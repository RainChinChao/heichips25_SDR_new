magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755684183
<< metal1 >>
rect 576 38576 99360 38600
rect 576 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 95072 38576
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95440 38536 99360 38576
rect 576 38512 99360 38536
rect 12739 38240 12797 38241
rect 12739 38200 12748 38240
rect 12788 38200 12797 38240
rect 12739 38199 12797 38200
rect 12067 37988 12125 37989
rect 12067 37948 12076 37988
rect 12116 37948 12125 37988
rect 12067 37947 12125 37948
rect 576 37820 99360 37844
rect 576 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 93832 37820
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 94200 37780 99360 37820
rect 576 37756 99360 37780
rect 13315 37652 13373 37653
rect 13315 37612 13324 37652
rect 13364 37612 13373 37652
rect 13315 37611 13373 37612
rect 18115 37484 18173 37485
rect 18115 37444 18124 37484
rect 18164 37444 18173 37484
rect 18115 37443 18173 37444
rect 25699 37484 25757 37485
rect 25699 37444 25708 37484
rect 25748 37444 25757 37484
rect 25699 37443 25757 37444
rect 26763 37484 26805 37493
rect 26763 37444 26764 37484
rect 26804 37444 26805 37484
rect 26763 37435 26805 37444
rect 39811 37484 39869 37485
rect 39811 37444 39820 37484
rect 39860 37444 39869 37484
rect 39811 37443 39869 37444
rect 11299 37400 11357 37401
rect 11299 37360 11308 37400
rect 11348 37360 11357 37400
rect 11299 37359 11357 37360
rect 12163 37400 12221 37401
rect 12163 37360 12172 37400
rect 12212 37360 12221 37400
rect 12163 37359 12221 37360
rect 19459 37400 19517 37401
rect 19459 37360 19468 37400
rect 19508 37360 19517 37400
rect 19459 37359 19517 37360
rect 22147 37400 22205 37401
rect 22147 37360 22156 37400
rect 22196 37360 22205 37400
rect 22147 37359 22205 37360
rect 22531 37400 22589 37401
rect 22531 37360 22540 37400
rect 22580 37360 22589 37400
rect 22531 37359 22589 37360
rect 27427 37400 27485 37401
rect 27427 37360 27436 37400
rect 27476 37360 27485 37400
rect 27427 37359 27485 37360
rect 39331 37400 39389 37401
rect 39331 37360 39340 37400
rect 39380 37360 39389 37400
rect 39331 37359 39389 37360
rect 40675 37400 40733 37401
rect 40675 37360 40684 37400
rect 40724 37360 40733 37400
rect 40675 37359 40733 37360
rect 10923 37316 10965 37325
rect 10923 37276 10924 37316
rect 10964 37276 10965 37316
rect 10923 37267 10965 37276
rect 17931 37232 17973 37241
rect 17931 37192 17932 37232
rect 17972 37192 17973 37232
rect 17931 37183 17973 37192
rect 18787 37232 18845 37233
rect 18787 37192 18796 37232
rect 18836 37192 18845 37232
rect 18787 37191 18845 37192
rect 22635 37232 22677 37241
rect 22635 37192 22636 37232
rect 22676 37192 22677 37232
rect 22635 37183 22677 37192
rect 25515 37232 25557 37241
rect 25515 37192 25516 37232
rect 25556 37192 25557 37232
rect 25515 37183 25557 37192
rect 38659 37232 38717 37233
rect 38659 37192 38668 37232
rect 38708 37192 38717 37232
rect 38659 37191 38717 37192
rect 39627 37232 39669 37241
rect 39627 37192 39628 37232
rect 39668 37192 39669 37232
rect 39627 37183 39669 37192
rect 40003 37232 40061 37233
rect 40003 37192 40012 37232
rect 40052 37192 40061 37232
rect 40003 37191 40061 37192
rect 576 37064 99360 37088
rect 576 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 95072 37064
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95440 37024 99360 37064
rect 576 37000 99360 37024
rect 10731 36896 10773 36905
rect 10731 36856 10732 36896
rect 10772 36856 10773 36896
rect 10731 36847 10773 36856
rect 19171 36896 19229 36897
rect 19171 36856 19180 36896
rect 19220 36856 19229 36896
rect 19171 36855 19229 36856
rect 27523 36896 27581 36897
rect 27523 36856 27532 36896
rect 27572 36856 27581 36896
rect 27523 36855 27581 36856
rect 39523 36896 39581 36897
rect 39523 36856 39532 36896
rect 39572 36856 39581 36896
rect 39523 36855 39581 36856
rect 42115 36896 42173 36897
rect 42115 36856 42124 36896
rect 42164 36856 42173 36896
rect 42115 36855 42173 36856
rect 16779 36812 16821 36821
rect 16779 36772 16780 36812
rect 16820 36772 16821 36812
rect 16779 36763 16821 36772
rect 21867 36812 21909 36821
rect 21867 36772 21868 36812
rect 21908 36772 21909 36812
rect 21867 36763 21909 36772
rect 25131 36812 25173 36821
rect 25131 36772 25132 36812
rect 25172 36772 25173 36812
rect 25131 36763 25173 36772
rect 39723 36812 39765 36821
rect 39723 36772 39724 36812
rect 39764 36772 39765 36812
rect 39723 36763 39765 36772
rect 7939 36728 7997 36729
rect 7939 36688 7948 36728
rect 7988 36688 7997 36728
rect 7939 36687 7997 36688
rect 10923 36728 10965 36737
rect 10923 36688 10924 36728
rect 10964 36688 10965 36728
rect 10923 36679 10965 36688
rect 11299 36728 11357 36729
rect 11299 36688 11308 36728
rect 11348 36688 11357 36728
rect 11299 36687 11357 36688
rect 12163 36728 12221 36729
rect 12163 36688 12172 36728
rect 12212 36688 12221 36728
rect 12163 36687 12221 36688
rect 17155 36728 17213 36729
rect 17155 36688 17164 36728
rect 17204 36688 17213 36728
rect 17155 36687 17213 36688
rect 18019 36728 18077 36729
rect 18019 36688 18028 36728
rect 18068 36688 18077 36728
rect 18019 36687 18077 36688
rect 22243 36728 22301 36729
rect 22243 36688 22252 36728
rect 22292 36688 22301 36728
rect 22243 36687 22301 36688
rect 23107 36728 23165 36729
rect 23107 36688 23116 36728
rect 23156 36688 23165 36728
rect 23107 36687 23165 36688
rect 25507 36728 25565 36729
rect 25507 36688 25516 36728
rect 25556 36688 25565 36728
rect 25507 36687 25565 36688
rect 26371 36728 26429 36729
rect 26371 36688 26380 36728
rect 26420 36688 26429 36728
rect 26371 36687 26429 36688
rect 29635 36728 29693 36729
rect 29635 36688 29644 36728
rect 29684 36688 29693 36728
rect 29635 36687 29693 36688
rect 35779 36728 35837 36729
rect 35779 36688 35788 36728
rect 35828 36688 35837 36728
rect 35779 36687 35837 36688
rect 37131 36728 37173 36737
rect 37131 36688 37132 36728
rect 37172 36688 37173 36728
rect 37131 36679 37173 36688
rect 37507 36728 37565 36729
rect 37507 36688 37516 36728
rect 37556 36688 37565 36728
rect 37507 36687 37565 36688
rect 38371 36728 38429 36729
rect 38371 36688 38380 36728
rect 38420 36688 38429 36728
rect 38371 36687 38429 36688
rect 40099 36728 40157 36729
rect 40099 36688 40108 36728
rect 40148 36688 40157 36728
rect 40099 36687 40157 36688
rect 40963 36728 41021 36729
rect 40963 36688 40972 36728
rect 41012 36688 41021 36728
rect 40963 36687 41021 36688
rect 10531 36644 10589 36645
rect 10531 36604 10540 36644
rect 10580 36604 10589 36644
rect 10531 36603 10589 36604
rect 34339 36644 34397 36645
rect 34339 36604 34348 36644
rect 34388 36604 34397 36644
rect 34339 36603 34397 36604
rect 7267 36560 7325 36561
rect 7267 36520 7276 36560
rect 7316 36520 7325 36560
rect 7267 36519 7325 36520
rect 13315 36560 13373 36561
rect 13315 36520 13324 36560
rect 13364 36520 13373 36560
rect 13315 36519 13373 36520
rect 34155 36560 34197 36569
rect 34155 36520 34156 36560
rect 34196 36520 34197 36560
rect 34155 36511 34197 36520
rect 35107 36560 35165 36561
rect 35107 36520 35116 36560
rect 35156 36520 35165 36560
rect 35107 36519 35165 36520
rect 24259 36476 24317 36477
rect 24259 36436 24268 36476
rect 24308 36436 24317 36476
rect 24259 36435 24317 36436
rect 28963 36476 29021 36477
rect 28963 36436 28972 36476
rect 29012 36436 29021 36476
rect 28963 36435 29021 36436
rect 576 36308 99360 36332
rect 576 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 93832 36308
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 94200 36268 99360 36308
rect 576 36244 99360 36268
rect 8131 36140 8189 36141
rect 8131 36100 8140 36140
rect 8180 36100 8189 36140
rect 8131 36099 8189 36100
rect 10827 36140 10869 36149
rect 10827 36100 10828 36140
rect 10868 36100 10869 36140
rect 10827 36091 10869 36100
rect 21867 36140 21909 36149
rect 21867 36100 21868 36140
rect 21908 36100 21909 36140
rect 21867 36091 21909 36100
rect 26283 36140 26325 36149
rect 26283 36100 26284 36140
rect 26324 36100 26325 36140
rect 26283 36091 26325 36100
rect 30211 36140 30269 36141
rect 30211 36100 30220 36140
rect 30260 36100 30269 36140
rect 30211 36099 30269 36100
rect 35587 36140 35645 36141
rect 35587 36100 35596 36140
rect 35636 36100 35645 36140
rect 35587 36099 35645 36100
rect 37419 36140 37461 36149
rect 37419 36100 37420 36140
rect 37460 36100 37461 36140
rect 37419 36091 37461 36100
rect 11011 35972 11069 35973
rect 11011 35932 11020 35972
rect 11060 35932 11069 35972
rect 11011 35931 11069 35932
rect 18219 35972 18261 35981
rect 18219 35932 18220 35972
rect 18260 35932 18261 35972
rect 18219 35923 18261 35932
rect 27427 35972 27485 35973
rect 27427 35932 27436 35972
rect 27476 35932 27485 35972
rect 27427 35931 27485 35932
rect 37603 35972 37661 35973
rect 37603 35932 37612 35972
rect 37652 35932 37661 35972
rect 37603 35931 37661 35932
rect 6115 35888 6173 35889
rect 6115 35848 6124 35888
rect 6164 35848 6173 35888
rect 6115 35847 6173 35848
rect 6979 35888 7037 35889
rect 6979 35848 6988 35888
rect 7028 35848 7037 35888
rect 6979 35847 7037 35848
rect 10435 35888 10493 35889
rect 10435 35848 10444 35888
rect 10484 35848 10493 35888
rect 10435 35847 10493 35848
rect 10635 35888 10677 35897
rect 10635 35848 10636 35888
rect 10676 35848 10677 35888
rect 10635 35839 10677 35848
rect 11875 35888 11933 35889
rect 11875 35848 11884 35888
rect 11924 35848 11933 35888
rect 11875 35847 11933 35848
rect 16195 35888 16253 35889
rect 16195 35848 16204 35888
rect 16244 35848 16253 35888
rect 16195 35847 16253 35848
rect 17059 35888 17117 35889
rect 17059 35848 17068 35888
rect 17108 35848 17117 35888
rect 17059 35847 17117 35848
rect 19075 35888 19133 35889
rect 19075 35848 19084 35888
rect 19124 35848 19133 35888
rect 19075 35847 19133 35848
rect 21771 35888 21813 35897
rect 21771 35848 21772 35888
rect 21812 35848 21813 35888
rect 21771 35839 21813 35848
rect 21955 35888 22013 35889
rect 21955 35848 21964 35888
rect 22004 35848 22013 35888
rect 21955 35847 22013 35848
rect 26179 35888 26237 35889
rect 26179 35848 26188 35888
rect 26228 35848 26237 35888
rect 26179 35847 26237 35848
rect 26379 35888 26421 35897
rect 26379 35848 26380 35888
rect 26420 35848 26421 35888
rect 26379 35839 26421 35848
rect 28195 35888 28253 35889
rect 28195 35848 28204 35888
rect 28244 35848 28253 35888
rect 28195 35847 28253 35848
rect 29059 35888 29117 35889
rect 29059 35848 29068 35888
rect 29108 35848 29117 35888
rect 29059 35847 29117 35848
rect 33195 35888 33237 35897
rect 33195 35848 33196 35888
rect 33236 35848 33237 35888
rect 33195 35839 33237 35848
rect 33571 35888 33629 35889
rect 33571 35848 33580 35888
rect 33620 35848 33629 35888
rect 33571 35847 33629 35848
rect 34435 35888 34493 35889
rect 34435 35848 34444 35888
rect 34484 35848 34493 35888
rect 34435 35847 34493 35848
rect 39619 35888 39677 35889
rect 39619 35848 39628 35888
rect 39668 35848 39677 35888
rect 39619 35847 39677 35848
rect 39819 35888 39861 35897
rect 39819 35848 39820 35888
rect 39860 35848 39861 35888
rect 39819 35839 39861 35848
rect 5739 35804 5781 35813
rect 5739 35764 5740 35804
rect 5780 35764 5781 35804
rect 5739 35755 5781 35764
rect 10539 35804 10581 35813
rect 10539 35764 10540 35804
rect 10580 35764 10581 35804
rect 10539 35755 10581 35764
rect 15819 35804 15861 35813
rect 15819 35764 15820 35804
rect 15860 35764 15861 35804
rect 15819 35755 15861 35764
rect 27819 35804 27861 35813
rect 27819 35764 27820 35804
rect 27860 35764 27861 35804
rect 27819 35755 27861 35764
rect 39723 35804 39765 35813
rect 39723 35764 39724 35804
rect 39764 35764 39765 35804
rect 39723 35755 39765 35764
rect 11203 35720 11261 35721
rect 11203 35680 11212 35720
rect 11252 35680 11261 35720
rect 11203 35679 11261 35680
rect 18403 35720 18461 35721
rect 18403 35680 18412 35720
rect 18452 35680 18461 35720
rect 18403 35679 18461 35680
rect 27627 35720 27669 35729
rect 27627 35680 27628 35720
rect 27668 35680 27669 35720
rect 27627 35671 27669 35680
rect 576 35552 99360 35576
rect 576 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 95072 35552
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95440 35512 99360 35552
rect 576 35488 99360 35512
rect 5931 35384 5973 35393
rect 5931 35344 5932 35384
rect 5972 35344 5973 35384
rect 5931 35335 5973 35344
rect 25795 35384 25853 35385
rect 25795 35344 25804 35384
rect 25844 35344 25853 35384
rect 25795 35343 25853 35344
rect 36931 35384 36989 35385
rect 36931 35344 36940 35384
rect 36980 35344 36989 35384
rect 36931 35343 36989 35344
rect 9003 35300 9045 35309
rect 9003 35260 9004 35300
rect 9044 35260 9045 35300
rect 9003 35251 9045 35260
rect 39523 35300 39581 35301
rect 39523 35260 39532 35300
rect 39572 35260 39581 35300
rect 39523 35259 39581 35260
rect 6315 35216 6357 35225
rect 6315 35176 6316 35216
rect 6356 35176 6357 35216
rect 6315 35167 6357 35176
rect 6691 35216 6749 35217
rect 6691 35176 6700 35216
rect 6740 35176 6749 35216
rect 6691 35175 6749 35176
rect 7555 35216 7613 35217
rect 7555 35176 7564 35216
rect 7604 35176 7613 35216
rect 7555 35175 7613 35176
rect 8907 35216 8949 35225
rect 8907 35176 8908 35216
rect 8948 35176 8949 35216
rect 8907 35167 8949 35176
rect 9091 35216 9149 35217
rect 9091 35176 9100 35216
rect 9140 35176 9149 35216
rect 9091 35175 9149 35176
rect 20515 35216 20573 35217
rect 20515 35176 20524 35216
rect 20564 35176 20573 35216
rect 20515 35175 20573 35176
rect 21475 35216 21533 35217
rect 21475 35176 21484 35216
rect 21524 35176 21533 35216
rect 21475 35175 21533 35176
rect 25699 35216 25757 35217
rect 25699 35176 25708 35216
rect 25748 35176 25757 35216
rect 25699 35175 25757 35176
rect 33195 35216 33237 35225
rect 33195 35176 33196 35216
rect 33236 35176 33237 35216
rect 33195 35167 33237 35176
rect 33571 35216 33629 35217
rect 33571 35176 33580 35216
rect 33620 35176 33629 35216
rect 33571 35175 33629 35176
rect 34435 35216 34493 35217
rect 34435 35176 34444 35216
rect 34484 35176 34493 35216
rect 34435 35175 34493 35176
rect 35779 35216 35837 35217
rect 35779 35176 35788 35216
rect 35828 35176 35837 35216
rect 35779 35175 35837 35176
rect 36835 35216 36893 35217
rect 36835 35176 36844 35216
rect 36884 35176 36893 35216
rect 36835 35175 36893 35176
rect 37131 35216 37173 35225
rect 37131 35176 37132 35216
rect 37172 35176 37173 35216
rect 37131 35167 37173 35176
rect 37227 35216 37269 35225
rect 37227 35176 37228 35216
rect 37268 35176 37269 35216
rect 37227 35167 37269 35176
rect 37315 35216 37373 35217
rect 37315 35176 37324 35216
rect 37364 35176 37373 35216
rect 37315 35175 37373 35176
rect 39043 35216 39101 35217
rect 39043 35176 39052 35216
rect 39092 35176 39101 35216
rect 39043 35175 39101 35176
rect 39427 35216 39485 35217
rect 39427 35176 39436 35216
rect 39476 35176 39485 35216
rect 39427 35175 39485 35176
rect 6115 35132 6173 35133
rect 6115 35092 6124 35132
rect 6164 35092 6173 35132
rect 6115 35091 6173 35092
rect 17059 35132 17117 35133
rect 17059 35092 17068 35132
rect 17108 35092 17117 35132
rect 17059 35091 17117 35092
rect 35595 35132 35637 35141
rect 35595 35092 35596 35132
rect 35636 35092 35637 35132
rect 35595 35083 35637 35092
rect 16875 35048 16917 35057
rect 16875 35008 16876 35048
rect 16916 35008 16917 35048
rect 16875 34999 16917 35008
rect 8707 34964 8765 34965
rect 8707 34924 8716 34964
rect 8756 34924 8765 34964
rect 8707 34923 8765 34924
rect 21195 34964 21237 34973
rect 21195 34924 21196 34964
rect 21236 34924 21237 34964
rect 21195 34915 21237 34924
rect 25507 34964 25565 34965
rect 25507 34924 25516 34964
rect 25556 34924 25565 34964
rect 25507 34923 25565 34924
rect 36451 34964 36509 34965
rect 36451 34924 36460 34964
rect 36500 34924 36509 34964
rect 36451 34923 36509 34924
rect 36643 34964 36701 34965
rect 36643 34924 36652 34964
rect 36692 34924 36701 34964
rect 36643 34923 36701 34924
rect 576 34796 99360 34820
rect 576 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 93832 34796
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 94200 34756 99360 34796
rect 576 34732 99360 34756
rect 7179 34628 7221 34637
rect 7179 34588 7180 34628
rect 7220 34588 7221 34628
rect 7179 34579 7221 34588
rect 34155 34628 34197 34637
rect 34155 34588 34156 34628
rect 34196 34588 34197 34628
rect 34155 34579 34197 34588
rect 12459 34544 12501 34553
rect 12459 34504 12460 34544
rect 12500 34504 12501 34544
rect 12459 34495 12501 34504
rect 7363 34460 7421 34461
rect 7363 34420 7372 34460
rect 7412 34420 7421 34460
rect 7363 34419 7421 34420
rect 23307 34460 23349 34469
rect 23307 34420 23308 34460
rect 23348 34420 23349 34460
rect 23307 34411 23349 34420
rect 34339 34460 34397 34461
rect 34339 34420 34348 34460
rect 34388 34420 34397 34460
rect 34339 34419 34397 34420
rect 8803 34376 8861 34377
rect 8803 34336 8812 34376
rect 8852 34336 8861 34376
rect 8803 34335 8861 34336
rect 9283 34376 9341 34377
rect 9283 34336 9292 34376
rect 9332 34336 9341 34376
rect 9283 34335 9341 34336
rect 9667 34376 9725 34377
rect 9667 34336 9676 34376
rect 9716 34336 9725 34376
rect 9667 34335 9725 34336
rect 10531 34376 10589 34377
rect 10531 34336 10540 34376
rect 10580 34336 10589 34376
rect 10531 34335 10589 34336
rect 11875 34376 11933 34377
rect 11875 34336 11884 34376
rect 11924 34336 11933 34376
rect 11875 34335 11933 34336
rect 12163 34376 12221 34377
rect 12163 34336 12172 34376
rect 12212 34336 12221 34376
rect 12163 34335 12221 34336
rect 13123 34376 13181 34377
rect 13123 34336 13132 34376
rect 13172 34336 13181 34376
rect 13123 34335 13181 34336
rect 21283 34376 21341 34377
rect 21283 34336 21292 34376
rect 21332 34336 21341 34376
rect 21283 34335 21341 34336
rect 22147 34376 22205 34377
rect 22147 34336 22156 34376
rect 22196 34336 22205 34376
rect 22147 34335 22205 34336
rect 24163 34376 24221 34377
rect 24163 34336 24172 34376
rect 24212 34336 24221 34376
rect 24163 34335 24221 34336
rect 24451 34376 24509 34377
rect 24451 34336 24460 34376
rect 24500 34336 24509 34376
rect 24451 34335 24509 34336
rect 25315 34376 25373 34377
rect 25315 34336 25324 34376
rect 25364 34336 25373 34376
rect 25315 34335 25373 34336
rect 26275 34376 26333 34377
rect 26275 34336 26284 34376
rect 26324 34336 26333 34376
rect 26275 34335 26333 34336
rect 20907 34292 20949 34301
rect 20907 34252 20908 34292
rect 20948 34252 20949 34292
rect 20907 34243 20949 34252
rect 8131 34208 8189 34209
rect 8131 34168 8140 34208
rect 8180 34168 8189 34208
rect 8131 34167 8189 34168
rect 9771 34208 9813 34217
rect 9771 34168 9772 34208
rect 9812 34168 9813 34208
rect 9771 34159 9813 34168
rect 10435 34208 10493 34209
rect 10435 34168 10444 34208
rect 10484 34168 10493 34208
rect 10435 34167 10493 34168
rect 10723 34208 10781 34209
rect 10723 34168 10732 34208
rect 10772 34168 10781 34208
rect 10723 34167 10781 34168
rect 24651 34208 24693 34217
rect 24651 34168 24652 34208
rect 24692 34168 24693 34208
rect 24651 34159 24693 34168
rect 576 34040 99360 34064
rect 576 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 95072 34040
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95440 34000 99360 34040
rect 576 33976 99360 34000
rect 6699 33872 6741 33881
rect 6699 33832 6700 33872
rect 6740 33832 6741 33872
rect 6699 33823 6741 33832
rect 19179 33872 19221 33881
rect 19179 33832 19180 33872
rect 19220 33832 19221 33872
rect 19179 33823 19221 33832
rect 18411 33788 18453 33797
rect 18411 33748 18412 33788
rect 18452 33748 18453 33788
rect 18411 33739 18453 33748
rect 25707 33788 25749 33797
rect 25707 33748 25708 33788
rect 25748 33748 25749 33788
rect 25707 33739 25749 33748
rect 40299 33788 40341 33797
rect 40299 33748 40300 33788
rect 40340 33748 40341 33788
rect 40299 33739 40341 33748
rect 7171 33704 7229 33705
rect 7171 33664 7180 33704
rect 7220 33664 7229 33704
rect 7171 33663 7229 33664
rect 17059 33704 17117 33705
rect 17059 33664 17068 33704
rect 17108 33664 17117 33704
rect 17059 33663 17117 33664
rect 18315 33704 18357 33713
rect 18315 33664 18316 33704
rect 18356 33664 18357 33704
rect 18315 33655 18357 33664
rect 18499 33704 18557 33705
rect 18499 33664 18508 33704
rect 18548 33664 18557 33704
rect 18499 33663 18557 33664
rect 18691 33704 18749 33705
rect 18691 33664 18700 33704
rect 18740 33664 18749 33704
rect 18691 33663 18749 33664
rect 18979 33704 19037 33705
rect 18979 33664 18988 33704
rect 19028 33664 19037 33704
rect 18979 33663 19037 33664
rect 25315 33704 25373 33705
rect 25315 33664 25324 33704
rect 25364 33664 25373 33704
rect 25315 33663 25373 33664
rect 26083 33704 26141 33705
rect 26083 33664 26092 33704
rect 26132 33664 26141 33704
rect 26083 33663 26141 33664
rect 26947 33704 27005 33705
rect 26947 33664 26956 33704
rect 26996 33664 27005 33704
rect 26947 33663 27005 33664
rect 40675 33704 40733 33705
rect 40675 33664 40684 33704
rect 40724 33664 40733 33704
rect 40675 33663 40733 33664
rect 41539 33704 41597 33705
rect 41539 33664 41548 33704
rect 41588 33664 41597 33704
rect 41539 33663 41597 33664
rect 6315 33620 6357 33629
rect 6315 33580 6316 33620
rect 6356 33580 6357 33620
rect 6315 33571 6357 33580
rect 15715 33620 15773 33621
rect 15715 33580 15724 33620
rect 15764 33580 15773 33620
rect 15715 33579 15773 33580
rect 15531 33452 15573 33461
rect 15531 33412 15532 33452
rect 15572 33412 15573 33452
rect 15531 33403 15573 33412
rect 16387 33452 16445 33453
rect 16387 33412 16396 33452
rect 16436 33412 16445 33452
rect 16387 33411 16445 33412
rect 28099 33452 28157 33453
rect 28099 33412 28108 33452
rect 28148 33412 28157 33452
rect 28099 33411 28157 33412
rect 42691 33452 42749 33453
rect 42691 33412 42700 33452
rect 42740 33412 42749 33452
rect 42691 33411 42749 33412
rect 576 33284 99360 33308
rect 576 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 18232 33284
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18600 33244 33352 33284
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33720 33244 48472 33284
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48840 33244 63592 33284
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63960 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 93832 33284
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 94200 33244 99360 33284
rect 576 33220 99360 33244
rect 16867 33116 16925 33117
rect 16867 33076 16876 33116
rect 16916 33076 16925 33116
rect 16867 33075 16925 33076
rect 4099 32864 4157 32865
rect 4099 32824 4108 32864
rect 4148 32824 4157 32864
rect 4099 32823 4157 32824
rect 14475 32864 14517 32873
rect 14475 32824 14476 32864
rect 14516 32824 14517 32864
rect 14475 32815 14517 32824
rect 14851 32864 14909 32865
rect 14851 32824 14860 32864
rect 14900 32824 14909 32864
rect 14851 32823 14909 32824
rect 15715 32864 15773 32865
rect 15715 32824 15724 32864
rect 15764 32824 15773 32864
rect 15715 32823 15773 32824
rect 18027 32864 18069 32873
rect 18027 32824 18028 32864
rect 18068 32824 18069 32864
rect 18027 32815 18069 32824
rect 18211 32864 18269 32865
rect 18211 32824 18220 32864
rect 18260 32824 18269 32864
rect 18211 32823 18269 32824
rect 27235 32864 27293 32865
rect 27235 32824 27244 32864
rect 27284 32824 27293 32864
rect 27235 32823 27293 32824
rect 27427 32864 27485 32865
rect 27427 32824 27436 32864
rect 27476 32824 27485 32864
rect 27427 32823 27485 32824
rect 3435 32780 3477 32789
rect 3435 32740 3436 32780
rect 3476 32740 3477 32780
rect 3435 32731 3477 32740
rect 18123 32780 18165 32789
rect 18123 32740 18124 32780
rect 18164 32740 18165 32780
rect 18123 32731 18165 32740
rect 26571 32780 26613 32789
rect 26571 32740 26572 32780
rect 26612 32740 26613 32780
rect 26571 32731 26613 32740
rect 28099 32696 28157 32697
rect 28099 32656 28108 32696
rect 28148 32656 28157 32696
rect 28099 32655 28157 32656
rect 576 32528 99360 32552
rect 576 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 19472 32528
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19840 32488 34592 32528
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34960 32488 49712 32528
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 50080 32488 64832 32528
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 65200 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 95072 32528
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95440 32488 99360 32528
rect 576 32464 99360 32488
rect 4291 32360 4349 32361
rect 4291 32320 4300 32360
rect 4340 32320 4349 32360
rect 4291 32319 4349 32320
rect 10059 32360 10101 32369
rect 10059 32320 10060 32360
rect 10100 32320 10101 32360
rect 10059 32311 10101 32320
rect 26571 32360 26613 32369
rect 26571 32320 26572 32360
rect 26612 32320 26613 32360
rect 26571 32311 26613 32320
rect 11019 32276 11061 32285
rect 11019 32236 11020 32276
rect 11060 32236 11061 32276
rect 11019 32227 11061 32236
rect 28107 32276 28149 32285
rect 28107 32236 28108 32276
rect 28148 32236 28149 32276
rect 28107 32227 28149 32236
rect 35499 32276 35541 32285
rect 35499 32236 35500 32276
rect 35540 32236 35541 32276
rect 35499 32227 35541 32236
rect 42883 32276 42941 32277
rect 42883 32236 42892 32276
rect 42932 32236 42941 32276
rect 42883 32235 42941 32236
rect 1899 32192 1941 32201
rect 1899 32152 1900 32192
rect 1940 32152 1941 32192
rect 1899 32143 1941 32152
rect 2275 32192 2333 32193
rect 2275 32152 2284 32192
rect 2324 32152 2333 32192
rect 2275 32151 2333 32152
rect 3139 32192 3197 32193
rect 3139 32152 3148 32192
rect 3188 32152 3197 32192
rect 3139 32151 3197 32152
rect 10443 32192 10485 32201
rect 10443 32152 10444 32192
rect 10484 32152 10485 32192
rect 10443 32143 10485 32152
rect 11395 32192 11453 32193
rect 11395 32152 11404 32192
rect 11444 32152 11453 32192
rect 11395 32151 11453 32152
rect 12259 32192 12317 32193
rect 12259 32152 12268 32192
rect 12308 32152 12317 32192
rect 12259 32151 12317 32152
rect 19843 32192 19901 32193
rect 19843 32152 19852 32192
rect 19892 32152 19901 32192
rect 19843 32151 19901 32152
rect 26187 32192 26229 32201
rect 26187 32152 26188 32192
rect 26228 32152 26229 32192
rect 26187 32143 26229 32152
rect 26275 32192 26333 32193
rect 26275 32152 26284 32192
rect 26324 32152 26333 32192
rect 26275 32151 26333 32152
rect 28483 32192 28541 32193
rect 28483 32152 28492 32192
rect 28532 32152 28541 32192
rect 28483 32151 28541 32152
rect 29347 32192 29405 32193
rect 29347 32152 29356 32192
rect 29396 32152 29405 32192
rect 29347 32151 29405 32152
rect 35875 32192 35933 32193
rect 35875 32152 35884 32192
rect 35924 32152 35933 32192
rect 35875 32151 35933 32152
rect 36739 32192 36797 32193
rect 36739 32152 36748 32192
rect 36788 32152 36797 32192
rect 36739 32151 36797 32152
rect 38371 32192 38429 32193
rect 38371 32152 38380 32192
rect 38420 32152 38429 32192
rect 38371 32151 38429 32152
rect 38475 32192 38517 32201
rect 38475 32152 38476 32192
rect 38516 32152 38517 32192
rect 38475 32143 38517 32152
rect 42979 32192 43037 32193
rect 42979 32152 42988 32192
rect 43028 32152 43037 32192
rect 42979 32151 43037 32152
rect 43363 32192 43421 32193
rect 43363 32152 43372 32192
rect 43412 32152 43421 32192
rect 43363 32151 43421 32152
rect 48931 32192 48989 32193
rect 48931 32152 48940 32192
rect 48980 32152 48989 32192
rect 48931 32151 48989 32152
rect 18211 32108 18269 32109
rect 18211 32068 18220 32108
rect 18260 32068 18269 32108
rect 18211 32067 18269 32068
rect 13411 31940 13469 31941
rect 13411 31900 13420 31940
rect 13460 31900 13469 31940
rect 13411 31899 13469 31900
rect 18027 31940 18069 31949
rect 18027 31900 18028 31940
rect 18068 31900 18069 31940
rect 18027 31891 18069 31900
rect 19171 31940 19229 31941
rect 19171 31900 19180 31940
rect 19220 31900 19229 31940
rect 19171 31899 19229 31900
rect 30499 31940 30557 31941
rect 30499 31900 30508 31940
rect 30548 31900 30557 31940
rect 30499 31899 30557 31900
rect 37891 31940 37949 31941
rect 37891 31900 37900 31940
rect 37940 31900 37949 31940
rect 37891 31899 37949 31900
rect 38187 31940 38229 31949
rect 38187 31900 38188 31940
rect 38228 31900 38229 31940
rect 38187 31891 38229 31900
rect 48259 31940 48317 31941
rect 48259 31900 48268 31940
rect 48308 31900 48317 31940
rect 48259 31899 48317 31900
rect 576 31772 99360 31796
rect 576 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 18232 31772
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18600 31732 33352 31772
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33720 31732 48472 31772
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48840 31732 63592 31772
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63960 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 93832 31772
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 94200 31732 99360 31772
rect 576 31708 99360 31732
rect 2187 31604 2229 31613
rect 2187 31564 2188 31604
rect 2228 31564 2229 31604
rect 2187 31555 2229 31564
rect 19843 31604 19901 31605
rect 19843 31564 19852 31604
rect 19892 31564 19901 31604
rect 19843 31563 19901 31564
rect 23115 31604 23157 31613
rect 23115 31564 23116 31604
rect 23156 31564 23157 31604
rect 23115 31555 23157 31564
rect 26283 31604 26325 31613
rect 26283 31564 26284 31604
rect 26324 31564 26325 31604
rect 26283 31555 26325 31564
rect 49507 31520 49565 31521
rect 49507 31480 49516 31520
rect 49556 31480 49565 31520
rect 49507 31479 49565 31480
rect 2371 31436 2429 31437
rect 2371 31396 2380 31436
rect 2420 31396 2429 31436
rect 2371 31395 2429 31396
rect 41547 31436 41589 31445
rect 41547 31396 41548 31436
rect 41588 31396 41589 31436
rect 41547 31387 41589 31396
rect 46723 31436 46781 31437
rect 46723 31396 46732 31436
rect 46772 31396 46781 31436
rect 46723 31395 46781 31396
rect 2947 31352 3005 31353
rect 2947 31312 2956 31352
rect 2996 31312 3005 31352
rect 2947 31311 3005 31312
rect 3811 31352 3869 31353
rect 3811 31312 3820 31352
rect 3860 31312 3869 31352
rect 3811 31311 3869 31312
rect 9291 31352 9333 31361
rect 9291 31312 9292 31352
rect 9332 31312 9333 31352
rect 9291 31303 9333 31312
rect 9667 31352 9725 31353
rect 9667 31312 9676 31352
rect 9716 31312 9725 31352
rect 9667 31311 9725 31312
rect 10531 31352 10589 31353
rect 10531 31312 10540 31352
rect 10580 31312 10589 31352
rect 10531 31311 10589 31312
rect 17451 31352 17493 31361
rect 17451 31312 17452 31352
rect 17492 31312 17493 31352
rect 17451 31303 17493 31312
rect 17827 31352 17885 31353
rect 17827 31312 17836 31352
rect 17876 31312 17885 31352
rect 17827 31311 17885 31312
rect 18691 31352 18749 31353
rect 18691 31312 18700 31352
rect 18740 31312 18749 31352
rect 18691 31311 18749 31312
rect 20131 31352 20189 31353
rect 20131 31312 20140 31352
rect 20180 31312 20189 31352
rect 20131 31311 20189 31312
rect 23307 31352 23349 31361
rect 23307 31312 23308 31352
rect 23348 31312 23349 31352
rect 23307 31303 23349 31312
rect 25315 31352 25373 31353
rect 25315 31312 25324 31352
rect 25364 31312 25373 31352
rect 25315 31311 25373 31312
rect 25995 31352 26037 31361
rect 25995 31312 25996 31352
rect 26036 31312 26037 31352
rect 25995 31303 26037 31312
rect 26179 31352 26237 31353
rect 26179 31312 26188 31352
rect 26228 31312 26237 31352
rect 26179 31311 26237 31312
rect 26379 31352 26421 31361
rect 26379 31312 26380 31352
rect 26420 31312 26421 31352
rect 26379 31303 26421 31312
rect 33475 31352 33533 31353
rect 33475 31312 33484 31352
rect 33524 31312 33533 31352
rect 33475 31311 33533 31312
rect 34339 31352 34397 31353
rect 34339 31312 34348 31352
rect 34388 31312 34397 31352
rect 34339 31311 34397 31312
rect 36931 31352 36989 31353
rect 36931 31312 36940 31352
rect 36980 31312 36989 31352
rect 36931 31311 36989 31312
rect 37123 31352 37181 31353
rect 37123 31312 37132 31352
rect 37172 31312 37181 31352
rect 37123 31311 37181 31312
rect 37987 31352 38045 31353
rect 37987 31312 37996 31352
rect 38036 31312 38045 31352
rect 37987 31311 38045 31312
rect 42403 31352 42461 31353
rect 42403 31312 42412 31352
rect 42452 31312 42461 31352
rect 42403 31311 42461 31312
rect 47491 31352 47549 31353
rect 47491 31312 47500 31352
rect 47540 31312 47549 31352
rect 47491 31311 47549 31312
rect 48355 31352 48413 31353
rect 48355 31312 48364 31352
rect 48404 31312 48413 31352
rect 48355 31311 48413 31312
rect 50947 31352 51005 31353
rect 50947 31312 50956 31352
rect 50996 31312 51005 31352
rect 50947 31311 51005 31312
rect 2571 31268 2613 31277
rect 2571 31228 2572 31268
rect 2612 31228 2613 31268
rect 2571 31219 2613 31228
rect 34731 31268 34773 31277
rect 34731 31228 34732 31268
rect 34772 31228 34773 31268
rect 34731 31219 34773 31228
rect 36267 31268 36309 31277
rect 36267 31228 36268 31268
rect 36308 31228 36309 31268
rect 36267 31219 36309 31228
rect 47115 31268 47157 31277
rect 47115 31228 47116 31268
rect 47156 31228 47157 31268
rect 47115 31219 47157 31228
rect 4963 31184 5021 31185
rect 4963 31144 4972 31184
rect 5012 31144 5021 31184
rect 4963 31143 5021 31144
rect 11683 31184 11741 31185
rect 11683 31144 11692 31184
rect 11732 31144 11741 31184
rect 11683 31143 11741 31144
rect 20035 31184 20093 31185
rect 20035 31144 20044 31184
rect 20084 31144 20093 31184
rect 20035 31143 20093 31144
rect 20323 31184 20381 31185
rect 20323 31144 20332 31184
rect 20372 31144 20381 31184
rect 20323 31143 20381 31144
rect 32323 31184 32381 31185
rect 32323 31144 32332 31184
rect 32372 31144 32381 31184
rect 32323 31143 32381 31144
rect 37795 31184 37853 31185
rect 37795 31144 37804 31184
rect 37844 31144 37853 31184
rect 37795 31143 37853 31144
rect 38659 31184 38717 31185
rect 38659 31144 38668 31184
rect 38708 31144 38717 31184
rect 38659 31143 38717 31144
rect 41931 31184 41973 31193
rect 41931 31144 41932 31184
rect 41972 31144 41973 31184
rect 41931 31135 41973 31144
rect 46923 31184 46965 31193
rect 46923 31144 46924 31184
rect 46964 31144 46965 31184
rect 46923 31135 46965 31144
rect 50275 31184 50333 31185
rect 50275 31144 50284 31184
rect 50324 31144 50333 31184
rect 50275 31143 50333 31144
rect 576 31016 99360 31040
rect 576 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 19472 31016
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19840 30976 34592 31016
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34960 30976 49712 31016
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 50080 30976 64832 31016
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 65200 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 95072 31016
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95440 30976 99360 31016
rect 576 30952 99360 30976
rect 3339 30848 3381 30857
rect 3339 30808 3340 30848
rect 3380 30808 3381 30848
rect 3339 30799 3381 30808
rect 25987 30848 26045 30849
rect 25987 30808 25996 30848
rect 26036 30808 26045 30848
rect 25987 30807 26045 30808
rect 35019 30848 35061 30857
rect 35019 30808 35020 30848
rect 35060 30808 35061 30848
rect 35019 30799 35061 30808
rect 37027 30848 37085 30849
rect 37027 30808 37036 30848
rect 37076 30808 37085 30848
rect 37027 30807 37085 30808
rect 42307 30848 42365 30849
rect 42307 30808 42316 30848
rect 42356 30808 42365 30848
rect 42307 30807 42365 30808
rect 48939 30848 48981 30857
rect 48939 30808 48940 30848
rect 48980 30808 48981 30848
rect 48939 30799 48981 30808
rect 51523 30848 51581 30849
rect 51523 30808 51532 30848
rect 51572 30808 51581 30848
rect 51523 30807 51581 30808
rect 21963 30764 22005 30773
rect 21963 30724 21964 30764
rect 22004 30724 22005 30764
rect 21963 30715 22005 30724
rect 26947 30764 27005 30765
rect 26947 30724 26956 30764
rect 26996 30724 27005 30764
rect 26947 30723 27005 30724
rect 31075 30764 31133 30765
rect 31075 30724 31084 30764
rect 31124 30724 31133 30764
rect 31075 30723 31133 30724
rect 41155 30764 41213 30765
rect 41155 30724 41164 30764
rect 41204 30724 41213 30764
rect 41155 30723 41213 30724
rect 49131 30764 49173 30773
rect 49131 30724 49132 30764
rect 49172 30724 49173 30764
rect 49131 30715 49173 30724
rect 4011 30680 4053 30689
rect 4011 30640 4012 30680
rect 4052 30640 4053 30680
rect 4011 30631 4053 30640
rect 4195 30680 4253 30681
rect 4195 30640 4204 30680
rect 4244 30640 4253 30680
rect 4195 30639 4253 30640
rect 5059 30680 5117 30681
rect 5059 30640 5068 30680
rect 5108 30640 5117 30680
rect 5059 30639 5117 30640
rect 7275 30680 7317 30689
rect 7275 30640 7276 30680
rect 7316 30640 7317 30680
rect 7275 30631 7317 30640
rect 7651 30680 7709 30681
rect 7651 30640 7660 30680
rect 7700 30640 7709 30680
rect 7651 30639 7709 30640
rect 8515 30680 8573 30681
rect 8515 30640 8524 30680
rect 8564 30640 8573 30680
rect 8515 30639 8573 30640
rect 13507 30680 13565 30681
rect 13507 30640 13516 30680
rect 13556 30640 13565 30680
rect 13507 30639 13565 30640
rect 17547 30680 17589 30689
rect 17547 30640 17548 30680
rect 17588 30640 17589 30680
rect 17547 30631 17589 30640
rect 17923 30680 17981 30681
rect 17923 30640 17932 30680
rect 17972 30640 17981 30680
rect 17923 30639 17981 30640
rect 18787 30680 18845 30681
rect 18787 30640 18796 30680
rect 18836 30640 18845 30680
rect 18787 30639 18845 30640
rect 22339 30680 22397 30681
rect 22339 30640 22348 30680
rect 22388 30640 22397 30680
rect 22339 30639 22397 30640
rect 23203 30680 23261 30681
rect 23203 30640 23212 30680
rect 23252 30640 23261 30680
rect 23203 30639 23261 30640
rect 25795 30680 25853 30681
rect 25795 30640 25804 30680
rect 25844 30640 25853 30680
rect 25795 30639 25853 30640
rect 26659 30680 26717 30681
rect 26659 30640 26668 30680
rect 26708 30640 26717 30680
rect 26659 30639 26717 30640
rect 27043 30680 27101 30681
rect 27043 30640 27052 30680
rect 27092 30640 27101 30680
rect 27043 30639 27101 30640
rect 27427 30680 27485 30681
rect 27427 30640 27436 30680
rect 27476 30640 27485 30680
rect 27427 30639 27485 30640
rect 30595 30680 30653 30681
rect 30595 30640 30604 30680
rect 30644 30640 30653 30680
rect 30595 30639 30653 30640
rect 30979 30680 31037 30681
rect 30979 30640 30988 30680
rect 31028 30640 31037 30680
rect 30979 30639 31037 30640
rect 34147 30680 34205 30681
rect 34147 30640 34156 30680
rect 34196 30640 34205 30680
rect 34147 30639 34205 30640
rect 34531 30680 34589 30681
rect 34531 30640 34540 30680
rect 34580 30640 34589 30680
rect 34531 30639 34589 30640
rect 36643 30680 36701 30681
rect 36643 30640 36652 30680
rect 36692 30640 36701 30680
rect 36643 30639 36701 30640
rect 38179 30680 38237 30681
rect 38179 30640 38188 30680
rect 38228 30640 38237 30680
rect 38179 30639 38237 30640
rect 39043 30680 39101 30681
rect 39043 30640 39052 30680
rect 39092 30640 39101 30680
rect 39043 30639 39101 30640
rect 39435 30680 39477 30689
rect 39435 30640 39436 30680
rect 39476 30640 39477 30680
rect 39435 30631 39477 30640
rect 42019 30680 42077 30681
rect 42019 30640 42028 30680
rect 42068 30640 42077 30680
rect 42019 30639 42077 30640
rect 43459 30680 43517 30681
rect 43459 30640 43468 30680
rect 43508 30640 43517 30680
rect 43459 30639 43517 30640
rect 44323 30680 44381 30681
rect 44323 30640 44332 30680
rect 44372 30640 44381 30680
rect 44323 30639 44381 30640
rect 44715 30680 44757 30689
rect 44715 30640 44716 30680
rect 44756 30640 44757 30680
rect 44715 30631 44757 30640
rect 46147 30680 46205 30681
rect 46147 30640 46156 30680
rect 46196 30640 46205 30680
rect 46147 30639 46205 30640
rect 48355 30680 48413 30681
rect 48355 30640 48364 30680
rect 48404 30640 48413 30680
rect 48355 30639 48413 30640
rect 48555 30680 48597 30689
rect 48555 30640 48556 30680
rect 48596 30640 48597 30680
rect 48555 30631 48597 30640
rect 49507 30680 49565 30681
rect 49507 30640 49516 30680
rect 49556 30640 49565 30680
rect 49507 30639 49565 30640
rect 50371 30680 50429 30681
rect 50371 30640 50380 30680
rect 50420 30640 50429 30680
rect 50371 30639 50429 30640
rect 3523 30596 3581 30597
rect 3523 30556 3532 30596
rect 3572 30556 3581 30596
rect 3523 30555 3581 30556
rect 24363 30596 24405 30605
rect 24363 30556 24364 30596
rect 24404 30556 24405 30596
rect 24363 30547 24405 30556
rect 48739 30596 48797 30597
rect 48739 30556 48748 30596
rect 48788 30556 48797 30596
rect 48739 30555 48797 30556
rect 4387 30512 4445 30513
rect 4387 30472 4396 30512
rect 4436 30472 4445 30512
rect 4387 30471 4445 30472
rect 4107 30428 4149 30437
rect 4107 30388 4108 30428
rect 4148 30388 4149 30428
rect 4107 30379 4149 30388
rect 9667 30428 9725 30429
rect 9667 30388 9676 30428
rect 9716 30388 9725 30428
rect 9667 30387 9725 30388
rect 14179 30428 14237 30429
rect 14179 30388 14188 30428
rect 14228 30388 14237 30428
rect 14179 30387 14237 30388
rect 19939 30428 19997 30429
rect 19939 30388 19948 30428
rect 19988 30388 19997 30428
rect 19939 30387 19997 30388
rect 25123 30428 25181 30429
rect 25123 30388 25132 30428
rect 25172 30388 25181 30428
rect 25123 30387 25181 30388
rect 25987 30428 26045 30429
rect 25987 30388 25996 30428
rect 26036 30388 26045 30428
rect 25987 30387 26045 30388
rect 35971 30428 36029 30429
rect 35971 30388 35980 30428
rect 36020 30388 36029 30428
rect 35971 30387 36029 30388
rect 48459 30428 48501 30437
rect 48459 30388 48460 30428
rect 48500 30388 48501 30428
rect 48459 30379 48501 30388
rect 576 30260 99360 30284
rect 576 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 18232 30260
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18600 30220 33352 30260
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33720 30220 48472 30260
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48840 30220 63592 30260
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63960 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 93832 30260
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 94200 30220 99360 30260
rect 576 30196 99360 30220
rect 16107 30092 16149 30101
rect 16107 30052 16108 30092
rect 16148 30052 16149 30092
rect 16107 30043 16149 30052
rect 17931 30092 17973 30101
rect 17931 30052 17932 30092
rect 17972 30052 17973 30092
rect 17931 30043 17973 30052
rect 19171 30092 19229 30093
rect 19171 30052 19180 30092
rect 19220 30052 19229 30092
rect 19171 30051 19229 30052
rect 37995 30092 38037 30101
rect 37995 30052 37996 30092
rect 38036 30052 38037 30092
rect 37995 30043 38037 30052
rect 43083 30092 43125 30101
rect 43083 30052 43084 30092
rect 43124 30052 43125 30092
rect 43083 30043 43125 30052
rect 45667 30092 45725 30093
rect 45667 30052 45676 30092
rect 45716 30052 45725 30092
rect 45667 30051 45725 30052
rect 46731 30092 46773 30101
rect 46731 30052 46732 30092
rect 46772 30052 46773 30092
rect 46731 30043 46773 30052
rect 18115 29924 18173 29925
rect 18115 29884 18124 29924
rect 18164 29884 18173 29924
rect 18115 29883 18173 29884
rect 5155 29840 5213 29841
rect 5155 29800 5164 29840
rect 5204 29800 5213 29840
rect 5155 29799 5213 29800
rect 5443 29840 5501 29841
rect 5443 29800 5452 29840
rect 5492 29800 5501 29840
rect 5443 29799 5501 29800
rect 11107 29840 11165 29841
rect 11107 29800 11116 29840
rect 11156 29800 11165 29840
rect 11107 29799 11165 29800
rect 11491 29840 11549 29841
rect 11491 29800 11500 29840
rect 11540 29800 11549 29840
rect 11491 29799 11549 29800
rect 15915 29840 15957 29849
rect 15915 29800 15916 29840
rect 15956 29800 15957 29840
rect 15915 29791 15957 29800
rect 19843 29840 19901 29841
rect 19843 29800 19852 29840
rect 19892 29800 19901 29840
rect 19843 29799 19901 29800
rect 25707 29840 25749 29849
rect 25707 29800 25708 29840
rect 25748 29800 25749 29840
rect 25707 29791 25749 29800
rect 26083 29840 26141 29841
rect 26083 29800 26092 29840
rect 26132 29800 26141 29840
rect 26083 29799 26141 29800
rect 26947 29840 27005 29841
rect 26947 29800 26956 29840
rect 26996 29800 27005 29840
rect 26947 29799 27005 29800
rect 28387 29840 28445 29841
rect 28387 29800 28396 29840
rect 28436 29800 28445 29840
rect 28387 29799 28445 29800
rect 37411 29840 37469 29841
rect 37411 29800 37420 29840
rect 37460 29800 37469 29840
rect 37411 29799 37469 29800
rect 37699 29840 37757 29841
rect 37699 29800 37708 29840
rect 37748 29800 37757 29840
rect 37699 29799 37757 29800
rect 37899 29840 37941 29849
rect 37899 29800 37900 29840
rect 37940 29800 37941 29840
rect 37899 29791 37941 29800
rect 38083 29840 38141 29841
rect 38083 29800 38092 29840
rect 38132 29800 38141 29840
rect 38083 29799 38141 29800
rect 42787 29840 42845 29841
rect 42787 29800 42796 29840
rect 42836 29800 42845 29840
rect 42787 29799 42845 29800
rect 45859 29840 45917 29841
rect 45859 29800 45868 29840
rect 45908 29800 45917 29840
rect 45859 29799 45917 29800
rect 46243 29840 46301 29841
rect 46243 29800 46252 29840
rect 46292 29800 46301 29840
rect 46243 29799 46301 29800
rect 47395 29840 47453 29841
rect 47395 29800 47404 29840
rect 47444 29800 47453 29840
rect 47395 29799 47453 29800
rect 47779 29840 47837 29841
rect 47779 29800 47788 29840
rect 47828 29800 47837 29840
rect 47779 29799 47837 29800
rect 5635 29756 5693 29757
rect 5635 29716 5644 29756
rect 5684 29716 5693 29756
rect 5635 29715 5693 29716
rect 37219 29756 37277 29757
rect 37219 29716 37228 29756
rect 37268 29716 37277 29756
rect 37219 29715 37277 29716
rect 47875 29756 47933 29757
rect 47875 29716 47884 29756
rect 47924 29716 47933 29756
rect 47875 29715 47933 29716
rect 11595 29672 11637 29681
rect 11595 29632 11596 29672
rect 11636 29632 11637 29672
rect 11595 29623 11637 29632
rect 28099 29672 28157 29673
rect 28099 29632 28108 29672
rect 28148 29632 28157 29672
rect 28099 29631 28157 29632
rect 29059 29672 29117 29673
rect 29059 29632 29068 29672
rect 29108 29632 29117 29672
rect 29059 29631 29117 29632
rect 43275 29672 43317 29681
rect 43275 29632 43276 29672
rect 43316 29632 43317 29672
rect 43275 29623 43317 29632
rect 45955 29672 46013 29673
rect 45955 29632 45964 29672
rect 46004 29632 46013 29672
rect 45955 29631 46013 29632
rect 576 29504 99360 29528
rect 576 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 19472 29504
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19840 29464 34592 29504
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34960 29464 49712 29504
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 50080 29464 64832 29504
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 65200 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 95072 29504
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95440 29464 99360 29504
rect 576 29440 99360 29464
rect 5163 29252 5205 29261
rect 5163 29212 5164 29252
rect 5204 29212 5205 29252
rect 5163 29203 5205 29212
rect 30411 29252 30453 29261
rect 30411 29212 30412 29252
rect 30452 29212 30453 29252
rect 30411 29203 30453 29212
rect 34539 29252 34581 29261
rect 34539 29212 34540 29252
rect 34580 29212 34581 29252
rect 34539 29203 34581 29212
rect 46923 29252 46965 29261
rect 46923 29212 46924 29252
rect 46964 29212 46965 29252
rect 46923 29203 46965 29212
rect 4867 29168 4925 29169
rect 4867 29128 4876 29168
rect 4916 29128 4925 29168
rect 4867 29127 4925 29128
rect 5067 29168 5109 29177
rect 5067 29128 5068 29168
rect 5108 29128 5109 29168
rect 5067 29119 5109 29128
rect 5251 29168 5309 29169
rect 5251 29128 5260 29168
rect 5300 29128 5309 29168
rect 5251 29127 5309 29128
rect 8803 29168 8861 29169
rect 8803 29128 8812 29168
rect 8852 29128 8861 29168
rect 8803 29127 8861 29128
rect 9763 29168 9821 29169
rect 9763 29128 9772 29168
rect 9812 29128 9821 29168
rect 9763 29127 9821 29128
rect 12363 29168 12405 29177
rect 12363 29128 12364 29168
rect 12404 29128 12405 29168
rect 12363 29119 12405 29128
rect 12451 29168 12509 29169
rect 12451 29128 12460 29168
rect 12500 29128 12509 29168
rect 12451 29127 12509 29128
rect 22147 29168 22205 29169
rect 22147 29128 22156 29168
rect 22196 29128 22205 29168
rect 22147 29127 22205 29128
rect 23019 29168 23061 29177
rect 23019 29128 23020 29168
rect 23060 29128 23061 29168
rect 23019 29119 23061 29128
rect 28491 29168 28533 29177
rect 28491 29128 28492 29168
rect 28532 29128 28533 29168
rect 28491 29119 28533 29128
rect 28675 29168 28733 29169
rect 28675 29128 28684 29168
rect 28724 29128 28733 29168
rect 28675 29127 28733 29128
rect 29155 29168 29213 29169
rect 29155 29128 29164 29168
rect 29204 29128 29213 29168
rect 29155 29127 29213 29128
rect 30115 29168 30173 29169
rect 30115 29128 30124 29168
rect 30164 29128 30173 29168
rect 30115 29127 30173 29128
rect 31075 29168 31133 29169
rect 31075 29128 31084 29168
rect 31124 29128 31133 29168
rect 31075 29127 31133 29128
rect 33283 29168 33341 29169
rect 33283 29128 33292 29168
rect 33332 29128 33341 29168
rect 33283 29127 33341 29128
rect 34147 29168 34205 29169
rect 34147 29128 34156 29168
rect 34196 29128 34205 29168
rect 34147 29127 34205 29128
rect 46819 29168 46877 29169
rect 46819 29128 46828 29168
rect 46868 29128 46877 29168
rect 46819 29127 46877 29128
rect 47019 29168 47061 29177
rect 47019 29128 47020 29168
rect 47060 29128 47061 29168
rect 47019 29119 47061 29128
rect 32139 29084 32181 29093
rect 32139 29044 32140 29084
rect 32180 29044 32181 29084
rect 32139 29035 32181 29044
rect 4195 29000 4253 29001
rect 4195 28960 4204 29000
rect 4244 28960 4253 29000
rect 4195 28959 4253 28960
rect 9483 29000 9525 29009
rect 9483 28960 9484 29000
rect 9524 28960 9525 29000
rect 9483 28951 9525 28960
rect 12651 28916 12693 28925
rect 12651 28876 12652 28916
rect 12692 28876 12693 28916
rect 12651 28867 12693 28876
rect 28587 28916 28629 28925
rect 28587 28876 28588 28916
rect 28628 28876 28629 28916
rect 28587 28867 28629 28876
rect 576 28748 99360 28772
rect 576 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 18232 28748
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18600 28708 33352 28748
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33720 28708 48472 28748
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48840 28708 63592 28748
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63960 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 93832 28748
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 94200 28708 99360 28748
rect 576 28684 99360 28708
rect 4675 28580 4733 28581
rect 4675 28540 4684 28580
rect 4724 28540 4733 28580
rect 4675 28539 4733 28540
rect 5835 28580 5877 28589
rect 5835 28540 5836 28580
rect 5876 28540 5877 28580
rect 5835 28531 5877 28540
rect 13035 28580 13077 28589
rect 13035 28540 13036 28580
rect 13076 28540 13077 28580
rect 13035 28531 13077 28540
rect 44899 28412 44957 28413
rect 44899 28372 44908 28412
rect 44948 28372 44957 28412
rect 44899 28371 44957 28372
rect 45675 28412 45717 28421
rect 45675 28372 45676 28412
rect 45716 28372 45717 28412
rect 45675 28363 45717 28372
rect 2659 28328 2717 28329
rect 2659 28288 2668 28328
rect 2708 28288 2717 28328
rect 2659 28287 2717 28288
rect 3523 28328 3581 28329
rect 3523 28288 3532 28328
rect 3572 28288 3581 28328
rect 3523 28287 3581 28288
rect 5155 28328 5213 28329
rect 5155 28288 5164 28328
rect 5204 28288 5213 28328
rect 5155 28287 5213 28288
rect 6115 28328 6173 28329
rect 6115 28288 6124 28328
rect 6164 28288 6173 28328
rect 6115 28287 6173 28288
rect 6499 28328 6557 28329
rect 6499 28288 6508 28328
rect 6548 28288 6557 28328
rect 6499 28287 6557 28288
rect 12067 28328 12125 28329
rect 12067 28288 12076 28328
rect 12116 28288 12125 28328
rect 12067 28287 12125 28288
rect 12747 28328 12789 28337
rect 12747 28288 12748 28328
rect 12788 28288 12789 28328
rect 12747 28279 12789 28288
rect 12931 28328 12989 28329
rect 12931 28288 12940 28328
rect 12980 28288 12989 28328
rect 12931 28287 12989 28288
rect 13131 28328 13173 28337
rect 13131 28288 13132 28328
rect 13172 28288 13173 28328
rect 13131 28279 13173 28288
rect 25123 28328 25181 28329
rect 25123 28288 25132 28328
rect 25172 28288 25181 28328
rect 25123 28287 25181 28288
rect 26083 28328 26141 28329
rect 26083 28288 26092 28328
rect 26132 28288 26141 28328
rect 26083 28287 26141 28288
rect 26947 28328 27005 28329
rect 26947 28288 26956 28328
rect 26996 28288 27005 28328
rect 26947 28287 27005 28288
rect 28003 28328 28061 28329
rect 28003 28288 28012 28328
rect 28052 28288 28061 28328
rect 28003 28287 28061 28288
rect 28291 28328 28349 28329
rect 28291 28288 28300 28328
rect 28340 28288 28349 28328
rect 28291 28287 28349 28288
rect 28771 28328 28829 28329
rect 28771 28288 28780 28328
rect 28820 28288 28829 28328
rect 28771 28287 28829 28288
rect 28867 28328 28925 28329
rect 28867 28288 28876 28328
rect 28916 28288 28925 28328
rect 28867 28287 28925 28288
rect 41731 28328 41789 28329
rect 41731 28288 41740 28328
rect 41780 28288 41789 28328
rect 41731 28287 41789 28288
rect 42603 28328 42645 28337
rect 42603 28288 42604 28328
rect 42644 28288 42645 28328
rect 42603 28279 42645 28288
rect 46339 28328 46397 28329
rect 46339 28288 46348 28328
rect 46388 28288 46397 28328
rect 46339 28287 46397 28288
rect 2283 28244 2325 28253
rect 2283 28204 2284 28244
rect 2324 28204 2325 28244
rect 2283 28195 2325 28204
rect 27811 28244 27869 28245
rect 27811 28204 27820 28244
rect 27860 28204 27869 28244
rect 27811 28203 27869 28204
rect 6403 28160 6461 28161
rect 6403 28120 6412 28160
rect 6452 28120 6461 28160
rect 6403 28119 6461 28120
rect 6691 28160 6749 28161
rect 6691 28120 6700 28160
rect 6740 28120 6749 28160
rect 6691 28119 6749 28120
rect 26275 28160 26333 28161
rect 26275 28120 26284 28160
rect 26324 28120 26333 28160
rect 26275 28119 26333 28120
rect 29067 28160 29109 28169
rect 29067 28120 29068 28160
rect 29108 28120 29109 28160
rect 29067 28111 29109 28120
rect 44715 28160 44757 28169
rect 44715 28120 44716 28160
rect 44756 28120 44757 28160
rect 44715 28111 44757 28120
rect 576 27992 99360 28016
rect 576 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 19472 27992
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19840 27952 34592 27992
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34960 27952 49712 27992
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 50080 27952 64832 27992
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 65200 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 95072 27992
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95440 27952 99360 27992
rect 576 27928 99360 27952
rect 46147 27824 46205 27825
rect 46147 27784 46156 27824
rect 46196 27784 46205 27824
rect 46147 27783 46205 27784
rect 8619 27740 8661 27749
rect 8619 27700 8620 27740
rect 8660 27700 8661 27740
rect 8619 27691 8661 27700
rect 14179 27740 14237 27741
rect 14179 27700 14188 27740
rect 14228 27700 14237 27740
rect 14179 27699 14237 27700
rect 43755 27740 43797 27749
rect 43755 27700 43756 27740
rect 43796 27700 43797 27740
rect 43755 27691 43797 27700
rect 47211 27740 47253 27749
rect 47211 27700 47212 27740
rect 47252 27700 47253 27740
rect 47211 27691 47253 27700
rect 3915 27656 3957 27665
rect 3915 27616 3916 27656
rect 3956 27616 3957 27656
rect 3915 27607 3957 27616
rect 4291 27656 4349 27657
rect 4291 27616 4300 27656
rect 4340 27616 4349 27656
rect 4291 27615 4349 27616
rect 5155 27656 5213 27657
rect 5155 27616 5164 27656
rect 5204 27616 5213 27656
rect 5155 27615 5213 27616
rect 8995 27656 9053 27657
rect 8995 27616 9004 27656
rect 9044 27616 9053 27656
rect 8995 27615 9053 27616
rect 9859 27656 9917 27657
rect 9859 27616 9868 27656
rect 9908 27616 9917 27656
rect 9859 27615 9917 27616
rect 13507 27656 13565 27657
rect 13507 27616 13516 27656
rect 13556 27616 13565 27656
rect 13507 27615 13565 27616
rect 13699 27656 13757 27657
rect 13699 27616 13708 27656
rect 13748 27616 13757 27656
rect 13699 27615 13757 27616
rect 14083 27656 14141 27657
rect 14083 27616 14092 27656
rect 14132 27616 14141 27656
rect 14083 27615 14141 27616
rect 14563 27656 14621 27657
rect 14563 27616 14572 27656
rect 14612 27616 14621 27656
rect 14563 27615 14621 27616
rect 22051 27656 22109 27657
rect 22051 27616 22060 27656
rect 22100 27616 22109 27656
rect 22051 27615 22109 27616
rect 22915 27656 22973 27657
rect 22915 27616 22924 27656
rect 22964 27616 22973 27656
rect 22915 27615 22973 27616
rect 23307 27656 23349 27665
rect 23307 27616 23308 27656
rect 23348 27616 23349 27656
rect 23307 27607 23349 27616
rect 29731 27656 29789 27657
rect 29731 27616 29740 27656
rect 29780 27616 29789 27656
rect 29731 27615 29789 27616
rect 42499 27656 42557 27657
rect 42499 27616 42508 27656
rect 42548 27616 42557 27656
rect 42499 27615 42557 27616
rect 43371 27656 43413 27665
rect 43371 27616 43372 27656
rect 43412 27616 43413 27656
rect 43371 27607 43413 27616
rect 44131 27656 44189 27657
rect 44131 27616 44140 27656
rect 44180 27616 44189 27656
rect 44131 27615 44189 27616
rect 44995 27656 45053 27657
rect 44995 27616 45004 27656
rect 45044 27616 45053 27656
rect 44995 27615 45053 27616
rect 47875 27656 47933 27657
rect 47875 27616 47884 27656
rect 47924 27616 47933 27656
rect 47875 27615 47933 27616
rect 3427 27572 3485 27573
rect 3427 27532 3436 27572
rect 3476 27532 3485 27572
rect 3427 27531 3485 27532
rect 11019 27572 11061 27581
rect 11019 27532 11020 27572
rect 11060 27532 11061 27572
rect 11019 27523 11061 27532
rect 47011 27572 47069 27573
rect 47011 27532 47020 27572
rect 47060 27532 47069 27572
rect 47011 27531 47069 27532
rect 3243 27488 3285 27497
rect 3243 27448 3244 27488
rect 3284 27448 3285 27488
rect 3243 27439 3285 27448
rect 6307 27404 6365 27405
rect 6307 27364 6316 27404
rect 6356 27364 6365 27404
rect 6307 27363 6365 27364
rect 12835 27404 12893 27405
rect 12835 27364 12844 27404
rect 12884 27364 12893 27404
rect 12835 27363 12893 27364
rect 15235 27404 15293 27405
rect 15235 27364 15244 27404
rect 15284 27364 15293 27404
rect 15235 27363 15293 27364
rect 20899 27404 20957 27405
rect 20899 27364 20908 27404
rect 20948 27364 20957 27404
rect 20899 27363 20957 27364
rect 30403 27404 30461 27405
rect 30403 27364 30412 27404
rect 30452 27364 30461 27404
rect 30403 27363 30461 27364
rect 46827 27404 46869 27413
rect 46827 27364 46828 27404
rect 46868 27364 46869 27404
rect 46827 27355 46869 27364
rect 576 27236 99360 27260
rect 576 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 18232 27236
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18600 27196 33352 27236
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33720 27196 48472 27236
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48840 27196 63592 27236
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63960 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 93832 27236
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 94200 27196 99360 27236
rect 576 27172 99360 27196
rect 4491 27068 4533 27077
rect 4491 27028 4492 27068
rect 4532 27028 4533 27068
rect 4491 27019 4533 27028
rect 5635 27068 5693 27069
rect 5635 27028 5644 27068
rect 5684 27028 5693 27068
rect 5635 27027 5693 27028
rect 44043 27068 44085 27077
rect 44043 27028 44044 27068
rect 44084 27028 44085 27068
rect 44043 27019 44085 27028
rect 49411 27068 49469 27069
rect 49411 27028 49420 27068
rect 49460 27028 49469 27068
rect 49411 27027 49469 27028
rect 4675 26900 4733 26901
rect 4675 26860 4684 26900
rect 4724 26860 4733 26900
rect 4675 26859 4733 26860
rect 39531 26900 39573 26909
rect 39531 26860 39532 26900
rect 39572 26860 39573 26900
rect 39531 26851 39573 26860
rect 6307 26816 6365 26817
rect 6307 26776 6316 26816
rect 6356 26776 6365 26816
rect 6307 26775 6365 26776
rect 9187 26816 9245 26817
rect 9187 26776 9196 26816
rect 9236 26776 9245 26816
rect 9187 26775 9245 26776
rect 10059 26816 10101 26825
rect 10059 26776 10060 26816
rect 10100 26776 10101 26816
rect 10059 26767 10101 26776
rect 12747 26816 12789 26825
rect 12747 26776 12748 26816
rect 12788 26776 12789 26816
rect 12747 26767 12789 26776
rect 13123 26816 13181 26817
rect 13123 26776 13132 26816
rect 13172 26776 13181 26816
rect 13123 26775 13181 26776
rect 13987 26816 14045 26817
rect 13987 26776 13996 26816
rect 14036 26776 14045 26816
rect 13987 26775 14045 26776
rect 15339 26816 15381 26825
rect 15339 26776 15340 26816
rect 15380 26776 15381 26816
rect 15339 26767 15381 26776
rect 15715 26816 15773 26817
rect 15715 26776 15724 26816
rect 15764 26776 15773 26816
rect 15715 26775 15773 26776
rect 16579 26816 16637 26817
rect 16579 26776 16588 26816
rect 16628 26776 16637 26816
rect 16579 26775 16637 26776
rect 19555 26816 19613 26817
rect 19555 26776 19564 26816
rect 19604 26776 19613 26816
rect 19555 26775 19613 26776
rect 20515 26816 20573 26817
rect 20515 26776 20524 26816
rect 20564 26776 20573 26816
rect 20515 26775 20573 26776
rect 28963 26816 29021 26817
rect 28963 26776 28972 26816
rect 29012 26776 29021 26816
rect 28963 26775 29021 26776
rect 29827 26816 29885 26817
rect 29827 26776 29836 26816
rect 29876 26776 29885 26816
rect 29827 26775 29885 26776
rect 30219 26816 30261 26825
rect 30219 26776 30220 26816
rect 30260 26776 30261 26816
rect 30219 26767 30261 26776
rect 32131 26816 32189 26817
rect 32131 26776 32140 26816
rect 32180 26776 32189 26816
rect 32131 26775 32189 26776
rect 37507 26816 37565 26817
rect 37507 26776 37516 26816
rect 37556 26776 37565 26816
rect 37507 26775 37565 26776
rect 38371 26816 38429 26817
rect 38371 26776 38380 26816
rect 38420 26776 38429 26816
rect 38371 26775 38429 26776
rect 40387 26816 40445 26817
rect 40387 26776 40396 26816
rect 40436 26776 40445 26816
rect 40387 26775 40445 26776
rect 44427 26816 44469 26825
rect 44427 26776 44428 26816
rect 44468 26776 44469 26816
rect 44427 26767 44469 26776
rect 47019 26816 47061 26825
rect 47019 26776 47020 26816
rect 47060 26776 47061 26816
rect 47019 26767 47061 26776
rect 47395 26816 47453 26817
rect 47395 26776 47404 26816
rect 47444 26776 47453 26816
rect 47395 26775 47453 26776
rect 48259 26816 48317 26817
rect 48259 26776 48268 26816
rect 48308 26776 48317 26816
rect 48259 26775 48317 26776
rect 37131 26732 37173 26741
rect 37131 26692 37132 26732
rect 37172 26692 37173 26732
rect 37131 26683 37173 26692
rect 15139 26648 15197 26649
rect 15139 26608 15148 26648
rect 15188 26608 15197 26648
rect 15139 26607 15197 26608
rect 17731 26648 17789 26649
rect 17731 26608 17740 26648
rect 17780 26608 17789 26648
rect 17731 26607 17789 26608
rect 27811 26648 27869 26649
rect 27811 26608 27820 26648
rect 27860 26608 27869 26648
rect 27811 26607 27869 26608
rect 31459 26648 31517 26649
rect 31459 26608 31468 26648
rect 31508 26608 31517 26648
rect 31459 26607 31517 26608
rect 39715 26648 39773 26649
rect 39715 26608 39724 26648
rect 39764 26608 39773 26648
rect 39715 26607 39773 26608
rect 576 26480 99360 26504
rect 576 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 19472 26480
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19840 26440 34592 26480
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34960 26440 49712 26480
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 50080 26440 64832 26480
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 65200 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 95072 26480
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95440 26440 99360 26480
rect 576 26416 99360 26440
rect 11787 26312 11829 26321
rect 11787 26272 11788 26312
rect 11828 26272 11829 26312
rect 11787 26263 11829 26272
rect 30219 26312 30261 26321
rect 30219 26272 30220 26312
rect 30260 26272 30261 26312
rect 30219 26263 30261 26272
rect 33283 26312 33341 26313
rect 33283 26272 33292 26312
rect 33332 26272 33341 26312
rect 33283 26271 33341 26272
rect 38187 26312 38229 26321
rect 38187 26272 38188 26312
rect 38228 26272 38229 26312
rect 38187 26263 38229 26272
rect 4867 26144 4925 26145
rect 4867 26104 4876 26144
rect 4916 26104 4925 26144
rect 4867 26103 4925 26104
rect 11403 26144 11445 26153
rect 11403 26104 11404 26144
rect 11444 26104 11445 26144
rect 11403 26095 11445 26104
rect 18979 26144 19037 26145
rect 18979 26104 18988 26144
rect 19028 26104 19037 26144
rect 18979 26103 19037 26104
rect 19659 26144 19701 26153
rect 19659 26104 19660 26144
rect 19700 26104 19701 26144
rect 19659 26095 19701 26104
rect 19851 26144 19893 26153
rect 19851 26104 19852 26144
rect 19892 26104 19893 26144
rect 19851 26095 19893 26104
rect 20227 26144 20285 26145
rect 20227 26104 20236 26144
rect 20276 26104 20285 26144
rect 20227 26103 20285 26104
rect 21091 26144 21149 26145
rect 21091 26104 21100 26144
rect 21140 26104 21149 26144
rect 21091 26103 21149 26104
rect 29835 26144 29877 26153
rect 29835 26104 29836 26144
rect 29876 26104 29877 26144
rect 29835 26095 29877 26104
rect 30691 26144 30749 26145
rect 30691 26104 30700 26144
rect 30740 26104 30749 26144
rect 30691 26103 30749 26104
rect 30891 26144 30933 26153
rect 30891 26104 30892 26144
rect 30932 26104 30933 26144
rect 30891 26095 30933 26104
rect 31267 26144 31325 26145
rect 31267 26104 31276 26144
rect 31316 26104 31325 26144
rect 31267 26103 31325 26104
rect 32131 26144 32189 26145
rect 32131 26104 32140 26144
rect 32180 26104 32189 26144
rect 32131 26103 32189 26104
rect 34539 26144 34581 26153
rect 34539 26104 34540 26144
rect 34580 26104 34581 26144
rect 34539 26095 34581 26104
rect 34915 26144 34973 26145
rect 34915 26104 34924 26144
rect 34964 26104 34973 26144
rect 34915 26103 34973 26104
rect 35779 26144 35837 26145
rect 35779 26104 35788 26144
rect 35828 26104 35837 26144
rect 35779 26103 35837 26104
rect 41355 26144 41397 26153
rect 41355 26104 41356 26144
rect 41396 26104 41397 26144
rect 41355 26095 41397 26104
rect 41731 26144 41789 26145
rect 41731 26104 41740 26144
rect 41780 26104 41789 26144
rect 41731 26103 41789 26104
rect 42595 26144 42653 26145
rect 42595 26104 42604 26144
rect 42644 26104 42653 26144
rect 42595 26103 42653 26104
rect 46627 26144 46685 26145
rect 46627 26104 46636 26144
rect 46676 26104 46685 26144
rect 46627 26103 46685 26104
rect 3427 26060 3485 26061
rect 3427 26020 3436 26060
rect 3476 26020 3485 26060
rect 3427 26019 3485 26020
rect 23779 26060 23837 26061
rect 23779 26020 23788 26060
rect 23828 26020 23837 26060
rect 23779 26019 23837 26020
rect 38371 26060 38429 26061
rect 38371 26020 38380 26060
rect 38420 26020 38429 26060
rect 38371 26019 38429 26020
rect 3243 25892 3285 25901
rect 3243 25852 3244 25892
rect 3284 25852 3285 25892
rect 3243 25843 3285 25852
rect 4195 25892 4253 25893
rect 4195 25852 4204 25892
rect 4244 25852 4253 25892
rect 4195 25851 4253 25852
rect 22243 25892 22301 25893
rect 22243 25852 22252 25892
rect 22292 25852 22301 25892
rect 22243 25851 22301 25852
rect 23595 25892 23637 25901
rect 23595 25852 23596 25892
rect 23636 25852 23637 25892
rect 23595 25843 23637 25852
rect 36931 25892 36989 25893
rect 36931 25852 36940 25892
rect 36980 25852 36989 25892
rect 36931 25851 36989 25852
rect 43747 25892 43805 25893
rect 43747 25852 43756 25892
rect 43796 25852 43805 25892
rect 43747 25851 43805 25852
rect 46347 25892 46389 25901
rect 46347 25852 46348 25892
rect 46388 25852 46389 25892
rect 46347 25843 46389 25852
rect 576 25724 99360 25748
rect 576 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 18232 25724
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18600 25684 33352 25724
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33720 25684 48472 25724
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48840 25684 63592 25724
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63960 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 93832 25724
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 94200 25684 99360 25724
rect 576 25660 99360 25684
rect 4771 25556 4829 25557
rect 4771 25516 4780 25556
rect 4820 25516 4829 25556
rect 4771 25515 4829 25516
rect 18123 25556 18165 25565
rect 18123 25516 18124 25556
rect 18164 25516 18165 25556
rect 18123 25507 18165 25516
rect 25995 25556 26037 25565
rect 25995 25516 25996 25556
rect 26036 25516 26037 25556
rect 25995 25507 26037 25516
rect 31851 25556 31893 25565
rect 31851 25516 31852 25556
rect 31892 25516 31893 25556
rect 31851 25507 31893 25516
rect 34347 25556 34389 25565
rect 34347 25516 34348 25556
rect 34388 25516 34389 25556
rect 34347 25507 34389 25516
rect 19459 25388 19517 25389
rect 19459 25348 19468 25388
rect 19508 25348 19517 25388
rect 19459 25347 19517 25348
rect 32035 25388 32093 25389
rect 32035 25348 32044 25388
rect 32084 25348 32093 25388
rect 32035 25347 32093 25348
rect 39627 25388 39669 25397
rect 39627 25348 39628 25388
rect 39668 25348 39669 25388
rect 39627 25339 39669 25348
rect 2379 25304 2421 25313
rect 2379 25264 2380 25304
rect 2420 25264 2421 25304
rect 2379 25255 2421 25264
rect 2755 25304 2813 25305
rect 2755 25264 2764 25304
rect 2804 25264 2813 25304
rect 2755 25263 2813 25264
rect 3619 25304 3677 25305
rect 3619 25264 3628 25304
rect 3668 25264 3677 25304
rect 3619 25263 3677 25264
rect 16771 25304 16829 25305
rect 16771 25264 16780 25304
rect 16820 25264 16829 25304
rect 16771 25263 16829 25264
rect 17059 25304 17117 25305
rect 17059 25264 17068 25304
rect 17108 25264 17117 25304
rect 17059 25263 17117 25264
rect 17835 25304 17877 25313
rect 17835 25264 17836 25304
rect 17876 25264 17877 25304
rect 17835 25255 17877 25264
rect 17923 25304 17981 25305
rect 17923 25264 17932 25304
rect 17972 25264 17981 25304
rect 17923 25263 17981 25264
rect 18403 25304 18461 25305
rect 18403 25264 18412 25304
rect 18452 25264 18461 25304
rect 18403 25263 18461 25264
rect 21859 25304 21917 25305
rect 21859 25264 21868 25304
rect 21908 25264 21917 25304
rect 21859 25263 21917 25264
rect 22819 25304 22877 25305
rect 22819 25264 22828 25304
rect 22868 25264 22877 25304
rect 22819 25263 22877 25264
rect 23203 25304 23261 25305
rect 23203 25264 23212 25304
rect 23252 25264 23261 25304
rect 23203 25263 23261 25264
rect 23595 25304 23637 25313
rect 23595 25264 23596 25304
rect 23636 25264 23637 25304
rect 23595 25255 23637 25264
rect 23971 25304 24029 25305
rect 23971 25264 23980 25304
rect 24020 25264 24029 25304
rect 23971 25263 24029 25264
rect 24835 25304 24893 25305
rect 24835 25264 24844 25304
rect 24884 25264 24893 25304
rect 24835 25263 24893 25264
rect 34051 25304 34109 25305
rect 34051 25264 34060 25304
rect 34100 25264 34109 25304
rect 34051 25263 34109 25264
rect 35011 25304 35069 25305
rect 35011 25264 35020 25304
rect 35060 25264 35069 25304
rect 35011 25263 35069 25264
rect 39523 25304 39581 25305
rect 39523 25264 39532 25304
rect 39572 25264 39581 25304
rect 39523 25263 39581 25264
rect 39723 25304 39765 25313
rect 39723 25264 39724 25304
rect 39764 25264 39765 25304
rect 39723 25255 39765 25264
rect 40291 25304 40349 25305
rect 40291 25264 40300 25304
rect 40340 25264 40349 25304
rect 40291 25263 40349 25264
rect 40675 25304 40733 25305
rect 40675 25264 40684 25304
rect 40724 25264 40733 25304
rect 40675 25263 40733 25264
rect 41251 25304 41309 25305
rect 41251 25264 41260 25304
rect 41300 25264 41309 25304
rect 41251 25263 41309 25264
rect 41635 25304 41693 25305
rect 41635 25264 41644 25304
rect 41684 25264 41693 25304
rect 41635 25263 41693 25264
rect 17251 25220 17309 25221
rect 17251 25180 17260 25220
rect 17300 25180 17309 25220
rect 17251 25179 17309 25180
rect 41731 25220 41789 25221
rect 41731 25180 41740 25220
rect 41780 25180 41789 25220
rect 41731 25179 41789 25180
rect 19075 25136 19133 25137
rect 19075 25096 19084 25136
rect 19124 25096 19133 25136
rect 19075 25095 19133 25096
rect 22531 25136 22589 25137
rect 22531 25096 22540 25136
rect 22580 25096 22589 25136
rect 22531 25095 22589 25096
rect 23307 25136 23349 25145
rect 23307 25096 23308 25136
rect 23348 25096 23349 25136
rect 23307 25087 23349 25096
rect 40779 25136 40821 25145
rect 40779 25096 40780 25136
rect 40820 25096 40821 25136
rect 40779 25087 40821 25096
rect 576 24968 99360 24992
rect 576 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 19472 24968
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19840 24928 34592 24968
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34960 24928 49712 24968
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 50080 24928 64832 24968
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 65200 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 95072 24968
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95440 24928 99360 24968
rect 576 24904 99360 24928
rect 32715 24800 32757 24809
rect 32715 24760 32716 24800
rect 32756 24760 32757 24800
rect 32715 24751 32757 24760
rect 38659 24800 38717 24801
rect 38659 24760 38668 24800
rect 38708 24760 38717 24800
rect 38659 24759 38717 24760
rect 31947 24716 31989 24725
rect 31947 24676 31948 24716
rect 31988 24676 31989 24716
rect 31947 24667 31989 24676
rect 33091 24716 33149 24717
rect 33091 24676 33100 24716
rect 33140 24676 33149 24716
rect 33091 24675 33149 24676
rect 18403 24632 18461 24633
rect 18403 24592 18412 24632
rect 18452 24592 18461 24632
rect 18403 24591 18461 24592
rect 18603 24632 18645 24641
rect 18603 24592 18604 24632
rect 18644 24592 18645 24632
rect 18603 24583 18645 24592
rect 31851 24632 31893 24641
rect 31851 24592 31852 24632
rect 31892 24592 31893 24632
rect 31851 24583 31893 24592
rect 32035 24632 32093 24633
rect 32035 24592 32044 24632
rect 32084 24592 32093 24632
rect 32035 24591 32093 24592
rect 32227 24632 32285 24633
rect 32227 24592 32236 24632
rect 32276 24592 32285 24632
rect 32227 24591 32285 24592
rect 32515 24632 32573 24633
rect 32515 24592 32524 24632
rect 32564 24592 32573 24632
rect 32515 24591 32573 24592
rect 33955 24632 34013 24633
rect 33955 24592 33964 24632
rect 34004 24592 34013 24632
rect 33955 24591 34013 24592
rect 39331 24632 39389 24633
rect 39331 24592 39340 24632
rect 39380 24592 39389 24632
rect 39331 24591 39389 24592
rect 42307 24632 42365 24633
rect 42307 24592 42316 24632
rect 42356 24592 42365 24632
rect 42307 24591 42365 24592
rect 43267 24632 43325 24633
rect 43267 24592 43276 24632
rect 43316 24592 43325 24632
rect 43267 24591 43325 24592
rect 37891 24548 37949 24549
rect 37891 24508 37900 24548
rect 37940 24508 37949 24548
rect 37891 24507 37949 24508
rect 18507 24464 18549 24473
rect 18507 24424 18508 24464
rect 18548 24424 18549 24464
rect 18507 24415 18549 24424
rect 37707 24380 37749 24389
rect 37707 24340 37708 24380
rect 37748 24340 37749 24380
rect 37707 24331 37749 24340
rect 576 24212 99360 24236
rect 576 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 18232 24212
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18600 24172 33352 24212
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33720 24172 48472 24212
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48840 24172 63592 24212
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63960 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 93832 24212
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 94200 24172 99360 24212
rect 576 24148 99360 24172
rect 18691 24044 18749 24045
rect 18691 24004 18700 24044
rect 18740 24004 18749 24044
rect 18691 24003 18749 24004
rect 39235 24044 39293 24045
rect 39235 24004 39244 24044
rect 39284 24004 39293 24044
rect 39235 24003 39293 24004
rect 16771 23960 16829 23961
rect 16771 23920 16780 23960
rect 16820 23920 16829 23960
rect 16771 23919 16829 23920
rect 3619 23876 3677 23877
rect 3619 23836 3628 23876
rect 3668 23836 3677 23876
rect 3619 23835 3677 23836
rect 42891 23876 42933 23885
rect 42891 23836 42892 23876
rect 42932 23836 42933 23876
rect 42891 23827 42933 23836
rect 43171 23876 43229 23877
rect 43171 23836 43180 23876
rect 43220 23836 43229 23876
rect 43171 23835 43229 23836
rect 4107 23792 4149 23801
rect 4107 23752 4108 23792
rect 4148 23752 4149 23792
rect 4107 23743 4149 23752
rect 4291 23792 4349 23793
rect 4291 23752 4300 23792
rect 4340 23752 4349 23792
rect 4291 23751 4349 23752
rect 5155 23792 5213 23793
rect 5155 23752 5164 23792
rect 5204 23752 5213 23792
rect 5155 23751 5213 23752
rect 9475 23792 9533 23793
rect 9475 23752 9484 23792
rect 9524 23752 9533 23792
rect 9475 23751 9533 23752
rect 10339 23792 10397 23793
rect 10339 23752 10348 23792
rect 10388 23752 10397 23792
rect 10339 23751 10397 23752
rect 13507 23792 13565 23793
rect 13507 23752 13516 23792
rect 13556 23752 13565 23792
rect 13507 23751 13565 23752
rect 14755 23792 14813 23793
rect 14755 23752 14764 23792
rect 14804 23752 14813 23792
rect 14755 23751 14813 23752
rect 15619 23792 15677 23793
rect 15619 23752 15628 23792
rect 15668 23752 15677 23792
rect 15619 23751 15677 23752
rect 19363 23792 19421 23793
rect 19363 23752 19372 23792
rect 19412 23752 19421 23792
rect 19363 23751 19421 23752
rect 36843 23792 36885 23801
rect 36843 23752 36844 23792
rect 36884 23752 36885 23792
rect 36843 23743 36885 23752
rect 37219 23792 37277 23793
rect 37219 23752 37228 23792
rect 37268 23752 37277 23792
rect 37219 23751 37277 23752
rect 38083 23792 38141 23793
rect 38083 23752 38092 23792
rect 38132 23752 38141 23792
rect 38083 23751 38141 23752
rect 42787 23792 42845 23793
rect 42787 23752 42796 23792
rect 42836 23752 42845 23792
rect 42787 23751 42845 23752
rect 42987 23792 43029 23801
rect 42987 23752 42988 23792
rect 43028 23752 43029 23792
rect 42987 23743 43029 23752
rect 43755 23792 43797 23801
rect 43755 23752 43756 23792
rect 43796 23752 43797 23792
rect 43755 23743 43797 23752
rect 44419 23792 44477 23793
rect 44419 23752 44428 23792
rect 44468 23752 44477 23792
rect 44419 23751 44477 23752
rect 4203 23708 4245 23717
rect 4203 23668 4204 23708
rect 4244 23668 4245 23708
rect 4203 23659 4245 23668
rect 9099 23708 9141 23717
rect 9099 23668 9100 23708
rect 9140 23668 9141 23708
rect 9099 23659 9141 23668
rect 14187 23708 14229 23717
rect 14187 23668 14188 23708
rect 14228 23668 14229 23708
rect 14187 23659 14229 23668
rect 14379 23708 14421 23717
rect 14379 23668 14380 23708
rect 14420 23668 14421 23708
rect 14379 23659 14421 23668
rect 3435 23624 3477 23633
rect 3435 23584 3436 23624
rect 3476 23584 3477 23624
rect 3435 23575 3477 23584
rect 4483 23624 4541 23625
rect 4483 23584 4492 23624
rect 4532 23584 4541 23624
rect 4483 23583 4541 23584
rect 11491 23624 11549 23625
rect 11491 23584 11500 23624
rect 11540 23584 11549 23624
rect 11491 23583 11549 23584
rect 43371 23624 43413 23633
rect 43371 23584 43372 23624
rect 43412 23584 43413 23624
rect 43371 23575 43413 23584
rect 576 23456 99360 23480
rect 576 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 19472 23456
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19840 23416 34592 23456
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34960 23416 49712 23456
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 50080 23416 64832 23456
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 65200 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 95072 23456
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95440 23416 99360 23456
rect 576 23392 99360 23416
rect 5059 23288 5117 23289
rect 5059 23248 5068 23288
rect 5108 23248 5117 23288
rect 5059 23247 5117 23248
rect 6019 23288 6077 23289
rect 6019 23248 6028 23288
rect 6068 23248 6077 23288
rect 6019 23247 6077 23248
rect 6307 23288 6365 23289
rect 6307 23248 6316 23288
rect 6356 23248 6365 23288
rect 6307 23247 6365 23248
rect 13707 23288 13749 23297
rect 13707 23248 13708 23288
rect 13748 23248 13749 23288
rect 13707 23239 13749 23248
rect 39043 23288 39101 23289
rect 39043 23248 39052 23288
rect 39092 23248 39101 23288
rect 39043 23247 39101 23248
rect 42691 23288 42749 23289
rect 42691 23248 42700 23288
rect 42740 23248 42749 23288
rect 42691 23247 42749 23248
rect 2667 23204 2709 23213
rect 2667 23164 2668 23204
rect 2708 23164 2709 23204
rect 2667 23155 2709 23164
rect 5731 23204 5789 23205
rect 5731 23164 5740 23204
rect 5780 23164 5789 23204
rect 5731 23163 5789 23164
rect 7563 23204 7605 23213
rect 7563 23164 7564 23204
rect 7604 23164 7605 23204
rect 7563 23155 7605 23164
rect 19075 23204 19133 23205
rect 19075 23164 19084 23204
rect 19124 23164 19133 23204
rect 19075 23163 19133 23164
rect 31755 23204 31797 23213
rect 31755 23164 31756 23204
rect 31796 23164 31797 23204
rect 31755 23155 31797 23164
rect 45963 23204 46005 23213
rect 45963 23164 45964 23204
rect 46004 23164 46005 23204
rect 45963 23155 46005 23164
rect 3043 23120 3101 23121
rect 3043 23080 3052 23120
rect 3092 23080 3101 23120
rect 3043 23079 3101 23080
rect 3907 23120 3965 23121
rect 3907 23080 3916 23120
rect 3956 23080 3965 23120
rect 3907 23079 3965 23080
rect 5251 23120 5309 23121
rect 5251 23080 5260 23120
rect 5300 23080 5309 23120
rect 5251 23079 5309 23080
rect 5539 23120 5597 23121
rect 5539 23080 5548 23120
rect 5588 23080 5597 23120
rect 5539 23079 5597 23080
rect 6115 23120 6173 23121
rect 6115 23080 6124 23120
rect 6164 23080 6173 23120
rect 6115 23079 6173 23080
rect 7939 23120 7997 23121
rect 7939 23080 7948 23120
rect 7988 23080 7997 23120
rect 7939 23079 7997 23080
rect 8803 23120 8861 23121
rect 8803 23080 8812 23120
rect 8852 23080 8861 23120
rect 8803 23079 8861 23080
rect 12835 23120 12893 23121
rect 12835 23080 12844 23120
rect 12884 23080 12893 23120
rect 12835 23079 12893 23080
rect 13987 23120 14045 23121
rect 13987 23080 13996 23120
rect 14036 23080 14045 23120
rect 13987 23079 14045 23080
rect 14091 23120 14133 23129
rect 14091 23080 14092 23120
rect 14132 23080 14133 23120
rect 14091 23071 14133 23080
rect 18595 23120 18653 23121
rect 18595 23080 18604 23120
rect 18644 23080 18653 23120
rect 18595 23079 18653 23080
rect 18979 23120 19037 23121
rect 18979 23080 18988 23120
rect 19028 23080 19037 23120
rect 18979 23079 19037 23080
rect 19555 23120 19613 23121
rect 19555 23080 19564 23120
rect 19604 23080 19613 23120
rect 19555 23079 19613 23080
rect 21859 23120 21917 23121
rect 21859 23080 21868 23120
rect 21908 23080 21917 23120
rect 21859 23079 21917 23080
rect 21963 23120 22005 23129
rect 21963 23080 21964 23120
rect 22004 23080 22005 23120
rect 21963 23071 22005 23080
rect 22339 23120 22397 23121
rect 22339 23080 22348 23120
rect 22388 23080 22397 23120
rect 22339 23079 22397 23080
rect 24835 23120 24893 23121
rect 24835 23080 24844 23120
rect 24884 23080 24893 23120
rect 24835 23079 24893 23080
rect 25707 23120 25749 23129
rect 25707 23080 25708 23120
rect 25748 23080 25749 23120
rect 25707 23071 25749 23080
rect 26179 23120 26237 23121
rect 26179 23080 26188 23120
rect 26228 23080 26237 23120
rect 26179 23079 26237 23080
rect 27139 23120 27197 23121
rect 27139 23080 27148 23120
rect 27188 23080 27197 23120
rect 27139 23079 27197 23080
rect 28771 23120 28829 23121
rect 28771 23080 28780 23120
rect 28820 23080 28829 23120
rect 28771 23079 28829 23080
rect 29451 23120 29493 23129
rect 29451 23080 29452 23120
rect 29492 23080 29493 23120
rect 29451 23071 29493 23080
rect 31659 23120 31701 23129
rect 31659 23080 31660 23120
rect 31700 23080 31701 23120
rect 31659 23071 31701 23080
rect 31843 23120 31901 23121
rect 31843 23080 31852 23120
rect 31892 23080 31901 23120
rect 31843 23079 31901 23080
rect 33667 23120 33725 23121
rect 33667 23080 33676 23120
rect 33716 23080 33725 23120
rect 33667 23079 33725 23080
rect 34627 23120 34685 23121
rect 34627 23080 34636 23120
rect 34676 23080 34685 23120
rect 34627 23079 34685 23080
rect 38947 23120 39005 23121
rect 38947 23080 38956 23120
rect 38996 23080 39005 23120
rect 38947 23079 39005 23080
rect 43363 23120 43421 23121
rect 43363 23080 43372 23120
rect 43412 23080 43421 23120
rect 43363 23079 43421 23080
rect 44707 23120 44765 23121
rect 44707 23080 44716 23120
rect 44756 23080 44765 23120
rect 44707 23079 44765 23080
rect 45571 23120 45629 23121
rect 45571 23080 45580 23120
rect 45620 23080 45629 23120
rect 45571 23079 45629 23080
rect 47883 23120 47925 23129
rect 47883 23080 47884 23120
rect 47924 23080 47925 23120
rect 47883 23071 47925 23080
rect 48259 23120 48317 23121
rect 48259 23080 48268 23120
rect 48308 23080 48317 23120
rect 48259 23079 48317 23080
rect 49123 23120 49181 23121
rect 49123 23080 49132 23120
rect 49172 23080 49181 23120
rect 49123 23079 49181 23080
rect 29635 23036 29693 23037
rect 29635 22996 29644 23036
rect 29684 22996 29693 23036
rect 29635 22995 29693 22996
rect 32515 23036 32573 23037
rect 32515 22996 32524 23036
rect 32564 22996 32573 23036
rect 32515 22995 32573 22996
rect 33963 23036 34005 23045
rect 33963 22996 33964 23036
rect 34004 22996 34005 23036
rect 33963 22987 34005 22996
rect 43563 23036 43605 23045
rect 43563 22996 43564 23036
rect 43604 22996 43605 23036
rect 43563 22987 43605 22996
rect 9955 22868 10013 22869
rect 9955 22828 9964 22868
rect 10004 22828 10013 22868
rect 9955 22827 10013 22828
rect 13507 22868 13565 22869
rect 13507 22828 13516 22868
rect 13556 22828 13565 22868
rect 13507 22827 13565 22828
rect 20227 22868 20285 22869
rect 20227 22828 20236 22868
rect 20276 22828 20285 22868
rect 20227 22827 20285 22828
rect 21675 22868 21717 22877
rect 21675 22828 21676 22868
rect 21716 22828 21717 22868
rect 21675 22819 21717 22828
rect 23011 22868 23069 22869
rect 23011 22828 23020 22868
rect 23060 22828 23069 22868
rect 23011 22827 23069 22828
rect 29835 22868 29877 22877
rect 29835 22828 29836 22868
rect 29876 22828 29877 22868
rect 29835 22819 29877 22828
rect 32331 22868 32373 22877
rect 32331 22828 32332 22868
rect 32372 22828 32373 22868
rect 32331 22819 32373 22828
rect 33195 22868 33237 22877
rect 33195 22828 33196 22868
rect 33236 22828 33237 22868
rect 33195 22819 33237 22828
rect 38755 22868 38813 22869
rect 38755 22828 38764 22868
rect 38804 22828 38813 22868
rect 38755 22827 38813 22828
rect 50275 22868 50333 22869
rect 50275 22828 50284 22868
rect 50324 22828 50333 22868
rect 50275 22827 50333 22828
rect 576 22700 99360 22724
rect 576 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 18232 22700
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18600 22660 33352 22700
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33720 22660 48472 22700
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48840 22660 63592 22700
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63960 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 93832 22700
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 94200 22660 99360 22700
rect 576 22636 99360 22660
rect 4203 22532 4245 22541
rect 4203 22492 4204 22532
rect 4244 22492 4245 22532
rect 4203 22483 4245 22492
rect 4483 22532 4541 22533
rect 4483 22492 4492 22532
rect 4532 22492 4541 22532
rect 4483 22491 4541 22492
rect 13995 22532 14037 22541
rect 13995 22492 13996 22532
rect 14036 22492 14037 22532
rect 13995 22483 14037 22492
rect 18499 22532 18557 22533
rect 18499 22492 18508 22532
rect 18548 22492 18557 22532
rect 18499 22491 18557 22492
rect 22147 22532 22205 22533
rect 22147 22492 22156 22532
rect 22196 22492 22205 22532
rect 22147 22491 22205 22492
rect 23019 22532 23061 22541
rect 23019 22492 23020 22532
rect 23060 22492 23061 22532
rect 23019 22483 23061 22492
rect 28195 22532 28253 22533
rect 28195 22492 28204 22532
rect 28244 22492 28253 22532
rect 28195 22491 28253 22492
rect 34531 22532 34589 22533
rect 34531 22492 34540 22532
rect 34580 22492 34589 22532
rect 34531 22491 34589 22492
rect 44995 22532 45053 22533
rect 44995 22492 45004 22532
rect 45044 22492 45053 22532
rect 44995 22491 45053 22492
rect 651 22448 693 22457
rect 651 22408 652 22448
rect 692 22408 693 22448
rect 651 22399 693 22408
rect 47979 22448 48021 22457
rect 47979 22408 47980 22448
rect 48020 22408 48021 22448
rect 47979 22399 48021 22408
rect 3619 22364 3677 22365
rect 3619 22324 3628 22364
rect 3668 22324 3677 22364
rect 3619 22323 3677 22324
rect 22443 22364 22485 22373
rect 22443 22324 22444 22364
rect 22484 22324 22485 22364
rect 22443 22315 22485 22324
rect 31075 22364 31133 22365
rect 31075 22324 31084 22364
rect 31124 22324 31133 22364
rect 31075 22323 31133 22324
rect 42211 22364 42269 22365
rect 42211 22324 42220 22364
rect 42260 22324 42269 22364
rect 42211 22323 42269 22324
rect 4107 22280 4149 22289
rect 4107 22240 4108 22280
rect 4148 22240 4149 22280
rect 4107 22231 4149 22240
rect 4291 22280 4349 22281
rect 4291 22240 4300 22280
rect 4340 22240 4349 22280
rect 4291 22239 4349 22240
rect 5155 22280 5213 22281
rect 5155 22240 5164 22280
rect 5204 22240 5213 22280
rect 5155 22239 5213 22240
rect 11107 22280 11165 22281
rect 11107 22240 11116 22280
rect 11156 22240 11165 22280
rect 11107 22239 11165 22240
rect 11395 22280 11453 22281
rect 11395 22240 11404 22280
rect 11444 22240 11453 22280
rect 11395 22239 11453 22240
rect 13891 22280 13949 22281
rect 13891 22240 13900 22280
rect 13940 22240 13949 22280
rect 13891 22239 13949 22240
rect 14091 22280 14133 22289
rect 14091 22240 14092 22280
rect 14132 22240 14133 22280
rect 14091 22231 14133 22240
rect 14467 22280 14525 22281
rect 14467 22240 14476 22280
rect 14516 22240 14525 22280
rect 14467 22239 14525 22240
rect 14851 22280 14909 22281
rect 14851 22240 14860 22280
rect 14900 22240 14909 22280
rect 14851 22239 14909 22240
rect 15235 22280 15293 22281
rect 15235 22240 15244 22280
rect 15284 22240 15293 22280
rect 15235 22239 15293 22240
rect 16483 22280 16541 22281
rect 16483 22240 16492 22280
rect 16532 22240 16541 22280
rect 16483 22239 16541 22240
rect 17347 22280 17405 22281
rect 17347 22240 17356 22280
rect 17396 22240 17405 22280
rect 17347 22239 17405 22240
rect 19755 22280 19797 22289
rect 19755 22240 19756 22280
rect 19796 22240 19797 22280
rect 19755 22231 19797 22240
rect 20131 22280 20189 22281
rect 20131 22240 20140 22280
rect 20180 22240 20189 22280
rect 20131 22239 20189 22240
rect 20995 22280 21053 22281
rect 20995 22240 21004 22280
rect 21044 22240 21053 22280
rect 20995 22239 21053 22240
rect 23211 22280 23253 22289
rect 23211 22240 23212 22280
rect 23252 22240 23253 22280
rect 23211 22231 23253 22240
rect 29347 22280 29405 22281
rect 29347 22240 29356 22280
rect 29396 22240 29405 22280
rect 29347 22239 29405 22240
rect 30211 22280 30269 22281
rect 30211 22240 30220 22280
rect 30260 22240 30269 22280
rect 30211 22239 30269 22240
rect 30603 22280 30645 22289
rect 30603 22240 30604 22280
rect 30644 22240 30645 22280
rect 30603 22231 30645 22240
rect 31939 22280 31997 22281
rect 31939 22240 31948 22280
rect 31988 22240 31997 22280
rect 31939 22239 31997 22240
rect 32139 22280 32181 22289
rect 32139 22240 32140 22280
rect 32180 22240 32181 22280
rect 32139 22231 32181 22240
rect 32515 22280 32573 22281
rect 32515 22240 32524 22280
rect 32564 22240 32573 22280
rect 32515 22239 32573 22240
rect 33379 22280 33437 22281
rect 33379 22240 33388 22280
rect 33428 22240 33437 22280
rect 33379 22239 33437 22240
rect 42979 22280 43037 22281
rect 42979 22240 42988 22280
rect 43028 22240 43037 22280
rect 42979 22239 43037 22240
rect 43843 22280 43901 22281
rect 43843 22240 43852 22280
rect 43892 22240 43901 22280
rect 43843 22239 43901 22240
rect 47299 22280 47357 22281
rect 47299 22240 47308 22280
rect 47348 22240 47357 22280
rect 47299 22239 47357 22240
rect 48835 22280 48893 22281
rect 48835 22240 48844 22280
rect 48884 22240 48893 22280
rect 48835 22239 48893 22240
rect 49699 22280 49757 22281
rect 49699 22240 49708 22280
rect 49748 22240 49757 22280
rect 49699 22239 49757 22240
rect 11587 22196 11645 22197
rect 11587 22156 11596 22196
rect 11636 22156 11645 22196
rect 11587 22155 11645 22156
rect 14947 22196 15005 22197
rect 14947 22156 14956 22196
rect 14996 22156 15005 22196
rect 14947 22155 15005 22156
rect 15915 22196 15957 22205
rect 15915 22156 15916 22196
rect 15956 22156 15957 22196
rect 15915 22147 15957 22156
rect 16107 22196 16149 22205
rect 16107 22156 16108 22196
rect 16148 22156 16149 22196
rect 16107 22147 16149 22156
rect 42603 22196 42645 22205
rect 42603 22156 42604 22196
rect 42644 22156 42645 22196
rect 42603 22147 42645 22156
rect 48459 22196 48501 22205
rect 48459 22156 48460 22196
rect 48500 22156 48501 22196
rect 48459 22147 48501 22156
rect 3435 22112 3477 22121
rect 3435 22072 3436 22112
rect 3476 22072 3477 22112
rect 3435 22063 3477 22072
rect 30891 22112 30933 22121
rect 30891 22072 30892 22112
rect 30932 22072 30933 22112
rect 30891 22063 30933 22072
rect 31267 22112 31325 22113
rect 31267 22072 31276 22112
rect 31316 22072 31325 22112
rect 31267 22071 31325 22072
rect 42411 22112 42453 22121
rect 42411 22072 42412 22112
rect 42452 22072 42453 22112
rect 42411 22063 42453 22072
rect 50851 22112 50909 22113
rect 50851 22072 50860 22112
rect 50900 22072 50909 22112
rect 50851 22071 50909 22072
rect 576 21944 99360 21968
rect 576 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 19472 21944
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19840 21904 34592 21944
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34960 21904 49712 21944
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 50080 21904 64832 21944
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 65200 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 95072 21944
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95440 21904 99360 21944
rect 576 21880 99360 21904
rect 5059 21776 5117 21777
rect 5059 21736 5068 21776
rect 5108 21736 5117 21776
rect 5059 21735 5117 21736
rect 15235 21776 15293 21777
rect 15235 21736 15244 21776
rect 15284 21736 15293 21776
rect 15235 21735 15293 21736
rect 32707 21776 32765 21777
rect 32707 21736 32716 21776
rect 32756 21736 32765 21776
rect 32707 21735 32765 21736
rect 33763 21776 33821 21777
rect 33763 21736 33772 21776
rect 33812 21736 33821 21776
rect 33763 21735 33821 21736
rect 48075 21776 48117 21785
rect 48075 21736 48076 21776
rect 48116 21736 48117 21776
rect 48075 21727 48117 21736
rect 49035 21776 49077 21785
rect 49035 21736 49036 21776
rect 49076 21736 49077 21776
rect 49035 21727 49077 21736
rect 2667 21692 2709 21701
rect 2667 21652 2668 21692
rect 2708 21652 2709 21692
rect 2667 21643 2709 21652
rect 21955 21692 22013 21693
rect 21955 21652 21964 21692
rect 22004 21652 22013 21692
rect 21955 21651 22013 21652
rect 22731 21692 22773 21701
rect 22731 21652 22732 21692
rect 22772 21652 22773 21692
rect 22731 21643 22773 21652
rect 30315 21692 30357 21701
rect 30315 21652 30316 21692
rect 30356 21652 30357 21692
rect 30315 21643 30357 21652
rect 37419 21692 37461 21701
rect 37419 21652 37420 21692
rect 37460 21652 37461 21692
rect 37419 21643 37461 21652
rect 3043 21608 3101 21609
rect 3043 21568 3052 21608
rect 3092 21568 3101 21608
rect 3043 21567 3101 21568
rect 3907 21608 3965 21609
rect 3907 21568 3916 21608
rect 3956 21568 3965 21608
rect 3907 21567 3965 21568
rect 15907 21608 15965 21609
rect 15907 21568 15916 21608
rect 15956 21568 15965 21608
rect 15907 21567 15965 21568
rect 21667 21608 21725 21609
rect 21667 21568 21676 21608
rect 21716 21568 21725 21608
rect 21667 21567 21725 21568
rect 22051 21608 22109 21609
rect 22051 21568 22060 21608
rect 22100 21568 22109 21608
rect 22051 21567 22109 21568
rect 22435 21608 22493 21609
rect 22435 21568 22444 21608
rect 22484 21568 22493 21608
rect 22435 21567 22493 21568
rect 22635 21608 22677 21617
rect 22635 21568 22636 21608
rect 22676 21568 22677 21608
rect 22635 21559 22677 21568
rect 22819 21608 22877 21609
rect 22819 21568 22828 21608
rect 22868 21568 22877 21608
rect 22819 21567 22877 21568
rect 30691 21608 30749 21609
rect 30691 21568 30700 21608
rect 30740 21568 30749 21608
rect 30691 21567 30749 21568
rect 31555 21608 31613 21609
rect 31555 21568 31564 21608
rect 31604 21568 31613 21608
rect 31555 21567 31613 21568
rect 33859 21608 33917 21609
rect 33859 21568 33868 21608
rect 33908 21568 33917 21608
rect 33859 21567 33917 21568
rect 37795 21608 37853 21609
rect 37795 21568 37804 21608
rect 37844 21568 37853 21608
rect 37795 21567 37853 21568
rect 38659 21608 38717 21609
rect 38659 21568 38668 21608
rect 38708 21568 38717 21608
rect 38659 21567 38717 21568
rect 50083 21608 50141 21609
rect 50083 21568 50092 21608
rect 50132 21568 50141 21608
rect 50083 21567 50141 21568
rect 50947 21608 51005 21609
rect 50947 21568 50956 21608
rect 50996 21568 51005 21608
rect 50947 21567 51005 21568
rect 48259 21524 48317 21525
rect 48259 21484 48268 21524
rect 48308 21484 48317 21524
rect 48259 21483 48317 21484
rect 49219 21524 49277 21525
rect 49219 21484 49228 21524
rect 49268 21484 49277 21524
rect 49219 21483 49277 21484
rect 50283 21524 50325 21533
rect 50283 21484 50284 21524
rect 50324 21484 50325 21524
rect 50283 21475 50325 21484
rect 20995 21440 21053 21441
rect 20995 21400 21004 21440
rect 21044 21400 21053 21440
rect 20995 21399 21053 21400
rect 39811 21440 39869 21441
rect 39811 21400 39820 21440
rect 39860 21400 39869 21440
rect 39811 21399 39869 21400
rect 49411 21440 49469 21441
rect 49411 21400 49420 21440
rect 49460 21400 49469 21440
rect 49411 21399 49469 21400
rect 34051 21356 34109 21357
rect 34051 21316 34060 21356
rect 34100 21316 34109 21356
rect 34051 21315 34109 21316
rect 576 21188 99360 21212
rect 576 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 18232 21188
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18600 21148 33352 21188
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33720 21148 48472 21188
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48840 21148 63592 21188
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63960 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 93832 21188
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 94200 21148 99360 21188
rect 576 21124 99360 21148
rect 10155 21020 10197 21029
rect 10155 20980 10156 21020
rect 10196 20980 10197 21020
rect 10155 20971 10197 20980
rect 651 20936 693 20945
rect 651 20896 652 20936
rect 692 20896 693 20936
rect 651 20887 693 20896
rect 26083 20852 26141 20853
rect 26083 20812 26092 20852
rect 26132 20812 26141 20852
rect 26083 20811 26141 20812
rect 26859 20852 26901 20861
rect 26859 20812 26860 20852
rect 26900 20812 26901 20852
rect 26859 20803 26901 20812
rect 9859 20768 9917 20769
rect 9859 20728 9868 20768
rect 9908 20728 9917 20768
rect 9859 20727 9917 20728
rect 14571 20768 14613 20777
rect 14571 20728 14572 20768
rect 14612 20728 14613 20768
rect 14571 20719 14613 20728
rect 27523 20768 27581 20769
rect 27523 20728 27532 20768
rect 27572 20728 27581 20768
rect 27523 20727 27581 20728
rect 38947 20768 39005 20769
rect 38947 20728 38956 20768
rect 38996 20728 39005 20768
rect 38947 20727 39005 20728
rect 39627 20768 39669 20777
rect 39627 20728 39628 20768
rect 39668 20728 39669 20768
rect 39627 20719 39669 20728
rect 40483 20768 40541 20769
rect 40483 20728 40492 20768
rect 40532 20728 40541 20768
rect 40483 20727 40541 20728
rect 14187 20600 14229 20609
rect 14187 20560 14188 20600
rect 14228 20560 14229 20600
rect 14187 20551 14229 20560
rect 25899 20600 25941 20609
rect 25899 20560 25900 20600
rect 25940 20560 25941 20600
rect 25899 20551 25941 20560
rect 39811 20600 39869 20601
rect 39811 20560 39820 20600
rect 39860 20560 39869 20600
rect 39811 20559 39869 20560
rect 576 20432 99360 20456
rect 576 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 19472 20432
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19840 20392 34592 20432
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34960 20392 49712 20432
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 50080 20392 64832 20432
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 65200 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 95072 20432
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95440 20392 99360 20432
rect 576 20368 99360 20392
rect 27331 20264 27389 20265
rect 27331 20224 27340 20264
rect 27380 20224 27389 20264
rect 27331 20223 27389 20224
rect 24939 20180 24981 20189
rect 24939 20140 24940 20180
rect 24980 20140 24981 20180
rect 24939 20131 24981 20140
rect 49803 20180 49845 20189
rect 49803 20140 49804 20180
rect 49844 20140 49845 20180
rect 49803 20131 49845 20140
rect 8715 20096 8757 20105
rect 8715 20056 8716 20096
rect 8756 20056 8757 20096
rect 8715 20047 8757 20056
rect 9091 20096 9149 20097
rect 9091 20056 9100 20096
rect 9140 20056 9149 20096
rect 9091 20055 9149 20056
rect 9955 20096 10013 20097
rect 9955 20056 9964 20096
rect 10004 20056 10013 20096
rect 9955 20055 10013 20056
rect 13035 20096 13077 20105
rect 13035 20056 13036 20096
rect 13076 20056 13077 20096
rect 13035 20047 13077 20056
rect 13411 20096 13469 20097
rect 13411 20056 13420 20096
rect 13460 20056 13469 20096
rect 13411 20055 13469 20056
rect 14275 20096 14333 20097
rect 14275 20056 14284 20096
rect 14324 20056 14333 20096
rect 14275 20055 14333 20056
rect 21091 20096 21149 20097
rect 21091 20056 21100 20096
rect 21140 20056 21149 20096
rect 21091 20055 21149 20056
rect 25315 20096 25373 20097
rect 25315 20056 25324 20096
rect 25364 20056 25373 20096
rect 25315 20055 25373 20056
rect 26179 20096 26237 20097
rect 26179 20056 26188 20096
rect 26228 20056 26237 20096
rect 26179 20055 26237 20056
rect 29155 20096 29213 20097
rect 29155 20056 29164 20096
rect 29204 20056 29213 20096
rect 29155 20055 29213 20056
rect 30115 20096 30173 20097
rect 30115 20056 30124 20096
rect 30164 20056 30173 20096
rect 30115 20055 30173 20056
rect 30499 20096 30557 20097
rect 30499 20056 30508 20096
rect 30548 20056 30557 20096
rect 30499 20055 30557 20056
rect 31459 20096 31517 20097
rect 31459 20056 31468 20096
rect 31508 20056 31517 20096
rect 31459 20055 31517 20056
rect 36075 20096 36117 20105
rect 36075 20056 36076 20096
rect 36116 20056 36117 20096
rect 36075 20047 36117 20056
rect 36451 20096 36509 20097
rect 36451 20056 36460 20096
rect 36500 20056 36509 20096
rect 36451 20055 36509 20056
rect 37315 20096 37373 20097
rect 37315 20056 37324 20096
rect 37364 20056 37373 20096
rect 37315 20055 37373 20056
rect 39723 20096 39765 20105
rect 39723 20056 39724 20096
rect 39764 20056 39765 20096
rect 39723 20047 39765 20056
rect 39819 20096 39861 20105
rect 39819 20056 39820 20096
rect 39860 20056 39861 20096
rect 39819 20047 39861 20056
rect 39907 20096 39965 20097
rect 39907 20056 39916 20096
rect 39956 20056 39965 20096
rect 39907 20055 39965 20056
rect 40579 20096 40637 20097
rect 40579 20056 40588 20096
rect 40628 20056 40637 20096
rect 40579 20055 40637 20056
rect 40675 20096 40733 20097
rect 40675 20056 40684 20096
rect 40724 20056 40733 20096
rect 40675 20055 40733 20056
rect 41731 20096 41789 20097
rect 41731 20056 41740 20096
rect 41780 20056 41789 20096
rect 41731 20055 41789 20056
rect 48171 20096 48213 20105
rect 48171 20056 48172 20096
rect 48212 20056 48213 20096
rect 48171 20047 48213 20056
rect 48835 20096 48893 20097
rect 48835 20056 48844 20096
rect 48884 20056 48893 20096
rect 48835 20055 48893 20056
rect 49315 20096 49373 20097
rect 49315 20056 49324 20096
rect 49364 20056 49373 20096
rect 49315 20055 49373 20056
rect 49515 20096 49557 20105
rect 49515 20056 49516 20096
rect 49556 20056 49557 20096
rect 49515 20047 49557 20056
rect 49699 20096 49757 20097
rect 49699 20056 49708 20096
rect 49748 20056 49757 20096
rect 49699 20055 49757 20056
rect 49899 20096 49941 20105
rect 49899 20056 49900 20096
rect 49940 20056 49941 20096
rect 49899 20047 49941 20056
rect 11115 20012 11157 20021
rect 11115 19972 11116 20012
rect 11156 19972 11157 20012
rect 11115 19963 11157 19972
rect 15435 20012 15477 20021
rect 15435 19972 15436 20012
rect 15476 19972 15477 20012
rect 15435 19963 15477 19972
rect 40867 20012 40925 20013
rect 40867 19972 40876 20012
rect 40916 19972 40925 20012
rect 40867 19971 40925 19972
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 20419 19844 20477 19845
rect 20419 19804 20428 19844
rect 20468 19804 20477 19844
rect 20419 19803 20477 19804
rect 29835 19844 29877 19853
rect 29835 19804 29836 19844
rect 29876 19804 29877 19844
rect 29835 19795 29877 19804
rect 30795 19844 30837 19853
rect 30795 19804 30796 19844
rect 30836 19804 30837 19844
rect 30795 19795 30837 19804
rect 38467 19844 38525 19845
rect 38467 19804 38476 19844
rect 38516 19804 38525 19844
rect 38467 19803 38525 19804
rect 41059 19844 41117 19845
rect 41059 19804 41068 19844
rect 41108 19804 41117 19844
rect 41059 19803 41117 19804
rect 49419 19844 49461 19853
rect 49419 19804 49420 19844
rect 49460 19804 49461 19844
rect 49419 19795 49461 19804
rect 576 19676 99360 19700
rect 576 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 18232 19676
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18600 19636 33352 19676
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33720 19636 48472 19676
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48840 19636 63592 19676
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63960 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 93832 19676
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 94200 19636 99360 19676
rect 576 19612 99360 19636
rect 3619 19508 3677 19509
rect 3619 19468 3628 19508
rect 3668 19468 3677 19508
rect 3619 19467 3677 19468
rect 48739 19508 48797 19509
rect 48739 19468 48748 19508
rect 48788 19468 48797 19508
rect 48739 19467 48797 19468
rect 651 19424 693 19433
rect 651 19384 652 19424
rect 692 19384 693 19424
rect 651 19375 693 19384
rect 2851 19340 2909 19341
rect 2851 19300 2860 19340
rect 2900 19300 2909 19340
rect 2851 19299 2909 19300
rect 4291 19256 4349 19257
rect 4291 19216 4300 19256
rect 4340 19216 4349 19256
rect 4291 19215 4349 19216
rect 26571 19256 26613 19265
rect 26571 19216 26572 19256
rect 26612 19216 26613 19256
rect 26571 19207 26613 19216
rect 26755 19256 26813 19257
rect 26755 19216 26764 19256
rect 26804 19216 26813 19256
rect 26755 19215 26813 19216
rect 27619 19256 27677 19257
rect 27619 19216 27628 19256
rect 27668 19216 27677 19256
rect 27619 19215 27677 19216
rect 34915 19256 34973 19257
rect 34915 19216 34924 19256
rect 34964 19216 34973 19256
rect 34915 19215 34973 19216
rect 39331 19256 39389 19257
rect 39331 19216 39340 19256
rect 39380 19216 39389 19256
rect 39331 19215 39389 19216
rect 39715 19256 39773 19257
rect 39715 19216 39724 19256
rect 39764 19216 39773 19256
rect 39715 19215 39773 19216
rect 46723 19256 46781 19257
rect 46723 19216 46732 19256
rect 46772 19216 46781 19256
rect 46723 19215 46781 19216
rect 47587 19256 47645 19257
rect 47587 19216 47596 19256
rect 47636 19216 47645 19256
rect 47587 19215 47645 19216
rect 50179 19256 50237 19257
rect 50179 19216 50188 19256
rect 50228 19216 50237 19256
rect 50179 19215 50237 19216
rect 50467 19256 50525 19257
rect 50467 19216 50476 19256
rect 50516 19216 50525 19256
rect 50467 19215 50525 19216
rect 26667 19172 26709 19181
rect 26667 19132 26668 19172
rect 26708 19132 26709 19172
rect 26667 19123 26709 19132
rect 46347 19172 46389 19181
rect 46347 19132 46348 19172
rect 46388 19132 46389 19172
rect 46347 19123 46389 19132
rect 2667 19088 2709 19097
rect 2667 19048 2668 19088
rect 2708 19048 2709 19088
rect 2667 19039 2709 19048
rect 26947 19088 27005 19089
rect 26947 19048 26956 19088
rect 26996 19048 27005 19088
rect 26947 19047 27005 19048
rect 35403 19088 35445 19097
rect 35403 19048 35404 19088
rect 35444 19048 35445 19088
rect 35403 19039 35445 19048
rect 39819 19088 39861 19097
rect 39819 19048 39820 19088
rect 39860 19048 39861 19088
rect 39819 19039 39861 19048
rect 50667 19088 50709 19097
rect 50667 19048 50668 19088
rect 50708 19048 50709 19088
rect 50667 19039 50709 19048
rect 576 18920 99360 18944
rect 576 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 19472 18920
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19840 18880 34592 18920
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34960 18880 49712 18920
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 50080 18880 64832 18920
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 65200 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 95072 18920
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95440 18880 99360 18920
rect 576 18856 99360 18880
rect 4099 18752 4157 18753
rect 4099 18712 4108 18752
rect 4148 18712 4157 18752
rect 4099 18711 4157 18712
rect 7467 18752 7509 18761
rect 7467 18712 7468 18752
rect 7508 18712 7509 18752
rect 7467 18703 7509 18712
rect 8715 18752 8757 18761
rect 8715 18712 8716 18752
rect 8756 18712 8757 18752
rect 8715 18703 8757 18712
rect 11779 18752 11837 18753
rect 11779 18712 11788 18752
rect 11828 18712 11837 18752
rect 11779 18711 11837 18712
rect 12067 18752 12125 18753
rect 12067 18712 12076 18752
rect 12116 18712 12125 18752
rect 12067 18711 12125 18712
rect 12259 18752 12317 18753
rect 12259 18712 12268 18752
rect 12308 18712 12317 18752
rect 12259 18711 12317 18712
rect 27523 18752 27581 18753
rect 27523 18712 27532 18752
rect 27572 18712 27581 18752
rect 27523 18711 27581 18712
rect 1707 18668 1749 18677
rect 1707 18628 1708 18668
rect 1748 18628 1749 18668
rect 1707 18619 1749 18628
rect 19755 18668 19797 18677
rect 19755 18628 19756 18668
rect 19796 18628 19797 18668
rect 19755 18619 19797 18628
rect 41067 18668 41109 18677
rect 41067 18628 41068 18668
rect 41108 18628 41109 18668
rect 41067 18619 41109 18628
rect 52011 18668 52053 18677
rect 52011 18628 52012 18668
rect 52052 18628 52053 18668
rect 52011 18619 52053 18628
rect 2083 18584 2141 18585
rect 2083 18544 2092 18584
rect 2132 18544 2141 18584
rect 2083 18543 2141 18544
rect 2947 18584 3005 18585
rect 2947 18544 2956 18584
rect 2996 18544 3005 18584
rect 2947 18543 3005 18544
rect 6979 18584 7037 18585
rect 6979 18544 6988 18584
rect 7028 18544 7037 18584
rect 6979 18543 7037 18544
rect 7939 18584 7997 18585
rect 7939 18544 7948 18584
rect 7988 18544 7997 18584
rect 7939 18543 7997 18544
rect 8227 18584 8285 18585
rect 8227 18544 8236 18584
rect 8276 18544 8285 18584
rect 8227 18543 8285 18544
rect 8611 18584 8669 18585
rect 8611 18544 8620 18584
rect 8660 18544 8669 18584
rect 8611 18543 8669 18544
rect 11875 18584 11933 18585
rect 11875 18544 11884 18584
rect 11924 18544 11933 18584
rect 11875 18543 11933 18544
rect 12931 18584 12989 18585
rect 12931 18544 12940 18584
rect 12980 18544 12989 18584
rect 12931 18543 12989 18544
rect 18499 18584 18557 18585
rect 18499 18544 18508 18584
rect 18548 18544 18557 18584
rect 18499 18543 18557 18544
rect 19363 18584 19421 18585
rect 19363 18544 19372 18584
rect 19412 18544 19421 18584
rect 19363 18543 19421 18544
rect 23491 18584 23549 18585
rect 23491 18544 23500 18584
rect 23540 18544 23549 18584
rect 23491 18543 23549 18544
rect 25131 18584 25173 18593
rect 25131 18544 25132 18584
rect 25172 18544 25173 18584
rect 25131 18535 25173 18544
rect 25507 18584 25565 18585
rect 25507 18544 25516 18584
rect 25556 18544 25565 18584
rect 25507 18543 25565 18544
rect 26371 18584 26429 18585
rect 26371 18544 26380 18584
rect 26420 18544 26429 18584
rect 26371 18543 26429 18544
rect 40675 18584 40733 18585
rect 40675 18544 40684 18584
rect 40724 18544 40733 18584
rect 40675 18543 40733 18544
rect 41443 18584 41501 18585
rect 41443 18544 41452 18584
rect 41492 18544 41501 18584
rect 41443 18543 41501 18544
rect 42307 18584 42365 18585
rect 42307 18544 42316 18584
rect 42356 18544 42365 18584
rect 42307 18543 42365 18544
rect 46731 18584 46773 18593
rect 46731 18544 46732 18584
rect 46772 18544 46773 18584
rect 46731 18535 46773 18544
rect 47107 18584 47165 18585
rect 47107 18544 47116 18584
rect 47156 18544 47165 18584
rect 47107 18543 47165 18544
rect 47971 18584 48029 18585
rect 47971 18544 47980 18584
rect 48020 18544 48029 18584
rect 47971 18543 48029 18544
rect 52387 18584 52445 18585
rect 52387 18544 52396 18584
rect 52436 18544 52445 18584
rect 52387 18543 52445 18544
rect 53251 18584 53309 18585
rect 53251 18544 53260 18584
rect 53300 18544 53309 18584
rect 53251 18543 53309 18544
rect 6787 18500 6845 18501
rect 6787 18460 6796 18500
rect 6836 18460 6845 18500
rect 6787 18459 6845 18460
rect 651 18416 693 18425
rect 651 18376 652 18416
rect 692 18376 693 18416
rect 651 18367 693 18376
rect 6603 18332 6645 18341
rect 6603 18292 6604 18332
rect 6644 18292 6645 18332
rect 6603 18283 6645 18292
rect 17347 18332 17405 18333
rect 17347 18292 17356 18332
rect 17396 18292 17405 18332
rect 17347 18291 17405 18292
rect 22819 18332 22877 18333
rect 22819 18292 22828 18332
rect 22868 18292 22877 18332
rect 22819 18291 22877 18292
rect 40003 18332 40061 18333
rect 40003 18292 40012 18332
rect 40052 18292 40061 18332
rect 40003 18291 40061 18292
rect 43459 18332 43517 18333
rect 43459 18292 43468 18332
rect 43508 18292 43517 18332
rect 43459 18291 43517 18292
rect 49123 18332 49181 18333
rect 49123 18292 49132 18332
rect 49172 18292 49181 18332
rect 49123 18291 49181 18292
rect 54403 18332 54461 18333
rect 54403 18292 54412 18332
rect 54452 18292 54461 18332
rect 54403 18291 54461 18292
rect 576 18164 99360 18188
rect 576 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 18232 18164
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18600 18124 33352 18164
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33720 18124 48472 18164
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48840 18124 63592 18164
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63960 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 93832 18164
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 94200 18124 99360 18164
rect 576 18100 99360 18124
rect 7651 17996 7709 17997
rect 7651 17956 7660 17996
rect 7700 17956 7709 17996
rect 7651 17955 7709 17956
rect 13315 17996 13373 17997
rect 13315 17956 13324 17996
rect 13364 17956 13373 17996
rect 13315 17955 13373 17956
rect 23395 17996 23453 17997
rect 23395 17956 23404 17996
rect 23444 17956 23453 17996
rect 23395 17955 23453 17956
rect 25899 17996 25941 18005
rect 25899 17956 25900 17996
rect 25940 17956 25941 17996
rect 25899 17947 25941 17956
rect 47211 17996 47253 18005
rect 47211 17956 47212 17996
rect 47252 17956 47253 17996
rect 47211 17947 47253 17956
rect 47595 17996 47637 18005
rect 47595 17956 47596 17996
rect 47636 17956 47637 17996
rect 47595 17947 47637 17956
rect 48547 17996 48605 17997
rect 48547 17956 48556 17996
rect 48596 17956 48605 17996
rect 48547 17955 48605 17956
rect 651 17912 693 17921
rect 651 17872 652 17912
rect 692 17872 693 17912
rect 651 17863 693 17872
rect 24643 17912 24701 17913
rect 24643 17872 24652 17912
rect 24692 17872 24701 17912
rect 24643 17871 24701 17872
rect 6507 17828 6549 17837
rect 6507 17788 6508 17828
rect 6548 17788 6549 17828
rect 6507 17779 6549 17788
rect 23971 17828 24029 17829
rect 23971 17788 23980 17828
rect 24020 17788 24029 17828
rect 23971 17787 24029 17788
rect 26083 17828 26141 17829
rect 26083 17788 26092 17828
rect 26132 17788 26141 17828
rect 26083 17787 26141 17788
rect 32331 17828 32373 17837
rect 32331 17788 32332 17828
rect 32372 17788 32373 17828
rect 32331 17779 32373 17788
rect 47395 17828 47453 17829
rect 47395 17788 47404 17828
rect 47444 17788 47453 17828
rect 47395 17787 47453 17788
rect 47779 17828 47837 17829
rect 47779 17788 47788 17828
rect 47828 17788 47837 17828
rect 47779 17787 47837 17788
rect 26678 17759 26720 17768
rect 4483 17744 4541 17745
rect 4483 17704 4492 17744
rect 4532 17704 4541 17744
rect 4483 17703 4541 17704
rect 5347 17744 5405 17745
rect 5347 17704 5356 17744
rect 5396 17704 5405 17744
rect 5347 17703 5405 17704
rect 6691 17744 6749 17745
rect 6691 17704 6700 17744
rect 6740 17704 6749 17744
rect 6691 17703 6749 17704
rect 8323 17744 8381 17745
rect 8323 17704 8332 17744
rect 8372 17704 8381 17744
rect 8323 17703 8381 17704
rect 8811 17744 8853 17753
rect 8811 17704 8812 17744
rect 8852 17704 8853 17744
rect 8811 17695 8853 17704
rect 8995 17744 9053 17745
rect 8995 17704 9004 17744
rect 9044 17704 9053 17744
rect 8995 17703 9053 17704
rect 11299 17744 11357 17745
rect 11299 17704 11308 17744
rect 11348 17704 11357 17744
rect 11299 17703 11357 17704
rect 12163 17744 12221 17745
rect 12163 17704 12172 17744
rect 12212 17704 12221 17744
rect 12163 17703 12221 17704
rect 18979 17744 19037 17745
rect 18979 17704 18988 17744
rect 19028 17704 19037 17744
rect 18979 17703 19037 17704
rect 21379 17744 21437 17745
rect 21379 17704 21388 17744
rect 21428 17704 21437 17744
rect 21379 17703 21437 17704
rect 22243 17744 22301 17745
rect 22243 17704 22252 17744
rect 22292 17704 22301 17744
rect 22243 17703 22301 17704
rect 25315 17744 25373 17745
rect 25315 17704 25324 17744
rect 25364 17704 25373 17744
rect 25315 17703 25373 17704
rect 26475 17744 26517 17753
rect 26475 17704 26476 17744
rect 26516 17704 26517 17744
rect 26475 17695 26517 17704
rect 26571 17744 26613 17753
rect 26571 17704 26572 17744
rect 26612 17704 26613 17744
rect 26678 17719 26679 17759
rect 26719 17719 26720 17759
rect 26678 17710 26720 17719
rect 27142 17744 27200 17745
rect 26571 17695 26613 17704
rect 27142 17704 27151 17744
rect 27191 17704 27200 17744
rect 27142 17703 27200 17704
rect 27523 17744 27581 17745
rect 27523 17704 27532 17744
rect 27572 17704 27581 17744
rect 27523 17703 27581 17704
rect 27811 17744 27869 17745
rect 27811 17704 27820 17744
rect 27860 17704 27869 17744
rect 27811 17703 27869 17704
rect 30307 17744 30365 17745
rect 30307 17704 30316 17744
rect 30356 17704 30365 17744
rect 30307 17703 30365 17704
rect 31171 17744 31229 17745
rect 31171 17704 31180 17744
rect 31220 17704 31229 17744
rect 31171 17703 31229 17704
rect 41443 17744 41501 17745
rect 41443 17704 41452 17744
rect 41492 17704 41501 17744
rect 41443 17703 41501 17704
rect 41827 17744 41885 17745
rect 41827 17704 41836 17744
rect 41876 17704 41885 17744
rect 41827 17703 41885 17704
rect 48163 17744 48221 17745
rect 48163 17704 48172 17744
rect 48212 17704 48221 17744
rect 48163 17703 48221 17704
rect 49219 17744 49277 17745
rect 49219 17704 49228 17744
rect 49268 17704 49277 17744
rect 49219 17703 49277 17704
rect 4107 17660 4149 17669
rect 4107 17620 4108 17660
rect 4148 17620 4149 17660
rect 4107 17611 4149 17620
rect 7371 17660 7413 17669
rect 7371 17620 7372 17660
rect 7412 17620 7413 17660
rect 7371 17611 7413 17620
rect 8907 17660 8949 17669
rect 8907 17620 8908 17660
rect 8948 17620 8949 17660
rect 8907 17611 8949 17620
rect 10923 17660 10965 17669
rect 10923 17620 10924 17660
rect 10964 17620 10965 17660
rect 10923 17611 10965 17620
rect 21003 17660 21045 17669
rect 21003 17620 21004 17660
rect 21044 17620 21045 17660
rect 21003 17611 21045 17620
rect 28003 17660 28061 17661
rect 28003 17620 28012 17660
rect 28052 17620 28061 17660
rect 28003 17619 28061 17620
rect 29931 17660 29973 17669
rect 29931 17620 29932 17660
rect 29972 17620 29973 17660
rect 29931 17611 29973 17620
rect 41923 17660 41981 17661
rect 41923 17620 41932 17660
rect 41972 17620 41981 17660
rect 41923 17619 41981 17620
rect 23787 17576 23829 17585
rect 23787 17536 23788 17576
rect 23828 17536 23829 17576
rect 23787 17527 23829 17536
rect 27043 17576 27101 17577
rect 27043 17536 27052 17576
rect 27092 17536 27101 17576
rect 27043 17535 27101 17536
rect 27331 17576 27389 17577
rect 27331 17536 27340 17576
rect 27380 17536 27389 17576
rect 27331 17535 27389 17536
rect 48067 17576 48125 17577
rect 48067 17536 48076 17576
rect 48116 17536 48125 17576
rect 48067 17535 48125 17536
rect 48355 17576 48413 17577
rect 48355 17536 48364 17576
rect 48404 17536 48413 17576
rect 48355 17535 48413 17536
rect 576 17408 99360 17432
rect 576 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 19472 17408
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19840 17368 34592 17408
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34960 17368 49712 17408
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 50080 17368 64832 17408
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 65200 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 95072 17408
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95440 17368 99360 17408
rect 576 17344 99360 17368
rect 5259 17240 5301 17249
rect 5259 17200 5260 17240
rect 5300 17200 5301 17240
rect 5259 17191 5301 17200
rect 8035 17240 8093 17241
rect 8035 17200 8044 17240
rect 8084 17200 8093 17240
rect 8035 17199 8093 17200
rect 10539 17240 10581 17249
rect 10539 17200 10540 17240
rect 10580 17200 10581 17240
rect 10539 17191 10581 17200
rect 21771 17240 21813 17249
rect 21771 17200 21772 17240
rect 21812 17200 21813 17240
rect 21771 17191 21813 17200
rect 25123 17240 25181 17241
rect 25123 17200 25132 17240
rect 25172 17200 25181 17240
rect 25123 17199 25181 17200
rect 39619 17240 39677 17241
rect 39619 17200 39628 17240
rect 39668 17200 39677 17240
rect 39619 17199 39677 17200
rect 54987 17240 55029 17249
rect 54987 17200 54988 17240
rect 55028 17200 55029 17240
rect 54987 17191 55029 17200
rect 5643 17156 5685 17165
rect 5643 17116 5644 17156
rect 5684 17116 5685 17156
rect 5643 17107 5685 17116
rect 8331 17156 8373 17165
rect 8331 17116 8332 17156
rect 8372 17116 8373 17156
rect 8331 17107 8373 17116
rect 10731 17156 10773 17165
rect 10731 17116 10732 17156
rect 10772 17116 10773 17156
rect 10731 17107 10773 17116
rect 18891 17156 18933 17165
rect 18891 17116 18892 17156
rect 18932 17116 18933 17156
rect 18891 17107 18933 17116
rect 22731 17156 22773 17165
rect 22731 17116 22732 17156
rect 22772 17116 22773 17156
rect 22731 17107 22773 17116
rect 30987 17156 31029 17165
rect 30987 17116 30988 17156
rect 31028 17116 31029 17156
rect 30987 17107 31029 17116
rect 34051 17156 34109 17157
rect 34051 17116 34060 17156
rect 34100 17116 34109 17156
rect 34051 17115 34109 17116
rect 40011 17156 40053 17165
rect 40011 17116 40012 17156
rect 40052 17116 40053 17156
rect 40011 17107 40053 17116
rect 6019 17072 6077 17073
rect 6019 17032 6028 17072
rect 6068 17032 6077 17072
rect 6019 17031 6077 17032
rect 6883 17072 6941 17073
rect 6883 17032 6892 17072
rect 6932 17032 6941 17072
rect 6883 17031 6941 17032
rect 8235 17072 8277 17081
rect 8235 17032 8236 17072
rect 8276 17032 8277 17072
rect 8235 17023 8277 17032
rect 8419 17072 8477 17073
rect 8419 17032 8428 17072
rect 8468 17032 8477 17072
rect 8419 17031 8477 17032
rect 11107 17072 11165 17073
rect 11107 17032 11116 17072
rect 11156 17032 11165 17072
rect 11107 17031 11165 17032
rect 11971 17072 12029 17073
rect 11971 17032 11980 17072
rect 12020 17032 12029 17072
rect 11971 17031 12029 17032
rect 17635 17072 17693 17073
rect 17635 17032 17644 17072
rect 17684 17032 17693 17072
rect 17635 17031 17693 17032
rect 18499 17072 18557 17073
rect 18499 17032 18508 17072
rect 18548 17032 18557 17072
rect 18499 17031 18557 17032
rect 19171 17072 19229 17073
rect 19171 17032 19180 17072
rect 19220 17032 19229 17072
rect 19171 17031 19229 17032
rect 23107 17072 23165 17073
rect 23107 17032 23116 17072
rect 23156 17032 23165 17072
rect 23107 17031 23165 17032
rect 23971 17072 24029 17073
rect 23971 17032 23980 17072
rect 24020 17032 24029 17072
rect 23971 17031 24029 17032
rect 31363 17072 31421 17073
rect 31363 17032 31372 17072
rect 31412 17032 31421 17072
rect 31363 17031 31421 17032
rect 32227 17072 32285 17073
rect 32227 17032 32236 17072
rect 32276 17032 32285 17072
rect 32227 17031 32285 17032
rect 33571 17072 33629 17073
rect 33571 17032 33580 17072
rect 33620 17032 33629 17072
rect 33571 17031 33629 17032
rect 33859 17072 33917 17073
rect 33859 17032 33868 17072
rect 33908 17032 33917 17072
rect 33859 17031 33917 17032
rect 36355 17072 36413 17073
rect 36355 17032 36364 17072
rect 36404 17032 36413 17072
rect 36355 17031 36413 17032
rect 37035 17072 37077 17081
rect 37035 17032 37036 17072
rect 37076 17032 37077 17072
rect 37035 17023 37077 17032
rect 37227 17072 37269 17081
rect 37227 17032 37228 17072
rect 37268 17032 37269 17072
rect 37227 17023 37269 17032
rect 37603 17072 37661 17073
rect 37603 17032 37612 17072
rect 37652 17032 37661 17072
rect 37603 17031 37661 17032
rect 38467 17072 38525 17073
rect 38467 17032 38476 17072
rect 38516 17032 38525 17072
rect 38467 17031 38525 17032
rect 40387 17072 40445 17073
rect 40387 17032 40396 17072
rect 40436 17032 40445 17072
rect 40387 17031 40445 17032
rect 41251 17072 41309 17073
rect 41251 17032 41260 17072
rect 41300 17032 41309 17072
rect 41251 17031 41309 17032
rect 54499 17072 54557 17073
rect 54499 17032 54508 17072
rect 54548 17032 54557 17072
rect 54499 17031 54557 17032
rect 54883 17072 54941 17073
rect 54883 17032 54892 17072
rect 54932 17032 54941 17072
rect 54883 17031 54941 17032
rect 56419 17072 56477 17073
rect 56419 17032 56428 17072
rect 56468 17032 56477 17072
rect 56419 17031 56477 17032
rect 57283 17072 57341 17073
rect 57283 17032 57292 17072
rect 57332 17032 57341 17072
rect 57283 17031 57341 17032
rect 57675 17072 57717 17081
rect 57675 17032 57676 17072
rect 57716 17032 57717 17072
rect 57675 17023 57717 17032
rect 5443 16988 5501 16989
rect 5443 16948 5452 16988
rect 5492 16948 5501 16988
rect 5443 16947 5501 16948
rect 10339 16988 10397 16989
rect 10339 16948 10348 16988
rect 10388 16948 10397 16988
rect 10339 16947 10397 16948
rect 21955 16988 22013 16989
rect 21955 16948 21964 16988
rect 22004 16948 22013 16988
rect 21955 16947 22013 16948
rect 55275 16988 55317 16997
rect 55275 16948 55276 16988
rect 55316 16948 55317 16988
rect 55275 16939 55317 16948
rect 651 16904 693 16913
rect 651 16864 652 16904
rect 692 16864 693 16904
rect 651 16855 693 16864
rect 19467 16904 19509 16913
rect 19467 16864 19468 16904
rect 19508 16864 19509 16904
rect 19467 16855 19509 16864
rect 13123 16820 13181 16821
rect 13123 16780 13132 16820
rect 13172 16780 13181 16820
rect 13123 16779 13181 16780
rect 16483 16820 16541 16821
rect 16483 16780 16492 16820
rect 16532 16780 16541 16820
rect 16483 16779 16541 16780
rect 33379 16820 33437 16821
rect 33379 16780 33388 16820
rect 33428 16780 33437 16820
rect 33379 16779 33437 16780
rect 42403 16820 42461 16821
rect 42403 16780 42412 16820
rect 42452 16780 42461 16820
rect 42403 16779 42461 16780
rect 576 16652 99360 16676
rect 576 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 18232 16652
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18600 16612 33352 16652
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33720 16612 48472 16652
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48840 16612 63592 16652
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63960 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 93832 16652
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 94200 16612 99360 16652
rect 576 16588 99360 16612
rect 651 16400 693 16409
rect 651 16360 652 16400
rect 692 16360 693 16400
rect 651 16351 693 16360
rect 10827 16400 10869 16409
rect 10827 16360 10828 16400
rect 10868 16360 10869 16400
rect 10827 16351 10869 16360
rect 11683 16400 11741 16401
rect 11683 16360 11692 16400
rect 11732 16360 11741 16400
rect 11683 16359 11741 16360
rect 12939 16400 12981 16409
rect 12939 16360 12940 16400
rect 12980 16360 12981 16400
rect 12939 16351 12981 16360
rect 11011 16316 11069 16317
rect 11011 16276 11020 16316
rect 11060 16276 11069 16316
rect 11011 16275 11069 16276
rect 36355 16316 36413 16317
rect 36355 16276 36364 16316
rect 36404 16276 36413 16316
rect 36355 16275 36413 16276
rect 12355 16232 12413 16233
rect 12355 16192 12364 16232
rect 12404 16192 12413 16232
rect 12355 16191 12413 16192
rect 12643 16232 12701 16233
rect 12643 16192 12652 16232
rect 12692 16192 12701 16232
rect 12643 16191 12701 16192
rect 34915 16232 34973 16233
rect 34915 16192 34924 16232
rect 34964 16192 34973 16232
rect 34915 16191 34973 16192
rect 36067 16232 36125 16233
rect 36067 16192 36076 16232
rect 36116 16192 36125 16232
rect 36067 16191 36125 16192
rect 36163 16232 36221 16233
rect 36163 16192 36172 16232
rect 36212 16192 36221 16232
rect 36163 16191 36221 16192
rect 13507 16148 13565 16149
rect 13507 16108 13516 16148
rect 13556 16108 13565 16148
rect 13507 16107 13565 16108
rect 35587 16064 35645 16065
rect 35587 16024 35596 16064
rect 35636 16024 35645 16064
rect 35587 16023 35645 16024
rect 576 15896 99360 15920
rect 576 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 19472 15896
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19840 15856 34592 15896
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34960 15856 49712 15896
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 50080 15856 64832 15896
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 65200 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 95072 15896
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95440 15856 99360 15896
rect 576 15832 99360 15856
rect 643 15728 701 15729
rect 643 15688 652 15728
rect 692 15688 701 15728
rect 643 15687 701 15688
rect 32995 15728 33053 15729
rect 32995 15688 33004 15728
rect 33044 15688 33053 15728
rect 32995 15687 33053 15688
rect 35787 15644 35829 15653
rect 35787 15604 35788 15644
rect 35828 15604 35829 15644
rect 35787 15595 35829 15604
rect 49227 15644 49269 15653
rect 49227 15604 49228 15644
rect 49268 15604 49269 15644
rect 49227 15595 49269 15604
rect 30603 15560 30645 15569
rect 30603 15520 30604 15560
rect 30644 15520 30645 15560
rect 30603 15511 30645 15520
rect 30979 15560 31037 15561
rect 30979 15520 30988 15560
rect 31028 15520 31037 15560
rect 30979 15519 31037 15520
rect 31843 15560 31901 15561
rect 31843 15520 31852 15560
rect 31892 15520 31901 15560
rect 31843 15519 31901 15520
rect 35691 15560 35733 15569
rect 35691 15520 35692 15560
rect 35732 15520 35733 15560
rect 35691 15511 35733 15520
rect 35875 15560 35933 15561
rect 35875 15520 35884 15560
rect 35924 15520 35933 15560
rect 35875 15519 35933 15520
rect 36075 15560 36117 15569
rect 36075 15520 36076 15560
rect 36116 15520 36117 15560
rect 36075 15511 36117 15520
rect 36739 15560 36797 15561
rect 36739 15520 36748 15560
rect 36788 15520 36797 15560
rect 36739 15519 36797 15520
rect 41539 15560 41597 15561
rect 41539 15520 41548 15560
rect 41588 15520 41597 15560
rect 41539 15519 41597 15520
rect 41731 15560 41789 15561
rect 41731 15520 41740 15560
rect 41780 15520 41789 15560
rect 41731 15519 41789 15520
rect 42603 15560 42645 15569
rect 42603 15520 42604 15560
rect 42644 15520 42645 15560
rect 42603 15511 42645 15520
rect 49603 15560 49661 15561
rect 49603 15520 49612 15560
rect 49652 15520 49661 15560
rect 49603 15519 49661 15520
rect 50467 15560 50525 15561
rect 50467 15520 50476 15560
rect 50516 15520 50525 15560
rect 50467 15519 50525 15520
rect 52771 15560 52829 15561
rect 52771 15520 52780 15560
rect 52820 15520 52829 15560
rect 52771 15519 52829 15520
rect 51627 15476 51669 15485
rect 51627 15436 51628 15476
rect 51668 15436 51669 15476
rect 51627 15427 51669 15436
rect 40867 15308 40925 15309
rect 40867 15268 40876 15308
rect 40916 15268 40925 15308
rect 40867 15267 40925 15268
rect 52099 15308 52157 15309
rect 52099 15268 52108 15308
rect 52148 15268 52157 15308
rect 52099 15267 52157 15268
rect 576 15140 99360 15164
rect 576 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 18232 15140
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18600 15100 33352 15140
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33720 15100 48472 15140
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48840 15100 63592 15140
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63960 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 93832 15140
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 94200 15100 99360 15140
rect 576 15076 99360 15100
rect 9483 14972 9525 14981
rect 9483 14932 9484 14972
rect 9524 14932 9525 14972
rect 9483 14923 9525 14932
rect 21867 14972 21909 14981
rect 21867 14932 21868 14972
rect 21908 14932 21909 14972
rect 21867 14923 21909 14932
rect 47115 14972 47157 14981
rect 47115 14932 47116 14972
rect 47156 14932 47157 14972
rect 47115 14923 47157 14932
rect 23115 14888 23157 14897
rect 23115 14848 23116 14888
rect 23156 14848 23157 14888
rect 23115 14839 23157 14848
rect 23499 14888 23541 14897
rect 23499 14848 23500 14888
rect 23540 14848 23541 14888
rect 23499 14839 23541 14848
rect 52579 14804 52637 14805
rect 52579 14764 52588 14804
rect 52628 14764 52637 14804
rect 52579 14763 52637 14764
rect 56995 14804 57053 14805
rect 56995 14764 57004 14804
rect 57044 14764 57053 14804
rect 56995 14763 57053 14764
rect 9763 14720 9821 14721
rect 9763 14680 9772 14720
rect 9812 14680 9821 14720
rect 9763 14679 9821 14680
rect 16483 14720 16541 14721
rect 16483 14680 16492 14720
rect 16532 14680 16541 14720
rect 16483 14679 16541 14680
rect 21675 14720 21717 14729
rect 21675 14680 21676 14720
rect 21716 14680 21717 14720
rect 21675 14671 21717 14680
rect 22923 14720 22965 14729
rect 22923 14680 22924 14720
rect 22964 14680 22965 14720
rect 22923 14671 22965 14680
rect 35971 14720 36029 14721
rect 35971 14680 35980 14720
rect 36020 14680 36029 14720
rect 35971 14679 36029 14680
rect 36259 14720 36317 14721
rect 36259 14680 36268 14720
rect 36308 14680 36317 14720
rect 36259 14679 36317 14680
rect 40779 14720 40821 14729
rect 40779 14680 40780 14720
rect 40820 14680 40821 14720
rect 40779 14671 40821 14680
rect 40875 14720 40917 14729
rect 40875 14680 40876 14720
rect 40916 14680 40917 14720
rect 40875 14671 40917 14680
rect 40963 14720 41021 14721
rect 40963 14680 40972 14720
rect 41012 14680 41021 14720
rect 40963 14679 41021 14680
rect 41443 14720 41501 14721
rect 41443 14680 41452 14720
rect 41492 14680 41501 14720
rect 41443 14679 41501 14680
rect 41539 14720 41597 14721
rect 41539 14680 41548 14720
rect 41588 14680 41597 14720
rect 41539 14679 41597 14680
rect 45091 14720 45149 14721
rect 45091 14680 45100 14720
rect 45140 14680 45149 14720
rect 45091 14679 45149 14680
rect 46051 14720 46109 14721
rect 46051 14680 46060 14720
rect 46100 14680 46109 14720
rect 46051 14679 46109 14680
rect 46627 14720 46685 14721
rect 46627 14680 46636 14720
rect 46676 14680 46685 14720
rect 46627 14679 46685 14680
rect 47587 14720 47645 14721
rect 47587 14680 47596 14720
rect 47636 14680 47645 14720
rect 47587 14679 47645 14680
rect 51243 14720 51285 14729
rect 51243 14680 51244 14720
rect 51284 14680 51285 14720
rect 51243 14671 51285 14680
rect 51427 14720 51485 14721
rect 51427 14680 51436 14720
rect 51476 14680 51485 14720
rect 51427 14679 51485 14680
rect 52291 14720 52349 14721
rect 52291 14680 52300 14720
rect 52340 14680 52349 14720
rect 52291 14679 52349 14680
rect 52771 14720 52829 14721
rect 52771 14680 52780 14720
rect 52820 14680 52829 14720
rect 52771 14679 52829 14680
rect 52867 14720 52925 14721
rect 52867 14680 52876 14720
rect 52916 14680 52925 14720
rect 52867 14679 52925 14680
rect 58627 14720 58685 14721
rect 58627 14680 58636 14720
rect 58676 14680 58685 14720
rect 58627 14679 58685 14680
rect 51339 14636 51381 14645
rect 51339 14596 51340 14636
rect 51380 14596 51381 14636
rect 51339 14587 51381 14596
rect 643 14552 701 14553
rect 643 14512 652 14552
rect 692 14512 701 14552
rect 643 14511 701 14512
rect 17155 14552 17213 14553
rect 17155 14512 17164 14552
rect 17204 14512 17213 14552
rect 17155 14511 17213 14512
rect 36459 14552 36501 14561
rect 36459 14512 36460 14552
rect 36500 14512 36501 14552
rect 36459 14503 36501 14512
rect 41259 14552 41301 14561
rect 41259 14512 41260 14552
rect 41300 14512 41301 14552
rect 41259 14503 41301 14512
rect 51619 14552 51677 14553
rect 51619 14512 51628 14552
rect 51668 14512 51677 14552
rect 51619 14511 51677 14512
rect 56811 14552 56853 14561
rect 56811 14512 56812 14552
rect 56852 14512 56853 14552
rect 56811 14503 56853 14512
rect 57955 14552 58013 14553
rect 57955 14512 57964 14552
rect 58004 14512 58013 14552
rect 57955 14511 58013 14512
rect 576 14384 99360 14408
rect 576 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 19472 14384
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19840 14344 34592 14384
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34960 14344 49712 14384
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 50080 14344 64832 14384
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 65200 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 95072 14384
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95440 14344 99360 14384
rect 576 14320 99360 14344
rect 36067 14216 36125 14217
rect 36067 14176 36076 14216
rect 36116 14176 36125 14216
rect 36067 14175 36125 14176
rect 40963 14216 41021 14217
rect 40963 14176 40972 14216
rect 41012 14176 41021 14216
rect 40963 14175 41021 14176
rect 52675 14216 52733 14217
rect 52675 14176 52684 14216
rect 52724 14176 52733 14216
rect 52675 14175 52733 14176
rect 55947 14216 55989 14225
rect 55947 14176 55948 14216
rect 55988 14176 55989 14216
rect 55947 14167 55989 14176
rect 58723 14216 58781 14217
rect 58723 14176 58732 14216
rect 58772 14176 58781 14216
rect 58723 14175 58781 14176
rect 50379 14132 50421 14141
rect 50379 14092 50380 14132
rect 50420 14092 50421 14132
rect 50379 14083 50421 14092
rect 52963 14132 53021 14133
rect 52963 14092 52972 14132
rect 53012 14092 53021 14132
rect 52963 14091 53021 14092
rect 56331 14132 56373 14141
rect 56331 14092 56332 14132
rect 56372 14092 56373 14132
rect 56331 14083 56373 14092
rect 4195 14048 4253 14049
rect 4195 14008 4204 14048
rect 4244 14008 4253 14048
rect 4195 14007 4253 14008
rect 12163 14048 12221 14049
rect 12163 14008 12172 14048
rect 12212 14008 12221 14048
rect 12163 14007 12221 14008
rect 13123 14048 13181 14049
rect 13123 14008 13132 14048
rect 13172 14008 13181 14048
rect 13123 14007 13181 14008
rect 13995 14048 14037 14057
rect 13995 14008 13996 14048
rect 14036 14008 14037 14048
rect 13995 13999 14037 14008
rect 15139 14048 15197 14049
rect 15139 14008 15148 14048
rect 15188 14008 15197 14048
rect 15139 14007 15197 14008
rect 15819 14048 15861 14057
rect 15819 14008 15820 14048
rect 15860 14008 15861 14048
rect 15819 13999 15861 14008
rect 16011 14048 16053 14057
rect 16011 14008 16012 14048
rect 16052 14008 16053 14048
rect 16011 13999 16053 14008
rect 16387 14048 16445 14049
rect 16387 14008 16396 14048
rect 16436 14008 16445 14048
rect 16387 14007 16445 14008
rect 17251 14048 17309 14049
rect 17251 14008 17260 14048
rect 17300 14008 17309 14048
rect 17251 14007 17309 14008
rect 18603 14048 18645 14057
rect 18603 14008 18604 14048
rect 18644 14008 18645 14048
rect 18603 13999 18645 14008
rect 18795 14048 18837 14057
rect 18795 14008 18796 14048
rect 18836 14008 18837 14048
rect 18795 13999 18837 14008
rect 18979 14048 19037 14049
rect 18979 14008 18988 14048
rect 19028 14008 19037 14048
rect 18979 14007 19037 14008
rect 19659 14048 19701 14057
rect 19659 14008 19660 14048
rect 19700 14008 19701 14048
rect 19659 13999 19701 14008
rect 26563 14048 26621 14049
rect 26563 14008 26572 14048
rect 26612 14008 26621 14048
rect 26563 14007 26621 14008
rect 33675 14048 33717 14057
rect 33675 14008 33676 14048
rect 33716 14008 33717 14048
rect 33675 13999 33717 14008
rect 34051 14048 34109 14049
rect 34051 14008 34060 14048
rect 34100 14008 34109 14048
rect 34051 14007 34109 14008
rect 34915 14048 34973 14049
rect 34915 14008 34924 14048
rect 34964 14008 34973 14048
rect 34915 14007 34973 14008
rect 36931 14048 36989 14049
rect 36931 14008 36940 14048
rect 36980 14008 36989 14048
rect 36931 14007 36989 14008
rect 38947 14048 39005 14049
rect 38947 14008 38956 14048
rect 38996 14008 39005 14048
rect 38947 14007 39005 14008
rect 39907 14048 39965 14049
rect 39907 14008 39916 14048
rect 39956 14008 39965 14048
rect 39907 14007 39965 14008
rect 40291 14048 40349 14049
rect 40291 14008 40300 14048
rect 40340 14008 40349 14048
rect 40291 14007 40349 14008
rect 42115 14048 42173 14049
rect 42115 14008 42124 14048
rect 42164 14008 42173 14048
rect 42115 14007 42173 14008
rect 49123 14048 49181 14049
rect 49123 14008 49132 14048
rect 49172 14008 49181 14048
rect 49123 14007 49181 14008
rect 49987 14048 50045 14049
rect 49987 14008 49996 14048
rect 50036 14008 50045 14048
rect 49987 14007 50045 14008
rect 51235 14048 51293 14049
rect 51235 14008 51244 14048
rect 51284 14008 51293 14048
rect 51235 14007 51293 14008
rect 52003 14048 52061 14049
rect 52003 14008 52012 14048
rect 52052 14008 52061 14048
rect 52003 14007 52061 14008
rect 53059 14048 53117 14049
rect 53059 14008 53068 14048
rect 53108 14008 53117 14048
rect 53059 14007 53117 14008
rect 53443 14048 53501 14049
rect 53443 14008 53452 14048
rect 53492 14008 53501 14048
rect 53443 14007 53501 14008
rect 54595 14048 54653 14049
rect 54595 14008 54604 14048
rect 54644 14008 54653 14048
rect 54595 14007 54653 14008
rect 55459 14048 55517 14049
rect 55459 14008 55468 14048
rect 55508 14008 55517 14048
rect 55459 14007 55517 14008
rect 55843 14048 55901 14049
rect 55843 14008 55852 14048
rect 55892 14008 55901 14048
rect 55843 14007 55901 14008
rect 56707 14048 56765 14049
rect 56707 14008 56716 14048
rect 56756 14008 56765 14048
rect 56707 14007 56765 14008
rect 57571 14048 57629 14049
rect 57571 14008 57580 14048
rect 57620 14008 57629 14048
rect 57571 14007 57629 14008
rect 18411 13964 18453 13973
rect 18411 13924 18412 13964
rect 18452 13924 18453 13964
rect 18411 13915 18453 13924
rect 25315 13964 25373 13965
rect 25315 13924 25324 13964
rect 25364 13924 25373 13964
rect 25315 13923 25373 13924
rect 12835 13880 12893 13881
rect 12835 13840 12844 13880
rect 12884 13840 12893 13880
rect 12835 13839 12893 13840
rect 25131 13880 25173 13889
rect 25131 13840 25132 13880
rect 25172 13840 25173 13880
rect 25131 13831 25173 13840
rect 25891 13880 25949 13881
rect 25891 13840 25900 13880
rect 25940 13840 25949 13880
rect 25891 13839 25949 13840
rect 47971 13880 48029 13881
rect 47971 13840 47980 13880
rect 48020 13840 48029 13880
rect 47971 13839 48029 13840
rect 3523 13796 3581 13797
rect 3523 13756 3532 13796
rect 3572 13756 3581 13796
rect 3523 13755 3581 13756
rect 18795 13796 18837 13805
rect 18795 13756 18796 13796
rect 18836 13756 18837 13796
rect 18795 13747 18837 13756
rect 37603 13796 37661 13797
rect 37603 13756 37612 13796
rect 37652 13756 37661 13796
rect 37603 13755 37661 13756
rect 39243 13796 39285 13805
rect 39243 13756 39244 13796
rect 39284 13756 39285 13796
rect 39243 13747 39285 13756
rect 41443 13796 41501 13797
rect 41443 13756 41452 13796
rect 41492 13756 41501 13796
rect 41443 13755 41501 13756
rect 50563 13796 50621 13797
rect 50563 13756 50572 13796
rect 50612 13756 50621 13796
rect 50563 13755 50621 13756
rect 576 13628 99360 13652
rect 576 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 18232 13628
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18600 13588 33352 13628
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33720 13588 48472 13628
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48840 13588 63592 13628
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63960 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 93832 13628
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 94200 13588 99360 13628
rect 576 13564 99360 13588
rect 4483 13460 4541 13461
rect 4483 13420 4492 13460
rect 4532 13420 4541 13460
rect 4483 13419 4541 13420
rect 14659 13460 14717 13461
rect 14659 13420 14668 13460
rect 14708 13420 14717 13460
rect 14659 13419 14717 13420
rect 26275 13460 26333 13461
rect 26275 13420 26284 13460
rect 26324 13420 26333 13460
rect 26275 13419 26333 13420
rect 32515 13460 32573 13461
rect 32515 13420 32524 13460
rect 32564 13420 32573 13460
rect 32515 13419 32573 13420
rect 39619 13460 39677 13461
rect 39619 13420 39628 13460
rect 39668 13420 39677 13460
rect 39619 13419 39677 13420
rect 49995 13460 50037 13469
rect 49995 13420 49996 13460
rect 50036 13420 50037 13460
rect 49995 13411 50037 13420
rect 51811 13460 51869 13461
rect 51811 13420 51820 13460
rect 51860 13420 51869 13460
rect 51811 13419 51869 13420
rect 54891 13460 54933 13469
rect 54891 13420 54892 13460
rect 54932 13420 54933 13460
rect 54891 13411 54933 13420
rect 23307 13376 23349 13385
rect 23307 13336 23308 13376
rect 23348 13336 23349 13376
rect 23307 13327 23349 13336
rect 28579 13292 28637 13293
rect 28579 13252 28588 13292
rect 28628 13252 28637 13292
rect 28579 13251 28637 13252
rect 2467 13208 2525 13209
rect 2467 13168 2476 13208
rect 2516 13168 2525 13208
rect 2467 13167 2525 13168
rect 3331 13208 3389 13209
rect 3331 13168 3340 13208
rect 3380 13168 3389 13208
rect 3331 13167 3389 13168
rect 8035 13208 8093 13209
rect 8035 13168 8044 13208
rect 8084 13168 8093 13208
rect 8035 13167 8093 13168
rect 9187 13208 9245 13209
rect 9187 13168 9196 13208
rect 9236 13168 9245 13208
rect 9187 13167 9245 13168
rect 11683 13208 11741 13209
rect 11683 13168 11692 13208
rect 11732 13168 11741 13208
rect 11683 13167 11741 13168
rect 12267 13208 12309 13217
rect 12267 13168 12268 13208
rect 12308 13168 12309 13208
rect 12267 13159 12309 13168
rect 12643 13208 12701 13209
rect 12643 13168 12652 13208
rect 12692 13168 12701 13208
rect 12643 13167 12701 13168
rect 13507 13208 13565 13209
rect 13507 13168 13516 13208
rect 13556 13168 13565 13208
rect 13507 13167 13565 13168
rect 18691 13208 18749 13209
rect 18691 13168 18700 13208
rect 18740 13168 18749 13208
rect 18691 13167 18749 13168
rect 19075 13208 19133 13209
rect 19075 13168 19084 13208
rect 19124 13168 19133 13208
rect 19075 13167 19133 13168
rect 19363 13208 19421 13209
rect 19363 13168 19372 13208
rect 19412 13168 19421 13208
rect 19363 13167 19421 13168
rect 20227 13208 20285 13209
rect 20227 13168 20236 13208
rect 20276 13168 20285 13208
rect 20227 13167 20285 13168
rect 20331 13208 20373 13217
rect 20331 13168 20332 13208
rect 20372 13168 20373 13208
rect 20331 13159 20373 13168
rect 20427 13208 20469 13217
rect 20427 13168 20428 13208
rect 20468 13168 20469 13208
rect 20427 13159 20469 13168
rect 23499 13208 23541 13217
rect 23499 13168 23500 13208
rect 23540 13168 23541 13208
rect 23499 13159 23541 13168
rect 23883 13208 23925 13217
rect 23883 13168 23884 13208
rect 23924 13168 23925 13208
rect 23883 13159 23925 13168
rect 24259 13208 24317 13209
rect 24259 13168 24268 13208
rect 24308 13168 24317 13208
rect 24259 13167 24317 13168
rect 25123 13208 25181 13209
rect 25123 13168 25132 13208
rect 25172 13168 25181 13208
rect 25123 13167 25181 13168
rect 28875 13208 28917 13217
rect 28875 13168 28876 13208
rect 28916 13168 28917 13208
rect 28875 13159 28917 13168
rect 28971 13208 29013 13217
rect 28971 13168 28972 13208
rect 29012 13168 29013 13208
rect 28971 13159 29013 13168
rect 29059 13208 29117 13209
rect 29059 13168 29068 13208
rect 29108 13168 29117 13208
rect 29059 13167 29117 13168
rect 30115 13208 30173 13209
rect 30115 13168 30124 13208
rect 30164 13168 30173 13208
rect 30115 13167 30173 13168
rect 30499 13208 30557 13209
rect 30499 13168 30508 13208
rect 30548 13168 30557 13208
rect 30499 13167 30557 13168
rect 30883 13208 30941 13209
rect 30883 13168 30892 13208
rect 30932 13168 30941 13208
rect 30883 13167 30941 13168
rect 32323 13208 32381 13209
rect 32323 13168 32332 13208
rect 32372 13168 32381 13208
rect 32323 13167 32381 13168
rect 37227 13208 37269 13217
rect 37227 13168 37228 13208
rect 37268 13168 37269 13208
rect 37227 13159 37269 13168
rect 37603 13208 37661 13209
rect 37603 13168 37612 13208
rect 37652 13168 37661 13208
rect 37603 13167 37661 13168
rect 38467 13208 38525 13209
rect 38467 13168 38476 13208
rect 38516 13168 38525 13208
rect 38467 13167 38525 13168
rect 39811 13208 39869 13209
rect 39811 13168 39820 13208
rect 39860 13168 39869 13208
rect 39811 13167 39869 13168
rect 40195 13208 40253 13209
rect 40195 13168 40204 13208
rect 40244 13168 40253 13208
rect 40195 13167 40253 13168
rect 41451 13208 41493 13217
rect 41451 13168 41452 13208
rect 41492 13168 41493 13208
rect 41451 13159 41493 13168
rect 41827 13208 41885 13209
rect 41827 13168 41836 13208
rect 41876 13168 41885 13208
rect 41827 13167 41885 13168
rect 42691 13208 42749 13209
rect 42691 13168 42700 13208
rect 42740 13168 42749 13208
rect 42691 13167 42749 13168
rect 47107 13208 47165 13209
rect 47107 13168 47116 13208
rect 47156 13168 47165 13208
rect 47107 13167 47165 13168
rect 47971 13208 48029 13209
rect 47971 13168 47980 13208
rect 48020 13168 48029 13208
rect 47971 13167 48029 13168
rect 48363 13208 48405 13217
rect 48363 13168 48364 13208
rect 48404 13168 48405 13208
rect 48363 13159 48405 13168
rect 49315 13208 49373 13209
rect 49315 13168 49324 13208
rect 49364 13168 49373 13208
rect 49315 13167 49373 13168
rect 50275 13208 50333 13209
rect 50275 13168 50284 13208
rect 50324 13168 50333 13208
rect 50275 13167 50333 13168
rect 52963 13208 53021 13209
rect 52963 13168 52972 13208
rect 53012 13168 53021 13208
rect 52963 13167 53021 13168
rect 53827 13208 53885 13209
rect 53827 13168 53836 13208
rect 53876 13168 53885 13208
rect 53827 13167 53885 13168
rect 54595 13208 54653 13209
rect 54595 13168 54604 13208
rect 54644 13168 54653 13208
rect 54595 13167 54653 13168
rect 56611 13208 56669 13209
rect 56611 13168 56620 13208
rect 56660 13168 56669 13208
rect 56611 13167 56669 13168
rect 57475 13208 57533 13209
rect 57475 13168 57484 13208
rect 57524 13168 57533 13208
rect 57475 13167 57533 13168
rect 2091 13124 2133 13133
rect 2091 13084 2092 13124
rect 2132 13084 2133 13124
rect 2091 13075 2133 13084
rect 7171 13124 7229 13125
rect 7171 13084 7180 13124
rect 7220 13084 7229 13124
rect 7171 13083 7229 13084
rect 30403 13124 30461 13125
rect 30403 13084 30412 13124
rect 30452 13084 30461 13124
rect 30403 13083 30461 13084
rect 54219 13124 54261 13133
rect 54219 13084 54220 13124
rect 54260 13084 54261 13124
rect 54219 13075 54261 13084
rect 56235 13124 56277 13133
rect 56235 13084 56236 13124
rect 56276 13084 56277 13124
rect 56235 13075 56277 13084
rect 643 13040 701 13041
rect 643 13000 652 13040
rect 692 13000 701 13040
rect 643 12999 701 13000
rect 9859 13040 9917 13041
rect 9859 13000 9868 13040
rect 9908 13000 9917 13040
rect 9859 12999 9917 13000
rect 11211 13040 11253 13049
rect 11211 13000 11212 13040
rect 11252 13000 11253 13040
rect 11211 12991 11253 13000
rect 18603 13040 18645 13049
rect 18603 13000 18604 13040
rect 18644 13000 18645 13040
rect 18603 12991 18645 13000
rect 20035 13040 20093 13041
rect 20035 13000 20044 13040
rect 20084 13000 20093 13040
rect 20035 12999 20093 13000
rect 28395 13040 28437 13049
rect 28395 13000 28396 13040
rect 28436 13000 28437 13040
rect 28395 12991 28437 13000
rect 29443 13040 29501 13041
rect 29443 13000 29452 13040
rect 29492 13000 29501 13040
rect 29443 12999 29501 13000
rect 32227 13040 32285 13041
rect 32227 13000 32236 13040
rect 32276 13000 32285 13040
rect 32227 12999 32285 13000
rect 40299 13040 40341 13049
rect 40299 13000 40300 13040
rect 40340 13000 40341 13040
rect 40299 12991 40341 13000
rect 43843 13040 43901 13041
rect 43843 13000 43852 13040
rect 43892 13000 43901 13040
rect 43843 12999 43901 13000
rect 45955 13040 46013 13041
rect 45955 13000 45964 13040
rect 46004 13000 46013 13040
rect 45955 12999 46013 13000
rect 55083 13040 55125 13049
rect 55083 13000 55084 13040
rect 55124 13000 55125 13040
rect 55083 12991 55125 13000
rect 58627 13040 58685 13041
rect 58627 13000 58636 13040
rect 58676 13000 58685 13040
rect 58627 12999 58685 13000
rect 576 12872 99360 12896
rect 576 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 19472 12872
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19840 12832 34592 12872
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34960 12832 49712 12872
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 50080 12832 64832 12872
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 65200 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 95072 12872
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95440 12832 99360 12872
rect 576 12808 99360 12832
rect 643 12704 701 12705
rect 643 12664 652 12704
rect 692 12664 701 12704
rect 643 12663 701 12664
rect 2187 12704 2229 12713
rect 2187 12664 2188 12704
rect 2228 12664 2229 12704
rect 2187 12655 2229 12664
rect 30019 12704 30077 12705
rect 30019 12664 30028 12704
rect 30068 12664 30077 12704
rect 30019 12663 30077 12664
rect 54883 12704 54941 12705
rect 54883 12664 54892 12704
rect 54932 12664 54941 12704
rect 54883 12663 54941 12664
rect 55171 12704 55229 12705
rect 55171 12664 55180 12704
rect 55220 12664 55229 12704
rect 55171 12663 55229 12664
rect 56235 12704 56277 12713
rect 56235 12664 56236 12704
rect 56276 12664 56277 12704
rect 56235 12655 56277 12664
rect 9483 12620 9525 12629
rect 9483 12580 9484 12620
rect 9524 12580 9525 12620
rect 9483 12571 9525 12580
rect 27627 12620 27669 12629
rect 27627 12580 27628 12620
rect 27668 12580 27669 12620
rect 27627 12571 27669 12580
rect 32611 12620 32669 12621
rect 32611 12580 32620 12620
rect 32660 12580 32669 12620
rect 32611 12579 32669 12580
rect 56715 12620 56757 12629
rect 56715 12580 56716 12620
rect 56756 12580 56757 12620
rect 56715 12571 56757 12580
rect 57675 12620 57717 12629
rect 57675 12580 57676 12620
rect 57716 12580 57717 12620
rect 57675 12571 57717 12580
rect 2571 12536 2613 12545
rect 2571 12496 2572 12536
rect 2612 12496 2613 12536
rect 2571 12487 2613 12496
rect 2947 12536 3005 12537
rect 2947 12496 2956 12536
rect 2996 12496 3005 12536
rect 2947 12495 3005 12496
rect 3811 12536 3869 12537
rect 3811 12496 3820 12536
rect 3860 12496 3869 12536
rect 3811 12495 3869 12496
rect 6219 12536 6261 12545
rect 6219 12496 6220 12536
rect 6260 12496 6261 12536
rect 6219 12487 6261 12496
rect 6595 12536 6653 12537
rect 6595 12496 6604 12536
rect 6644 12496 6653 12536
rect 6595 12495 6653 12496
rect 7459 12536 7517 12537
rect 7459 12496 7468 12536
rect 7508 12496 7517 12536
rect 7459 12495 7517 12496
rect 9859 12536 9917 12537
rect 9859 12496 9868 12536
rect 9908 12496 9917 12536
rect 9859 12495 9917 12496
rect 10723 12536 10781 12537
rect 10723 12496 10732 12536
rect 10772 12496 10781 12536
rect 10723 12495 10781 12496
rect 18499 12536 18557 12537
rect 18499 12496 18508 12536
rect 18548 12496 18557 12536
rect 18499 12495 18557 12496
rect 18595 12536 18653 12537
rect 18595 12496 18604 12536
rect 18644 12496 18653 12536
rect 18595 12495 18653 12496
rect 19651 12536 19709 12537
rect 19651 12496 19660 12536
rect 19700 12496 19709 12536
rect 19651 12495 19709 12496
rect 19851 12536 19893 12545
rect 19851 12496 19852 12536
rect 19892 12496 19893 12536
rect 19851 12487 19893 12496
rect 19947 12536 19989 12545
rect 19947 12496 19948 12536
rect 19988 12496 19989 12536
rect 19947 12487 19989 12496
rect 20043 12536 20085 12545
rect 20043 12496 20044 12536
rect 20084 12496 20085 12536
rect 20043 12487 20085 12496
rect 20139 12536 20181 12545
rect 20139 12496 20140 12536
rect 20180 12496 20181 12536
rect 20139 12487 20181 12496
rect 21283 12536 21341 12537
rect 21283 12496 21292 12536
rect 21332 12496 21341 12536
rect 21283 12495 21341 12496
rect 28003 12536 28061 12537
rect 28003 12496 28012 12536
rect 28052 12496 28061 12536
rect 28003 12495 28061 12496
rect 28867 12536 28925 12537
rect 28867 12496 28876 12536
rect 28916 12496 28925 12536
rect 28867 12495 28925 12496
rect 33475 12536 33533 12537
rect 33475 12496 33484 12536
rect 33524 12496 33533 12536
rect 33475 12495 33533 12496
rect 34435 12536 34493 12537
rect 34435 12496 34444 12536
rect 34484 12496 34493 12536
rect 34435 12495 34493 12496
rect 55075 12536 55133 12537
rect 55075 12496 55084 12536
rect 55124 12496 55133 12536
rect 55075 12495 55133 12496
rect 56611 12536 56669 12537
rect 56611 12496 56620 12536
rect 56660 12496 56669 12536
rect 56611 12495 56669 12496
rect 56811 12536 56853 12545
rect 56811 12496 56812 12536
rect 56852 12496 56853 12536
rect 56811 12487 56853 12496
rect 58339 12536 58397 12537
rect 58339 12496 58348 12536
rect 58388 12496 58397 12536
rect 58339 12495 58397 12496
rect 2371 12452 2429 12453
rect 2371 12412 2380 12452
rect 2420 12412 2429 12452
rect 2371 12411 2429 12412
rect 8619 12452 8661 12461
rect 8619 12412 8620 12452
rect 8660 12412 8661 12452
rect 8619 12403 8661 12412
rect 11883 12452 11925 12461
rect 11883 12412 11884 12452
rect 11924 12412 11925 12452
rect 11883 12403 11925 12412
rect 18787 12452 18845 12453
rect 18787 12412 18796 12452
rect 18836 12412 18845 12452
rect 18787 12411 18845 12412
rect 32227 12452 32285 12453
rect 32227 12412 32236 12452
rect 32276 12412 32285 12452
rect 32227 12411 32285 12412
rect 33771 12452 33813 12461
rect 33771 12412 33772 12452
rect 33812 12412 33813 12452
rect 33771 12403 33813 12412
rect 56419 12452 56477 12453
rect 56419 12412 56428 12452
rect 56468 12412 56477 12452
rect 56419 12411 56477 12412
rect 4963 12284 5021 12285
rect 4963 12244 4972 12284
rect 5012 12244 5021 12284
rect 4963 12243 5021 12244
rect 18979 12284 19037 12285
rect 18979 12244 18988 12284
rect 19028 12244 19037 12284
rect 18979 12243 19037 12244
rect 21955 12284 22013 12285
rect 21955 12244 21964 12284
rect 22004 12244 22013 12284
rect 21955 12243 22013 12244
rect 32043 12284 32085 12293
rect 32043 12244 32044 12284
rect 32084 12244 32085 12284
rect 32043 12235 32085 12244
rect 32811 12284 32853 12293
rect 32811 12244 32812 12284
rect 32852 12244 32853 12284
rect 32811 12235 32853 12244
rect 576 12116 99360 12140
rect 576 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 18232 12116
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18600 12076 33352 12116
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33720 12076 48472 12116
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48840 12076 63592 12116
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63960 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 93832 12116
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 94200 12076 99360 12116
rect 576 12052 99360 12076
rect 3243 11948 3285 11957
rect 3243 11908 3244 11948
rect 3284 11908 3285 11948
rect 3243 11899 3285 11908
rect 17259 11948 17301 11957
rect 17259 11908 17260 11948
rect 17300 11908 17301 11948
rect 17259 11899 17301 11908
rect 19179 11948 19221 11957
rect 19179 11908 19180 11948
rect 19220 11908 19221 11948
rect 19179 11899 19221 11908
rect 31275 11948 31317 11957
rect 31275 11908 31276 11948
rect 31316 11908 31317 11948
rect 31275 11899 31317 11908
rect 33955 11948 34013 11949
rect 33955 11908 33964 11948
rect 34004 11908 34013 11948
rect 33955 11907 34013 11908
rect 3427 11780 3485 11781
rect 3427 11740 3436 11780
rect 3476 11740 3485 11780
rect 3427 11739 3485 11740
rect 3915 11696 3957 11705
rect 3915 11656 3916 11696
rect 3956 11656 3957 11696
rect 3915 11647 3957 11656
rect 4011 11696 4053 11705
rect 4011 11656 4012 11696
rect 4052 11656 4053 11696
rect 4011 11647 4053 11656
rect 4099 11696 4157 11697
rect 4099 11656 4108 11696
rect 4148 11656 4157 11696
rect 4099 11655 4157 11656
rect 4963 11696 5021 11697
rect 4963 11656 4972 11696
rect 5012 11656 5021 11696
rect 4963 11655 5021 11656
rect 5155 11696 5213 11697
rect 5155 11656 5164 11696
rect 5204 11656 5213 11696
rect 5155 11655 5213 11656
rect 5443 11696 5501 11697
rect 5443 11656 5452 11696
rect 5492 11656 5501 11696
rect 5443 11655 5501 11656
rect 16675 11696 16733 11697
rect 16675 11656 16684 11696
rect 16724 11656 16733 11696
rect 16675 11655 16733 11656
rect 17163 11696 17205 11705
rect 17163 11656 17164 11696
rect 17204 11656 17205 11696
rect 17163 11647 17205 11656
rect 17347 11696 17405 11697
rect 17347 11656 17356 11696
rect 17396 11656 17405 11696
rect 17347 11655 17405 11656
rect 18883 11696 18941 11697
rect 18883 11656 18892 11696
rect 18932 11656 18941 11696
rect 18883 11655 18941 11656
rect 31171 11696 31229 11697
rect 31171 11656 31180 11696
rect 31220 11656 31229 11696
rect 31171 11655 31229 11656
rect 31371 11696 31413 11705
rect 31371 11656 31372 11696
rect 31412 11656 31413 11696
rect 31371 11647 31413 11656
rect 31563 11696 31605 11705
rect 31563 11656 31564 11696
rect 31604 11656 31605 11696
rect 31563 11647 31605 11656
rect 31939 11696 31997 11697
rect 31939 11656 31948 11696
rect 31988 11656 31997 11696
rect 31939 11655 31997 11656
rect 32803 11696 32861 11697
rect 32803 11656 32812 11696
rect 32852 11656 32861 11696
rect 32803 11655 32861 11656
rect 40675 11696 40733 11697
rect 40675 11656 40684 11696
rect 40724 11656 40733 11696
rect 40675 11655 40733 11656
rect 46819 11696 46877 11697
rect 46819 11656 46828 11696
rect 46868 11656 46877 11696
rect 46819 11655 46877 11656
rect 5635 11612 5693 11613
rect 5635 11572 5644 11612
rect 5684 11572 5693 11612
rect 5635 11571 5693 11572
rect 643 11528 701 11529
rect 643 11488 652 11528
rect 692 11488 701 11528
rect 643 11487 701 11488
rect 4291 11528 4349 11529
rect 4291 11488 4300 11528
rect 4340 11488 4349 11528
rect 4291 11487 4349 11488
rect 16003 11528 16061 11529
rect 16003 11488 16012 11528
rect 16052 11488 16061 11528
rect 16003 11487 16061 11488
rect 19371 11528 19413 11537
rect 19371 11488 19372 11528
rect 19412 11488 19413 11528
rect 19371 11479 19413 11488
rect 41347 11528 41405 11529
rect 41347 11488 41356 11528
rect 41396 11488 41405 11528
rect 41347 11487 41405 11488
rect 47491 11528 47549 11529
rect 47491 11488 47500 11528
rect 47540 11488 47549 11528
rect 47491 11487 47549 11488
rect 576 11360 99360 11384
rect 576 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 19472 11360
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19840 11320 34592 11360
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34960 11320 49712 11360
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 50080 11320 64832 11360
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 65200 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 95072 11360
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95440 11320 99360 11360
rect 576 11296 99360 11320
rect 643 11192 701 11193
rect 643 11152 652 11192
rect 692 11152 701 11192
rect 643 11151 701 11152
rect 16579 11192 16637 11193
rect 16579 11152 16588 11192
rect 16628 11152 16637 11192
rect 16579 11151 16637 11152
rect 32803 11192 32861 11193
rect 32803 11152 32812 11192
rect 32852 11152 32861 11192
rect 32803 11151 32861 11152
rect 54691 11192 54749 11193
rect 54691 11152 54700 11192
rect 54740 11152 54749 11192
rect 54691 11151 54749 11152
rect 23019 11108 23061 11117
rect 23019 11068 23020 11108
rect 23060 11068 23061 11108
rect 23019 11059 23061 11068
rect 36163 11108 36221 11109
rect 36163 11068 36172 11108
rect 36212 11068 36221 11108
rect 36163 11067 36221 11068
rect 43651 11108 43709 11109
rect 43651 11068 43660 11108
rect 43700 11068 43709 11108
rect 43651 11067 43709 11068
rect 55851 11108 55893 11117
rect 55851 11068 55852 11108
rect 55892 11068 55893 11108
rect 55851 11059 55893 11068
rect 15907 11024 15965 11025
rect 15907 10984 15916 11024
rect 15956 10984 15965 11024
rect 15907 10983 15965 10984
rect 23395 11024 23453 11025
rect 23395 10984 23404 11024
rect 23444 10984 23453 11024
rect 23395 10983 23453 10984
rect 24259 11024 24317 11025
rect 24259 10984 24268 11024
rect 24308 10984 24317 11024
rect 24259 10983 24317 10984
rect 33475 11024 33533 11025
rect 33475 10984 33484 11024
rect 33524 10984 33533 11024
rect 33475 10983 33533 10984
rect 37027 11024 37085 11025
rect 37027 10984 37036 11024
rect 37076 10984 37085 11024
rect 37027 10983 37085 10984
rect 39907 11024 39965 11025
rect 39907 10984 39916 11024
rect 39956 10984 39965 11024
rect 39907 10983 39965 10984
rect 43843 11024 43901 11025
rect 43843 10984 43852 11024
rect 43892 10984 43901 11024
rect 43843 10983 43901 10984
rect 44131 11024 44189 11025
rect 44131 10984 44140 11024
rect 44180 10984 44189 11024
rect 44131 10983 44189 10984
rect 44995 11024 45053 11025
rect 44995 10984 45004 11024
rect 45044 10984 45053 11024
rect 44995 10983 45053 10984
rect 55363 11024 55421 11025
rect 55363 10984 55372 11024
rect 55412 10984 55421 11024
rect 55363 10983 55421 10984
rect 55747 11024 55805 11025
rect 55747 10984 55756 11024
rect 55796 10984 55805 11024
rect 55747 10983 55805 10984
rect 55947 11024 55989 11033
rect 55947 10984 55948 11024
rect 55988 10984 55989 11024
rect 55947 10975 55989 10984
rect 31843 10940 31901 10941
rect 31843 10900 31852 10940
rect 31892 10900 31901 10940
rect 31843 10899 31901 10900
rect 54019 10940 54077 10941
rect 54019 10900 54028 10940
rect 54068 10900 54077 10940
rect 54019 10899 54077 10900
rect 25411 10772 25469 10773
rect 25411 10732 25420 10772
rect 25460 10732 25469 10772
rect 25411 10731 25469 10732
rect 31659 10772 31701 10781
rect 31659 10732 31660 10772
rect 31700 10732 31701 10772
rect 31659 10723 31701 10732
rect 40579 10772 40637 10773
rect 40579 10732 40588 10772
rect 40628 10732 40637 10772
rect 40579 10731 40637 10732
rect 44323 10772 44381 10773
rect 44323 10732 44332 10772
rect 44372 10732 44381 10772
rect 44323 10731 44381 10732
rect 53835 10772 53877 10781
rect 53835 10732 53836 10772
rect 53876 10732 53877 10772
rect 53835 10723 53877 10732
rect 576 10604 99360 10628
rect 576 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 18232 10604
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18600 10564 33352 10604
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33720 10564 48472 10604
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48840 10564 63592 10604
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63960 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 93832 10604
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 94200 10564 99360 10604
rect 576 10540 99360 10564
rect 3627 10436 3669 10445
rect 3627 10396 3628 10436
rect 3668 10396 3669 10436
rect 3627 10387 3669 10396
rect 33475 10436 33533 10437
rect 33475 10396 33484 10436
rect 33524 10396 33533 10436
rect 33475 10395 33533 10396
rect 38371 10436 38429 10437
rect 38371 10396 38380 10436
rect 38420 10396 38429 10436
rect 38371 10395 38429 10396
rect 44131 10436 44189 10437
rect 44131 10396 44140 10436
rect 44180 10396 44189 10436
rect 44131 10395 44189 10396
rect 52299 10436 52341 10445
rect 52299 10396 52300 10436
rect 52340 10396 52341 10436
rect 52299 10387 52341 10396
rect 55171 10436 55229 10437
rect 55171 10396 55180 10436
rect 55220 10396 55229 10436
rect 55171 10395 55229 10396
rect 55563 10352 55605 10361
rect 55563 10312 55564 10352
rect 55604 10312 55605 10352
rect 55563 10303 55605 10312
rect 25411 10268 25469 10269
rect 25411 10228 25420 10268
rect 25460 10228 25469 10268
rect 25411 10227 25469 10228
rect 47019 10268 47061 10277
rect 47019 10228 47020 10268
rect 47060 10228 47061 10268
rect 47019 10219 47061 10228
rect 48163 10268 48221 10269
rect 48163 10228 48172 10268
rect 48212 10228 48221 10268
rect 48163 10227 48221 10228
rect 55747 10268 55805 10269
rect 55747 10228 55756 10268
rect 55796 10228 55805 10268
rect 55747 10227 55805 10228
rect 56619 10268 56661 10277
rect 56619 10228 56620 10268
rect 56660 10228 56661 10268
rect 56619 10219 56661 10228
rect 4203 10184 4245 10193
rect 4203 10144 4204 10184
rect 4244 10144 4245 10184
rect 4203 10135 4245 10144
rect 12931 10184 12989 10185
rect 12931 10144 12940 10184
rect 12980 10144 12989 10184
rect 12931 10143 12989 10144
rect 16003 10184 16061 10185
rect 16003 10144 16012 10184
rect 16052 10144 16061 10184
rect 16003 10143 16061 10144
rect 16291 10184 16349 10185
rect 16291 10144 16300 10184
rect 16340 10144 16349 10184
rect 16291 10143 16349 10144
rect 18987 10184 19029 10193
rect 18987 10144 18988 10184
rect 19028 10144 19029 10184
rect 18987 10135 19029 10144
rect 19363 10184 19421 10185
rect 19363 10144 19372 10184
rect 19412 10144 19421 10184
rect 19363 10143 19421 10144
rect 20227 10184 20285 10185
rect 20227 10144 20236 10184
rect 20276 10144 20285 10184
rect 20227 10143 20285 10144
rect 25603 10184 25661 10185
rect 25603 10144 25612 10184
rect 25652 10144 25661 10184
rect 25603 10143 25661 10144
rect 25699 10184 25757 10185
rect 25699 10144 25708 10184
rect 25748 10144 25757 10184
rect 25699 10143 25757 10144
rect 31083 10184 31125 10193
rect 31083 10144 31084 10184
rect 31124 10144 31125 10184
rect 31083 10135 31125 10144
rect 31459 10184 31517 10185
rect 31459 10144 31468 10184
rect 31508 10144 31517 10184
rect 31459 10143 31517 10144
rect 32323 10184 32381 10185
rect 32323 10144 32332 10184
rect 32372 10144 32381 10184
rect 32323 10143 32381 10144
rect 39523 10184 39581 10185
rect 39523 10144 39532 10184
rect 39572 10144 39581 10184
rect 39523 10143 39581 10144
rect 40387 10184 40445 10185
rect 40387 10144 40396 10184
rect 40436 10144 40445 10184
rect 40387 10143 40445 10144
rect 40779 10184 40821 10193
rect 40779 10144 40780 10184
rect 40820 10144 40821 10184
rect 40779 10135 40821 10144
rect 45283 10184 45341 10185
rect 45283 10144 45292 10184
rect 45332 10144 45341 10184
rect 45283 10143 45341 10144
rect 46147 10184 46205 10185
rect 46147 10144 46156 10184
rect 46196 10144 46205 10184
rect 46147 10143 46205 10144
rect 46923 10184 46965 10193
rect 46923 10144 46924 10184
rect 46964 10144 46965 10184
rect 46923 10135 46965 10144
rect 47107 10184 47165 10185
rect 47107 10144 47116 10184
rect 47156 10144 47165 10184
rect 47107 10143 47165 10144
rect 47971 10184 48029 10185
rect 47971 10144 47980 10184
rect 48020 10144 48029 10184
rect 47971 10143 48029 10144
rect 48451 10184 48509 10185
rect 48451 10144 48460 10184
rect 48500 10144 48509 10184
rect 48451 10143 48509 10144
rect 48555 10184 48597 10193
rect 48555 10144 48556 10184
rect 48596 10144 48597 10184
rect 48555 10135 48597 10144
rect 49891 10184 49949 10185
rect 49891 10144 49900 10184
rect 49940 10144 49949 10184
rect 49891 10143 49949 10144
rect 50275 10184 50333 10185
rect 50275 10144 50284 10184
rect 50324 10144 50333 10184
rect 50275 10143 50333 10144
rect 51723 10184 51765 10193
rect 51723 10144 51724 10184
rect 51764 10144 51765 10184
rect 51723 10135 51765 10144
rect 52779 10184 52821 10193
rect 52779 10144 52780 10184
rect 52820 10144 52821 10184
rect 52779 10135 52821 10144
rect 53155 10184 53213 10185
rect 53155 10144 53164 10184
rect 53204 10144 53213 10184
rect 53155 10143 53213 10144
rect 54019 10184 54077 10185
rect 54019 10144 54028 10184
rect 54068 10144 54077 10184
rect 54019 10143 54077 10144
rect 57283 10184 57341 10185
rect 57283 10144 57292 10184
rect 57332 10144 57341 10184
rect 57283 10143 57341 10144
rect 16483 10100 16541 10101
rect 16483 10060 16492 10100
rect 16532 10060 16541 10100
rect 16483 10059 16541 10060
rect 46539 10100 46581 10109
rect 46539 10060 46540 10100
rect 46580 10060 46581 10100
rect 46539 10051 46581 10060
rect 47307 10100 47349 10109
rect 47307 10060 47308 10100
rect 47348 10060 47349 10100
rect 47307 10051 47349 10060
rect 49795 10100 49853 10101
rect 49795 10060 49804 10100
rect 49844 10060 49853 10100
rect 49795 10059 49853 10060
rect 643 10016 701 10017
rect 643 9976 652 10016
rect 692 9976 701 10016
rect 643 9975 701 9976
rect 12259 10016 12317 10017
rect 12259 9976 12268 10016
rect 12308 9976 12317 10016
rect 12259 9975 12317 9976
rect 21379 10016 21437 10017
rect 21379 9976 21388 10016
rect 21428 9976 21437 10016
rect 21379 9975 21437 9976
rect 576 9848 99360 9872
rect 576 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 19472 9848
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19840 9808 34592 9848
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34960 9808 49712 9848
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 50080 9808 64832 9848
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 65200 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 95072 9848
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95440 9808 99360 9848
rect 576 9784 99360 9808
rect 643 9680 701 9681
rect 643 9640 652 9680
rect 692 9640 701 9680
rect 643 9639 701 9640
rect 4387 9680 4445 9681
rect 4387 9640 4396 9680
rect 4436 9640 4445 9680
rect 4387 9639 4445 9640
rect 5251 9680 5309 9681
rect 5251 9640 5260 9680
rect 5300 9640 5309 9680
rect 5251 9639 5309 9640
rect 14275 9680 14333 9681
rect 14275 9640 14284 9680
rect 14324 9640 14333 9680
rect 14275 9639 14333 9640
rect 26467 9680 26525 9681
rect 26467 9640 26476 9680
rect 26516 9640 26525 9680
rect 26467 9639 26525 9640
rect 47211 9680 47253 9689
rect 47211 9640 47212 9680
rect 47252 9640 47253 9680
rect 47211 9631 47253 9640
rect 47875 9680 47933 9681
rect 47875 9640 47884 9680
rect 47924 9640 47933 9680
rect 47875 9639 47933 9640
rect 51819 9680 51861 9689
rect 51819 9640 51820 9680
rect 51860 9640 51861 9680
rect 51819 9631 51861 9640
rect 57283 9680 57341 9681
rect 57283 9640 57292 9680
rect 57332 9640 57341 9680
rect 57283 9639 57341 9640
rect 3243 9596 3285 9605
rect 3243 9556 3244 9596
rect 3284 9556 3285 9596
rect 3243 9547 3285 9556
rect 11883 9596 11925 9605
rect 11883 9556 11884 9596
rect 11924 9556 11925 9596
rect 11883 9547 11925 9556
rect 15915 9596 15957 9605
rect 15915 9556 15916 9596
rect 15956 9556 15957 9596
rect 15915 9547 15957 9556
rect 41163 9596 41205 9605
rect 41163 9556 41164 9596
rect 41204 9556 41205 9596
rect 41163 9547 41205 9556
rect 54891 9596 54933 9605
rect 54891 9556 54892 9596
rect 54932 9556 54933 9596
rect 54891 9547 54933 9556
rect 3147 9512 3189 9521
rect 3147 9472 3148 9512
rect 3188 9472 3189 9512
rect 3147 9463 3189 9472
rect 3331 9512 3389 9513
rect 3331 9472 3340 9512
rect 3380 9472 3389 9512
rect 3331 9471 3389 9472
rect 3531 9512 3573 9521
rect 3531 9472 3532 9512
rect 3572 9472 3573 9512
rect 3531 9463 3573 9472
rect 4195 9512 4253 9513
rect 4195 9472 4204 9512
rect 4244 9472 4253 9512
rect 4195 9471 4253 9472
rect 5059 9512 5117 9513
rect 5059 9472 5068 9512
rect 5108 9472 5117 9512
rect 5059 9471 5117 9472
rect 5347 9512 5405 9513
rect 5347 9472 5356 9512
rect 5396 9472 5405 9512
rect 5347 9471 5405 9472
rect 8035 9512 8093 9513
rect 8035 9472 8044 9512
rect 8084 9472 8093 9512
rect 8035 9471 8093 9472
rect 10627 9512 10685 9513
rect 10627 9472 10636 9512
rect 10676 9472 10685 9512
rect 10627 9471 10685 9472
rect 12259 9512 12317 9513
rect 12259 9472 12268 9512
rect 12308 9472 12317 9512
rect 12259 9471 12317 9472
rect 13123 9512 13181 9513
rect 13123 9472 13132 9512
rect 13172 9472 13181 9512
rect 13123 9471 13181 9472
rect 16291 9512 16349 9513
rect 16291 9472 16300 9512
rect 16340 9472 16349 9512
rect 16291 9471 16349 9472
rect 17155 9512 17213 9513
rect 17155 9472 17164 9512
rect 17204 9472 17213 9512
rect 17155 9471 17213 9472
rect 19659 9512 19701 9521
rect 19659 9472 19660 9512
rect 19700 9472 19701 9512
rect 19659 9463 19701 9472
rect 25899 9507 25941 9516
rect 25795 9470 25853 9471
rect 2947 9428 3005 9429
rect 2947 9388 2956 9428
rect 2996 9388 3005 9428
rect 2947 9387 3005 9388
rect 18891 9428 18933 9437
rect 25795 9430 25804 9470
rect 25844 9430 25853 9470
rect 25899 9467 25900 9507
rect 25940 9467 25941 9507
rect 25987 9512 26045 9513
rect 25987 9472 25996 9512
rect 26036 9472 26045 9512
rect 25987 9471 26045 9472
rect 26371 9512 26429 9513
rect 26371 9472 26380 9512
rect 26420 9472 26429 9512
rect 26371 9471 26429 9472
rect 26859 9512 26901 9521
rect 26859 9472 26860 9512
rect 26900 9472 26901 9512
rect 25899 9458 25941 9467
rect 26859 9463 26901 9472
rect 39907 9512 39965 9513
rect 39907 9472 39916 9512
rect 39956 9472 39965 9512
rect 39907 9471 39965 9472
rect 40771 9512 40829 9513
rect 40771 9472 40780 9512
rect 40820 9472 40829 9512
rect 40771 9471 40829 9472
rect 41347 9512 41405 9513
rect 41347 9472 41356 9512
rect 41396 9472 41405 9512
rect 41347 9471 41405 9472
rect 41547 9512 41589 9521
rect 41547 9472 41548 9512
rect 41588 9472 41589 9512
rect 41547 9463 41589 9472
rect 47299 9512 47357 9513
rect 47299 9472 47308 9512
rect 47348 9472 47357 9512
rect 47299 9471 47357 9472
rect 47683 9512 47741 9513
rect 47683 9472 47692 9512
rect 47732 9472 47741 9512
rect 47683 9471 47741 9472
rect 48547 9512 48605 9513
rect 48547 9472 48556 9512
rect 48596 9472 48605 9512
rect 48547 9471 48605 9472
rect 52291 9512 52349 9513
rect 52291 9472 52300 9512
rect 52340 9472 52349 9512
rect 52291 9471 52349 9472
rect 52867 9512 52925 9513
rect 52867 9472 52876 9512
rect 52916 9472 52925 9512
rect 52867 9471 52925 9472
rect 53059 9512 53117 9513
rect 53059 9472 53068 9512
rect 53108 9472 53117 9512
rect 53059 9471 53117 9472
rect 55267 9512 55325 9513
rect 55267 9472 55276 9512
rect 55316 9472 55325 9512
rect 55267 9471 55325 9472
rect 56131 9512 56189 9513
rect 56131 9472 56140 9512
rect 56180 9472 56189 9512
rect 56131 9471 56189 9472
rect 25795 9429 25853 9430
rect 18891 9388 18892 9428
rect 18932 9388 18933 9428
rect 18891 9379 18933 9388
rect 26179 9344 26237 9345
rect 26179 9304 26188 9344
rect 26228 9304 26237 9344
rect 26179 9303 26237 9304
rect 26859 9344 26901 9353
rect 26859 9304 26860 9344
rect 26900 9304 26901 9344
rect 26859 9295 26901 9304
rect 2763 9260 2805 9269
rect 2763 9220 2764 9260
rect 2804 9220 2805 9260
rect 2763 9211 2805 9220
rect 5539 9260 5597 9261
rect 5539 9220 5548 9260
rect 5588 9220 5597 9260
rect 5539 9219 5597 9220
rect 7363 9260 7421 9261
rect 7363 9220 7372 9260
rect 7412 9220 7421 9260
rect 7363 9219 7421 9220
rect 9955 9260 10013 9261
rect 9955 9220 9964 9260
rect 10004 9220 10013 9260
rect 9955 9219 10013 9220
rect 18307 9260 18365 9261
rect 18307 9220 18316 9260
rect 18356 9220 18365 9260
rect 18307 9219 18365 9220
rect 25515 9260 25557 9269
rect 25515 9220 25516 9260
rect 25556 9220 25557 9260
rect 25515 9211 25557 9220
rect 26667 9260 26709 9269
rect 26667 9220 26668 9260
rect 26708 9220 26709 9260
rect 26667 9211 26709 9220
rect 38755 9260 38813 9261
rect 38755 9220 38764 9260
rect 38804 9220 38813 9260
rect 38755 9219 38813 9220
rect 41451 9260 41493 9269
rect 41451 9220 41452 9260
rect 41492 9220 41493 9260
rect 41451 9211 41493 9220
rect 51819 9260 51861 9269
rect 51819 9220 51820 9260
rect 51860 9220 51861 9260
rect 51819 9211 51861 9220
rect 576 9092 99360 9116
rect 576 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 18232 9092
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18600 9052 33352 9092
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33720 9052 48472 9092
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48840 9052 63592 9092
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63960 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 93832 9092
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 94200 9052 99360 9092
rect 576 9028 99360 9052
rect 4387 8924 4445 8925
rect 4387 8884 4396 8924
rect 4436 8884 4445 8924
rect 4387 8883 4445 8884
rect 47875 8924 47933 8925
rect 47875 8884 47884 8924
rect 47924 8884 47933 8924
rect 47875 8883 47933 8884
rect 7171 8840 7229 8841
rect 7171 8800 7180 8840
rect 7220 8800 7229 8840
rect 7171 8799 7229 8800
rect 9763 8840 9821 8841
rect 9763 8800 9772 8840
rect 9812 8800 9821 8840
rect 9763 8799 9821 8800
rect 12355 8840 12413 8841
rect 12355 8800 12364 8840
rect 12404 8800 12413 8840
rect 12355 8799 12413 8800
rect 19179 8840 19221 8849
rect 19179 8800 19180 8840
rect 19220 8800 19221 8840
rect 19179 8791 19221 8800
rect 30027 8840 30069 8849
rect 30027 8800 30028 8840
rect 30068 8800 30069 8840
rect 30027 8791 30069 8800
rect 40195 8840 40253 8841
rect 40195 8800 40204 8840
rect 40244 8800 40253 8840
rect 40195 8799 40253 8800
rect 40579 8756 40637 8757
rect 40579 8716 40588 8756
rect 40628 8716 40637 8756
rect 40579 8715 40637 8716
rect 2371 8672 2429 8673
rect 2371 8632 2380 8672
rect 2420 8632 2429 8672
rect 2371 8631 2429 8632
rect 3235 8672 3293 8673
rect 3235 8632 3244 8672
rect 3284 8632 3293 8672
rect 3235 8631 3293 8632
rect 4779 8672 4821 8681
rect 4779 8632 4780 8672
rect 4820 8632 4821 8672
rect 4779 8623 4821 8632
rect 5155 8672 5213 8673
rect 5155 8632 5164 8672
rect 5204 8632 5213 8672
rect 5155 8631 5213 8632
rect 6019 8672 6077 8673
rect 6019 8632 6028 8672
rect 6068 8632 6077 8672
rect 6019 8631 6077 8632
rect 7371 8672 7413 8681
rect 7371 8632 7372 8672
rect 7412 8632 7413 8672
rect 7371 8623 7413 8632
rect 7747 8672 7805 8673
rect 7747 8632 7756 8672
rect 7796 8632 7805 8672
rect 7747 8631 7805 8632
rect 8611 8672 8669 8673
rect 8611 8632 8620 8672
rect 8660 8632 8669 8672
rect 8611 8631 8669 8632
rect 9963 8672 10005 8681
rect 9963 8632 9964 8672
rect 10004 8632 10005 8672
rect 9963 8623 10005 8632
rect 10339 8672 10397 8673
rect 10339 8632 10348 8672
rect 10388 8632 10397 8672
rect 10339 8631 10397 8632
rect 11203 8672 11261 8673
rect 11203 8632 11212 8672
rect 11252 8632 11261 8672
rect 11203 8631 11261 8632
rect 19371 8672 19413 8681
rect 19371 8632 19372 8672
rect 19412 8632 19413 8672
rect 19371 8623 19413 8632
rect 19755 8672 19797 8681
rect 19755 8632 19756 8672
rect 19796 8632 19797 8672
rect 19755 8623 19797 8632
rect 19939 8672 19997 8673
rect 19939 8632 19948 8672
rect 19988 8632 19997 8672
rect 19939 8631 19997 8632
rect 20907 8672 20949 8681
rect 20907 8632 20908 8672
rect 20948 8632 20949 8672
rect 20907 8623 20949 8632
rect 21099 8672 21141 8681
rect 21099 8632 21100 8672
rect 21140 8632 21141 8672
rect 21099 8623 21141 8632
rect 21571 8672 21629 8673
rect 21571 8632 21580 8672
rect 21620 8632 21629 8672
rect 21571 8631 21629 8632
rect 21675 8672 21717 8681
rect 21675 8632 21676 8672
rect 21716 8632 21717 8672
rect 21675 8623 21717 8632
rect 22059 8672 22101 8681
rect 22059 8632 22060 8672
rect 22100 8632 22101 8672
rect 22059 8623 22101 8632
rect 22243 8672 22301 8673
rect 22243 8632 22252 8672
rect 22292 8632 22301 8672
rect 22243 8631 22301 8632
rect 25995 8672 26037 8681
rect 25995 8632 25996 8672
rect 26036 8632 26037 8672
rect 25995 8623 26037 8632
rect 26091 8672 26133 8681
rect 26091 8632 26092 8672
rect 26132 8632 26133 8672
rect 26091 8623 26133 8632
rect 29347 8672 29405 8673
rect 29347 8632 29356 8672
rect 29396 8632 29405 8672
rect 29347 8631 29405 8632
rect 30027 8672 30069 8681
rect 30027 8632 30028 8672
rect 30068 8632 30069 8672
rect 30027 8623 30069 8632
rect 30219 8672 30261 8681
rect 30219 8632 30220 8672
rect 30260 8632 30261 8672
rect 30219 8623 30261 8632
rect 39043 8672 39101 8673
rect 39043 8632 39052 8672
rect 39092 8632 39101 8672
rect 39043 8631 39101 8632
rect 39523 8672 39581 8673
rect 39523 8632 39532 8672
rect 39572 8632 39581 8672
rect 39523 8631 39581 8632
rect 40771 8672 40829 8673
rect 40771 8632 40780 8672
rect 40820 8632 40829 8672
rect 40771 8631 40829 8632
rect 40867 8672 40925 8673
rect 40867 8632 40876 8672
rect 40916 8632 40925 8672
rect 40867 8631 40925 8632
rect 45859 8672 45917 8673
rect 45859 8632 45868 8672
rect 45908 8632 45917 8672
rect 45859 8631 45917 8632
rect 46723 8672 46781 8673
rect 46723 8632 46732 8672
rect 46772 8632 46781 8672
rect 46723 8631 46781 8632
rect 1995 8588 2037 8597
rect 1995 8548 1996 8588
rect 2036 8548 2037 8588
rect 1995 8539 2037 8548
rect 19851 8588 19893 8597
rect 19851 8548 19852 8588
rect 19892 8548 19893 8588
rect 19851 8539 19893 8548
rect 22155 8588 22197 8597
rect 22155 8548 22156 8588
rect 22196 8548 22197 8588
rect 22155 8539 22197 8548
rect 45483 8588 45525 8597
rect 45483 8548 45484 8588
rect 45524 8548 45525 8588
rect 45483 8539 45525 8548
rect 643 8504 701 8505
rect 643 8464 652 8504
rect 692 8464 701 8504
rect 643 8463 701 8464
rect 21003 8504 21045 8513
rect 21003 8464 21004 8504
rect 21044 8464 21045 8504
rect 21003 8455 21045 8464
rect 21291 8504 21333 8513
rect 21291 8464 21292 8504
rect 21332 8464 21333 8504
rect 21291 8455 21333 8464
rect 25795 8504 25853 8505
rect 25795 8464 25804 8504
rect 25844 8464 25853 8504
rect 25795 8463 25853 8464
rect 28675 8504 28733 8505
rect 28675 8464 28684 8504
rect 28724 8464 28733 8504
rect 28675 8463 28733 8464
rect 38371 8504 38429 8505
rect 38371 8464 38380 8504
rect 38420 8464 38429 8504
rect 38371 8463 38429 8464
rect 576 8336 99360 8360
rect 576 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 19472 8336
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19840 8296 34592 8336
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34960 8296 49712 8336
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 50080 8296 64832 8336
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 65200 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 95072 8336
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95440 8296 99360 8336
rect 576 8272 99360 8296
rect 643 8168 701 8169
rect 643 8128 652 8168
rect 692 8128 701 8168
rect 643 8127 701 8128
rect 2283 8168 2325 8177
rect 2283 8128 2284 8168
rect 2324 8128 2325 8168
rect 2283 8119 2325 8128
rect 5059 8168 5117 8169
rect 5059 8128 5068 8168
rect 5108 8128 5117 8168
rect 5059 8127 5117 8128
rect 9099 8168 9141 8177
rect 9099 8128 9100 8168
rect 9140 8128 9141 8168
rect 9099 8119 9141 8128
rect 21867 8168 21909 8177
rect 21867 8128 21868 8168
rect 21908 8128 21909 8168
rect 21867 8119 21909 8128
rect 23203 8168 23261 8169
rect 23203 8128 23212 8168
rect 23252 8128 23261 8168
rect 23203 8127 23261 8128
rect 24931 8168 24989 8169
rect 24931 8128 24940 8168
rect 24980 8128 24989 8168
rect 24931 8127 24989 8128
rect 29539 8168 29597 8169
rect 29539 8128 29548 8168
rect 29588 8128 29597 8168
rect 29539 8127 29597 8128
rect 45571 8168 45629 8169
rect 45571 8128 45580 8168
rect 45620 8128 45629 8168
rect 45571 8127 45629 8128
rect 2667 8084 2709 8093
rect 2667 8044 2668 8084
rect 2708 8044 2709 8084
rect 2667 8035 2709 8044
rect 18691 8084 18749 8085
rect 18691 8044 18700 8084
rect 18740 8044 18749 8084
rect 18691 8043 18749 8044
rect 27339 8084 27381 8093
rect 27339 8044 27340 8084
rect 27380 8044 27381 8084
rect 27339 8035 27381 8044
rect 39907 8084 39965 8085
rect 39907 8044 39916 8084
rect 39956 8044 39965 8084
rect 39907 8043 39965 8044
rect 3043 8000 3101 8001
rect 3043 7960 3052 8000
rect 3092 7960 3101 8000
rect 3043 7959 3101 7960
rect 3907 8000 3965 8001
rect 3907 7960 3916 8000
rect 3956 7960 3965 8000
rect 3907 7959 3965 7960
rect 8715 8000 8757 8009
rect 8715 7960 8716 8000
rect 8756 7960 8757 8000
rect 8715 7951 8757 7960
rect 18787 8000 18845 8001
rect 18787 7960 18796 8000
rect 18836 7960 18845 8000
rect 18787 7959 18845 7960
rect 19171 8000 19229 8001
rect 19171 7960 19180 8000
rect 19220 7960 19229 8000
rect 19171 7959 19229 7960
rect 22051 8000 22109 8001
rect 22051 7960 22060 8000
rect 22100 7960 22109 8000
rect 22051 7959 22109 7960
rect 22339 8000 22397 8001
rect 22339 7960 22348 8000
rect 22388 7960 22397 8000
rect 22339 7959 22397 7960
rect 22923 8000 22965 8009
rect 22923 7960 22924 8000
rect 22964 7960 22965 8000
rect 22923 7951 22965 7960
rect 23019 8000 23061 8009
rect 23019 7960 23020 8000
rect 23060 7960 23061 8000
rect 23019 7951 23061 7960
rect 23115 8000 23157 8009
rect 23115 7960 23116 8000
rect 23156 7960 23157 8000
rect 23115 7951 23157 7960
rect 26083 8000 26141 8001
rect 26083 7960 26092 8000
rect 26132 7960 26141 8000
rect 26083 7959 26141 7960
rect 26947 8000 27005 8001
rect 26947 7960 26956 8000
rect 26996 7960 27005 8000
rect 26947 7959 27005 7960
rect 29643 8000 29685 8009
rect 29643 7960 29644 8000
rect 29684 7960 29685 8000
rect 29643 7951 29685 7960
rect 29739 8000 29781 8009
rect 29739 7960 29740 8000
rect 29780 7960 29781 8000
rect 29739 7951 29781 7960
rect 29835 8000 29877 8009
rect 29835 7960 29836 8000
rect 29876 7960 29877 8000
rect 29835 7951 29877 7960
rect 30315 8000 30357 8009
rect 30315 7960 30316 8000
rect 30356 7960 30357 8000
rect 30315 7951 30357 7960
rect 30979 8000 31037 8001
rect 30979 7960 30988 8000
rect 31028 7960 31037 8000
rect 30979 7959 31037 7960
rect 32899 8000 32957 8001
rect 32899 7960 32908 8000
rect 32948 7960 32957 8000
rect 32899 7959 32957 7960
rect 33475 8000 33533 8001
rect 33475 7960 33484 8000
rect 33524 7960 33533 8000
rect 33475 7959 33533 7960
rect 34723 8000 34781 8001
rect 34723 7960 34732 8000
rect 34772 7960 34781 8000
rect 34723 7959 34781 7960
rect 35587 8000 35645 8001
rect 35587 7960 35596 8000
rect 35636 7960 35645 8000
rect 35587 7959 35645 7960
rect 35979 8000 36021 8009
rect 35979 7960 35980 8000
rect 36020 7960 36021 8000
rect 35979 7951 36021 7960
rect 37219 8000 37277 8001
rect 37219 7960 37228 8000
rect 37268 7960 37277 8000
rect 37219 7959 37277 7960
rect 37899 8000 37941 8009
rect 37899 7960 37900 8000
rect 37940 7960 37941 8000
rect 37899 7951 37941 7960
rect 38755 8000 38813 8001
rect 38755 7960 38764 8000
rect 38804 7960 38813 8000
rect 38755 7959 38813 7960
rect 40099 8000 40157 8001
rect 40099 7960 40108 8000
rect 40148 7960 40157 8000
rect 40099 7959 40157 7960
rect 40387 8000 40445 8001
rect 40387 7960 40396 8000
rect 40436 7960 40445 8000
rect 40387 7959 40445 7960
rect 46243 8000 46301 8001
rect 46243 7960 46252 8000
rect 46292 7960 46301 8000
rect 46243 7959 46301 7960
rect 50955 8000 50997 8009
rect 50955 7960 50956 8000
rect 50996 7960 50997 8000
rect 50955 7951 50997 7960
rect 2467 7916 2525 7917
rect 2467 7876 2476 7916
rect 2516 7876 2525 7916
rect 2467 7875 2525 7876
rect 38091 7832 38133 7841
rect 38091 7792 38092 7832
rect 38132 7792 38133 7832
rect 38091 7783 38133 7792
rect 32227 7748 32285 7749
rect 32227 7708 32236 7748
rect 32276 7708 32285 7748
rect 32227 7707 32285 7708
rect 36555 7748 36597 7757
rect 36555 7708 36556 7748
rect 36596 7708 36597 7748
rect 36555 7699 36597 7708
rect 51147 7748 51189 7757
rect 51147 7708 51148 7748
rect 51188 7708 51189 7748
rect 51147 7699 51189 7708
rect 576 7580 99360 7604
rect 576 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 18232 7580
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18600 7540 33352 7580
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33720 7540 48472 7580
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48840 7540 63592 7580
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63960 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 93832 7580
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 94200 7540 99360 7580
rect 576 7516 99360 7540
rect 18595 7412 18653 7413
rect 18595 7372 18604 7412
rect 18644 7372 18653 7412
rect 18595 7371 18653 7372
rect 20323 7412 20381 7413
rect 20323 7372 20332 7412
rect 20372 7372 20381 7412
rect 20323 7371 20381 7372
rect 30699 7412 30741 7421
rect 30699 7372 30700 7412
rect 30740 7372 30741 7412
rect 30699 7363 30741 7372
rect 50755 7412 50813 7413
rect 50755 7372 50764 7412
rect 50804 7372 50813 7412
rect 50755 7371 50813 7372
rect 29059 7244 29117 7245
rect 29059 7204 29068 7244
rect 29108 7204 29117 7244
rect 29059 7203 29117 7204
rect 10915 7160 10973 7161
rect 10915 7120 10924 7160
rect 10964 7120 10973 7160
rect 10915 7119 10973 7120
rect 11787 7160 11829 7169
rect 11787 7120 11788 7160
rect 11828 7120 11829 7160
rect 11787 7111 11829 7120
rect 16203 7160 16245 7169
rect 16203 7120 16204 7160
rect 16244 7120 16245 7160
rect 16203 7111 16245 7120
rect 16579 7160 16637 7161
rect 16579 7120 16588 7160
rect 16628 7120 16637 7160
rect 16579 7119 16637 7120
rect 17443 7160 17501 7161
rect 17443 7120 17452 7160
rect 17492 7120 17501 7160
rect 17443 7119 17501 7120
rect 21475 7160 21533 7161
rect 21475 7120 21484 7160
rect 21524 7120 21533 7160
rect 21475 7119 21533 7120
rect 22339 7160 22397 7161
rect 22339 7120 22348 7160
rect 22388 7120 22397 7160
rect 22339 7119 22397 7120
rect 22923 7160 22965 7169
rect 22923 7120 22924 7160
rect 22964 7120 22965 7160
rect 22923 7111 22965 7120
rect 23587 7160 23645 7161
rect 23587 7120 23596 7160
rect 23636 7120 23645 7160
rect 23587 7119 23645 7120
rect 26659 7160 26717 7161
rect 26659 7120 26668 7160
rect 26708 7120 26717 7160
rect 26659 7119 26717 7120
rect 28579 7160 28637 7161
rect 28579 7120 28588 7160
rect 28628 7120 28637 7160
rect 28579 7119 28637 7120
rect 28867 7160 28925 7161
rect 28867 7120 28876 7160
rect 28916 7120 28925 7160
rect 28867 7119 28925 7120
rect 29347 7160 29405 7161
rect 29347 7120 29356 7160
rect 29396 7120 29405 7160
rect 29347 7119 29405 7120
rect 29451 7160 29493 7169
rect 29451 7120 29452 7160
rect 29492 7120 29493 7160
rect 29451 7111 29493 7120
rect 30019 7160 30077 7161
rect 30019 7120 30028 7160
rect 30068 7120 30077 7160
rect 30019 7119 30077 7120
rect 30403 7160 30461 7161
rect 30403 7120 30412 7160
rect 30452 7120 30461 7160
rect 30403 7119 30461 7120
rect 30603 7160 30645 7169
rect 30603 7120 30604 7160
rect 30644 7120 30645 7160
rect 30603 7111 30645 7120
rect 30787 7160 30845 7161
rect 30787 7120 30796 7160
rect 30836 7120 30845 7160
rect 30787 7119 30845 7120
rect 32323 7160 32381 7161
rect 32323 7120 32332 7160
rect 32372 7120 32381 7160
rect 32323 7119 32381 7120
rect 34627 7160 34685 7161
rect 34627 7120 34636 7160
rect 34676 7120 34685 7160
rect 34627 7119 34685 7120
rect 35491 7160 35549 7161
rect 35491 7120 35500 7160
rect 35540 7120 35549 7160
rect 35491 7119 35549 7120
rect 38659 7160 38717 7161
rect 38659 7120 38668 7160
rect 38708 7120 38717 7160
rect 38659 7119 38717 7120
rect 40195 7160 40253 7161
rect 40195 7120 40204 7160
rect 40244 7120 40253 7160
rect 40195 7119 40253 7120
rect 48739 7160 48797 7161
rect 48739 7120 48748 7160
rect 48788 7120 48797 7160
rect 48739 7119 48797 7120
rect 49603 7160 49661 7161
rect 49603 7120 49612 7160
rect 49652 7120 49661 7160
rect 49603 7119 49661 7120
rect 22731 7076 22773 7085
rect 22731 7036 22732 7076
rect 22772 7036 22773 7076
rect 22731 7027 22773 7036
rect 25995 7076 26037 7085
rect 25995 7036 25996 7076
rect 26036 7036 26037 7076
rect 25995 7027 26037 7036
rect 35883 7076 35925 7085
rect 35883 7036 35884 7076
rect 35924 7036 35925 7076
rect 35883 7027 35925 7036
rect 37995 7076 38037 7085
rect 37995 7036 37996 7076
rect 38036 7036 38037 7076
rect 37995 7027 38037 7036
rect 48363 7076 48405 7085
rect 48363 7036 48364 7076
rect 48404 7036 48405 7076
rect 48363 7027 48405 7036
rect 643 6992 701 6993
rect 643 6952 652 6992
rect 692 6952 701 6992
rect 643 6951 701 6952
rect 28395 6992 28437 7001
rect 28395 6952 28396 6992
rect 28436 6952 28437 6992
rect 28395 6943 28437 6952
rect 29931 6992 29973 7001
rect 29931 6952 29932 6992
rect 29972 6952 29973 6992
rect 29931 6943 29973 6952
rect 31651 6992 31709 6993
rect 31651 6952 31660 6992
rect 31700 6952 31709 6992
rect 31651 6951 31709 6952
rect 33475 6992 33533 6993
rect 33475 6952 33484 6992
rect 33524 6952 33533 6992
rect 33475 6951 33533 6952
rect 39523 6992 39581 6993
rect 39523 6952 39532 6992
rect 39572 6952 39581 6992
rect 39523 6951 39581 6952
rect 576 6824 99360 6848
rect 576 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 19472 6824
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19840 6784 34592 6824
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34960 6784 49712 6824
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 50080 6784 64832 6824
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 65200 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 95072 6824
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95440 6784 99360 6824
rect 576 6760 99360 6784
rect 29443 6656 29501 6657
rect 29443 6616 29452 6656
rect 29492 6616 29501 6656
rect 29443 6615 29501 6616
rect 39819 6656 39861 6665
rect 39819 6616 39820 6656
rect 39860 6616 39861 6656
rect 39819 6607 39861 6616
rect 45291 6656 45333 6665
rect 45291 6616 45292 6656
rect 45332 6616 45333 6656
rect 45291 6607 45333 6616
rect 48643 6656 48701 6657
rect 48643 6616 48652 6656
rect 48692 6616 48701 6656
rect 48643 6615 48701 6616
rect 29739 6572 29781 6581
rect 29739 6532 29740 6572
rect 29780 6532 29781 6572
rect 29739 6523 29781 6532
rect 21571 6488 21629 6489
rect 21571 6448 21580 6488
rect 21620 6448 21629 6488
rect 21571 6447 21629 6448
rect 22531 6488 22589 6489
rect 22531 6448 22540 6488
rect 22580 6448 22589 6488
rect 22531 6447 22589 6448
rect 28771 6488 28829 6489
rect 28771 6448 28780 6488
rect 28820 6448 28829 6488
rect 28771 6447 28829 6448
rect 29643 6488 29685 6497
rect 29643 6448 29644 6488
rect 29684 6448 29685 6488
rect 29643 6439 29685 6448
rect 29827 6488 29885 6489
rect 29827 6448 29836 6488
rect 29876 6448 29885 6488
rect 29827 6447 29885 6448
rect 39331 6488 39389 6489
rect 39331 6448 39340 6488
rect 39380 6448 39389 6488
rect 39331 6447 39389 6448
rect 44803 6488 44861 6489
rect 44803 6448 44812 6488
rect 44852 6448 44861 6488
rect 44803 6447 44861 6448
rect 45187 6488 45245 6489
rect 45187 6448 45196 6488
rect 45236 6448 45245 6488
rect 45187 6447 45245 6448
rect 45571 6488 45629 6489
rect 45571 6448 45580 6488
rect 45620 6448 45629 6488
rect 45571 6447 45629 6448
rect 46251 6488 46293 6497
rect 46251 6448 46252 6488
rect 46292 6448 46293 6488
rect 46251 6439 46293 6448
rect 47971 6488 48029 6489
rect 47971 6448 47980 6488
rect 48020 6448 48029 6488
rect 47971 6447 48029 6448
rect 53731 6488 53789 6489
rect 53731 6448 53740 6488
rect 53780 6448 53789 6488
rect 53731 6447 53789 6448
rect 54019 6488 54077 6489
rect 54019 6448 54028 6488
rect 54068 6448 54077 6488
rect 54019 6447 54077 6448
rect 38755 6404 38813 6405
rect 38755 6364 38764 6404
rect 38804 6364 38813 6404
rect 38755 6363 38813 6364
rect 21867 6320 21909 6329
rect 21867 6280 21868 6320
rect 21908 6280 21909 6320
rect 21867 6271 21909 6280
rect 38571 6320 38613 6329
rect 38571 6280 38572 6320
rect 38612 6280 38613 6320
rect 38571 6271 38613 6280
rect 39627 6320 39669 6329
rect 39627 6280 39628 6320
rect 39668 6280 39669 6320
rect 39627 6271 39669 6280
rect 53059 6320 53117 6321
rect 53059 6280 53068 6320
rect 53108 6280 53117 6320
rect 53059 6279 53117 6280
rect 54315 6320 54357 6329
rect 54315 6280 54316 6320
rect 54356 6280 54357 6320
rect 54315 6271 54357 6280
rect 576 6068 99360 6092
rect 576 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 18232 6068
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18600 6028 33352 6068
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33720 6028 48472 6068
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48840 6028 63592 6068
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63960 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 93832 6068
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 94200 6028 99360 6068
rect 576 6004 99360 6028
rect 40099 5900 40157 5901
rect 40099 5860 40108 5900
rect 40148 5860 40157 5900
rect 40099 5859 40157 5860
rect 47403 5900 47445 5909
rect 47403 5860 47404 5900
rect 47444 5860 47445 5900
rect 47403 5851 47445 5860
rect 48363 5900 48405 5909
rect 48363 5860 48364 5900
rect 48404 5860 48405 5900
rect 48363 5851 48405 5860
rect 54979 5900 55037 5901
rect 54979 5860 54988 5900
rect 55028 5860 55037 5900
rect 54979 5859 55037 5860
rect 52195 5732 52253 5733
rect 52195 5692 52204 5732
rect 52244 5692 52253 5732
rect 52195 5691 52253 5692
rect 13027 5648 13085 5649
rect 13027 5608 13036 5648
rect 13076 5608 13085 5648
rect 13027 5607 13085 5608
rect 15139 5648 15197 5649
rect 15139 5608 15148 5648
rect 15188 5608 15197 5648
rect 15139 5607 15197 5608
rect 16099 5648 16157 5649
rect 16099 5608 16108 5648
rect 16148 5608 16157 5648
rect 16099 5607 16157 5608
rect 18115 5648 18173 5649
rect 18115 5608 18124 5648
rect 18164 5608 18173 5648
rect 18115 5607 18173 5608
rect 33859 5648 33917 5649
rect 33859 5608 33868 5648
rect 33908 5608 33917 5648
rect 33859 5607 33917 5608
rect 37707 5648 37749 5657
rect 37707 5608 37708 5648
rect 37748 5608 37749 5648
rect 37707 5599 37749 5608
rect 38083 5648 38141 5649
rect 38083 5608 38092 5648
rect 38132 5608 38141 5648
rect 38083 5607 38141 5608
rect 38947 5648 39005 5649
rect 38947 5608 38956 5648
rect 38996 5608 39005 5648
rect 38947 5607 39005 5608
rect 45283 5648 45341 5649
rect 45283 5608 45292 5648
rect 45332 5608 45341 5648
rect 45283 5607 45341 5608
rect 46443 5648 46485 5657
rect 46443 5608 46444 5648
rect 46484 5608 46485 5648
rect 46443 5599 46485 5608
rect 46539 5648 46581 5657
rect 46539 5608 46540 5648
rect 46580 5608 46581 5648
rect 46539 5599 46581 5608
rect 46627 5648 46685 5649
rect 46627 5608 46636 5648
rect 46676 5608 46685 5648
rect 46627 5607 46685 5608
rect 47203 5648 47261 5649
rect 47203 5608 47212 5648
rect 47252 5608 47261 5648
rect 47203 5607 47261 5608
rect 47299 5648 47357 5649
rect 47299 5608 47308 5648
rect 47348 5608 47357 5648
rect 47299 5607 47357 5608
rect 48643 5648 48701 5649
rect 48643 5608 48652 5648
rect 48692 5608 48701 5648
rect 48643 5607 48701 5608
rect 52963 5648 53021 5649
rect 52963 5608 52972 5648
rect 53012 5608 53021 5648
rect 52963 5607 53021 5608
rect 53827 5648 53885 5649
rect 53827 5608 53836 5648
rect 53876 5608 53885 5648
rect 53827 5607 53885 5608
rect 56611 5648 56669 5649
rect 56611 5608 56620 5648
rect 56660 5608 56669 5648
rect 56611 5607 56669 5608
rect 17251 5564 17309 5565
rect 17251 5524 17260 5564
rect 17300 5524 17309 5564
rect 17251 5523 17309 5524
rect 45963 5564 46005 5573
rect 45963 5524 45964 5564
rect 46004 5524 46005 5564
rect 45963 5515 46005 5524
rect 52587 5564 52629 5573
rect 52587 5524 52588 5564
rect 52628 5524 52629 5564
rect 52587 5515 52629 5524
rect 643 5480 701 5481
rect 643 5440 652 5480
rect 692 5440 701 5480
rect 643 5439 701 5440
rect 12355 5480 12413 5481
rect 12355 5440 12364 5480
rect 12404 5440 12413 5480
rect 12355 5439 12413 5440
rect 15627 5480 15669 5489
rect 15627 5440 15628 5480
rect 15668 5440 15669 5480
rect 15627 5431 15669 5440
rect 33387 5480 33429 5489
rect 33387 5440 33388 5480
rect 33428 5440 33429 5480
rect 33387 5431 33429 5440
rect 48171 5480 48213 5489
rect 48171 5440 48172 5480
rect 48212 5440 48213 5480
rect 48171 5431 48213 5440
rect 52395 5480 52437 5489
rect 52395 5440 52396 5480
rect 52436 5440 52437 5480
rect 52395 5431 52437 5440
rect 55939 5480 55997 5481
rect 55939 5440 55948 5480
rect 55988 5440 55997 5480
rect 55939 5439 55997 5440
rect 576 5312 99360 5336
rect 576 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 95072 5312
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95440 5272 99360 5312
rect 576 5248 99360 5272
rect 43651 5144 43709 5145
rect 43651 5104 43660 5144
rect 43700 5104 43709 5144
rect 43651 5103 43709 5104
rect 52195 5144 52253 5145
rect 52195 5104 52204 5144
rect 52244 5104 52253 5144
rect 52195 5103 52253 5104
rect 47691 5060 47733 5069
rect 47691 5020 47692 5060
rect 47732 5020 47733 5060
rect 47691 5011 47733 5020
rect 51907 5060 51965 5061
rect 51907 5020 51916 5060
rect 51956 5020 51965 5060
rect 51907 5019 51965 5020
rect 11499 4976 11541 4985
rect 11499 4936 11500 4976
rect 11540 4936 11541 4976
rect 11499 4927 11541 4936
rect 11875 4976 11933 4977
rect 11875 4936 11884 4976
rect 11924 4936 11933 4976
rect 11875 4935 11933 4936
rect 12739 4976 12797 4977
rect 12739 4936 12748 4976
rect 12788 4936 12797 4976
rect 12739 4935 12797 4936
rect 25603 4976 25661 4977
rect 25603 4936 25612 4976
rect 25652 4936 25661 4976
rect 25603 4935 25661 4936
rect 26283 4976 26325 4985
rect 26283 4936 26284 4976
rect 26324 4936 26325 4976
rect 26283 4927 26325 4936
rect 26475 4976 26517 4985
rect 26475 4936 26476 4976
rect 26516 4936 26517 4976
rect 26475 4927 26517 4936
rect 26851 4976 26909 4977
rect 26851 4936 26860 4976
rect 26900 4936 26909 4976
rect 26851 4935 26909 4936
rect 27715 4976 27773 4977
rect 27715 4936 27724 4976
rect 27764 4936 27773 4976
rect 27715 4935 27773 4936
rect 41259 4976 41301 4985
rect 41259 4936 41260 4976
rect 41300 4936 41301 4976
rect 41259 4927 41301 4936
rect 41635 4976 41693 4977
rect 41635 4936 41644 4976
rect 41684 4936 41693 4976
rect 41635 4935 41693 4936
rect 42499 4976 42557 4977
rect 42499 4936 42508 4976
rect 42548 4936 42557 4976
rect 42499 4935 42557 4936
rect 46435 4976 46493 4977
rect 46435 4936 46444 4976
rect 46484 4936 46493 4976
rect 46435 4935 46493 4936
rect 47299 4976 47357 4977
rect 47299 4936 47308 4976
rect 47348 4936 47357 4976
rect 47299 4935 47357 4936
rect 52099 4976 52157 4977
rect 52099 4936 52108 4976
rect 52148 4936 52157 4976
rect 52099 4935 52157 4936
rect 54795 4976 54837 4985
rect 54795 4936 54796 4976
rect 54836 4936 54837 4976
rect 54795 4927 54837 4936
rect 55171 4976 55229 4977
rect 55171 4936 55180 4976
rect 55220 4936 55229 4976
rect 55171 4935 55229 4936
rect 56035 4976 56093 4977
rect 56035 4936 56044 4976
rect 56084 4936 56093 4976
rect 56035 4935 56093 4936
rect 835 4892 893 4893
rect 835 4852 844 4892
rect 884 4852 893 4892
rect 835 4851 893 4852
rect 28875 4892 28917 4901
rect 28875 4852 28876 4892
rect 28916 4852 28917 4892
rect 28875 4843 28917 4852
rect 39235 4892 39293 4893
rect 39235 4852 39244 4892
rect 39284 4852 39293 4892
rect 39235 4851 39293 4852
rect 45291 4892 45333 4901
rect 45291 4852 45292 4892
rect 45332 4852 45333 4892
rect 45291 4843 45333 4852
rect 54403 4892 54461 4893
rect 54403 4852 54412 4892
rect 54452 4852 54461 4892
rect 54403 4851 54461 4852
rect 57195 4892 57237 4901
rect 57195 4852 57196 4892
rect 57236 4852 57237 4892
rect 57195 4843 57237 4852
rect 651 4808 693 4817
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 54603 4808 54645 4817
rect 54603 4768 54604 4808
rect 54644 4768 54645 4808
rect 54603 4759 54645 4768
rect 13891 4724 13949 4725
rect 13891 4684 13900 4724
rect 13940 4684 13949 4724
rect 13891 4683 13949 4684
rect 576 4556 99360 4580
rect 576 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 93832 4556
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 94200 4516 99360 4556
rect 576 4492 99360 4516
rect 13603 4388 13661 4389
rect 13603 4348 13612 4388
rect 13652 4348 13661 4388
rect 13603 4347 13661 4348
rect 30307 4388 30365 4389
rect 30307 4348 30316 4388
rect 30356 4348 30365 4388
rect 30307 4347 30365 4348
rect 40675 4388 40733 4389
rect 40675 4348 40684 4388
rect 40724 4348 40733 4388
rect 40675 4347 40733 4348
rect 835 4220 893 4221
rect 835 4180 844 4220
rect 884 4180 893 4220
rect 835 4179 893 4180
rect 10819 4220 10877 4221
rect 10819 4180 10828 4220
rect 10868 4180 10877 4220
rect 10819 4179 10877 4180
rect 23787 4220 23829 4229
rect 23787 4180 23788 4220
rect 23828 4180 23829 4220
rect 23787 4171 23829 4180
rect 34435 4220 34493 4221
rect 34435 4180 34444 4220
rect 34484 4180 34493 4220
rect 34435 4179 34493 4180
rect 38955 4220 38997 4229
rect 38955 4180 38956 4220
rect 38996 4180 38997 4220
rect 38955 4171 38997 4180
rect 11587 4136 11645 4137
rect 11587 4096 11596 4136
rect 11636 4096 11645 4136
rect 11587 4095 11645 4096
rect 12451 4136 12509 4137
rect 12451 4096 12460 4136
rect 12500 4096 12509 4136
rect 12451 4095 12509 4096
rect 20515 4136 20573 4137
rect 20515 4096 20524 4136
rect 20564 4096 20573 4136
rect 20515 4095 20573 4096
rect 21763 4136 21821 4137
rect 21763 4096 21772 4136
rect 21812 4096 21821 4136
rect 21763 4095 21821 4096
rect 22627 4136 22685 4137
rect 22627 4096 22636 4136
rect 22676 4096 22685 4136
rect 22627 4095 22685 4096
rect 24355 4136 24413 4137
rect 24355 4096 24364 4136
rect 24404 4096 24413 4136
rect 24355 4095 24413 4096
rect 27043 4136 27101 4137
rect 27043 4096 27052 4136
rect 27092 4096 27101 4136
rect 27043 4095 27101 4096
rect 28291 4136 28349 4137
rect 28291 4096 28300 4136
rect 28340 4096 28349 4136
rect 28291 4095 28349 4096
rect 29155 4136 29213 4137
rect 29155 4096 29164 4136
rect 29204 4096 29213 4136
rect 29155 4095 29213 4096
rect 38275 4136 38333 4137
rect 38275 4096 38284 4136
rect 38324 4096 38333 4136
rect 38275 4095 38333 4096
rect 40011 4136 40053 4145
rect 40011 4096 40012 4136
rect 40052 4096 40053 4136
rect 40011 4087 40053 4096
rect 40107 4136 40149 4145
rect 40107 4096 40108 4136
rect 40148 4096 40149 4136
rect 40107 4087 40149 4096
rect 40195 4136 40253 4137
rect 40195 4096 40204 4136
rect 40244 4096 40253 4136
rect 40195 4095 40253 4096
rect 40483 4136 40541 4137
rect 40483 4096 40492 4136
rect 40532 4096 40541 4136
rect 40483 4095 40541 4096
rect 41059 4136 41117 4137
rect 41059 4096 41068 4136
rect 41108 4096 41117 4136
rect 41059 4095 41117 4096
rect 41347 4136 41405 4137
rect 41347 4096 41356 4136
rect 41396 4096 41405 4136
rect 41347 4095 41405 4096
rect 54019 4136 54077 4137
rect 54019 4096 54028 4136
rect 54068 4096 54077 4136
rect 54019 4095 54077 4096
rect 54219 4136 54261 4145
rect 54219 4096 54220 4136
rect 54260 4096 54261 4136
rect 54219 4087 54261 4096
rect 56515 4136 56573 4137
rect 56515 4096 56524 4136
rect 56564 4096 56573 4136
rect 56515 4095 56573 4096
rect 11211 4052 11253 4061
rect 11211 4012 11212 4052
rect 11252 4012 11253 4052
rect 11211 4003 11253 4012
rect 21195 4052 21237 4061
rect 21195 4012 21196 4052
rect 21236 4012 21237 4052
rect 21195 4003 21237 4012
rect 21387 4052 21429 4061
rect 21387 4012 21388 4052
rect 21428 4012 21429 4052
rect 21387 4003 21429 4012
rect 27915 4052 27957 4061
rect 27915 4012 27916 4052
rect 27956 4012 27957 4052
rect 27915 4003 27957 4012
rect 54123 4052 54165 4061
rect 54123 4012 54124 4052
rect 54164 4012 54165 4052
rect 54123 4003 54165 4012
rect 651 3968 693 3977
rect 651 3928 652 3968
rect 692 3928 693 3968
rect 651 3919 693 3928
rect 11019 3968 11061 3977
rect 11019 3928 11020 3968
rect 11060 3928 11061 3968
rect 11019 3919 11061 3928
rect 25027 3968 25085 3969
rect 25027 3928 25036 3968
rect 25076 3928 25085 3968
rect 25027 3927 25085 3928
rect 27715 3968 27773 3969
rect 27715 3928 27724 3968
rect 27764 3928 27773 3968
rect 27715 3927 27773 3928
rect 34251 3968 34293 3977
rect 34251 3928 34252 3968
rect 34292 3928 34293 3968
rect 34251 3919 34293 3928
rect 40387 3968 40445 3969
rect 40387 3928 40396 3968
rect 40436 3928 40445 3968
rect 40387 3927 40445 3928
rect 41547 3968 41589 3977
rect 41547 3928 41548 3968
rect 41588 3928 41589 3968
rect 41547 3919 41589 3928
rect 55843 3968 55901 3969
rect 55843 3928 55852 3968
rect 55892 3928 55901 3968
rect 55843 3927 55901 3928
rect 576 3800 99360 3824
rect 576 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 95072 3800
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95440 3760 99360 3800
rect 576 3736 99360 3760
rect 11787 3632 11829 3641
rect 11787 3592 11788 3632
rect 11828 3592 11829 3632
rect 11787 3583 11829 3592
rect 12547 3632 12605 3633
rect 12547 3592 12556 3632
rect 12596 3592 12605 3632
rect 12547 3591 12605 3592
rect 20035 3632 20093 3633
rect 20035 3592 20044 3632
rect 20084 3592 20093 3632
rect 20035 3591 20093 3592
rect 24547 3632 24605 3633
rect 24547 3592 24556 3632
rect 24596 3592 24605 3632
rect 24547 3591 24605 3592
rect 27139 3632 27197 3633
rect 27139 3592 27148 3632
rect 27188 3592 27197 3632
rect 27139 3591 27197 3592
rect 35779 3632 35837 3633
rect 35779 3592 35788 3632
rect 35828 3592 35837 3632
rect 35779 3591 35837 3592
rect 47595 3632 47637 3641
rect 47595 3592 47596 3632
rect 47636 3592 47637 3632
rect 47595 3583 47637 3592
rect 52291 3632 52349 3633
rect 52291 3592 52300 3632
rect 52340 3592 52349 3632
rect 52291 3591 52349 3592
rect 53643 3632 53685 3641
rect 53643 3592 53644 3632
rect 53684 3592 53685 3632
rect 53643 3583 53685 3592
rect 56803 3632 56861 3633
rect 56803 3592 56812 3632
rect 56852 3592 56861 3632
rect 56803 3591 56861 3592
rect 13035 3548 13077 3557
rect 13035 3508 13036 3548
rect 13076 3508 13077 3548
rect 13035 3499 13077 3508
rect 24747 3548 24789 3557
rect 24747 3508 24748 3548
rect 24788 3508 24789 3548
rect 24747 3499 24789 3508
rect 33387 3548 33429 3557
rect 33387 3508 33388 3548
rect 33428 3508 33429 3548
rect 33387 3499 33429 3508
rect 40299 3548 40341 3557
rect 40299 3508 40300 3548
rect 40340 3508 40341 3548
rect 40299 3499 40341 3508
rect 52011 3548 52053 3557
rect 52011 3508 52012 3548
rect 52052 3508 52053 3548
rect 52011 3499 52053 3508
rect 7083 3464 7125 3473
rect 7083 3424 7084 3464
rect 7124 3424 7125 3464
rect 7083 3415 7125 3424
rect 7459 3464 7517 3465
rect 7459 3424 7468 3464
rect 7508 3424 7517 3464
rect 7459 3423 7517 3424
rect 8323 3464 8381 3465
rect 8323 3424 8332 3464
rect 8372 3424 8381 3464
rect 8323 3423 8381 3424
rect 10923 3464 10965 3473
rect 10923 3424 10924 3464
rect 10964 3424 10965 3464
rect 10923 3415 10965 3424
rect 11107 3464 11165 3465
rect 11107 3424 11116 3464
rect 11156 3424 11165 3464
rect 11107 3423 11165 3424
rect 11307 3464 11349 3473
rect 11307 3424 11308 3464
rect 11348 3424 11349 3464
rect 11307 3415 11349 3424
rect 11491 3464 11549 3465
rect 11491 3424 11500 3464
rect 11540 3424 11549 3464
rect 11491 3423 11549 3424
rect 12643 3464 12701 3465
rect 12643 3424 12652 3464
rect 12692 3424 12701 3464
rect 12643 3423 12701 3424
rect 13699 3464 13757 3465
rect 13699 3424 13708 3464
rect 13748 3424 13757 3464
rect 13699 3423 13757 3424
rect 17643 3464 17685 3473
rect 17643 3424 17644 3464
rect 17684 3424 17685 3464
rect 17643 3415 17685 3424
rect 18019 3464 18077 3465
rect 18019 3424 18028 3464
rect 18068 3424 18077 3464
rect 18019 3423 18077 3424
rect 18883 3464 18941 3465
rect 18883 3424 18892 3464
rect 18932 3424 18941 3464
rect 18883 3423 18941 3424
rect 21091 3464 21149 3465
rect 21091 3424 21100 3464
rect 21140 3424 21149 3464
rect 21091 3423 21149 3424
rect 21771 3464 21813 3473
rect 21771 3424 21772 3464
rect 21812 3424 21813 3464
rect 21771 3415 21813 3424
rect 22155 3464 22197 3473
rect 22155 3424 22156 3464
rect 22196 3424 22197 3464
rect 22155 3415 22197 3424
rect 22531 3464 22589 3465
rect 22531 3424 22540 3464
rect 22580 3424 22589 3464
rect 22531 3423 22589 3424
rect 23395 3464 23453 3465
rect 23395 3424 23404 3464
rect 23444 3424 23453 3464
rect 23395 3423 23453 3424
rect 25123 3464 25181 3465
rect 25123 3424 25132 3464
rect 25172 3424 25181 3464
rect 25123 3423 25181 3424
rect 25987 3464 26045 3465
rect 25987 3424 25996 3464
rect 26036 3424 26045 3464
rect 25987 3423 26045 3424
rect 33763 3464 33821 3465
rect 33763 3424 33772 3464
rect 33812 3424 33821 3464
rect 33763 3423 33821 3424
rect 34627 3464 34685 3465
rect 34627 3424 34636 3464
rect 34676 3424 34685 3464
rect 34627 3423 34685 3424
rect 38851 3464 38909 3465
rect 38851 3424 38860 3464
rect 38900 3424 38909 3464
rect 38851 3423 38909 3424
rect 40203 3464 40245 3473
rect 40203 3424 40204 3464
rect 40244 3424 40245 3464
rect 40203 3415 40245 3424
rect 40387 3464 40445 3465
rect 40387 3424 40396 3464
rect 40436 3424 40445 3464
rect 40387 3423 40445 3424
rect 40971 3464 41013 3473
rect 40971 3424 40972 3464
rect 41012 3424 41013 3464
rect 40971 3415 41013 3424
rect 41635 3464 41693 3465
rect 41635 3424 41644 3464
rect 41684 3424 41693 3464
rect 41635 3423 41693 3424
rect 47683 3464 47741 3465
rect 47683 3424 47692 3464
rect 47732 3424 47741 3464
rect 47683 3423 47741 3424
rect 48067 3464 48125 3465
rect 48067 3424 48076 3464
rect 48116 3424 48125 3464
rect 48067 3423 48125 3424
rect 51907 3464 51965 3465
rect 51907 3424 51916 3464
rect 51956 3424 51965 3464
rect 51907 3423 51965 3424
rect 52107 3464 52149 3473
rect 52107 3424 52108 3464
rect 52148 3424 52149 3464
rect 52107 3415 52149 3424
rect 52963 3464 53021 3465
rect 52963 3424 52972 3464
rect 53012 3424 53021 3464
rect 52963 3423 53021 3424
rect 53155 3464 53213 3465
rect 53155 3424 53164 3464
rect 53204 3424 53213 3464
rect 53155 3423 53213 3424
rect 53539 3464 53597 3465
rect 53539 3424 53548 3464
rect 53588 3424 53597 3464
rect 53539 3423 53597 3424
rect 54411 3464 54453 3473
rect 54411 3424 54412 3464
rect 54452 3424 54453 3464
rect 54411 3415 54453 3424
rect 54787 3464 54845 3465
rect 54787 3424 54796 3464
rect 54836 3424 54845 3464
rect 54787 3423 54845 3424
rect 55651 3464 55709 3465
rect 55651 3424 55660 3464
rect 55700 3424 55709 3464
rect 55651 3423 55709 3424
rect 835 3380 893 3381
rect 835 3340 844 3380
rect 884 3340 893 3380
rect 835 3339 893 3340
rect 11971 3380 12029 3381
rect 11971 3340 11980 3380
rect 12020 3340 12029 3380
rect 11971 3339 12029 3340
rect 38371 3380 38429 3381
rect 38371 3340 38380 3380
rect 38420 3340 38429 3380
rect 38371 3339 38429 3340
rect 39531 3380 39573 3389
rect 39531 3340 39532 3380
rect 39572 3340 39573 3380
rect 39531 3331 39573 3340
rect 40003 3380 40061 3381
rect 40003 3340 40012 3380
rect 40052 3340 40061 3380
rect 40003 3339 40061 3340
rect 51427 3380 51485 3381
rect 51427 3340 51436 3380
rect 51476 3340 51485 3380
rect 51427 3339 51485 3340
rect 651 3212 693 3221
rect 651 3172 652 3212
rect 692 3172 693 3212
rect 651 3163 693 3172
rect 9475 3212 9533 3213
rect 9475 3172 9484 3212
rect 9524 3172 9533 3212
rect 9475 3171 9533 3172
rect 11019 3212 11061 3221
rect 11019 3172 11020 3212
rect 11060 3172 11061 3212
rect 11019 3163 11061 3172
rect 11403 3212 11445 3221
rect 11403 3172 11404 3212
rect 11444 3172 11445 3212
rect 11403 3163 11445 3172
rect 12835 3212 12893 3213
rect 12835 3172 12844 3212
rect 12884 3172 12893 3212
rect 12835 3171 12893 3172
rect 38187 3212 38229 3221
rect 38187 3172 38188 3212
rect 38228 3172 38229 3212
rect 38187 3163 38229 3172
rect 39819 3212 39861 3221
rect 39819 3172 39820 3212
rect 39860 3172 39861 3212
rect 39819 3163 39861 3172
rect 51243 3212 51285 3221
rect 51243 3172 51244 3212
rect 51284 3172 51285 3212
rect 51243 3163 51285 3172
rect 576 3044 99360 3068
rect 576 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 93832 3044
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 94200 3004 99360 3044
rect 576 2980 99360 3004
rect 19843 2876 19901 2877
rect 19843 2836 19852 2876
rect 19892 2836 19901 2876
rect 19843 2835 19901 2836
rect 39139 2876 39197 2877
rect 39139 2836 39148 2876
rect 39188 2836 39197 2876
rect 39139 2835 39197 2836
rect 41731 2876 41789 2877
rect 41731 2836 41740 2876
rect 41780 2836 41789 2876
rect 41731 2835 41789 2836
rect 46435 2876 46493 2877
rect 46435 2836 46444 2876
rect 46484 2836 46493 2876
rect 46435 2835 46493 2836
rect 47107 2876 47165 2877
rect 47107 2836 47116 2876
rect 47156 2836 47165 2876
rect 47107 2835 47165 2836
rect 52867 2876 52925 2877
rect 52867 2836 52876 2876
rect 52916 2836 52925 2876
rect 52867 2835 52925 2836
rect 54507 2876 54549 2885
rect 54507 2836 54508 2876
rect 54548 2836 54549 2876
rect 54507 2827 54549 2836
rect 835 2708 893 2709
rect 835 2668 844 2708
rect 884 2668 893 2708
rect 835 2667 893 2668
rect 9675 2708 9717 2717
rect 9675 2668 9676 2708
rect 9716 2668 9717 2708
rect 9675 2659 9717 2668
rect 54691 2708 54749 2709
rect 54691 2668 54700 2708
rect 54740 2668 54749 2708
rect 54691 2667 54749 2668
rect 7651 2624 7709 2625
rect 7651 2584 7660 2624
rect 7700 2584 7709 2624
rect 7651 2583 7709 2584
rect 8515 2624 8573 2625
rect 8515 2584 8524 2624
rect 8564 2584 8573 2624
rect 8515 2583 8573 2584
rect 9859 2624 9917 2625
rect 9859 2584 9868 2624
rect 9908 2584 9917 2624
rect 9859 2583 9917 2584
rect 11683 2624 11741 2625
rect 11683 2584 11692 2624
rect 11732 2584 11741 2624
rect 11683 2583 11741 2584
rect 11971 2624 12029 2625
rect 11971 2584 11980 2624
rect 12020 2584 12029 2624
rect 11971 2583 12029 2584
rect 14091 2624 14133 2633
rect 14091 2584 14092 2624
rect 14132 2584 14133 2624
rect 14091 2575 14133 2584
rect 14467 2624 14525 2625
rect 14467 2584 14476 2624
rect 14516 2584 14525 2624
rect 14467 2583 14525 2584
rect 15331 2624 15389 2625
rect 15331 2584 15340 2624
rect 15380 2584 15389 2624
rect 15331 2583 15389 2584
rect 17827 2624 17885 2625
rect 17827 2584 17836 2624
rect 17876 2584 17885 2624
rect 17827 2583 17885 2584
rect 18691 2624 18749 2625
rect 18691 2584 18700 2624
rect 18740 2584 18749 2624
rect 18691 2583 18749 2584
rect 36747 2624 36789 2633
rect 36747 2584 36748 2624
rect 36788 2584 36789 2624
rect 36747 2575 36789 2584
rect 37123 2624 37181 2625
rect 37123 2584 37132 2624
rect 37172 2584 37181 2624
rect 37123 2583 37181 2584
rect 37987 2624 38045 2625
rect 37987 2584 37996 2624
rect 38036 2584 38045 2624
rect 37987 2583 38045 2584
rect 39339 2624 39381 2633
rect 39339 2584 39340 2624
rect 39380 2584 39381 2624
rect 39339 2575 39381 2584
rect 39715 2624 39773 2625
rect 39715 2584 39724 2624
rect 39764 2584 39773 2624
rect 39715 2583 39773 2584
rect 40579 2624 40637 2625
rect 40579 2584 40588 2624
rect 40628 2584 40637 2624
rect 40579 2583 40637 2584
rect 44043 2624 44085 2633
rect 44043 2584 44044 2624
rect 44084 2584 44085 2624
rect 44043 2575 44085 2584
rect 44419 2624 44477 2625
rect 44419 2584 44428 2624
rect 44468 2584 44477 2624
rect 44419 2583 44477 2584
rect 45283 2624 45341 2625
rect 45283 2584 45292 2624
rect 45332 2584 45341 2624
rect 45283 2583 45341 2584
rect 48259 2624 48317 2625
rect 48259 2584 48268 2624
rect 48308 2584 48317 2624
rect 48259 2583 48317 2584
rect 49123 2624 49181 2625
rect 49123 2584 49132 2624
rect 49172 2584 49181 2624
rect 49123 2583 49181 2584
rect 49515 2624 49557 2633
rect 49515 2584 49516 2624
rect 49556 2584 49557 2624
rect 49515 2575 49557 2584
rect 50475 2624 50517 2633
rect 50475 2584 50476 2624
rect 50516 2584 50517 2624
rect 50475 2575 50517 2584
rect 50851 2624 50909 2625
rect 50851 2584 50860 2624
rect 50900 2584 50909 2624
rect 50851 2583 50909 2584
rect 51715 2624 51773 2625
rect 51715 2584 51724 2624
rect 51764 2584 51773 2624
rect 51715 2583 51773 2584
rect 7275 2540 7317 2549
rect 7275 2500 7276 2540
rect 7316 2500 7317 2540
rect 7275 2491 7317 2500
rect 10539 2540 10581 2549
rect 10539 2500 10540 2540
rect 10580 2500 10581 2540
rect 10539 2491 10581 2500
rect 12163 2540 12221 2541
rect 12163 2500 12172 2540
rect 12212 2500 12221 2540
rect 12163 2499 12221 2500
rect 17451 2540 17493 2549
rect 17451 2500 17452 2540
rect 17492 2500 17493 2540
rect 17451 2491 17493 2500
rect 651 2456 693 2465
rect 651 2416 652 2456
rect 692 2416 693 2456
rect 651 2407 693 2416
rect 16483 2456 16541 2457
rect 16483 2416 16492 2456
rect 16532 2416 16541 2456
rect 16483 2415 16541 2416
rect 576 2288 99360 2312
rect 576 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 95072 2288
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95440 2248 99360 2288
rect 576 2224 99360 2248
rect 7851 2120 7893 2129
rect 7851 2080 7852 2120
rect 7892 2080 7893 2120
rect 7851 2071 7893 2080
rect 8235 2120 8277 2129
rect 8235 2080 8236 2120
rect 8276 2080 8277 2120
rect 8235 2071 8277 2080
rect 8899 2120 8957 2121
rect 8899 2080 8908 2120
rect 8948 2080 8957 2120
rect 8899 2079 8957 2080
rect 17731 2120 17789 2121
rect 17731 2080 17740 2120
rect 17780 2080 17789 2120
rect 17731 2079 17789 2080
rect 9571 1952 9629 1953
rect 9571 1912 9580 1952
rect 9620 1912 9629 1952
rect 9571 1911 9629 1912
rect 17059 1952 17117 1953
rect 17059 1912 17068 1952
rect 17108 1912 17117 1952
rect 17059 1911 17117 1912
rect 8035 1868 8093 1869
rect 8035 1828 8044 1868
rect 8084 1828 8093 1868
rect 8035 1827 8093 1828
rect 8419 1868 8477 1869
rect 8419 1828 8428 1868
rect 8468 1828 8477 1868
rect 8419 1827 8477 1828
rect 576 1532 99360 1556
rect 576 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 93832 1532
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 94200 1492 99360 1532
rect 576 1468 99360 1492
rect 576 776 99360 800
rect 576 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 95072 776
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95440 736 99360 776
rect 576 712 99360 736
<< via1 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 12748 38200 12788 38240
rect 12076 37948 12116 37988
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 13324 37612 13364 37652
rect 18124 37444 18164 37484
rect 25708 37444 25748 37484
rect 26764 37444 26804 37484
rect 39820 37444 39860 37484
rect 11308 37360 11348 37400
rect 12172 37360 12212 37400
rect 19468 37360 19508 37400
rect 22156 37360 22196 37400
rect 22540 37360 22580 37400
rect 27436 37360 27476 37400
rect 39340 37360 39380 37400
rect 40684 37360 40724 37400
rect 10924 37276 10964 37316
rect 17932 37192 17972 37232
rect 18796 37192 18836 37232
rect 22636 37192 22676 37232
rect 25516 37192 25556 37232
rect 38668 37192 38708 37232
rect 39628 37192 39668 37232
rect 40012 37192 40052 37232
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 10732 36856 10772 36896
rect 19180 36856 19220 36896
rect 27532 36856 27572 36896
rect 39532 36856 39572 36896
rect 42124 36856 42164 36896
rect 16780 36772 16820 36812
rect 21868 36772 21908 36812
rect 25132 36772 25172 36812
rect 39724 36772 39764 36812
rect 7948 36688 7988 36728
rect 10924 36688 10964 36728
rect 11308 36688 11348 36728
rect 12172 36688 12212 36728
rect 17164 36688 17204 36728
rect 18028 36688 18068 36728
rect 22252 36688 22292 36728
rect 23116 36688 23156 36728
rect 25516 36688 25556 36728
rect 26380 36688 26420 36728
rect 29644 36688 29684 36728
rect 35788 36688 35828 36728
rect 37132 36688 37172 36728
rect 37516 36688 37556 36728
rect 38380 36688 38420 36728
rect 40108 36688 40148 36728
rect 40972 36688 41012 36728
rect 10540 36604 10580 36644
rect 34348 36604 34388 36644
rect 7276 36520 7316 36560
rect 13324 36520 13364 36560
rect 34156 36520 34196 36560
rect 35116 36520 35156 36560
rect 24268 36436 24308 36476
rect 28972 36436 29012 36476
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 8140 36100 8180 36140
rect 10828 36100 10868 36140
rect 21868 36100 21908 36140
rect 26284 36100 26324 36140
rect 30220 36100 30260 36140
rect 35596 36100 35636 36140
rect 37420 36100 37460 36140
rect 11020 35932 11060 35972
rect 18220 35932 18260 35972
rect 27436 35932 27476 35972
rect 37612 35932 37652 35972
rect 6124 35848 6164 35888
rect 6988 35848 7028 35888
rect 10444 35848 10484 35888
rect 10636 35848 10676 35888
rect 11884 35848 11924 35888
rect 16204 35848 16244 35888
rect 17068 35848 17108 35888
rect 19084 35848 19124 35888
rect 21772 35848 21812 35888
rect 21964 35848 22004 35888
rect 26188 35848 26228 35888
rect 26380 35848 26420 35888
rect 28204 35848 28244 35888
rect 29068 35848 29108 35888
rect 33196 35848 33236 35888
rect 33580 35848 33620 35888
rect 34444 35848 34484 35888
rect 39628 35848 39668 35888
rect 39820 35848 39860 35888
rect 5740 35764 5780 35804
rect 10540 35764 10580 35804
rect 15820 35764 15860 35804
rect 27820 35764 27860 35804
rect 39724 35764 39764 35804
rect 11212 35680 11252 35720
rect 18412 35680 18452 35720
rect 27628 35680 27668 35720
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 5932 35344 5972 35384
rect 25804 35344 25844 35384
rect 36940 35344 36980 35384
rect 9004 35260 9044 35300
rect 39532 35260 39572 35300
rect 6316 35176 6356 35216
rect 6700 35176 6740 35216
rect 7564 35176 7604 35216
rect 8908 35176 8948 35216
rect 9100 35176 9140 35216
rect 20524 35176 20564 35216
rect 21484 35176 21524 35216
rect 25708 35176 25748 35216
rect 33196 35176 33236 35216
rect 33580 35176 33620 35216
rect 34444 35176 34484 35216
rect 35788 35176 35828 35216
rect 36844 35176 36884 35216
rect 37132 35176 37172 35216
rect 37228 35176 37268 35216
rect 37324 35176 37364 35216
rect 39052 35176 39092 35216
rect 39436 35176 39476 35216
rect 6124 35092 6164 35132
rect 17068 35092 17108 35132
rect 35596 35092 35636 35132
rect 16876 35008 16916 35048
rect 8716 34924 8756 34964
rect 21196 34924 21236 34964
rect 25516 34924 25556 34964
rect 36460 34924 36500 34964
rect 36652 34924 36692 34964
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 7180 34588 7220 34628
rect 34156 34588 34196 34628
rect 12460 34504 12500 34544
rect 7372 34420 7412 34460
rect 23308 34420 23348 34460
rect 34348 34420 34388 34460
rect 8812 34336 8852 34376
rect 9292 34336 9332 34376
rect 9676 34336 9716 34376
rect 10540 34336 10580 34376
rect 11884 34336 11924 34376
rect 12172 34336 12212 34376
rect 13132 34336 13172 34376
rect 21292 34336 21332 34376
rect 22156 34336 22196 34376
rect 24172 34336 24212 34376
rect 24460 34336 24500 34376
rect 25324 34336 25364 34376
rect 26284 34336 26324 34376
rect 20908 34252 20948 34292
rect 8140 34168 8180 34208
rect 9772 34168 9812 34208
rect 10444 34168 10484 34208
rect 10732 34168 10772 34208
rect 24652 34168 24692 34208
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 6700 33832 6740 33872
rect 19180 33832 19220 33872
rect 18412 33748 18452 33788
rect 25708 33748 25748 33788
rect 40300 33748 40340 33788
rect 7180 33664 7220 33704
rect 17068 33664 17108 33704
rect 18316 33664 18356 33704
rect 18508 33664 18548 33704
rect 18700 33664 18740 33704
rect 18988 33664 19028 33704
rect 25324 33664 25364 33704
rect 26092 33664 26132 33704
rect 26956 33664 26996 33704
rect 40684 33664 40724 33704
rect 41548 33664 41588 33704
rect 6316 33580 6356 33620
rect 15724 33580 15764 33620
rect 15532 33412 15572 33452
rect 16396 33412 16436 33452
rect 28108 33412 28148 33452
rect 42700 33412 42740 33452
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 16876 33076 16916 33116
rect 4108 32824 4148 32864
rect 14476 32824 14516 32864
rect 14860 32824 14900 32864
rect 15724 32824 15764 32864
rect 18028 32824 18068 32864
rect 18220 32824 18260 32864
rect 27244 32824 27284 32864
rect 27436 32824 27476 32864
rect 3436 32740 3476 32780
rect 18124 32740 18164 32780
rect 26572 32740 26612 32780
rect 28108 32656 28148 32696
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 4300 32320 4340 32360
rect 10060 32320 10100 32360
rect 26572 32320 26612 32360
rect 11020 32236 11060 32276
rect 28108 32236 28148 32276
rect 35500 32236 35540 32276
rect 42892 32236 42932 32276
rect 1900 32152 1940 32192
rect 2284 32152 2324 32192
rect 3148 32152 3188 32192
rect 10444 32152 10484 32192
rect 11404 32152 11444 32192
rect 12268 32152 12308 32192
rect 19852 32152 19892 32192
rect 26188 32152 26228 32192
rect 26284 32152 26324 32192
rect 28492 32152 28532 32192
rect 29356 32152 29396 32192
rect 35884 32152 35924 32192
rect 36748 32152 36788 32192
rect 38380 32152 38420 32192
rect 38476 32152 38516 32192
rect 42988 32152 43028 32192
rect 43372 32152 43412 32192
rect 48940 32152 48980 32192
rect 18220 32068 18260 32108
rect 13420 31900 13460 31940
rect 18028 31900 18068 31940
rect 19180 31900 19220 31940
rect 30508 31900 30548 31940
rect 37900 31900 37940 31940
rect 38188 31900 38228 31940
rect 48268 31900 48308 31940
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 2188 31564 2228 31604
rect 19852 31564 19892 31604
rect 23116 31564 23156 31604
rect 26284 31564 26324 31604
rect 49516 31480 49556 31520
rect 2380 31396 2420 31436
rect 41548 31396 41588 31436
rect 46732 31396 46772 31436
rect 2956 31312 2996 31352
rect 3820 31312 3860 31352
rect 9292 31312 9332 31352
rect 9676 31312 9716 31352
rect 10540 31312 10580 31352
rect 17452 31312 17492 31352
rect 17836 31312 17876 31352
rect 18700 31312 18740 31352
rect 20140 31312 20180 31352
rect 23308 31312 23348 31352
rect 25324 31312 25364 31352
rect 25996 31312 26036 31352
rect 26188 31312 26228 31352
rect 26380 31312 26420 31352
rect 33484 31312 33524 31352
rect 34348 31312 34388 31352
rect 36940 31312 36980 31352
rect 37132 31312 37172 31352
rect 37996 31312 38036 31352
rect 42412 31312 42452 31352
rect 47500 31312 47540 31352
rect 48364 31312 48404 31352
rect 50956 31312 50996 31352
rect 2572 31228 2612 31268
rect 34732 31228 34772 31268
rect 36268 31228 36308 31268
rect 47116 31228 47156 31268
rect 4972 31144 5012 31184
rect 11692 31144 11732 31184
rect 20044 31144 20084 31184
rect 20332 31144 20372 31184
rect 32332 31144 32372 31184
rect 37804 31144 37844 31184
rect 38668 31144 38708 31184
rect 41932 31144 41972 31184
rect 46924 31144 46964 31184
rect 50284 31144 50324 31184
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 3340 30808 3380 30848
rect 25996 30808 26036 30848
rect 35020 30808 35060 30848
rect 37036 30808 37076 30848
rect 42316 30808 42356 30848
rect 48940 30808 48980 30848
rect 51532 30808 51572 30848
rect 21964 30724 22004 30764
rect 26956 30724 26996 30764
rect 31084 30724 31124 30764
rect 41164 30724 41204 30764
rect 49132 30724 49172 30764
rect 4012 30640 4052 30680
rect 4204 30640 4244 30680
rect 5068 30640 5108 30680
rect 7276 30640 7316 30680
rect 7660 30640 7700 30680
rect 8524 30640 8564 30680
rect 13516 30640 13556 30680
rect 17548 30640 17588 30680
rect 17932 30640 17972 30680
rect 18796 30640 18836 30680
rect 22348 30640 22388 30680
rect 23212 30640 23252 30680
rect 25804 30640 25844 30680
rect 26668 30640 26708 30680
rect 27052 30640 27092 30680
rect 27436 30640 27476 30680
rect 30604 30640 30644 30680
rect 30988 30640 31028 30680
rect 34156 30640 34196 30680
rect 34540 30640 34580 30680
rect 36652 30640 36692 30680
rect 38188 30640 38228 30680
rect 39052 30640 39092 30680
rect 39436 30640 39476 30680
rect 42028 30640 42068 30680
rect 43468 30640 43508 30680
rect 44332 30640 44372 30680
rect 44716 30640 44756 30680
rect 46156 30640 46196 30680
rect 48364 30640 48404 30680
rect 48556 30640 48596 30680
rect 49516 30640 49556 30680
rect 50380 30640 50420 30680
rect 3532 30556 3572 30596
rect 24364 30556 24404 30596
rect 48748 30556 48788 30596
rect 4396 30472 4436 30512
rect 4108 30388 4148 30428
rect 9676 30388 9716 30428
rect 14188 30388 14228 30428
rect 19948 30388 19988 30428
rect 25132 30388 25172 30428
rect 25996 30388 26036 30428
rect 35980 30388 36020 30428
rect 48460 30388 48500 30428
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 16108 30052 16148 30092
rect 17932 30052 17972 30092
rect 19180 30052 19220 30092
rect 37996 30052 38036 30092
rect 43084 30052 43124 30092
rect 45676 30052 45716 30092
rect 46732 30052 46772 30092
rect 18124 29884 18164 29924
rect 5164 29800 5204 29840
rect 5452 29800 5492 29840
rect 11116 29800 11156 29840
rect 11500 29800 11540 29840
rect 15916 29800 15956 29840
rect 19852 29800 19892 29840
rect 25708 29800 25748 29840
rect 26092 29800 26132 29840
rect 26956 29800 26996 29840
rect 28396 29800 28436 29840
rect 37420 29800 37460 29840
rect 37708 29800 37748 29840
rect 37900 29800 37940 29840
rect 38092 29800 38132 29840
rect 42796 29800 42836 29840
rect 45868 29800 45908 29840
rect 46252 29800 46292 29840
rect 47404 29800 47444 29840
rect 47788 29800 47828 29840
rect 5644 29716 5684 29756
rect 37228 29716 37268 29756
rect 47884 29716 47924 29756
rect 11596 29632 11636 29672
rect 28108 29632 28148 29672
rect 29068 29632 29108 29672
rect 43276 29632 43316 29672
rect 45964 29632 46004 29672
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 5164 29212 5204 29252
rect 30412 29212 30452 29252
rect 34540 29212 34580 29252
rect 46924 29212 46964 29252
rect 4876 29128 4916 29168
rect 5068 29128 5108 29168
rect 5260 29128 5300 29168
rect 8812 29128 8852 29168
rect 9772 29128 9812 29168
rect 12364 29128 12404 29168
rect 12460 29128 12500 29168
rect 22156 29128 22196 29168
rect 23020 29128 23060 29168
rect 28492 29128 28532 29168
rect 28684 29128 28724 29168
rect 29164 29128 29204 29168
rect 30124 29128 30164 29168
rect 31084 29128 31124 29168
rect 33292 29128 33332 29168
rect 34156 29128 34196 29168
rect 46828 29128 46868 29168
rect 47020 29128 47060 29168
rect 32140 29044 32180 29084
rect 4204 28960 4244 29000
rect 9484 28960 9524 29000
rect 12652 28876 12692 28916
rect 28588 28876 28628 28916
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 4684 28540 4724 28580
rect 5836 28540 5876 28580
rect 13036 28540 13076 28580
rect 44908 28372 44948 28412
rect 45676 28372 45716 28412
rect 2668 28288 2708 28328
rect 3532 28288 3572 28328
rect 5164 28288 5204 28328
rect 6124 28288 6164 28328
rect 6508 28288 6548 28328
rect 12076 28288 12116 28328
rect 12748 28288 12788 28328
rect 12940 28288 12980 28328
rect 13132 28288 13172 28328
rect 25132 28288 25172 28328
rect 26092 28288 26132 28328
rect 26956 28288 26996 28328
rect 28012 28288 28052 28328
rect 28300 28288 28340 28328
rect 28780 28288 28820 28328
rect 28876 28288 28916 28328
rect 41740 28288 41780 28328
rect 42604 28288 42644 28328
rect 46348 28288 46388 28328
rect 2284 28204 2324 28244
rect 27820 28204 27860 28244
rect 6412 28120 6452 28160
rect 6700 28120 6740 28160
rect 26284 28120 26324 28160
rect 29068 28120 29108 28160
rect 44716 28120 44756 28160
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 46156 27784 46196 27824
rect 8620 27700 8660 27740
rect 14188 27700 14228 27740
rect 43756 27700 43796 27740
rect 47212 27700 47252 27740
rect 3916 27616 3956 27656
rect 4300 27616 4340 27656
rect 5164 27616 5204 27656
rect 9004 27616 9044 27656
rect 9868 27616 9908 27656
rect 13516 27616 13556 27656
rect 13708 27616 13748 27656
rect 14092 27616 14132 27656
rect 14572 27616 14612 27656
rect 22060 27616 22100 27656
rect 22924 27616 22964 27656
rect 23308 27616 23348 27656
rect 29740 27616 29780 27656
rect 42508 27616 42548 27656
rect 43372 27616 43412 27656
rect 44140 27616 44180 27656
rect 45004 27616 45044 27656
rect 47884 27616 47924 27656
rect 3436 27532 3476 27572
rect 11020 27532 11060 27572
rect 47020 27532 47060 27572
rect 3244 27448 3284 27488
rect 6316 27364 6356 27404
rect 12844 27364 12884 27404
rect 15244 27364 15284 27404
rect 20908 27364 20948 27404
rect 30412 27364 30452 27404
rect 46828 27364 46868 27404
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 4492 27028 4532 27068
rect 5644 27028 5684 27068
rect 44044 27028 44084 27068
rect 49420 27028 49460 27068
rect 4684 26860 4724 26900
rect 39532 26860 39572 26900
rect 6316 26776 6356 26816
rect 9196 26776 9236 26816
rect 10060 26776 10100 26816
rect 12748 26776 12788 26816
rect 13132 26776 13172 26816
rect 13996 26776 14036 26816
rect 15340 26776 15380 26816
rect 15724 26776 15764 26816
rect 16588 26776 16628 26816
rect 19564 26776 19604 26816
rect 20524 26776 20564 26816
rect 28972 26776 29012 26816
rect 29836 26776 29876 26816
rect 30220 26776 30260 26816
rect 32140 26776 32180 26816
rect 37516 26776 37556 26816
rect 38380 26776 38420 26816
rect 40396 26776 40436 26816
rect 44428 26776 44468 26816
rect 47020 26776 47060 26816
rect 47404 26776 47444 26816
rect 48268 26776 48308 26816
rect 37132 26692 37172 26732
rect 15148 26608 15188 26648
rect 17740 26608 17780 26648
rect 27820 26608 27860 26648
rect 31468 26608 31508 26648
rect 39724 26608 39764 26648
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 11788 26272 11828 26312
rect 30220 26272 30260 26312
rect 33292 26272 33332 26312
rect 38188 26272 38228 26312
rect 4876 26104 4916 26144
rect 11404 26104 11444 26144
rect 18988 26104 19028 26144
rect 19660 26104 19700 26144
rect 19852 26104 19892 26144
rect 20236 26104 20276 26144
rect 21100 26104 21140 26144
rect 29836 26104 29876 26144
rect 30700 26104 30740 26144
rect 30892 26104 30932 26144
rect 31276 26104 31316 26144
rect 32140 26104 32180 26144
rect 34540 26104 34580 26144
rect 34924 26104 34964 26144
rect 35788 26104 35828 26144
rect 41356 26104 41396 26144
rect 41740 26104 41780 26144
rect 42604 26104 42644 26144
rect 46636 26104 46676 26144
rect 3436 26020 3476 26060
rect 23788 26020 23828 26060
rect 38380 26020 38420 26060
rect 3244 25852 3284 25892
rect 4204 25852 4244 25892
rect 22252 25852 22292 25892
rect 23596 25852 23636 25892
rect 36940 25852 36980 25892
rect 43756 25852 43796 25892
rect 46348 25852 46388 25892
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 4780 25516 4820 25556
rect 18124 25516 18164 25556
rect 25996 25516 26036 25556
rect 31852 25516 31892 25556
rect 34348 25516 34388 25556
rect 19468 25348 19508 25388
rect 32044 25348 32084 25388
rect 39628 25348 39668 25388
rect 2380 25264 2420 25304
rect 2764 25264 2804 25304
rect 3628 25264 3668 25304
rect 16780 25264 16820 25304
rect 17068 25264 17108 25304
rect 17836 25264 17876 25304
rect 17932 25264 17972 25304
rect 18412 25264 18452 25304
rect 21868 25264 21908 25304
rect 22828 25264 22868 25304
rect 23212 25264 23252 25304
rect 23596 25264 23636 25304
rect 23980 25264 24020 25304
rect 24844 25264 24884 25304
rect 34060 25264 34100 25304
rect 35020 25264 35060 25304
rect 39532 25264 39572 25304
rect 39724 25264 39764 25304
rect 40300 25264 40340 25304
rect 40684 25264 40724 25304
rect 41260 25264 41300 25304
rect 41644 25264 41684 25304
rect 17260 25180 17300 25220
rect 41740 25180 41780 25220
rect 19084 25096 19124 25136
rect 22540 25096 22580 25136
rect 23308 25096 23348 25136
rect 40780 25096 40820 25136
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 32716 24760 32756 24800
rect 38668 24760 38708 24800
rect 31948 24676 31988 24716
rect 33100 24676 33140 24716
rect 18412 24592 18452 24632
rect 18604 24592 18644 24632
rect 31852 24592 31892 24632
rect 32044 24592 32084 24632
rect 32236 24592 32276 24632
rect 32524 24592 32564 24632
rect 33964 24592 34004 24632
rect 39340 24592 39380 24632
rect 42316 24592 42356 24632
rect 43276 24592 43316 24632
rect 37900 24508 37940 24548
rect 18508 24424 18548 24464
rect 37708 24340 37748 24380
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 18700 24004 18740 24044
rect 39244 24004 39284 24044
rect 16780 23920 16820 23960
rect 3628 23836 3668 23876
rect 42892 23836 42932 23876
rect 43180 23836 43220 23876
rect 4108 23752 4148 23792
rect 4300 23752 4340 23792
rect 5164 23752 5204 23792
rect 9484 23752 9524 23792
rect 10348 23752 10388 23792
rect 13516 23752 13556 23792
rect 14764 23752 14804 23792
rect 15628 23752 15668 23792
rect 19372 23752 19412 23792
rect 36844 23752 36884 23792
rect 37228 23752 37268 23792
rect 38092 23752 38132 23792
rect 42796 23752 42836 23792
rect 42988 23752 43028 23792
rect 43756 23752 43796 23792
rect 44428 23752 44468 23792
rect 4204 23668 4244 23708
rect 9100 23668 9140 23708
rect 14188 23668 14228 23708
rect 14380 23668 14420 23708
rect 3436 23584 3476 23624
rect 4492 23584 4532 23624
rect 11500 23584 11540 23624
rect 43372 23584 43412 23624
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 5068 23248 5108 23288
rect 6028 23248 6068 23288
rect 6316 23248 6356 23288
rect 13708 23248 13748 23288
rect 39052 23248 39092 23288
rect 42700 23248 42740 23288
rect 2668 23164 2708 23204
rect 5740 23164 5780 23204
rect 7564 23164 7604 23204
rect 19084 23164 19124 23204
rect 31756 23164 31796 23204
rect 45964 23164 46004 23204
rect 3052 23080 3092 23120
rect 3916 23080 3956 23120
rect 5260 23080 5300 23120
rect 5548 23080 5588 23120
rect 6124 23080 6164 23120
rect 7948 23080 7988 23120
rect 8812 23080 8852 23120
rect 12844 23080 12884 23120
rect 13996 23080 14036 23120
rect 14092 23080 14132 23120
rect 18604 23080 18644 23120
rect 18988 23080 19028 23120
rect 19564 23080 19604 23120
rect 21868 23080 21908 23120
rect 21964 23080 22004 23120
rect 22348 23080 22388 23120
rect 24844 23080 24884 23120
rect 25708 23080 25748 23120
rect 26188 23080 26228 23120
rect 27148 23080 27188 23120
rect 28780 23080 28820 23120
rect 29452 23080 29492 23120
rect 31660 23080 31700 23120
rect 31852 23080 31892 23120
rect 33676 23080 33716 23120
rect 34636 23080 34676 23120
rect 38956 23080 38996 23120
rect 43372 23080 43412 23120
rect 44716 23080 44756 23120
rect 45580 23080 45620 23120
rect 47884 23080 47924 23120
rect 48268 23080 48308 23120
rect 49132 23080 49172 23120
rect 29644 22996 29684 23036
rect 32524 22996 32564 23036
rect 33964 22996 34004 23036
rect 43564 22996 43604 23036
rect 9964 22828 10004 22868
rect 13516 22828 13556 22868
rect 20236 22828 20276 22868
rect 21676 22828 21716 22868
rect 23020 22828 23060 22868
rect 29836 22828 29876 22868
rect 32332 22828 32372 22868
rect 33196 22828 33236 22868
rect 38764 22828 38804 22868
rect 50284 22828 50324 22868
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 4204 22492 4244 22532
rect 4492 22492 4532 22532
rect 13996 22492 14036 22532
rect 18508 22492 18548 22532
rect 22156 22492 22196 22532
rect 23020 22492 23060 22532
rect 28204 22492 28244 22532
rect 34540 22492 34580 22532
rect 45004 22492 45044 22532
rect 652 22408 692 22448
rect 47980 22408 48020 22448
rect 3628 22324 3668 22364
rect 22444 22324 22484 22364
rect 31084 22324 31124 22364
rect 42220 22324 42260 22364
rect 4108 22240 4148 22280
rect 4300 22240 4340 22280
rect 5164 22240 5204 22280
rect 11116 22240 11156 22280
rect 11404 22240 11444 22280
rect 13900 22240 13940 22280
rect 14092 22240 14132 22280
rect 14476 22240 14516 22280
rect 14860 22240 14900 22280
rect 15244 22240 15284 22280
rect 16492 22240 16532 22280
rect 17356 22240 17396 22280
rect 19756 22240 19796 22280
rect 20140 22240 20180 22280
rect 21004 22240 21044 22280
rect 23212 22240 23252 22280
rect 29356 22240 29396 22280
rect 30220 22240 30260 22280
rect 30604 22240 30644 22280
rect 31948 22240 31988 22280
rect 32140 22240 32180 22280
rect 32524 22240 32564 22280
rect 33388 22240 33428 22280
rect 42988 22240 43028 22280
rect 43852 22240 43892 22280
rect 47308 22240 47348 22280
rect 48844 22240 48884 22280
rect 49708 22240 49748 22280
rect 11596 22156 11636 22196
rect 14956 22156 14996 22196
rect 15916 22156 15956 22196
rect 16108 22156 16148 22196
rect 42604 22156 42644 22196
rect 48460 22156 48500 22196
rect 3436 22072 3476 22112
rect 30892 22072 30932 22112
rect 31276 22072 31316 22112
rect 42412 22072 42452 22112
rect 50860 22072 50900 22112
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 5068 21736 5108 21776
rect 15244 21736 15284 21776
rect 32716 21736 32756 21776
rect 33772 21736 33812 21776
rect 48076 21736 48116 21776
rect 49036 21736 49076 21776
rect 2668 21652 2708 21692
rect 21964 21652 22004 21692
rect 22732 21652 22772 21692
rect 30316 21652 30356 21692
rect 37420 21652 37460 21692
rect 3052 21568 3092 21608
rect 3916 21568 3956 21608
rect 15916 21568 15956 21608
rect 21676 21568 21716 21608
rect 22060 21568 22100 21608
rect 22444 21568 22484 21608
rect 22636 21568 22676 21608
rect 22828 21568 22868 21608
rect 30700 21568 30740 21608
rect 31564 21568 31604 21608
rect 33868 21568 33908 21608
rect 37804 21568 37844 21608
rect 38668 21568 38708 21608
rect 50092 21568 50132 21608
rect 50956 21568 50996 21608
rect 48268 21484 48308 21524
rect 49228 21484 49268 21524
rect 50284 21484 50324 21524
rect 21004 21400 21044 21440
rect 39820 21400 39860 21440
rect 49420 21400 49460 21440
rect 34060 21316 34100 21356
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 10156 20980 10196 21020
rect 652 20896 692 20936
rect 26092 20812 26132 20852
rect 26860 20812 26900 20852
rect 9868 20728 9908 20768
rect 14572 20728 14612 20768
rect 27532 20728 27572 20768
rect 38956 20728 38996 20768
rect 39628 20728 39668 20768
rect 40492 20728 40532 20768
rect 14188 20560 14228 20600
rect 25900 20560 25940 20600
rect 39820 20560 39860 20600
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 27340 20224 27380 20264
rect 24940 20140 24980 20180
rect 49804 20140 49844 20180
rect 8716 20056 8756 20096
rect 9100 20056 9140 20096
rect 9964 20056 10004 20096
rect 13036 20056 13076 20096
rect 13420 20056 13460 20096
rect 14284 20056 14324 20096
rect 21100 20056 21140 20096
rect 25324 20056 25364 20096
rect 26188 20056 26228 20096
rect 29164 20056 29204 20096
rect 30124 20056 30164 20096
rect 30508 20056 30548 20096
rect 31468 20056 31508 20096
rect 36076 20056 36116 20096
rect 36460 20056 36500 20096
rect 37324 20056 37364 20096
rect 39724 20056 39764 20096
rect 39820 20056 39860 20096
rect 39916 20056 39956 20096
rect 40588 20056 40628 20096
rect 40684 20056 40724 20096
rect 41740 20056 41780 20096
rect 48172 20056 48212 20096
rect 48844 20056 48884 20096
rect 49324 20056 49364 20096
rect 49516 20056 49556 20096
rect 49708 20056 49748 20096
rect 49900 20056 49940 20096
rect 11116 19972 11156 20012
rect 15436 19972 15476 20012
rect 40876 19972 40916 20012
rect 652 19888 692 19928
rect 20428 19804 20468 19844
rect 29836 19804 29876 19844
rect 30796 19804 30836 19844
rect 38476 19804 38516 19844
rect 41068 19804 41108 19844
rect 49420 19804 49460 19844
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 3628 19468 3668 19508
rect 48748 19468 48788 19508
rect 652 19384 692 19424
rect 2860 19300 2900 19340
rect 4300 19216 4340 19256
rect 26572 19216 26612 19256
rect 26764 19216 26804 19256
rect 27628 19216 27668 19256
rect 34924 19216 34964 19256
rect 39340 19216 39380 19256
rect 39724 19216 39764 19256
rect 46732 19216 46772 19256
rect 47596 19216 47636 19256
rect 50188 19216 50228 19256
rect 50476 19216 50516 19256
rect 26668 19132 26708 19172
rect 46348 19132 46388 19172
rect 2668 19048 2708 19088
rect 26956 19048 26996 19088
rect 35404 19048 35444 19088
rect 39820 19048 39860 19088
rect 50668 19048 50708 19088
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 4108 18712 4148 18752
rect 7468 18712 7508 18752
rect 8716 18712 8756 18752
rect 11788 18712 11828 18752
rect 12076 18712 12116 18752
rect 12268 18712 12308 18752
rect 27532 18712 27572 18752
rect 1708 18628 1748 18668
rect 19756 18628 19796 18668
rect 41068 18628 41108 18668
rect 52012 18628 52052 18668
rect 2092 18544 2132 18584
rect 2956 18544 2996 18584
rect 6988 18544 7028 18584
rect 7948 18544 7988 18584
rect 8236 18544 8276 18584
rect 8620 18544 8660 18584
rect 11884 18544 11924 18584
rect 12940 18544 12980 18584
rect 18508 18544 18548 18584
rect 19372 18544 19412 18584
rect 23500 18544 23540 18584
rect 25132 18544 25172 18584
rect 25516 18544 25556 18584
rect 26380 18544 26420 18584
rect 40684 18544 40724 18584
rect 41452 18544 41492 18584
rect 42316 18544 42356 18584
rect 46732 18544 46772 18584
rect 47116 18544 47156 18584
rect 47980 18544 48020 18584
rect 52396 18544 52436 18584
rect 53260 18544 53300 18584
rect 6796 18460 6836 18500
rect 652 18376 692 18416
rect 6604 18292 6644 18332
rect 17356 18292 17396 18332
rect 22828 18292 22868 18332
rect 40012 18292 40052 18332
rect 43468 18292 43508 18332
rect 49132 18292 49172 18332
rect 54412 18292 54452 18332
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 7660 17956 7700 17996
rect 13324 17956 13364 17996
rect 23404 17956 23444 17996
rect 25900 17956 25940 17996
rect 47212 17956 47252 17996
rect 47596 17956 47636 17996
rect 48556 17956 48596 17996
rect 652 17872 692 17912
rect 24652 17872 24692 17912
rect 6508 17788 6548 17828
rect 23980 17788 24020 17828
rect 26092 17788 26132 17828
rect 32332 17788 32372 17828
rect 47404 17788 47444 17828
rect 47788 17788 47828 17828
rect 4492 17704 4532 17744
rect 5356 17704 5396 17744
rect 6700 17704 6740 17744
rect 8332 17704 8372 17744
rect 8812 17704 8852 17744
rect 9004 17704 9044 17744
rect 11308 17704 11348 17744
rect 12172 17704 12212 17744
rect 18988 17704 19028 17744
rect 21388 17704 21428 17744
rect 22252 17704 22292 17744
rect 25324 17704 25364 17744
rect 26476 17704 26516 17744
rect 26572 17704 26612 17744
rect 26679 17719 26719 17759
rect 27151 17704 27191 17744
rect 27532 17704 27572 17744
rect 27820 17704 27860 17744
rect 30316 17704 30356 17744
rect 31180 17704 31220 17744
rect 41452 17704 41492 17744
rect 41836 17704 41876 17744
rect 48172 17704 48212 17744
rect 49228 17704 49268 17744
rect 4108 17620 4148 17660
rect 7372 17620 7412 17660
rect 8908 17620 8948 17660
rect 10924 17620 10964 17660
rect 21004 17620 21044 17660
rect 28012 17620 28052 17660
rect 29932 17620 29972 17660
rect 41932 17620 41972 17660
rect 23788 17536 23828 17576
rect 27052 17536 27092 17576
rect 27340 17536 27380 17576
rect 48076 17536 48116 17576
rect 48364 17536 48404 17576
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 5260 17200 5300 17240
rect 8044 17200 8084 17240
rect 10540 17200 10580 17240
rect 21772 17200 21812 17240
rect 25132 17200 25172 17240
rect 39628 17200 39668 17240
rect 54988 17200 55028 17240
rect 5644 17116 5684 17156
rect 8332 17116 8372 17156
rect 10732 17116 10772 17156
rect 18892 17116 18932 17156
rect 22732 17116 22772 17156
rect 30988 17116 31028 17156
rect 34060 17116 34100 17156
rect 40012 17116 40052 17156
rect 6028 17032 6068 17072
rect 6892 17032 6932 17072
rect 8236 17032 8276 17072
rect 8428 17032 8468 17072
rect 11116 17032 11156 17072
rect 11980 17032 12020 17072
rect 17644 17032 17684 17072
rect 18508 17032 18548 17072
rect 19180 17032 19220 17072
rect 23116 17032 23156 17072
rect 23980 17032 24020 17072
rect 31372 17032 31412 17072
rect 32236 17032 32276 17072
rect 33580 17032 33620 17072
rect 33868 17032 33908 17072
rect 36364 17032 36404 17072
rect 37036 17032 37076 17072
rect 37228 17032 37268 17072
rect 37612 17032 37652 17072
rect 38476 17032 38516 17072
rect 40396 17032 40436 17072
rect 41260 17032 41300 17072
rect 54508 17032 54548 17072
rect 54892 17032 54932 17072
rect 56428 17032 56468 17072
rect 57292 17032 57332 17072
rect 57676 17032 57716 17072
rect 5452 16948 5492 16988
rect 10348 16948 10388 16988
rect 21964 16948 22004 16988
rect 55276 16948 55316 16988
rect 652 16864 692 16904
rect 19468 16864 19508 16904
rect 13132 16780 13172 16820
rect 16492 16780 16532 16820
rect 33388 16780 33428 16820
rect 42412 16780 42452 16820
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 652 16360 692 16400
rect 10828 16360 10868 16400
rect 11692 16360 11732 16400
rect 12940 16360 12980 16400
rect 11020 16276 11060 16316
rect 36364 16276 36404 16316
rect 12364 16192 12404 16232
rect 12652 16192 12692 16232
rect 34924 16192 34964 16232
rect 36076 16192 36116 16232
rect 36172 16192 36212 16232
rect 13516 16108 13556 16148
rect 35596 16024 35636 16064
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 652 15688 692 15728
rect 33004 15688 33044 15728
rect 35788 15604 35828 15644
rect 49228 15604 49268 15644
rect 30604 15520 30644 15560
rect 30988 15520 31028 15560
rect 31852 15520 31892 15560
rect 35692 15520 35732 15560
rect 35884 15520 35924 15560
rect 36076 15520 36116 15560
rect 36748 15520 36788 15560
rect 41548 15520 41588 15560
rect 41740 15520 41780 15560
rect 42604 15520 42644 15560
rect 49612 15520 49652 15560
rect 50476 15520 50516 15560
rect 52780 15520 52820 15560
rect 51628 15436 51668 15476
rect 40876 15268 40916 15308
rect 52108 15268 52148 15308
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 9484 14932 9524 14972
rect 21868 14932 21908 14972
rect 47116 14932 47156 14972
rect 23116 14848 23156 14888
rect 23500 14848 23540 14888
rect 52588 14764 52628 14804
rect 57004 14764 57044 14804
rect 9772 14680 9812 14720
rect 16492 14680 16532 14720
rect 21676 14680 21716 14720
rect 22924 14680 22964 14720
rect 35980 14680 36020 14720
rect 36268 14680 36308 14720
rect 40780 14680 40820 14720
rect 40876 14680 40916 14720
rect 40972 14680 41012 14720
rect 41452 14680 41492 14720
rect 41548 14680 41588 14720
rect 45100 14680 45140 14720
rect 46060 14680 46100 14720
rect 46636 14680 46676 14720
rect 47596 14680 47636 14720
rect 51244 14680 51284 14720
rect 51436 14680 51476 14720
rect 52300 14680 52340 14720
rect 52780 14680 52820 14720
rect 52876 14680 52916 14720
rect 58636 14680 58676 14720
rect 51340 14596 51380 14636
rect 652 14512 692 14552
rect 17164 14512 17204 14552
rect 36460 14512 36500 14552
rect 41260 14512 41300 14552
rect 51628 14512 51668 14552
rect 56812 14512 56852 14552
rect 57964 14512 58004 14552
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 36076 14176 36116 14216
rect 40972 14176 41012 14216
rect 52684 14176 52724 14216
rect 55948 14176 55988 14216
rect 58732 14176 58772 14216
rect 50380 14092 50420 14132
rect 52972 14092 53012 14132
rect 56332 14092 56372 14132
rect 4204 14008 4244 14048
rect 12172 14008 12212 14048
rect 13132 14008 13172 14048
rect 13996 14008 14036 14048
rect 15148 14008 15188 14048
rect 15820 14008 15860 14048
rect 16012 14008 16052 14048
rect 16396 14008 16436 14048
rect 17260 14008 17300 14048
rect 18604 14008 18644 14048
rect 18796 14008 18836 14048
rect 18988 14008 19028 14048
rect 19660 14008 19700 14048
rect 26572 14008 26612 14048
rect 33676 14008 33716 14048
rect 34060 14008 34100 14048
rect 34924 14008 34964 14048
rect 36940 14008 36980 14048
rect 38956 14008 38996 14048
rect 39916 14008 39956 14048
rect 40300 14008 40340 14048
rect 42124 14008 42164 14048
rect 49132 14008 49172 14048
rect 49996 14008 50036 14048
rect 51244 14008 51284 14048
rect 52012 14008 52052 14048
rect 53068 14008 53108 14048
rect 53452 14008 53492 14048
rect 54604 14008 54644 14048
rect 55468 14008 55508 14048
rect 55852 14008 55892 14048
rect 56716 14008 56756 14048
rect 57580 14008 57620 14048
rect 18412 13924 18452 13964
rect 25324 13924 25364 13964
rect 12844 13840 12884 13880
rect 25132 13840 25172 13880
rect 25900 13840 25940 13880
rect 47980 13840 48020 13880
rect 3532 13756 3572 13796
rect 18796 13756 18836 13796
rect 37612 13756 37652 13796
rect 39244 13756 39284 13796
rect 41452 13756 41492 13796
rect 50572 13756 50612 13796
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 4492 13420 4532 13460
rect 14668 13420 14708 13460
rect 26284 13420 26324 13460
rect 32524 13420 32564 13460
rect 39628 13420 39668 13460
rect 49996 13420 50036 13460
rect 51820 13420 51860 13460
rect 54892 13420 54932 13460
rect 23308 13336 23348 13376
rect 28588 13252 28628 13292
rect 2476 13168 2516 13208
rect 3340 13168 3380 13208
rect 8044 13168 8084 13208
rect 9196 13168 9236 13208
rect 11692 13168 11732 13208
rect 12268 13168 12308 13208
rect 12652 13168 12692 13208
rect 13516 13168 13556 13208
rect 18700 13168 18740 13208
rect 19084 13168 19124 13208
rect 19372 13168 19412 13208
rect 20236 13168 20276 13208
rect 20332 13168 20372 13208
rect 20428 13168 20468 13208
rect 23500 13168 23540 13208
rect 23884 13168 23924 13208
rect 24268 13168 24308 13208
rect 25132 13168 25172 13208
rect 28876 13168 28916 13208
rect 28972 13168 29012 13208
rect 29068 13168 29108 13208
rect 30124 13168 30164 13208
rect 30508 13168 30548 13208
rect 30892 13168 30932 13208
rect 32332 13168 32372 13208
rect 37228 13168 37268 13208
rect 37612 13168 37652 13208
rect 38476 13168 38516 13208
rect 39820 13168 39860 13208
rect 40204 13168 40244 13208
rect 41452 13168 41492 13208
rect 41836 13168 41876 13208
rect 42700 13168 42740 13208
rect 47116 13168 47156 13208
rect 47980 13168 48020 13208
rect 48364 13168 48404 13208
rect 49324 13168 49364 13208
rect 50284 13168 50324 13208
rect 52972 13168 53012 13208
rect 53836 13168 53876 13208
rect 54604 13168 54644 13208
rect 56620 13168 56660 13208
rect 57484 13168 57524 13208
rect 2092 13084 2132 13124
rect 7180 13084 7220 13124
rect 30412 13084 30452 13124
rect 54220 13084 54260 13124
rect 56236 13084 56276 13124
rect 652 13000 692 13040
rect 9868 13000 9908 13040
rect 11212 13000 11252 13040
rect 18604 13000 18644 13040
rect 20044 13000 20084 13040
rect 28396 13000 28436 13040
rect 29452 13000 29492 13040
rect 32236 13000 32276 13040
rect 40300 13000 40340 13040
rect 43852 13000 43892 13040
rect 45964 13000 46004 13040
rect 55084 13000 55124 13040
rect 58636 13000 58676 13040
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 652 12664 692 12704
rect 2188 12664 2228 12704
rect 30028 12664 30068 12704
rect 54892 12664 54932 12704
rect 55180 12664 55220 12704
rect 56236 12664 56276 12704
rect 9484 12580 9524 12620
rect 27628 12580 27668 12620
rect 32620 12580 32660 12620
rect 56716 12580 56756 12620
rect 57676 12580 57716 12620
rect 2572 12496 2612 12536
rect 2956 12496 2996 12536
rect 3820 12496 3860 12536
rect 6220 12496 6260 12536
rect 6604 12496 6644 12536
rect 7468 12496 7508 12536
rect 9868 12496 9908 12536
rect 10732 12496 10772 12536
rect 18508 12496 18548 12536
rect 18604 12496 18644 12536
rect 19660 12496 19700 12536
rect 19852 12496 19892 12536
rect 19948 12496 19988 12536
rect 20044 12496 20084 12536
rect 20140 12496 20180 12536
rect 21292 12496 21332 12536
rect 28012 12496 28052 12536
rect 28876 12496 28916 12536
rect 33484 12496 33524 12536
rect 34444 12496 34484 12536
rect 55084 12496 55124 12536
rect 56620 12496 56660 12536
rect 56812 12496 56852 12536
rect 58348 12496 58388 12536
rect 2380 12412 2420 12452
rect 8620 12412 8660 12452
rect 11884 12412 11924 12452
rect 18796 12412 18836 12452
rect 32236 12412 32276 12452
rect 33772 12412 33812 12452
rect 56428 12412 56468 12452
rect 4972 12244 5012 12284
rect 18988 12244 19028 12284
rect 21964 12244 22004 12284
rect 32044 12244 32084 12284
rect 32812 12244 32852 12284
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 3244 11908 3284 11948
rect 17260 11908 17300 11948
rect 19180 11908 19220 11948
rect 31276 11908 31316 11948
rect 33964 11908 34004 11948
rect 3436 11740 3476 11780
rect 3916 11656 3956 11696
rect 4012 11656 4052 11696
rect 4108 11656 4148 11696
rect 4972 11656 5012 11696
rect 5164 11656 5204 11696
rect 5452 11656 5492 11696
rect 16684 11656 16724 11696
rect 17164 11656 17204 11696
rect 17356 11656 17396 11696
rect 18892 11656 18932 11696
rect 31180 11656 31220 11696
rect 31372 11656 31412 11696
rect 31564 11656 31604 11696
rect 31948 11656 31988 11696
rect 32812 11656 32852 11696
rect 40684 11656 40724 11696
rect 46828 11656 46868 11696
rect 5644 11572 5684 11612
rect 652 11488 692 11528
rect 4300 11488 4340 11528
rect 16012 11488 16052 11528
rect 19372 11488 19412 11528
rect 41356 11488 41396 11528
rect 47500 11488 47540 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 652 11152 692 11192
rect 16588 11152 16628 11192
rect 32812 11152 32852 11192
rect 54700 11152 54740 11192
rect 23020 11068 23060 11108
rect 36172 11068 36212 11108
rect 43660 11068 43700 11108
rect 55852 11068 55892 11108
rect 15916 10984 15956 11024
rect 23404 10984 23444 11024
rect 24268 10984 24308 11024
rect 33484 10984 33524 11024
rect 37036 10984 37076 11024
rect 39916 10984 39956 11024
rect 43852 10984 43892 11024
rect 44140 10984 44180 11024
rect 45004 10984 45044 11024
rect 55372 10984 55412 11024
rect 55756 10984 55796 11024
rect 55948 10984 55988 11024
rect 31852 10900 31892 10940
rect 54028 10900 54068 10940
rect 25420 10732 25460 10772
rect 31660 10732 31700 10772
rect 40588 10732 40628 10772
rect 44332 10732 44372 10772
rect 53836 10732 53876 10772
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 3628 10396 3668 10436
rect 33484 10396 33524 10436
rect 38380 10396 38420 10436
rect 44140 10396 44180 10436
rect 52300 10396 52340 10436
rect 55180 10396 55220 10436
rect 55564 10312 55604 10352
rect 25420 10228 25460 10268
rect 47020 10228 47060 10268
rect 48172 10228 48212 10268
rect 55756 10228 55796 10268
rect 56620 10228 56660 10268
rect 4204 10144 4244 10184
rect 12940 10144 12980 10184
rect 16012 10144 16052 10184
rect 16300 10144 16340 10184
rect 18988 10144 19028 10184
rect 19372 10144 19412 10184
rect 20236 10144 20276 10184
rect 25612 10144 25652 10184
rect 25708 10144 25748 10184
rect 31084 10144 31124 10184
rect 31468 10144 31508 10184
rect 32332 10144 32372 10184
rect 39532 10144 39572 10184
rect 40396 10144 40436 10184
rect 40780 10144 40820 10184
rect 45292 10144 45332 10184
rect 46156 10144 46196 10184
rect 46924 10144 46964 10184
rect 47116 10144 47156 10184
rect 47980 10144 48020 10184
rect 48460 10144 48500 10184
rect 48556 10144 48596 10184
rect 49900 10144 49940 10184
rect 50284 10144 50324 10184
rect 51724 10144 51764 10184
rect 52780 10144 52820 10184
rect 53164 10144 53204 10184
rect 54028 10144 54068 10184
rect 57292 10144 57332 10184
rect 16492 10060 16532 10100
rect 46540 10060 46580 10100
rect 47308 10060 47348 10100
rect 49804 10060 49844 10100
rect 652 9976 692 10016
rect 12268 9976 12308 10016
rect 21388 9976 21428 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 652 9640 692 9680
rect 4396 9640 4436 9680
rect 5260 9640 5300 9680
rect 14284 9640 14324 9680
rect 26476 9640 26516 9680
rect 47212 9640 47252 9680
rect 47884 9640 47924 9680
rect 51820 9640 51860 9680
rect 57292 9640 57332 9680
rect 3244 9556 3284 9596
rect 11884 9556 11924 9596
rect 15916 9556 15956 9596
rect 41164 9556 41204 9596
rect 54892 9556 54932 9596
rect 3148 9472 3188 9512
rect 3340 9472 3380 9512
rect 3532 9472 3572 9512
rect 4204 9472 4244 9512
rect 5068 9472 5108 9512
rect 5356 9472 5396 9512
rect 8044 9472 8084 9512
rect 10636 9472 10676 9512
rect 12268 9472 12308 9512
rect 13132 9472 13172 9512
rect 16300 9472 16340 9512
rect 17164 9472 17204 9512
rect 19660 9472 19700 9512
rect 2956 9388 2996 9428
rect 25804 9430 25844 9470
rect 25900 9467 25940 9507
rect 25996 9472 26036 9512
rect 26380 9472 26420 9512
rect 26860 9472 26900 9512
rect 39916 9472 39956 9512
rect 40780 9472 40820 9512
rect 41356 9472 41396 9512
rect 41548 9472 41588 9512
rect 47308 9472 47348 9512
rect 47692 9472 47732 9512
rect 48556 9472 48596 9512
rect 52300 9472 52340 9512
rect 52876 9472 52916 9512
rect 53068 9472 53108 9512
rect 55276 9472 55316 9512
rect 56140 9472 56180 9512
rect 18892 9388 18932 9428
rect 26188 9304 26228 9344
rect 26860 9304 26900 9344
rect 2764 9220 2804 9260
rect 5548 9220 5588 9260
rect 7372 9220 7412 9260
rect 9964 9220 10004 9260
rect 18316 9220 18356 9260
rect 25516 9220 25556 9260
rect 26668 9220 26708 9260
rect 38764 9220 38804 9260
rect 41452 9220 41492 9260
rect 51820 9220 51860 9260
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 4396 8884 4436 8924
rect 47884 8884 47924 8924
rect 7180 8800 7220 8840
rect 9772 8800 9812 8840
rect 12364 8800 12404 8840
rect 19180 8800 19220 8840
rect 30028 8800 30068 8840
rect 40204 8800 40244 8840
rect 40588 8716 40628 8756
rect 2380 8632 2420 8672
rect 3244 8632 3284 8672
rect 4780 8632 4820 8672
rect 5164 8632 5204 8672
rect 6028 8632 6068 8672
rect 7372 8632 7412 8672
rect 7756 8632 7796 8672
rect 8620 8632 8660 8672
rect 9964 8632 10004 8672
rect 10348 8632 10388 8672
rect 11212 8632 11252 8672
rect 19372 8632 19412 8672
rect 19756 8632 19796 8672
rect 19948 8632 19988 8672
rect 20908 8632 20948 8672
rect 21100 8632 21140 8672
rect 21580 8632 21620 8672
rect 21676 8632 21716 8672
rect 22060 8632 22100 8672
rect 22252 8632 22292 8672
rect 25996 8632 26036 8672
rect 26092 8632 26132 8672
rect 29356 8632 29396 8672
rect 30028 8632 30068 8672
rect 30220 8632 30260 8672
rect 39052 8632 39092 8672
rect 39532 8632 39572 8672
rect 40780 8632 40820 8672
rect 40876 8632 40916 8672
rect 45868 8632 45908 8672
rect 46732 8632 46772 8672
rect 1996 8548 2036 8588
rect 19852 8548 19892 8588
rect 22156 8548 22196 8588
rect 45484 8548 45524 8588
rect 652 8464 692 8504
rect 21004 8464 21044 8504
rect 21292 8464 21332 8504
rect 25804 8464 25844 8504
rect 28684 8464 28724 8504
rect 38380 8464 38420 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 652 8128 692 8168
rect 2284 8128 2324 8168
rect 5068 8128 5108 8168
rect 9100 8128 9140 8168
rect 21868 8128 21908 8168
rect 23212 8128 23252 8168
rect 24940 8128 24980 8168
rect 29548 8128 29588 8168
rect 45580 8128 45620 8168
rect 2668 8044 2708 8084
rect 18700 8044 18740 8084
rect 27340 8044 27380 8084
rect 39916 8044 39956 8084
rect 3052 7960 3092 8000
rect 3916 7960 3956 8000
rect 8716 7960 8756 8000
rect 18796 7960 18836 8000
rect 19180 7960 19220 8000
rect 22060 7960 22100 8000
rect 22348 7960 22388 8000
rect 22924 7960 22964 8000
rect 23020 7960 23060 8000
rect 23116 7960 23156 8000
rect 26092 7960 26132 8000
rect 26956 7960 26996 8000
rect 29644 7960 29684 8000
rect 29740 7960 29780 8000
rect 29836 7960 29876 8000
rect 30316 7960 30356 8000
rect 30988 7960 31028 8000
rect 32908 7960 32948 8000
rect 33484 7960 33524 8000
rect 34732 7960 34772 8000
rect 35596 7960 35636 8000
rect 35980 7960 36020 8000
rect 37228 7960 37268 8000
rect 37900 7960 37940 8000
rect 38764 7960 38804 8000
rect 40108 7960 40148 8000
rect 40396 7960 40436 8000
rect 46252 7960 46292 8000
rect 50956 7960 50996 8000
rect 2476 7876 2516 7916
rect 38092 7792 38132 7832
rect 32236 7708 32276 7748
rect 36556 7708 36596 7748
rect 51148 7708 51188 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 18604 7372 18644 7412
rect 20332 7372 20372 7412
rect 30700 7372 30740 7412
rect 50764 7372 50804 7412
rect 29068 7204 29108 7244
rect 10924 7120 10964 7160
rect 11788 7120 11828 7160
rect 16204 7120 16244 7160
rect 16588 7120 16628 7160
rect 17452 7120 17492 7160
rect 21484 7120 21524 7160
rect 22348 7120 22388 7160
rect 22924 7120 22964 7160
rect 23596 7120 23636 7160
rect 26668 7120 26708 7160
rect 28588 7120 28628 7160
rect 28876 7120 28916 7160
rect 29356 7120 29396 7160
rect 29452 7120 29492 7160
rect 30028 7120 30068 7160
rect 30412 7120 30452 7160
rect 30604 7120 30644 7160
rect 30796 7120 30836 7160
rect 32332 7120 32372 7160
rect 34636 7120 34676 7160
rect 35500 7120 35540 7160
rect 38668 7120 38708 7160
rect 40204 7120 40244 7160
rect 48748 7120 48788 7160
rect 49612 7120 49652 7160
rect 22732 7036 22772 7076
rect 25996 7036 26036 7076
rect 35884 7036 35924 7076
rect 37996 7036 38036 7076
rect 48364 7036 48404 7076
rect 652 6952 692 6992
rect 28396 6952 28436 6992
rect 29932 6952 29972 6992
rect 31660 6952 31700 6992
rect 33484 6952 33524 6992
rect 39532 6952 39572 6992
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 29452 6616 29492 6656
rect 39820 6616 39860 6656
rect 45292 6616 45332 6656
rect 48652 6616 48692 6656
rect 29740 6532 29780 6572
rect 21580 6448 21620 6488
rect 22540 6448 22580 6488
rect 28780 6448 28820 6488
rect 29644 6448 29684 6488
rect 29836 6448 29876 6488
rect 39340 6448 39380 6488
rect 44812 6448 44852 6488
rect 45196 6448 45236 6488
rect 45580 6448 45620 6488
rect 46252 6448 46292 6488
rect 47980 6448 48020 6488
rect 53740 6448 53780 6488
rect 54028 6448 54068 6488
rect 38764 6364 38804 6404
rect 21868 6280 21908 6320
rect 38572 6280 38612 6320
rect 39628 6280 39668 6320
rect 53068 6280 53108 6320
rect 54316 6280 54356 6320
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 40108 5860 40148 5900
rect 47404 5860 47444 5900
rect 48364 5860 48404 5900
rect 54988 5860 55028 5900
rect 52204 5692 52244 5732
rect 13036 5608 13076 5648
rect 15148 5608 15188 5648
rect 16108 5608 16148 5648
rect 18124 5608 18164 5648
rect 33868 5608 33908 5648
rect 37708 5608 37748 5648
rect 38092 5608 38132 5648
rect 38956 5608 38996 5648
rect 45292 5608 45332 5648
rect 46444 5608 46484 5648
rect 46540 5608 46580 5648
rect 46636 5608 46676 5648
rect 47212 5608 47252 5648
rect 47308 5608 47348 5648
rect 48652 5608 48692 5648
rect 52972 5608 53012 5648
rect 53836 5608 53876 5648
rect 56620 5608 56660 5648
rect 17260 5524 17300 5564
rect 45964 5524 46004 5564
rect 52588 5524 52628 5564
rect 652 5440 692 5480
rect 12364 5440 12404 5480
rect 15628 5440 15668 5480
rect 33388 5440 33428 5480
rect 48172 5440 48212 5480
rect 52396 5440 52436 5480
rect 55948 5440 55988 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 43660 5104 43700 5144
rect 52204 5104 52244 5144
rect 47692 5020 47732 5060
rect 51916 5020 51956 5060
rect 11500 4936 11540 4976
rect 11884 4936 11924 4976
rect 12748 4936 12788 4976
rect 25612 4936 25652 4976
rect 26284 4936 26324 4976
rect 26476 4936 26516 4976
rect 26860 4936 26900 4976
rect 27724 4936 27764 4976
rect 41260 4936 41300 4976
rect 41644 4936 41684 4976
rect 42508 4936 42548 4976
rect 46444 4936 46484 4976
rect 47308 4936 47348 4976
rect 52108 4936 52148 4976
rect 54796 4936 54836 4976
rect 55180 4936 55220 4976
rect 56044 4936 56084 4976
rect 844 4852 884 4892
rect 28876 4852 28916 4892
rect 39244 4852 39284 4892
rect 45292 4852 45332 4892
rect 54412 4852 54452 4892
rect 57196 4852 57236 4892
rect 652 4768 692 4808
rect 54604 4768 54644 4808
rect 13900 4684 13940 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 13612 4348 13652 4388
rect 30316 4348 30356 4388
rect 40684 4348 40724 4388
rect 844 4180 884 4220
rect 10828 4180 10868 4220
rect 23788 4180 23828 4220
rect 34444 4180 34484 4220
rect 38956 4180 38996 4220
rect 11596 4096 11636 4136
rect 12460 4096 12500 4136
rect 20524 4096 20564 4136
rect 21772 4096 21812 4136
rect 22636 4096 22676 4136
rect 24364 4096 24404 4136
rect 27052 4096 27092 4136
rect 28300 4096 28340 4136
rect 29164 4096 29204 4136
rect 38284 4096 38324 4136
rect 40012 4096 40052 4136
rect 40108 4096 40148 4136
rect 40204 4096 40244 4136
rect 40492 4096 40532 4136
rect 41068 4096 41108 4136
rect 41356 4096 41396 4136
rect 54028 4096 54068 4136
rect 54220 4096 54260 4136
rect 56524 4096 56564 4136
rect 11212 4012 11252 4052
rect 21196 4012 21236 4052
rect 21388 4012 21428 4052
rect 27916 4012 27956 4052
rect 54124 4012 54164 4052
rect 652 3928 692 3968
rect 11020 3928 11060 3968
rect 25036 3928 25076 3968
rect 27724 3928 27764 3968
rect 34252 3928 34292 3968
rect 40396 3928 40436 3968
rect 41548 3928 41588 3968
rect 55852 3928 55892 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 11788 3592 11828 3632
rect 12556 3592 12596 3632
rect 20044 3592 20084 3632
rect 24556 3592 24596 3632
rect 27148 3592 27188 3632
rect 35788 3592 35828 3632
rect 47596 3592 47636 3632
rect 52300 3592 52340 3632
rect 53644 3592 53684 3632
rect 56812 3592 56852 3632
rect 13036 3508 13076 3548
rect 24748 3508 24788 3548
rect 33388 3508 33428 3548
rect 40300 3508 40340 3548
rect 52012 3508 52052 3548
rect 7084 3424 7124 3464
rect 7468 3424 7508 3464
rect 8332 3424 8372 3464
rect 10924 3424 10964 3464
rect 11116 3424 11156 3464
rect 11308 3424 11348 3464
rect 11500 3424 11540 3464
rect 12652 3424 12692 3464
rect 13708 3424 13748 3464
rect 17644 3424 17684 3464
rect 18028 3424 18068 3464
rect 18892 3424 18932 3464
rect 21100 3424 21140 3464
rect 21772 3424 21812 3464
rect 22156 3424 22196 3464
rect 22540 3424 22580 3464
rect 23404 3424 23444 3464
rect 25132 3424 25172 3464
rect 25996 3424 26036 3464
rect 33772 3424 33812 3464
rect 34636 3424 34676 3464
rect 38860 3424 38900 3464
rect 40204 3424 40244 3464
rect 40396 3424 40436 3464
rect 40972 3424 41012 3464
rect 41644 3424 41684 3464
rect 47692 3424 47732 3464
rect 48076 3424 48116 3464
rect 51916 3424 51956 3464
rect 52108 3424 52148 3464
rect 52972 3424 53012 3464
rect 53164 3424 53204 3464
rect 53548 3424 53588 3464
rect 54412 3424 54452 3464
rect 54796 3424 54836 3464
rect 55660 3424 55700 3464
rect 844 3340 884 3380
rect 11980 3340 12020 3380
rect 38380 3340 38420 3380
rect 39532 3340 39572 3380
rect 40012 3340 40052 3380
rect 51436 3340 51476 3380
rect 652 3172 692 3212
rect 9484 3172 9524 3212
rect 11020 3172 11060 3212
rect 11404 3172 11444 3212
rect 12844 3172 12884 3212
rect 38188 3172 38228 3212
rect 39820 3172 39860 3212
rect 51244 3172 51284 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 19852 2836 19892 2876
rect 39148 2836 39188 2876
rect 41740 2836 41780 2876
rect 46444 2836 46484 2876
rect 47116 2836 47156 2876
rect 52876 2836 52916 2876
rect 54508 2836 54548 2876
rect 844 2668 884 2708
rect 9676 2668 9716 2708
rect 54700 2668 54740 2708
rect 7660 2584 7700 2624
rect 8524 2584 8564 2624
rect 9868 2584 9908 2624
rect 11692 2584 11732 2624
rect 11980 2584 12020 2624
rect 14092 2584 14132 2624
rect 14476 2584 14516 2624
rect 15340 2584 15380 2624
rect 17836 2584 17876 2624
rect 18700 2584 18740 2624
rect 36748 2584 36788 2624
rect 37132 2584 37172 2624
rect 37996 2584 38036 2624
rect 39340 2584 39380 2624
rect 39724 2584 39764 2624
rect 40588 2584 40628 2624
rect 44044 2584 44084 2624
rect 44428 2584 44468 2624
rect 45292 2584 45332 2624
rect 48268 2584 48308 2624
rect 49132 2584 49172 2624
rect 49516 2584 49556 2624
rect 50476 2584 50516 2624
rect 50860 2584 50900 2624
rect 51724 2584 51764 2624
rect 7276 2500 7316 2540
rect 10540 2500 10580 2540
rect 12172 2500 12212 2540
rect 17452 2500 17492 2540
rect 652 2416 692 2456
rect 16492 2416 16532 2456
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 7852 2080 7892 2120
rect 8236 2080 8276 2120
rect 8908 2080 8948 2120
rect 17740 2080 17780 2120
rect 9580 1912 9620 1952
rect 17068 1912 17108 1952
rect 8044 1828 8084 1868
rect 8428 1828 8468 1868
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal2 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 95072 38576 95440 38585
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95072 38527 95440 38536
rect 12748 38240 12788 38249
rect 12788 38200 13364 38240
rect 12748 38191 12788 38200
rect 12076 37988 12116 37997
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 267 37568 309 37577
rect 267 37528 268 37568
rect 308 37528 309 37568
rect 267 37519 309 37528
rect 75 36728 117 36737
rect 75 36688 76 36728
rect 116 36688 117 36728
rect 75 36679 117 36688
rect 76 20105 116 36679
rect 268 23297 308 37519
rect 11308 37400 11348 37409
rect 10924 37316 10964 37325
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 10732 36896 10772 36905
rect 10924 36896 10964 37276
rect 10772 36856 10964 36896
rect 10732 36847 10772 36856
rect 7948 36728 7988 36737
rect 7276 36560 7316 36569
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 6123 35888 6165 35897
rect 6123 35848 6124 35888
rect 6164 35848 6165 35888
rect 6123 35839 6165 35848
rect 6699 35888 6741 35897
rect 6699 35848 6700 35888
rect 6740 35848 6741 35888
rect 6699 35839 6741 35848
rect 6988 35888 7028 35897
rect 5740 35804 5780 35813
rect 5780 35764 5972 35804
rect 5740 35755 5780 35764
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 5932 35384 5972 35764
rect 6124 35754 6164 35839
rect 5932 35335 5972 35344
rect 6700 35225 6740 35839
rect 6316 35216 6356 35225
rect 6123 35132 6165 35141
rect 6123 35092 6124 35132
rect 6164 35092 6165 35132
rect 6123 35083 6165 35092
rect 6124 34998 6164 35083
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 6316 34637 6356 35176
rect 6699 35216 6741 35225
rect 6699 35176 6700 35216
rect 6740 35176 6741 35216
rect 6699 35167 6741 35176
rect 6988 35057 7028 35848
rect 7276 35141 7316 36520
rect 7948 36140 7988 36688
rect 10924 36728 10964 36737
rect 10539 36644 10581 36653
rect 10539 36604 10540 36644
rect 10580 36604 10581 36644
rect 10539 36595 10581 36604
rect 8140 36140 8180 36149
rect 7948 36100 8140 36140
rect 10540 36140 10580 36595
rect 10828 36140 10868 36149
rect 10924 36140 10964 36688
rect 11308 36728 11348 37360
rect 11348 36688 11444 36728
rect 11308 36679 11348 36688
rect 10540 36100 10676 36140
rect 8140 36091 8180 36100
rect 10444 35888 10484 35897
rect 9675 35804 9717 35813
rect 9675 35764 9676 35804
rect 9716 35764 9717 35804
rect 9675 35755 9717 35764
rect 9004 35344 9332 35384
rect 9004 35300 9044 35344
rect 9004 35251 9044 35260
rect 7564 35216 7604 35225
rect 7275 35132 7317 35141
rect 7275 35092 7276 35132
rect 7316 35092 7317 35132
rect 7275 35083 7317 35092
rect 7564 35057 7604 35176
rect 8811 35216 8853 35225
rect 8811 35176 8812 35216
rect 8852 35176 8853 35216
rect 8811 35167 8853 35176
rect 8908 35216 8948 35227
rect 6699 35048 6741 35057
rect 6699 35008 6700 35048
rect 6740 35008 6741 35048
rect 6699 34999 6741 35008
rect 6987 35048 7029 35057
rect 6987 35008 6988 35048
rect 7028 35008 7029 35048
rect 6987 34999 7029 35008
rect 7563 35048 7605 35057
rect 7563 35008 7564 35048
rect 7604 35008 7605 35048
rect 7563 34999 7605 35008
rect 6315 34628 6357 34637
rect 6315 34588 6316 34628
rect 6356 34588 6357 34628
rect 6315 34579 6357 34588
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 6700 33872 6740 34999
rect 8716 34964 8756 34973
rect 8812 34964 8852 35167
rect 8908 35141 8948 35176
rect 9100 35216 9140 35225
rect 8907 35132 8949 35141
rect 8907 35092 8908 35132
rect 8948 35092 8949 35132
rect 8907 35083 8949 35092
rect 8812 34924 8948 34964
rect 7179 34628 7221 34637
rect 7179 34588 7180 34628
rect 7220 34588 7221 34628
rect 7179 34579 7221 34588
rect 7180 34494 7220 34579
rect 7372 34460 7412 34469
rect 7372 34217 7412 34420
rect 8716 34376 8756 34924
rect 8812 34376 8852 34385
rect 8716 34336 8812 34376
rect 8812 34327 8852 34336
rect 7371 34208 7413 34217
rect 7371 34168 7372 34208
rect 7412 34168 7413 34208
rect 7371 34159 7413 34168
rect 8139 34208 8181 34217
rect 8139 34168 8140 34208
rect 8180 34168 8181 34208
rect 8139 34159 8181 34168
rect 8140 34074 8180 34159
rect 6700 33823 6740 33832
rect 7180 33704 7220 33715
rect 7180 33629 7220 33664
rect 6316 33620 6356 33629
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 4108 32864 4148 32873
rect 3436 32780 3476 32789
rect 3476 32740 3572 32780
rect 3436 32731 3476 32740
rect 1900 32192 1940 32201
rect 2284 32192 2324 32201
rect 1940 32152 2228 32192
rect 1900 32143 1940 32152
rect 2188 31604 2228 32152
rect 2188 31555 2228 31564
rect 2284 31361 2324 32152
rect 3147 32192 3189 32201
rect 3147 32152 3148 32192
rect 3188 32152 3189 32192
rect 3147 32143 3189 32152
rect 3148 32058 3188 32143
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 3532 31445 3572 32740
rect 4108 32360 4148 32824
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 4300 32360 4340 32369
rect 4108 32320 4300 32360
rect 4300 32311 4340 32320
rect 6316 32201 6356 33580
rect 7179 33620 7221 33629
rect 7179 33580 7180 33620
rect 7220 33580 7221 33620
rect 7179 33571 7221 33580
rect 3819 32192 3861 32201
rect 3819 32152 3820 32192
rect 3860 32152 3861 32192
rect 3819 32143 3861 32152
rect 6315 32192 6357 32201
rect 6315 32152 6316 32192
rect 6356 32152 6357 32192
rect 6315 32143 6357 32152
rect 2379 31436 2421 31445
rect 2379 31396 2380 31436
rect 2420 31396 2421 31436
rect 2379 31387 2421 31396
rect 3531 31436 3573 31445
rect 3531 31396 3532 31436
rect 3572 31396 3573 31436
rect 3531 31387 3573 31396
rect 2283 31352 2325 31361
rect 2283 31312 2284 31352
rect 2324 31312 2325 31352
rect 2283 31303 2325 31312
rect 2380 31302 2420 31387
rect 2955 31352 2997 31361
rect 2955 31312 2956 31352
rect 2996 31312 2997 31352
rect 2955 31303 2997 31312
rect 3820 31352 3860 32143
rect 4011 31436 4053 31445
rect 4011 31396 4012 31436
rect 4052 31396 4053 31436
rect 4011 31387 4053 31396
rect 3820 31303 3860 31312
rect 2572 31268 2612 31277
rect 2612 31228 2900 31268
rect 2572 31219 2612 31228
rect 2667 31100 2709 31109
rect 2667 31060 2668 31100
rect 2708 31060 2709 31100
rect 2667 31051 2709 31060
rect 2668 28328 2708 31051
rect 2860 30848 2900 31228
rect 2956 31218 2996 31303
rect 3340 30848 3380 30857
rect 2860 30808 3340 30848
rect 3340 30799 3380 30808
rect 3531 30680 3573 30689
rect 3531 30640 3532 30680
rect 3572 30640 3573 30680
rect 3531 30631 3573 30640
rect 4012 30680 4052 31387
rect 7659 31352 7701 31361
rect 7659 31312 7660 31352
rect 7700 31312 7701 31352
rect 7659 31303 7701 31312
rect 4972 31184 5012 31193
rect 5012 31144 5108 31184
rect 4972 31135 5012 31144
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 4204 30689 4244 30774
rect 4012 30631 4052 30640
rect 4203 30680 4245 30689
rect 5068 30680 5108 31144
rect 4203 30640 4204 30680
rect 4244 30640 4340 30680
rect 4203 30631 4245 30640
rect 3532 30596 3572 30631
rect 3532 30545 3572 30556
rect 4300 30512 4340 30640
rect 5068 30631 5108 30640
rect 5643 30680 5685 30689
rect 5643 30640 5644 30680
rect 5684 30640 5685 30680
rect 5643 30631 5685 30640
rect 7275 30680 7317 30689
rect 7275 30640 7276 30680
rect 7316 30640 7317 30680
rect 7275 30631 7317 30640
rect 7660 30680 7700 31303
rect 7660 30631 7700 30640
rect 8524 30680 8564 30689
rect 4396 30512 4436 30521
rect 4300 30472 4396 30512
rect 4436 30472 4532 30512
rect 4396 30463 4436 30472
rect 4107 30428 4149 30437
rect 4107 30388 4108 30428
rect 4148 30388 4149 30428
rect 4107 30379 4149 30388
rect 4108 30294 4148 30379
rect 4492 30353 4532 30472
rect 5163 30428 5205 30437
rect 5163 30388 5164 30428
rect 5204 30388 5205 30428
rect 5163 30379 5205 30388
rect 4491 30344 4533 30353
rect 4491 30304 4492 30344
rect 4532 30304 4533 30344
rect 4491 30295 4533 30304
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 5164 29840 5204 30379
rect 5452 29840 5492 29849
rect 5164 29791 5204 29800
rect 5260 29800 5452 29840
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 5260 29336 5300 29800
rect 5452 29791 5492 29800
rect 5644 29756 5684 30631
rect 7276 30546 7316 30631
rect 6507 30344 6549 30353
rect 6507 30304 6508 30344
rect 6548 30304 6549 30344
rect 6507 30295 6549 30304
rect 5644 29707 5684 29716
rect 5164 29296 5300 29336
rect 5164 29252 5204 29296
rect 5164 29203 5204 29212
rect 4876 29168 4916 29177
rect 4684 29128 4876 29168
rect 3531 29000 3573 29009
rect 3531 28960 3532 29000
rect 3572 28960 3573 29000
rect 3531 28951 3573 28960
rect 4203 29000 4245 29009
rect 4203 28960 4204 29000
rect 4244 28960 4245 29000
rect 4203 28951 4245 28960
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 3532 28580 3572 28951
rect 4204 28866 4244 28951
rect 2284 28244 2324 28253
rect 2284 27497 2324 28204
rect 2668 27665 2708 28288
rect 3436 28540 3572 28580
rect 4684 28580 4724 29128
rect 4876 29119 4916 29128
rect 5068 29168 5108 29177
rect 5068 29009 5108 29128
rect 5260 29168 5300 29177
rect 5067 29000 5109 29009
rect 5067 28960 5068 29000
rect 5108 28960 5109 29000
rect 5067 28951 5109 28960
rect 2667 27656 2709 27665
rect 2667 27616 2668 27656
rect 2708 27616 2709 27656
rect 2667 27607 2709 27616
rect 2283 27488 2325 27497
rect 2283 27448 2284 27488
rect 2324 27448 2325 27488
rect 2283 27439 2325 27448
rect 2379 25892 2421 25901
rect 2379 25852 2380 25892
rect 2420 25852 2421 25892
rect 2379 25843 2421 25852
rect 2380 25304 2420 25843
rect 2668 25304 2708 27607
rect 3244 27497 3284 27582
rect 3436 27572 3476 28540
rect 4684 28531 4724 28540
rect 3532 28328 3572 28337
rect 5164 28328 5204 28337
rect 3572 28288 3668 28328
rect 3532 28279 3572 28288
rect 3628 27749 3668 28288
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 5164 27749 5204 28288
rect 5260 28169 5300 29128
rect 5835 28580 5877 28589
rect 5835 28540 5836 28580
rect 5876 28540 5877 28580
rect 5835 28531 5877 28540
rect 5836 28446 5876 28531
rect 6123 28328 6165 28337
rect 6123 28288 6124 28328
rect 6164 28288 6165 28328
rect 6123 28279 6165 28288
rect 6508 28328 6548 30295
rect 8524 28589 8564 30640
rect 8812 29168 8852 29177
rect 8523 28580 8565 28589
rect 8523 28540 8524 28580
rect 8564 28540 8565 28580
rect 8523 28531 8565 28540
rect 8812 28337 8852 29128
rect 6508 28279 6548 28288
rect 8811 28328 8853 28337
rect 8811 28288 8812 28328
rect 8852 28288 8853 28328
rect 8811 28279 8853 28288
rect 6124 28194 6164 28279
rect 5259 28160 5301 28169
rect 5259 28120 5260 28160
rect 5300 28120 5301 28160
rect 5259 28111 5301 28120
rect 6411 28160 6453 28169
rect 6411 28120 6412 28160
rect 6452 28120 6453 28160
rect 6411 28111 6453 28120
rect 6700 28160 6740 28169
rect 3627 27740 3669 27749
rect 3627 27700 3628 27740
rect 3668 27700 3669 27740
rect 3627 27691 3669 27700
rect 5163 27740 5205 27749
rect 5163 27700 5164 27740
rect 5204 27700 5205 27740
rect 5163 27691 5205 27700
rect 3436 27523 3476 27532
rect 3243 27488 3285 27497
rect 3243 27448 3244 27488
rect 3284 27448 3285 27488
rect 3243 27439 3285 27448
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 3435 26060 3477 26069
rect 3435 26020 3436 26060
rect 3476 26020 3477 26060
rect 3435 26011 3477 26020
rect 3244 25901 3284 25986
rect 3436 25926 3476 26011
rect 3243 25892 3285 25901
rect 3243 25852 3244 25892
rect 3284 25852 3285 25892
rect 3243 25843 3285 25852
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 2764 25304 2804 25313
rect 2668 25264 2764 25304
rect 2380 25255 2420 25264
rect 2764 25255 2804 25264
rect 3628 25304 3668 27691
rect 3916 27656 3956 27665
rect 4299 27656 4341 27665
rect 3956 27616 4148 27656
rect 3916 27607 3956 27616
rect 4108 27068 4148 27616
rect 4299 27616 4300 27656
rect 4340 27616 4341 27656
rect 4299 27607 4341 27616
rect 5164 27656 5204 27691
rect 4300 27522 4340 27607
rect 5164 27605 5204 27616
rect 5260 27077 5300 28111
rect 6412 28026 6452 28111
rect 6700 27749 6740 28120
rect 6699 27740 6741 27749
rect 6699 27700 6700 27740
rect 6740 27700 6741 27740
rect 6699 27691 6741 27700
rect 8619 27740 8661 27749
rect 8619 27700 8620 27740
rect 8660 27700 8661 27740
rect 8619 27691 8661 27700
rect 8620 27606 8660 27691
rect 6316 27404 6356 27413
rect 4492 27068 4532 27077
rect 4108 27028 4492 27068
rect 4492 27019 4532 27028
rect 4683 27068 4725 27077
rect 4683 27028 4684 27068
rect 4724 27028 4725 27068
rect 4683 27019 4725 27028
rect 5259 27068 5301 27077
rect 5259 27028 5260 27068
rect 5300 27028 5301 27068
rect 5259 27019 5301 27028
rect 5643 27068 5685 27077
rect 5643 27028 5644 27068
rect 5684 27028 5685 27068
rect 5643 27019 5685 27028
rect 4684 26900 4724 27019
rect 5644 26934 5684 27019
rect 4684 26851 4724 26860
rect 6316 26816 6356 27364
rect 8908 26825 8948 34924
rect 9100 34217 9140 35176
rect 9292 34376 9332 35344
rect 9292 34327 9332 34336
rect 9676 34376 9716 35755
rect 10444 35552 10484 35848
rect 10636 35888 10676 36100
rect 10868 36100 10964 36140
rect 10828 36091 10868 36100
rect 10636 35839 10676 35848
rect 11020 35972 11060 35981
rect 10539 35804 10581 35813
rect 10539 35764 10540 35804
rect 10580 35764 10581 35804
rect 10539 35755 10581 35764
rect 10540 35670 10580 35755
rect 11020 35720 11060 35932
rect 11212 35720 11252 35729
rect 11020 35680 11212 35720
rect 11020 35552 11060 35680
rect 11212 35671 11252 35680
rect 10444 35512 11060 35552
rect 10444 34376 10484 35512
rect 10540 34376 10580 34385
rect 10444 34336 10540 34376
rect 9676 34327 9716 34336
rect 10540 34327 10580 34336
rect 9099 34208 9141 34217
rect 9099 34168 9100 34208
rect 9140 34168 9141 34208
rect 9099 34159 9141 34168
rect 9772 34208 9812 34217
rect 9772 32780 9812 34168
rect 10443 34208 10485 34217
rect 10443 34168 10444 34208
rect 10484 34168 10485 34208
rect 10443 34159 10485 34168
rect 10732 34208 10772 34217
rect 10444 34074 10484 34159
rect 10059 33620 10101 33629
rect 10059 33580 10060 33620
rect 10100 33580 10101 33620
rect 10059 33571 10101 33580
rect 9292 32740 9812 32780
rect 9003 31352 9045 31361
rect 9003 31312 9004 31352
rect 9044 31312 9045 31352
rect 9003 31303 9045 31312
rect 9292 31352 9332 32740
rect 10060 32360 10100 33571
rect 10732 32780 10772 34168
rect 10732 32740 11060 32780
rect 10060 32311 10100 32320
rect 11020 32276 11060 32740
rect 11404 32705 11444 36688
rect 12076 36653 12116 37948
rect 13324 37652 13364 38200
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 93832 37820 94200 37829
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 93832 37771 94200 37780
rect 13324 37603 13364 37612
rect 18124 37484 18164 37493
rect 12172 37400 12212 37409
rect 12172 36728 12212 37360
rect 18124 37241 18164 37444
rect 25707 37484 25749 37493
rect 25707 37444 25708 37484
rect 25748 37444 25749 37484
rect 25707 37435 25749 37444
rect 26187 37484 26229 37493
rect 26187 37444 26188 37484
rect 26228 37444 26229 37484
rect 26187 37435 26229 37444
rect 26763 37484 26805 37493
rect 26763 37444 26764 37484
rect 26804 37444 26805 37484
rect 26763 37435 26805 37444
rect 39820 37484 39860 37493
rect 19468 37400 19508 37409
rect 22156 37400 22196 37409
rect 19180 37360 19468 37400
rect 17932 37232 17972 37241
rect 17932 36821 17972 37192
rect 18123 37232 18165 37241
rect 18123 37192 18124 37232
rect 18164 37192 18165 37232
rect 18123 37183 18165 37192
rect 18795 37232 18837 37241
rect 18795 37192 18796 37232
rect 18836 37192 18837 37232
rect 18795 37183 18837 37192
rect 18796 37098 18836 37183
rect 19180 36896 19220 37360
rect 19468 37351 19508 37360
rect 21964 37360 22156 37400
rect 21771 37232 21813 37241
rect 21771 37192 21772 37232
rect 21812 37192 21813 37232
rect 21771 37183 21813 37192
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 19180 36847 19220 36856
rect 16779 36812 16821 36821
rect 16779 36772 16780 36812
rect 16820 36772 16821 36812
rect 16779 36763 16821 36772
rect 17931 36812 17973 36821
rect 17931 36772 17932 36812
rect 17972 36772 17973 36812
rect 17931 36763 17973 36772
rect 12212 36688 12308 36728
rect 12172 36679 12212 36688
rect 12075 36644 12117 36653
rect 12075 36604 12076 36644
rect 12116 36604 12117 36644
rect 12075 36595 12117 36604
rect 11883 36560 11925 36569
rect 11883 36520 11884 36560
rect 11924 36520 11925 36560
rect 11883 36511 11925 36520
rect 11884 35888 11924 36511
rect 11884 35839 11924 35848
rect 12268 34385 12308 36688
rect 16780 36678 16820 36763
rect 17164 36728 17204 36737
rect 17164 36569 17204 36688
rect 18028 36728 18068 36737
rect 13323 36560 13365 36569
rect 13323 36520 13324 36560
rect 13364 36520 13365 36560
rect 13323 36511 13365 36520
rect 16203 36560 16245 36569
rect 16203 36520 16204 36560
rect 16244 36520 16245 36560
rect 16203 36511 16245 36520
rect 17163 36560 17205 36569
rect 17163 36520 17164 36560
rect 17204 36520 17205 36560
rect 17163 36511 17205 36520
rect 13324 36426 13364 36511
rect 16204 35888 16244 36511
rect 18028 35897 18068 36688
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 18219 35972 18261 35981
rect 18219 35932 18220 35972
rect 18260 35932 18261 35972
rect 18219 35923 18261 35932
rect 19083 35972 19125 35981
rect 19083 35932 19084 35972
rect 19124 35932 19125 35972
rect 19083 35923 19125 35932
rect 15819 35804 15861 35813
rect 15819 35764 15820 35804
rect 15860 35764 15861 35804
rect 15819 35755 15861 35764
rect 15820 35670 15860 35755
rect 12460 34544 12500 34553
rect 12460 34385 12500 34504
rect 11883 34376 11925 34385
rect 11883 34336 11884 34376
rect 11924 34336 11925 34376
rect 11883 34327 11925 34336
rect 12172 34376 12212 34385
rect 11884 34242 11924 34327
rect 12172 33629 12212 34336
rect 12267 34376 12309 34385
rect 12267 34336 12268 34376
rect 12308 34336 12309 34376
rect 12267 34327 12309 34336
rect 12459 34376 12501 34385
rect 12459 34336 12460 34376
rect 12500 34336 12501 34376
rect 12459 34327 12501 34336
rect 13132 34376 13172 34385
rect 12171 33620 12213 33629
rect 12171 33580 12172 33620
rect 12212 33580 12213 33620
rect 12171 33571 12213 33580
rect 11403 32696 11445 32705
rect 11403 32656 11404 32696
rect 11444 32656 11445 32696
rect 11403 32647 11445 32656
rect 11020 32227 11060 32236
rect 10444 32192 10484 32201
rect 9292 31303 9332 31312
rect 9675 31352 9717 31361
rect 9675 31312 9676 31352
rect 9716 31312 9717 31352
rect 9675 31303 9717 31312
rect 9004 27656 9044 31303
rect 9676 31218 9716 31303
rect 9675 30428 9717 30437
rect 9675 30388 9676 30428
rect 9716 30388 9717 30428
rect 9675 30379 9717 30388
rect 9676 30294 9716 30379
rect 10444 29177 10484 32152
rect 10539 32192 10581 32201
rect 10539 32152 10540 32192
rect 10580 32152 10581 32192
rect 10539 32143 10581 32152
rect 11404 32192 11444 32647
rect 11404 32143 11444 32152
rect 12268 32192 12308 34327
rect 13132 34049 13172 34336
rect 13131 34040 13173 34049
rect 13131 34000 13132 34040
rect 13172 34000 13173 34040
rect 13131 33991 13173 34000
rect 15627 34040 15669 34049
rect 15627 34000 15628 34040
rect 15668 34000 15669 34040
rect 15627 33991 15669 34000
rect 15532 33452 15572 33461
rect 14476 32873 14516 32958
rect 15532 32873 15572 33412
rect 14475 32864 14517 32873
rect 14475 32824 14476 32864
rect 14516 32824 14517 32864
rect 14475 32815 14517 32824
rect 14860 32864 14900 32873
rect 14860 32705 14900 32824
rect 15531 32864 15573 32873
rect 15531 32824 15532 32864
rect 15572 32824 15573 32864
rect 15628 32864 15668 33991
rect 15723 33620 15765 33629
rect 15723 33580 15724 33620
rect 15764 33580 15765 33620
rect 15723 33571 15765 33580
rect 15724 33486 15764 33571
rect 15724 32864 15764 32873
rect 15628 32824 15724 32864
rect 15531 32815 15573 32824
rect 15724 32815 15764 32824
rect 16204 32705 16244 35848
rect 17067 35888 17109 35897
rect 17067 35848 17068 35888
rect 17108 35848 17109 35888
rect 17067 35839 17109 35848
rect 18027 35888 18069 35897
rect 18027 35848 18028 35888
rect 18068 35848 18069 35888
rect 18027 35839 18069 35848
rect 16875 35804 16917 35813
rect 16875 35764 16876 35804
rect 16916 35764 16917 35804
rect 16875 35755 16917 35764
rect 16876 35048 16916 35755
rect 17068 35754 17108 35839
rect 18028 35225 18068 35839
rect 18220 35838 18260 35923
rect 19084 35888 19124 35923
rect 19084 35837 19124 35848
rect 21772 35888 21812 37183
rect 21867 36812 21909 36821
rect 21867 36772 21868 36812
rect 21908 36772 21909 36812
rect 21867 36763 21909 36772
rect 21868 36678 21908 36763
rect 21868 36140 21908 36149
rect 21964 36140 22004 37360
rect 22156 37351 22196 37360
rect 22540 37400 22580 37409
rect 22251 36728 22293 36737
rect 22251 36688 22252 36728
rect 22292 36688 22293 36728
rect 22251 36679 22293 36688
rect 22252 36594 22292 36679
rect 22540 36653 22580 37360
rect 25708 37350 25748 37435
rect 22636 37232 22676 37241
rect 22636 36821 22676 37192
rect 25131 37232 25173 37241
rect 25131 37192 25132 37232
rect 25172 37192 25173 37232
rect 25131 37183 25173 37192
rect 25515 37232 25557 37241
rect 25515 37192 25516 37232
rect 25556 37192 25557 37232
rect 25515 37183 25557 37192
rect 22635 36812 22677 36821
rect 22635 36772 22636 36812
rect 22676 36772 22677 36812
rect 22635 36763 22677 36772
rect 25132 36812 25172 37183
rect 25516 37098 25556 37183
rect 25132 36763 25172 36772
rect 23116 36728 23156 36737
rect 22539 36644 22581 36653
rect 22539 36604 22540 36644
rect 22580 36604 22581 36644
rect 22539 36595 22581 36604
rect 21908 36100 22004 36140
rect 21868 36091 21908 36100
rect 21772 35839 21812 35848
rect 21963 35888 22005 35897
rect 21963 35848 21964 35888
rect 22004 35848 22005 35888
rect 21963 35839 22005 35848
rect 21964 35754 22004 35839
rect 18412 35720 18452 35729
rect 18027 35216 18069 35225
rect 18027 35176 18028 35216
rect 18068 35176 18069 35216
rect 18027 35167 18069 35176
rect 18412 35141 18452 35680
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 18795 35216 18837 35225
rect 18795 35176 18796 35216
rect 18836 35176 18837 35216
rect 18795 35167 18837 35176
rect 20523 35216 20565 35225
rect 20523 35176 20524 35216
rect 20564 35176 20565 35216
rect 20523 35167 20565 35176
rect 21484 35216 21524 35225
rect 17067 35132 17109 35141
rect 17067 35092 17068 35132
rect 17108 35092 17109 35132
rect 17067 35083 17109 35092
rect 18123 35132 18165 35141
rect 18123 35092 18124 35132
rect 18164 35092 18165 35132
rect 18123 35083 18165 35092
rect 18411 35132 18453 35141
rect 18411 35092 18412 35132
rect 18452 35092 18453 35132
rect 18411 35083 18453 35092
rect 16876 34999 16916 35008
rect 17068 34998 17108 35083
rect 17068 33704 17108 33713
rect 16876 33664 17068 33704
rect 18124 33704 18164 35083
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 18412 33832 18740 33872
rect 18412 33788 18452 33832
rect 18412 33739 18452 33748
rect 18316 33704 18356 33713
rect 18124 33664 18316 33704
rect 16395 33620 16437 33629
rect 16395 33580 16396 33620
rect 16436 33580 16437 33620
rect 16395 33571 16437 33580
rect 16396 33452 16436 33571
rect 16396 32873 16436 33412
rect 16876 33116 16916 33664
rect 17068 33655 17108 33664
rect 18316 33655 18356 33664
rect 18508 33704 18548 33713
rect 18508 33452 18548 33664
rect 18700 33704 18740 33832
rect 18700 33655 18740 33664
rect 18508 33412 18740 33452
rect 18232 33284 18600 33293
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18232 33235 18600 33244
rect 16876 33067 16916 33076
rect 18028 32873 18068 32958
rect 18123 32948 18165 32957
rect 18123 32908 18124 32948
rect 18164 32908 18165 32948
rect 18123 32899 18165 32908
rect 16395 32864 16437 32873
rect 16395 32824 16396 32864
rect 16436 32824 16437 32864
rect 16395 32815 16437 32824
rect 18027 32864 18069 32873
rect 18027 32824 18028 32864
rect 18068 32824 18069 32864
rect 18027 32815 18069 32824
rect 18124 32780 18164 32899
rect 18124 32731 18164 32740
rect 18220 32864 18260 32873
rect 14859 32696 14901 32705
rect 14859 32656 14860 32696
rect 14900 32656 14901 32696
rect 14859 32647 14901 32656
rect 16203 32696 16245 32705
rect 16203 32656 16204 32696
rect 16244 32656 16245 32696
rect 16203 32647 16245 32656
rect 12268 32143 12308 32152
rect 10540 31352 10580 32143
rect 10540 31303 10580 31312
rect 13420 31940 13460 31949
rect 11692 31184 11732 31193
rect 11500 31144 11692 31184
rect 11115 30428 11157 30437
rect 11115 30388 11116 30428
rect 11156 30388 11157 30428
rect 11115 30379 11157 30388
rect 11116 29840 11156 30379
rect 11116 29791 11156 29800
rect 11500 29840 11540 31144
rect 11692 31135 11732 31144
rect 13420 30680 13460 31900
rect 13516 30680 13556 30689
rect 13420 30640 13516 30680
rect 13516 30631 13556 30640
rect 14188 30428 14228 30437
rect 11500 29791 11540 29800
rect 14092 30388 14188 30428
rect 11596 29672 11636 29681
rect 9771 29168 9813 29177
rect 9771 29128 9772 29168
rect 9812 29128 9813 29168
rect 9771 29119 9813 29128
rect 10443 29168 10485 29177
rect 10443 29128 10444 29168
rect 10484 29128 10485 29168
rect 11596 29168 11636 29632
rect 12364 29168 12404 29177
rect 11596 29128 12364 29168
rect 10443 29119 10485 29128
rect 12364 29119 12404 29128
rect 12460 29168 12500 29177
rect 9772 29034 9812 29119
rect 12460 29009 12500 29128
rect 9483 29000 9525 29009
rect 9483 28960 9484 29000
rect 9524 28960 9525 29000
rect 9483 28951 9525 28960
rect 11403 29000 11445 29009
rect 11403 28960 11404 29000
rect 11444 28960 11445 29000
rect 11403 28951 11445 28960
rect 12459 29000 12501 29009
rect 12459 28960 12460 29000
rect 12500 28960 12501 29000
rect 12459 28951 12501 28960
rect 13035 29000 13077 29009
rect 13035 28960 13036 29000
rect 13076 28960 13077 29000
rect 13035 28951 13077 28960
rect 9484 28866 9524 28951
rect 9868 27656 9908 27665
rect 9044 27616 9236 27656
rect 9004 27607 9044 27616
rect 6316 26767 6356 26776
rect 8907 26816 8949 26825
rect 8907 26776 8908 26816
rect 8948 26776 8949 26816
rect 8907 26767 8949 26776
rect 9196 26816 9236 27616
rect 9196 26767 9236 26776
rect 9483 26816 9525 26825
rect 9483 26776 9484 26816
rect 9524 26776 9525 26816
rect 9483 26767 9525 26776
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 4876 26144 4916 26153
rect 4107 26060 4149 26069
rect 4107 26020 4108 26060
rect 4148 26020 4149 26060
rect 4107 26011 4149 26020
rect 4108 25892 4148 26011
rect 4204 25892 4244 25901
rect 4108 25852 4204 25892
rect 3668 25264 3860 25304
rect 3628 25255 3668 25264
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 3820 23960 3860 25264
rect 3820 23920 3956 23960
rect 3628 23876 3668 23885
rect 3628 23633 3668 23836
rect 3436 23624 3476 23633
rect 2668 23584 3436 23624
rect 267 23288 309 23297
rect 267 23248 268 23288
rect 308 23248 309 23288
rect 267 23239 309 23248
rect 2668 23204 2708 23584
rect 3436 23575 3476 23584
rect 3627 23624 3669 23633
rect 3627 23584 3628 23624
rect 3668 23584 3669 23624
rect 3627 23575 3669 23584
rect 2668 23155 2708 23164
rect 3052 23120 3092 23131
rect 3052 23045 3092 23080
rect 3916 23120 3956 23920
rect 4108 23792 4148 25852
rect 4204 25843 4244 25852
rect 4780 25556 4820 25565
rect 4876 25556 4916 26104
rect 4820 25516 4916 25556
rect 4780 25507 4820 25516
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 4108 23743 4148 23752
rect 4300 23792 4340 23801
rect 4204 23708 4244 23717
rect 4204 23129 4244 23668
rect 4300 23633 4340 23752
rect 5164 23792 5204 23801
rect 4492 23633 4532 23718
rect 4299 23624 4341 23633
rect 4299 23584 4300 23624
rect 4340 23584 4341 23624
rect 4299 23575 4341 23584
rect 4491 23624 4533 23633
rect 4491 23584 4492 23624
rect 4532 23584 4533 23624
rect 4491 23575 4533 23584
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 5068 23288 5108 23297
rect 5164 23288 5204 23752
rect 8811 23792 8853 23801
rect 8811 23752 8812 23792
rect 8852 23752 8853 23792
rect 8811 23743 8853 23752
rect 9484 23792 9524 26767
rect 9868 26321 9908 27616
rect 11019 27572 11061 27581
rect 11019 27532 11020 27572
rect 11060 27532 11061 27572
rect 11019 27523 11061 27532
rect 11020 27438 11060 27523
rect 10059 26816 10101 26825
rect 10059 26776 10060 26816
rect 10100 26776 10101 26816
rect 10059 26767 10101 26776
rect 10060 26682 10100 26767
rect 9867 26312 9909 26321
rect 9867 26272 9868 26312
rect 9908 26272 9909 26312
rect 9867 26263 9909 26272
rect 10059 26312 10101 26321
rect 10059 26272 10060 26312
rect 10100 26272 10101 26312
rect 10059 26263 10101 26272
rect 10060 23801 10100 26263
rect 11404 26144 11444 28951
rect 12652 28916 12692 28925
rect 12076 28328 12116 28337
rect 12076 27581 12116 28288
rect 12652 27656 12692 28876
rect 13036 28580 13076 28951
rect 13036 28531 13076 28540
rect 14092 28337 14132 30388
rect 14188 30379 14228 30388
rect 15915 30176 15957 30185
rect 15915 30136 15916 30176
rect 15956 30136 15957 30176
rect 15915 30127 15957 30136
rect 15916 29840 15956 30127
rect 15916 29791 15956 29800
rect 16108 30092 16148 30101
rect 16204 30092 16244 32647
rect 18220 32276 18260 32824
rect 18124 32236 18260 32276
rect 17451 31940 17493 31949
rect 17451 31900 17452 31940
rect 17492 31900 17493 31940
rect 17451 31891 17493 31900
rect 18027 31940 18069 31949
rect 18027 31900 18028 31940
rect 18068 31900 18069 31940
rect 18027 31891 18069 31900
rect 17452 31352 17492 31891
rect 18028 31806 18068 31891
rect 17452 31303 17492 31312
rect 17836 31352 17876 31361
rect 17876 31312 17972 31352
rect 17836 31303 17876 31312
rect 17548 30680 17588 30689
rect 17548 30269 17588 30640
rect 17932 30680 17972 31312
rect 17972 30640 18068 30680
rect 17932 30631 17972 30640
rect 17547 30260 17589 30269
rect 17547 30220 17548 30260
rect 17588 30220 17589 30260
rect 17547 30211 17589 30220
rect 17931 30260 17973 30269
rect 17931 30220 17932 30260
rect 17972 30220 17973 30260
rect 17931 30211 17973 30220
rect 16148 30052 16244 30092
rect 17932 30092 17972 30211
rect 18028 30185 18068 30640
rect 18027 30176 18069 30185
rect 18027 30136 18028 30176
rect 18068 30136 18069 30176
rect 18027 30127 18069 30136
rect 18124 30101 18164 32236
rect 18220 32108 18260 32117
rect 18220 31949 18260 32068
rect 18700 31949 18740 33412
rect 18219 31940 18261 31949
rect 18219 31900 18220 31940
rect 18260 31900 18261 31940
rect 18219 31891 18261 31900
rect 18699 31940 18741 31949
rect 18699 31900 18700 31940
rect 18740 31900 18741 31940
rect 18699 31891 18741 31900
rect 18232 31772 18600 31781
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18232 31723 18600 31732
rect 18700 31352 18740 31361
rect 18796 31352 18836 35167
rect 20524 35082 20564 35167
rect 21196 34964 21236 34973
rect 21196 34553 21236 34924
rect 21195 34544 21237 34553
rect 21195 34504 21196 34544
rect 21236 34504 21237 34544
rect 21195 34495 21237 34504
rect 21484 34385 21524 35176
rect 23116 34553 23156 36688
rect 25515 36728 25557 36737
rect 25515 36688 25516 36728
rect 25556 36688 25557 36728
rect 25515 36679 25557 36688
rect 25516 36594 25556 36679
rect 24268 36476 24308 36485
rect 24308 36436 24500 36476
rect 24268 36427 24308 36436
rect 22155 34544 22197 34553
rect 22155 34504 22156 34544
rect 22196 34504 22197 34544
rect 22155 34495 22197 34504
rect 23115 34544 23157 34553
rect 23115 34504 23116 34544
rect 23156 34504 23157 34544
rect 23115 34495 23157 34504
rect 21292 34376 21332 34385
rect 19179 34292 19221 34301
rect 19179 34252 19180 34292
rect 19220 34252 19221 34292
rect 19179 34243 19221 34252
rect 20907 34292 20949 34301
rect 20907 34252 20908 34292
rect 20948 34252 20949 34292
rect 20907 34243 20949 34252
rect 19180 33872 19220 34243
rect 20908 34158 20948 34243
rect 21292 34049 21332 34336
rect 21483 34376 21525 34385
rect 21483 34336 21484 34376
rect 21524 34336 21525 34376
rect 21483 34327 21525 34336
rect 22156 34376 22196 34495
rect 23307 34460 23349 34469
rect 23307 34420 23308 34460
rect 23348 34420 23349 34460
rect 23307 34411 23349 34420
rect 24075 34460 24117 34469
rect 24075 34420 24076 34460
rect 24116 34420 24212 34460
rect 24075 34411 24117 34420
rect 22156 34327 22196 34336
rect 23115 34376 23157 34385
rect 23115 34336 23116 34376
rect 23156 34336 23157 34376
rect 23115 34327 23157 34336
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 21291 34040 21333 34049
rect 21291 34000 21292 34040
rect 21332 34000 21333 34040
rect 21291 33991 21333 34000
rect 22347 34040 22389 34049
rect 22347 34000 22348 34040
rect 22388 34000 22389 34040
rect 22347 33991 22389 34000
rect 19180 33823 19220 33832
rect 18988 33704 19028 33713
rect 18988 32957 19028 33664
rect 18987 32948 19029 32957
rect 18987 32908 18988 32948
rect 19028 32908 19029 32948
rect 18987 32899 19029 32908
rect 19472 32528 19840 32537
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19472 32479 19840 32488
rect 19852 32192 19892 32201
rect 19179 31940 19221 31949
rect 19179 31900 19180 31940
rect 19220 31900 19221 31940
rect 19179 31891 19221 31900
rect 19180 31806 19220 31891
rect 19852 31604 19892 32152
rect 20139 31940 20181 31949
rect 20139 31900 20140 31940
rect 20180 31900 20181 31940
rect 20139 31891 20181 31900
rect 19852 31555 19892 31564
rect 18740 31312 18836 31352
rect 20140 31352 20180 31891
rect 22348 31529 22388 33991
rect 23116 31604 23156 34327
rect 23308 34326 23348 34411
rect 24172 34376 24212 34420
rect 24172 34327 24212 34336
rect 24460 34376 24500 36436
rect 25707 35888 25749 35897
rect 26188 35888 26228 37435
rect 26764 37350 26804 37435
rect 27436 37400 27476 37409
rect 27436 36896 27476 37360
rect 39340 37400 39380 37409
rect 39380 37360 39572 37400
rect 39340 37351 39380 37360
rect 38668 37232 38708 37241
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 27532 36896 27572 36905
rect 27436 36856 27532 36896
rect 27532 36847 27572 36856
rect 26380 36728 26420 36737
rect 26283 36644 26325 36653
rect 26283 36604 26284 36644
rect 26324 36604 26325 36644
rect 26283 36595 26325 36604
rect 26284 36140 26324 36595
rect 26380 36140 26420 36688
rect 28203 36728 28245 36737
rect 28203 36688 28204 36728
rect 28244 36688 28245 36728
rect 28203 36679 28245 36688
rect 29643 36728 29685 36737
rect 29643 36688 29644 36728
rect 29684 36688 29685 36728
rect 29643 36679 29685 36688
rect 30219 36728 30261 36737
rect 35788 36728 35828 36737
rect 30219 36688 30220 36728
rect 30260 36688 30261 36728
rect 30219 36679 30261 36688
rect 35596 36688 35788 36728
rect 26380 36100 26516 36140
rect 26284 36091 26324 36100
rect 26380 35897 26420 35982
rect 25707 35848 25708 35888
rect 25748 35848 25749 35888
rect 25707 35839 25749 35848
rect 25804 35848 26188 35888
rect 25708 35216 25748 35839
rect 25804 35384 25844 35848
rect 26188 35839 26228 35848
rect 26379 35888 26421 35897
rect 26379 35848 26380 35888
rect 26420 35848 26421 35888
rect 26379 35839 26421 35848
rect 26476 35720 26516 36100
rect 27435 35972 27477 35981
rect 27435 35932 27436 35972
rect 27476 35932 27477 35972
rect 27435 35923 27477 35932
rect 27436 35838 27476 35923
rect 28204 35888 28244 36679
rect 29644 36594 29684 36679
rect 28972 36476 29012 36485
rect 28972 35981 29012 36436
rect 30220 36140 30260 36679
rect 34348 36644 34388 36655
rect 34348 36569 34388 36604
rect 33195 36560 33237 36569
rect 33195 36520 33196 36560
rect 33236 36520 33237 36560
rect 33195 36511 33237 36520
rect 34155 36560 34197 36569
rect 34155 36520 34156 36560
rect 34196 36520 34197 36560
rect 34155 36511 34197 36520
rect 34347 36560 34389 36569
rect 34347 36520 34348 36560
rect 34388 36520 34389 36560
rect 34347 36511 34389 36520
rect 35115 36560 35157 36569
rect 35115 36520 35116 36560
rect 35156 36520 35157 36560
rect 35115 36511 35157 36520
rect 30220 36091 30260 36100
rect 28971 35972 29013 35981
rect 28971 35932 28972 35972
rect 29012 35932 29013 35972
rect 28971 35923 29013 35932
rect 27820 35804 27860 35813
rect 25804 35335 25844 35344
rect 26284 35680 26516 35720
rect 27628 35720 27668 35729
rect 27820 35720 27860 35764
rect 27668 35680 27860 35720
rect 25748 35176 25940 35216
rect 25708 35167 25748 35176
rect 25516 34964 25556 34973
rect 25556 34924 25748 34964
rect 25516 34915 25556 34924
rect 24460 34327 24500 34336
rect 25323 34376 25365 34385
rect 25323 34336 25324 34376
rect 25364 34336 25365 34376
rect 25323 34327 25365 34336
rect 25324 34242 25364 34327
rect 24652 34208 24692 34217
rect 24652 32201 24692 34168
rect 25708 33788 25748 34924
rect 25708 33739 25748 33748
rect 25323 33704 25365 33713
rect 25323 33664 25324 33704
rect 25364 33664 25365 33704
rect 25323 33655 25365 33664
rect 25324 33570 25364 33655
rect 24651 32192 24693 32201
rect 24651 32152 24652 32192
rect 24692 32152 24693 32192
rect 24651 32143 24693 32152
rect 23116 31555 23156 31564
rect 22347 31520 22389 31529
rect 22347 31480 22348 31520
rect 22388 31480 22389 31520
rect 22347 31471 22389 31480
rect 18700 31303 18740 31312
rect 20140 31303 20180 31312
rect 20044 31184 20084 31193
rect 19472 31016 19840 31025
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19472 30967 19840 30976
rect 18796 30680 18836 30689
rect 18232 30260 18600 30269
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18232 30211 18600 30220
rect 12748 28328 12788 28337
rect 12940 28328 12980 28337
rect 12788 28288 12940 28328
rect 12748 28279 12788 28288
rect 12940 28279 12980 28288
rect 13131 28328 13173 28337
rect 13131 28288 13132 28328
rect 13172 28288 13173 28328
rect 13131 28279 13173 28288
rect 14091 28328 14133 28337
rect 14091 28288 14092 28328
rect 14132 28288 14133 28328
rect 14091 28279 14133 28288
rect 13132 28194 13172 28279
rect 13516 27656 13556 27665
rect 12652 27616 13516 27656
rect 13516 27607 13556 27616
rect 13708 27656 13748 27667
rect 13708 27581 13748 27616
rect 14092 27656 14132 28279
rect 14188 27740 14228 27749
rect 14228 27700 14612 27740
rect 14188 27691 14228 27700
rect 14092 27607 14132 27616
rect 14572 27656 14612 27700
rect 14572 27607 14612 27616
rect 12075 27572 12117 27581
rect 12075 27532 12076 27572
rect 12116 27532 12117 27572
rect 12075 27523 12117 27532
rect 13707 27572 13749 27581
rect 13707 27532 13708 27572
rect 13748 27532 13749 27572
rect 13707 27523 13749 27532
rect 12844 27404 12884 27413
rect 12748 26816 12788 26825
rect 12844 26816 12884 27364
rect 15244 27404 15284 27413
rect 12788 26776 12884 26816
rect 13131 26816 13173 26825
rect 13131 26776 13132 26816
rect 13172 26776 13173 26816
rect 12748 26767 12788 26776
rect 13131 26767 13173 26776
rect 13996 26816 14036 26825
rect 15244 26816 15284 27364
rect 16108 26825 16148 30052
rect 17932 30043 17972 30052
rect 18123 30092 18165 30101
rect 18123 30052 18124 30092
rect 18164 30052 18165 30092
rect 18123 30043 18165 30052
rect 18124 29924 18164 30043
rect 18124 29875 18164 29884
rect 18232 28748 18600 28757
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18232 28699 18600 28708
rect 18232 27236 18600 27245
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18232 27187 18600 27196
rect 18796 26825 18836 30640
rect 19948 30428 19988 30437
rect 19179 30092 19221 30101
rect 19179 30052 19180 30092
rect 19220 30052 19221 30092
rect 19179 30043 19221 30052
rect 19180 29958 19220 30043
rect 19852 29840 19892 29849
rect 19948 29840 19988 30388
rect 20044 30101 20084 31144
rect 20332 31184 20372 31193
rect 20332 30773 20372 31144
rect 20331 30764 20373 30773
rect 20331 30724 20332 30764
rect 20372 30724 20373 30764
rect 20331 30715 20373 30724
rect 21963 30764 22005 30773
rect 21963 30724 21964 30764
rect 22004 30724 22005 30764
rect 21963 30715 22005 30724
rect 21964 30630 22004 30715
rect 22348 30680 22388 31471
rect 23308 31352 23348 31361
rect 22348 30631 22388 30640
rect 23212 30680 23252 30689
rect 20139 30176 20181 30185
rect 20139 30136 20140 30176
rect 20180 30136 20181 30176
rect 20139 30127 20181 30136
rect 20043 30092 20085 30101
rect 20043 30052 20044 30092
rect 20084 30052 20085 30092
rect 20043 30043 20085 30052
rect 19892 29800 19988 29840
rect 19852 29791 19892 29800
rect 19472 29504 19840 29513
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19472 29455 19840 29464
rect 19472 27992 19840 28001
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19472 27943 19840 27952
rect 15340 26816 15380 26825
rect 15244 26776 15340 26816
rect 13132 26682 13172 26767
rect 13996 26321 14036 26776
rect 15340 26767 15380 26776
rect 15723 26816 15765 26825
rect 15723 26776 15724 26816
rect 15764 26776 15765 26816
rect 15723 26767 15765 26776
rect 16107 26816 16149 26825
rect 16107 26776 16108 26816
rect 16148 26776 16149 26816
rect 16107 26767 16149 26776
rect 16587 26816 16629 26825
rect 16587 26776 16588 26816
rect 16628 26776 16629 26816
rect 16587 26767 16629 26776
rect 18795 26816 18837 26825
rect 18795 26776 18796 26816
rect 18836 26776 18837 26816
rect 18795 26767 18837 26776
rect 19371 26816 19413 26825
rect 19371 26776 19372 26816
rect 19412 26776 19413 26816
rect 19371 26767 19413 26776
rect 19563 26816 19605 26825
rect 19563 26776 19564 26816
rect 19604 26776 19605 26816
rect 19563 26767 19605 26776
rect 15724 26682 15764 26767
rect 16588 26682 16628 26767
rect 15147 26648 15189 26657
rect 15147 26608 15148 26648
rect 15188 26608 15189 26648
rect 15147 26599 15189 26608
rect 17067 26648 17109 26657
rect 17067 26608 17068 26648
rect 17108 26608 17109 26648
rect 17067 26599 17109 26608
rect 17740 26648 17780 26657
rect 17780 26608 18068 26648
rect 17740 26599 17780 26608
rect 15148 26514 15188 26599
rect 11787 26312 11829 26321
rect 11787 26272 11788 26312
rect 11828 26272 11829 26312
rect 11787 26263 11829 26272
rect 13995 26312 14037 26321
rect 13995 26272 13996 26312
rect 14036 26272 14037 26312
rect 13995 26263 14037 26272
rect 11788 26178 11828 26263
rect 11404 26095 11444 26104
rect 13996 25229 14036 26263
rect 16780 25304 16820 25313
rect 13995 25220 14037 25229
rect 13995 25180 13996 25220
rect 14036 25180 14037 25220
rect 13995 25171 14037 25180
rect 15627 25220 15669 25229
rect 15627 25180 15628 25220
rect 15668 25180 15669 25220
rect 15627 25171 15669 25180
rect 6315 23708 6357 23717
rect 6315 23668 6316 23708
rect 6356 23668 6357 23708
rect 6315 23659 6357 23668
rect 6123 23624 6165 23633
rect 6123 23584 6124 23624
rect 6164 23584 6165 23624
rect 6123 23575 6165 23584
rect 5108 23248 5204 23288
rect 6028 23288 6068 23297
rect 5068 23239 5108 23248
rect 5739 23204 5781 23213
rect 5739 23164 5740 23204
rect 5780 23164 5781 23204
rect 5739 23155 5781 23164
rect 3916 23071 3956 23080
rect 4203 23120 4245 23129
rect 4203 23080 4204 23120
rect 4244 23080 4245 23120
rect 4203 23071 4245 23080
rect 5259 23120 5301 23129
rect 5259 23080 5260 23120
rect 5300 23080 5301 23120
rect 5259 23071 5301 23080
rect 5548 23120 5588 23129
rect 3051 23036 3093 23045
rect 2956 22996 3052 23036
rect 3092 22996 3093 23036
rect 652 22448 692 22457
rect 652 21617 692 22408
rect 2667 21692 2709 21701
rect 2667 21652 2668 21692
rect 2708 21652 2709 21692
rect 2667 21643 2709 21652
rect 651 21608 693 21617
rect 651 21568 652 21608
rect 692 21568 693 21608
rect 651 21559 693 21568
rect 2668 21558 2708 21643
rect 2956 21608 2996 22996
rect 3051 22987 3093 22996
rect 5260 22986 5300 23071
rect 5548 22709 5588 23080
rect 5740 23070 5780 23155
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 4203 22700 4245 22709
rect 4203 22660 4204 22700
rect 4244 22660 4245 22700
rect 4203 22651 4245 22660
rect 5547 22700 5589 22709
rect 5547 22660 5548 22700
rect 5588 22660 5589 22700
rect 5547 22651 5589 22660
rect 3627 22532 3669 22541
rect 3627 22492 3628 22532
rect 3668 22492 3669 22532
rect 3627 22483 3669 22492
rect 4204 22532 4244 22651
rect 6028 22541 6068 23248
rect 6124 23120 6164 23575
rect 6316 23288 6356 23659
rect 6316 23239 6356 23248
rect 7563 23204 7605 23213
rect 7563 23164 7564 23204
rect 7604 23164 7605 23204
rect 7563 23155 7605 23164
rect 6124 23071 6164 23080
rect 7564 23070 7604 23155
rect 7948 23120 7988 23131
rect 7948 23045 7988 23080
rect 8812 23120 8852 23743
rect 9099 23708 9141 23717
rect 9099 23668 9100 23708
rect 9140 23668 9141 23708
rect 9099 23659 9141 23668
rect 9100 23574 9140 23659
rect 8812 23071 8852 23080
rect 7947 23036 7989 23045
rect 7947 22996 7948 23036
rect 7988 22996 7989 23036
rect 7947 22987 7989 22996
rect 4204 22483 4244 22492
rect 4299 22532 4341 22541
rect 4299 22492 4300 22532
rect 4340 22492 4341 22532
rect 4299 22483 4341 22492
rect 4491 22532 4533 22541
rect 4491 22492 4492 22532
rect 4532 22492 4533 22532
rect 4491 22483 4533 22492
rect 6027 22532 6069 22541
rect 6027 22492 6028 22532
rect 6068 22492 6069 22532
rect 6027 22483 6069 22492
rect 3628 22364 3668 22483
rect 3628 22315 3668 22324
rect 4108 22280 4148 22289
rect 3436 22112 3476 22121
rect 3436 21701 3476 22072
rect 3435 21692 3477 21701
rect 3435 21652 3436 21692
rect 3476 21652 3477 21692
rect 3435 21643 3477 21652
rect 3052 21608 3092 21617
rect 2956 21568 3052 21608
rect 3052 21559 3092 21568
rect 3916 21608 3956 21617
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 652 20936 692 20945
rect 652 20777 692 20896
rect 651 20768 693 20777
rect 651 20728 652 20768
rect 692 20728 693 20768
rect 651 20719 693 20728
rect 2859 20180 2901 20189
rect 2859 20140 2860 20180
rect 2900 20140 2901 20180
rect 2859 20131 2901 20140
rect 3627 20180 3669 20189
rect 3627 20140 3628 20180
rect 3668 20140 3669 20180
rect 3627 20131 3669 20140
rect 75 20096 117 20105
rect 75 20056 76 20096
rect 116 20056 117 20096
rect 75 20047 117 20056
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 652 19794 692 19879
rect 652 19424 692 19433
rect 652 19097 692 19384
rect 2860 19340 2900 20131
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 3628 19508 3668 20131
rect 3628 19459 3668 19468
rect 2860 19291 2900 19300
rect 651 19088 693 19097
rect 651 19048 652 19088
rect 692 19048 693 19088
rect 651 19039 693 19048
rect 1707 19088 1749 19097
rect 1707 19048 1708 19088
rect 1748 19048 1749 19088
rect 1707 19039 1749 19048
rect 2667 19088 2709 19097
rect 2667 19048 2668 19088
rect 2708 19048 2709 19088
rect 2667 19039 2709 19048
rect 1708 18668 1748 19039
rect 2668 18954 2708 19039
rect 1708 18619 1748 18628
rect 3916 18593 3956 21568
rect 4108 20189 4148 22240
rect 4300 22280 4340 22483
rect 4492 22398 4532 22483
rect 4300 22231 4340 22240
rect 5164 22280 5204 22289
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 5068 21776 5108 21785
rect 5164 21776 5204 22240
rect 5108 21736 5204 21776
rect 5068 21727 5108 21736
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 9484 20189 9524 23752
rect 10059 23792 10101 23801
rect 10059 23752 10060 23792
rect 10100 23752 10101 23792
rect 10059 23743 10101 23752
rect 10347 23792 10389 23801
rect 10347 23752 10348 23792
rect 10388 23752 10389 23792
rect 10347 23743 10389 23752
rect 13516 23792 13556 23801
rect 14763 23792 14805 23801
rect 13556 23752 13748 23792
rect 13516 23743 13556 23752
rect 10348 23658 10388 23743
rect 11499 23624 11541 23633
rect 11499 23584 11500 23624
rect 11540 23584 11541 23624
rect 11499 23575 11541 23584
rect 12843 23624 12885 23633
rect 12843 23584 12844 23624
rect 12884 23584 12885 23624
rect 12843 23575 12885 23584
rect 11500 23490 11540 23575
rect 12844 23129 12884 23575
rect 13708 23288 13748 23752
rect 14763 23752 14764 23792
rect 14804 23752 14805 23792
rect 14763 23743 14805 23752
rect 15628 23792 15668 25171
rect 16780 23960 16820 25264
rect 17068 25304 17108 26599
rect 17068 25255 17108 25264
rect 17259 25304 17301 25313
rect 17259 25264 17260 25304
rect 17300 25264 17301 25304
rect 17259 25255 17301 25264
rect 17835 25304 17877 25313
rect 17835 25264 17836 25304
rect 17876 25264 17877 25304
rect 17835 25255 17877 25264
rect 17932 25304 17972 25313
rect 18028 25304 18068 26608
rect 19372 26153 19412 26767
rect 19564 26682 19604 26767
rect 19472 26480 19840 26489
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19472 26431 19840 26440
rect 18988 26144 19028 26153
rect 18232 25724 18600 25733
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18232 25675 18600 25684
rect 18988 25565 19028 26104
rect 19371 26144 19413 26153
rect 19371 26104 19372 26144
rect 19412 26104 19413 26144
rect 19371 26095 19413 26104
rect 19660 26144 19700 26153
rect 19852 26144 19892 26153
rect 19700 26104 19852 26144
rect 19660 26095 19700 26104
rect 19852 26095 19892 26104
rect 20140 26144 20180 30127
rect 22156 29168 22196 29177
rect 22059 27740 22101 27749
rect 22059 27700 22060 27740
rect 22100 27700 22101 27740
rect 22059 27691 22101 27700
rect 22060 27656 22100 27691
rect 22060 27605 22100 27616
rect 22156 27581 22196 29128
rect 23019 29168 23061 29177
rect 23019 29128 23020 29168
rect 23060 29128 23061 29168
rect 23019 29119 23061 29128
rect 22924 27656 22964 27665
rect 22155 27572 22197 27581
rect 22155 27532 22156 27572
rect 22196 27532 22197 27572
rect 22155 27523 22197 27532
rect 20907 27404 20949 27413
rect 20907 27364 20908 27404
rect 20948 27364 20949 27404
rect 20907 27355 20949 27364
rect 21867 27404 21909 27413
rect 21867 27364 21868 27404
rect 21908 27364 21909 27404
rect 21867 27355 21909 27364
rect 20908 27270 20948 27355
rect 20523 26816 20565 26825
rect 20523 26776 20524 26816
rect 20564 26776 20565 26816
rect 20523 26767 20565 26776
rect 20524 26682 20564 26767
rect 20236 26144 20276 26153
rect 20140 26104 20236 26144
rect 18123 25556 18165 25565
rect 18123 25516 18124 25556
rect 18164 25516 18165 25556
rect 18123 25507 18165 25516
rect 18987 25556 19029 25565
rect 18987 25516 18988 25556
rect 19028 25516 19029 25556
rect 18987 25507 19029 25516
rect 18124 25422 18164 25507
rect 19372 25388 19412 26095
rect 19468 25388 19508 25397
rect 19372 25348 19468 25388
rect 19468 25339 19508 25348
rect 18412 25304 18452 25313
rect 18028 25264 18412 25304
rect 17260 25220 17300 25255
rect 17260 25169 17300 25180
rect 17836 25170 17876 25255
rect 17932 24464 17972 25264
rect 18412 25255 18452 25264
rect 19084 25136 19124 25145
rect 18412 24760 18740 24800
rect 18412 24632 18452 24760
rect 18412 24583 18452 24592
rect 18603 24632 18645 24641
rect 18603 24592 18604 24632
rect 18644 24592 18645 24632
rect 18603 24583 18645 24592
rect 18604 24498 18644 24583
rect 18508 24464 18548 24473
rect 17932 24424 18508 24464
rect 18508 24415 18548 24424
rect 18232 24212 18600 24221
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18232 24163 18600 24172
rect 18700 24044 18740 24760
rect 19084 24641 19124 25096
rect 19472 24968 19840 24977
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19472 24919 19840 24928
rect 19083 24632 19125 24641
rect 19083 24592 19084 24632
rect 19124 24592 19125 24632
rect 19083 24583 19125 24592
rect 18700 23995 18740 24004
rect 19084 23960 19124 24583
rect 16780 23911 16820 23920
rect 18988 23920 19124 23960
rect 15628 23743 15668 23752
rect 16491 23792 16533 23801
rect 16491 23752 16492 23792
rect 16532 23752 16533 23792
rect 16491 23743 16533 23752
rect 18603 23792 18645 23801
rect 18603 23752 18604 23792
rect 18644 23752 18645 23792
rect 18603 23743 18645 23752
rect 14188 23708 14228 23717
rect 14380 23708 14420 23717
rect 14228 23668 14380 23708
rect 14188 23659 14228 23668
rect 14380 23659 14420 23668
rect 14764 23658 14804 23743
rect 13708 23239 13748 23248
rect 12843 23120 12885 23129
rect 12843 23080 12844 23120
rect 12884 23080 12885 23120
rect 12843 23071 12885 23080
rect 13996 23120 14036 23129
rect 10155 23036 10197 23045
rect 10155 22996 10156 23036
rect 10196 22996 10197 23036
rect 10155 22987 10197 22996
rect 9963 22868 10005 22877
rect 9963 22828 9964 22868
rect 10004 22828 10005 22868
rect 9963 22819 10005 22828
rect 9964 22734 10004 22819
rect 10156 21020 10196 22987
rect 12844 22986 12884 23071
rect 11115 22868 11157 22877
rect 11115 22828 11116 22868
rect 11156 22828 11157 22868
rect 11115 22819 11157 22828
rect 13515 22868 13557 22877
rect 13515 22828 13516 22868
rect 13556 22828 13557 22868
rect 13515 22819 13557 22828
rect 13899 22868 13941 22877
rect 13899 22828 13900 22868
rect 13940 22828 13941 22868
rect 13899 22819 13941 22828
rect 11116 22280 11156 22819
rect 13516 22734 13556 22819
rect 11595 22448 11637 22457
rect 11595 22408 11596 22448
rect 11636 22408 11637 22448
rect 11595 22399 11637 22408
rect 11116 22231 11156 22240
rect 11404 22280 11444 22289
rect 9868 20768 9908 20777
rect 9868 20189 9908 20728
rect 4107 20180 4149 20189
rect 4107 20140 4108 20180
rect 4148 20140 4149 20180
rect 4107 20131 4149 20140
rect 9099 20180 9141 20189
rect 9099 20140 9100 20180
rect 9140 20140 9141 20180
rect 9099 20131 9141 20140
rect 9483 20180 9525 20189
rect 9483 20140 9484 20180
rect 9524 20140 9525 20180
rect 9483 20131 9525 20140
rect 9867 20180 9909 20189
rect 9867 20140 9868 20180
rect 9908 20140 9909 20180
rect 9867 20131 9909 20140
rect 8716 20096 8756 20105
rect 4300 19256 4340 19265
rect 4108 19216 4300 19256
rect 4108 18752 4148 19216
rect 4300 19207 4340 19216
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 4108 18703 4148 18712
rect 7467 18752 7509 18761
rect 7467 18712 7468 18752
rect 7508 18712 7509 18752
rect 7467 18703 7509 18712
rect 8716 18752 8756 20056
rect 9100 20096 9140 20131
rect 9100 20045 9140 20056
rect 9964 20096 10004 20105
rect 9964 18761 10004 20056
rect 8716 18703 8756 18712
rect 9963 18752 10005 18761
rect 9963 18712 9964 18752
rect 10004 18712 10005 18752
rect 9963 18703 10005 18712
rect 7468 18618 7508 18703
rect 2092 18584 2132 18593
rect 652 18416 692 18425
rect 652 18257 692 18376
rect 651 18248 693 18257
rect 651 18208 652 18248
rect 692 18208 693 18248
rect 651 18199 693 18208
rect 652 17912 692 17921
rect 652 17417 692 17872
rect 2092 17753 2132 18544
rect 2955 18584 2997 18593
rect 2955 18544 2956 18584
rect 2996 18544 2997 18584
rect 2955 18535 2997 18544
rect 3915 18584 3957 18593
rect 3915 18544 3916 18584
rect 3956 18544 3957 18584
rect 3915 18535 3957 18544
rect 5355 18584 5397 18593
rect 5355 18544 5356 18584
rect 5396 18544 5397 18584
rect 5355 18535 5397 18544
rect 6988 18584 7028 18593
rect 2956 18450 2996 18535
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 5356 17753 5396 18535
rect 6795 18500 6837 18509
rect 6795 18460 6796 18500
rect 6836 18460 6837 18500
rect 6795 18451 6837 18460
rect 6796 18366 6836 18451
rect 5643 18332 5685 18341
rect 5643 18292 5644 18332
rect 5684 18292 5685 18332
rect 5643 18283 5685 18292
rect 6603 18332 6645 18341
rect 6603 18292 6604 18332
rect 6644 18292 6645 18332
rect 6603 18283 6645 18292
rect 2091 17744 2133 17753
rect 2091 17704 2092 17744
rect 2132 17704 2133 17744
rect 2091 17695 2133 17704
rect 4491 17744 4533 17753
rect 4491 17704 4492 17744
rect 4532 17704 4533 17744
rect 4491 17695 4533 17704
rect 5355 17744 5397 17753
rect 5355 17704 5356 17744
rect 5396 17704 5397 17744
rect 5355 17695 5397 17704
rect 4107 17660 4149 17669
rect 4107 17620 4108 17660
rect 4148 17620 4149 17660
rect 4107 17611 4149 17620
rect 4108 17526 4148 17611
rect 4492 17610 4532 17695
rect 5259 17660 5301 17669
rect 5259 17620 5260 17660
rect 5300 17620 5301 17660
rect 5259 17611 5301 17620
rect 651 17408 693 17417
rect 651 17368 652 17408
rect 692 17368 693 17408
rect 651 17359 693 17368
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 5260 17240 5300 17611
rect 5356 17610 5396 17695
rect 5260 17191 5300 17200
rect 5644 17156 5684 18283
rect 6604 18198 6644 18283
rect 6027 17828 6069 17837
rect 6027 17788 6028 17828
rect 6068 17788 6069 17828
rect 6027 17779 6069 17788
rect 6508 17828 6548 17837
rect 6548 17788 6740 17828
rect 6508 17779 6548 17788
rect 6028 17165 6068 17779
rect 6700 17744 6740 17788
rect 6988 17753 7028 18544
rect 7947 18584 7989 18593
rect 7947 18544 7948 18584
rect 7988 18544 7989 18584
rect 7947 18535 7989 18544
rect 8236 18584 8276 18593
rect 7659 18500 7701 18509
rect 7659 18460 7660 18500
rect 7700 18460 7701 18500
rect 7659 18451 7701 18460
rect 7660 18005 7700 18451
rect 7948 18450 7988 18535
rect 7659 17996 7701 18005
rect 7659 17956 7660 17996
rect 7700 17956 7701 17996
rect 7659 17947 7701 17956
rect 7660 17862 7700 17947
rect 6700 17695 6740 17704
rect 6987 17744 7029 17753
rect 6987 17704 6988 17744
rect 7028 17704 7029 17744
rect 6987 17695 7029 17704
rect 8043 17744 8085 17753
rect 8043 17704 8044 17744
rect 8084 17704 8085 17744
rect 8043 17695 8085 17704
rect 5644 17107 5684 17116
rect 6027 17156 6069 17165
rect 6027 17116 6028 17156
rect 6068 17116 6069 17156
rect 6027 17107 6069 17116
rect 6028 17072 6068 17107
rect 6028 17022 6068 17032
rect 6892 17072 6932 17081
rect 6988 17072 7028 17695
rect 6932 17032 7028 17072
rect 7372 17660 7412 17669
rect 6892 17023 6932 17032
rect 7372 16997 7412 17620
rect 8044 17240 8084 17695
rect 8236 17576 8276 18544
rect 8620 18584 8660 18593
rect 9483 18584 9525 18593
rect 8660 18544 8948 18584
rect 8620 18535 8660 18544
rect 8811 17996 8853 18005
rect 8811 17956 8812 17996
rect 8852 17956 8853 17996
rect 8811 17947 8853 17956
rect 8332 17753 8372 17838
rect 8331 17744 8373 17753
rect 8331 17704 8332 17744
rect 8372 17704 8373 17744
rect 8331 17695 8373 17704
rect 8812 17744 8852 17947
rect 8812 17695 8852 17704
rect 8908 17660 8948 18544
rect 9483 18544 9484 18584
rect 9524 18544 9525 18584
rect 9483 18535 9525 18544
rect 9003 17744 9045 17753
rect 9003 17704 9004 17744
rect 9044 17704 9045 17744
rect 9003 17695 9045 17704
rect 8908 17611 8948 17620
rect 9004 17610 9044 17695
rect 8236 17536 8372 17576
rect 8044 17191 8084 17200
rect 8332 17156 8372 17536
rect 8332 17107 8372 17116
rect 8236 17072 8276 17083
rect 8236 16997 8276 17032
rect 8428 17072 8468 17083
rect 8428 16997 8468 17032
rect 5451 16988 5493 16997
rect 5451 16948 5452 16988
rect 5492 16948 5493 16988
rect 5451 16939 5493 16948
rect 7371 16988 7413 16997
rect 7371 16948 7372 16988
rect 7412 16948 7413 16988
rect 7371 16939 7413 16948
rect 8235 16988 8277 16997
rect 8235 16948 8236 16988
rect 8276 16948 8277 16988
rect 8235 16939 8277 16948
rect 8427 16988 8469 16997
rect 8427 16948 8428 16988
rect 8468 16948 8469 16988
rect 8427 16939 8469 16948
rect 652 16904 692 16913
rect 652 16577 692 16864
rect 5452 16854 5492 16939
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 651 16568 693 16577
rect 651 16528 652 16568
rect 692 16528 693 16568
rect 651 16519 693 16528
rect 652 16400 692 16409
rect 556 16360 652 16400
rect 556 15737 596 16360
rect 652 16351 692 16360
rect 9484 16241 9524 18535
rect 10156 17165 10196 20980
rect 11404 20180 11444 22240
rect 11596 22196 11636 22399
rect 13900 22280 13940 22819
rect 13996 22532 14036 23080
rect 13996 22483 14036 22492
rect 14092 23120 14132 23129
rect 14092 22457 14132 23080
rect 14475 23120 14517 23129
rect 14475 23080 14476 23120
rect 14516 23080 14517 23120
rect 14475 23071 14517 23080
rect 14091 22448 14133 22457
rect 14091 22408 14092 22448
rect 14132 22408 14133 22448
rect 14091 22399 14133 22408
rect 13900 22231 13940 22240
rect 14091 22280 14133 22289
rect 14091 22240 14092 22280
rect 14132 22240 14133 22280
rect 14091 22231 14133 22240
rect 14476 22280 14516 23071
rect 16492 22373 16532 23743
rect 18604 23120 18644 23743
rect 18988 23120 19028 23920
rect 19371 23792 19413 23801
rect 19371 23752 19372 23792
rect 19412 23752 19413 23792
rect 19371 23743 19413 23752
rect 19372 23658 19412 23743
rect 19472 23456 19840 23465
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19472 23407 19840 23416
rect 19084 23204 19124 23213
rect 19124 23164 19604 23204
rect 19084 23155 19124 23164
rect 18644 23080 18740 23120
rect 18604 23071 18644 23080
rect 18232 22700 18600 22709
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18232 22651 18600 22660
rect 18508 22532 18548 22541
rect 18700 22532 18740 23080
rect 18988 23071 19028 23080
rect 19564 23120 19604 23164
rect 19564 23071 19604 23080
rect 19755 22868 19797 22877
rect 19755 22828 19756 22868
rect 19796 22828 19797 22868
rect 19755 22819 19797 22828
rect 18548 22492 18740 22532
rect 18508 22483 18548 22492
rect 16491 22364 16533 22373
rect 16491 22324 16492 22364
rect 16532 22324 16533 22364
rect 16491 22315 16533 22324
rect 14476 22231 14516 22240
rect 14859 22280 14901 22289
rect 15244 22280 15284 22289
rect 14859 22240 14860 22280
rect 14900 22240 14901 22280
rect 14859 22231 14901 22240
rect 14956 22240 15244 22280
rect 11596 22147 11636 22156
rect 14092 22146 14132 22231
rect 14860 21785 14900 22231
rect 14956 22196 14996 22240
rect 15244 22231 15284 22240
rect 16492 22280 16532 22315
rect 16492 22230 16532 22240
rect 17355 22280 17397 22289
rect 17355 22240 17356 22280
rect 17396 22240 17397 22280
rect 17355 22231 17397 22240
rect 19756 22280 19796 22819
rect 20140 22373 20180 26104
rect 20236 26095 20276 26104
rect 20331 26144 20373 26153
rect 20331 26104 20332 26144
rect 20372 26104 20373 26144
rect 20331 26095 20373 26104
rect 21099 26144 21141 26153
rect 21099 26104 21100 26144
rect 21140 26104 21141 26144
rect 21099 26095 21141 26104
rect 20235 22868 20277 22877
rect 20235 22828 20236 22868
rect 20276 22828 20277 22868
rect 20235 22819 20277 22828
rect 20236 22734 20276 22819
rect 20139 22364 20181 22373
rect 20139 22324 20140 22364
rect 20180 22324 20181 22364
rect 20139 22315 20181 22324
rect 19756 22231 19796 22240
rect 20140 22280 20180 22315
rect 20332 22289 20372 26095
rect 21100 26010 21140 26095
rect 21868 25304 21908 27355
rect 22156 26825 22196 27523
rect 22155 26816 22197 26825
rect 22155 26776 22156 26816
rect 22196 26776 22197 26816
rect 22155 26767 22197 26776
rect 22252 25892 22292 25901
rect 22252 25313 22292 25852
rect 22251 25304 22293 25313
rect 21908 25264 22100 25304
rect 21868 25255 21908 25264
rect 21963 25136 22005 25145
rect 21963 25096 21964 25136
rect 22004 25096 22005 25136
rect 21963 25087 22005 25096
rect 21867 23120 21909 23129
rect 21867 23080 21868 23120
rect 21908 23080 21909 23120
rect 21867 23071 21909 23080
rect 21964 23120 22004 25087
rect 21964 23071 22004 23080
rect 21868 22986 21908 23071
rect 21676 22868 21716 22877
rect 14956 22147 14996 22156
rect 15916 22196 15956 22205
rect 16108 22196 16148 22205
rect 15956 22156 16108 22196
rect 15916 22147 15956 22156
rect 16108 22147 16148 22156
rect 17356 22146 17396 22231
rect 20140 22229 20180 22240
rect 20331 22280 20373 22289
rect 20331 22240 20332 22280
rect 20372 22240 20373 22280
rect 20331 22231 20373 22240
rect 21003 22280 21045 22289
rect 21003 22240 21004 22280
rect 21044 22240 21045 22280
rect 21003 22231 21045 22240
rect 21004 22146 21044 22231
rect 19472 21944 19840 21953
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19472 21895 19840 21904
rect 14859 21776 14901 21785
rect 14859 21736 14860 21776
rect 14900 21736 14901 21776
rect 14859 21727 14901 21736
rect 15243 21776 15285 21785
rect 15243 21736 15244 21776
rect 15284 21736 15285 21776
rect 15243 21727 15285 21736
rect 15244 21642 15284 21727
rect 15916 21608 15956 21617
rect 15436 21568 15916 21608
rect 13995 20768 14037 20777
rect 13995 20728 13996 20768
rect 14036 20728 14037 20768
rect 13995 20719 14037 20728
rect 14571 20768 14613 20777
rect 14571 20728 14572 20768
rect 14612 20728 14613 20768
rect 14571 20719 14613 20728
rect 11116 20140 11444 20180
rect 13419 20180 13461 20189
rect 13419 20140 13420 20180
rect 13460 20140 13461 20180
rect 11116 20012 11156 20140
rect 13419 20131 13461 20140
rect 11116 19963 11156 19972
rect 13036 20096 13076 20105
rect 13036 19013 13076 20056
rect 13420 20096 13460 20131
rect 13420 20045 13460 20056
rect 12075 19004 12117 19013
rect 12075 18964 12076 19004
rect 12116 18964 12117 19004
rect 12075 18955 12117 18964
rect 13035 19004 13077 19013
rect 13035 18964 13036 19004
rect 13076 18964 13077 19004
rect 13035 18955 13077 18964
rect 11019 18752 11061 18761
rect 11019 18712 11020 18752
rect 11060 18712 11061 18752
rect 11019 18703 11061 18712
rect 11787 18752 11829 18761
rect 11787 18712 11788 18752
rect 11828 18712 11829 18752
rect 11787 18703 11829 18712
rect 12076 18752 12116 18955
rect 12076 18703 12116 18712
rect 12267 18752 12309 18761
rect 12267 18712 12268 18752
rect 12308 18712 12309 18752
rect 12267 18703 12309 18712
rect 11020 17753 11060 18703
rect 11788 18618 11828 18703
rect 12268 18618 12308 18703
rect 11884 18584 11924 18593
rect 11019 17744 11061 17753
rect 11019 17704 11020 17744
rect 11060 17704 11061 17744
rect 11019 17695 11061 17704
rect 11308 17744 11348 17753
rect 10924 17660 10964 17669
rect 10540 17240 10580 17249
rect 10580 17200 10772 17240
rect 10540 17191 10580 17200
rect 10155 17156 10197 17165
rect 10155 17116 10156 17156
rect 10196 17116 10197 17156
rect 10155 17107 10197 17116
rect 10732 17156 10772 17200
rect 10732 17107 10772 17116
rect 10347 16988 10389 16997
rect 10347 16948 10348 16988
rect 10388 16948 10389 16988
rect 10347 16939 10389 16948
rect 10348 16854 10388 16939
rect 10828 16400 10868 16409
rect 10924 16400 10964 17620
rect 10868 16360 10964 16400
rect 10828 16351 10868 16360
rect 11020 16316 11060 17695
rect 11308 17165 11348 17704
rect 11115 17156 11157 17165
rect 11115 17116 11116 17156
rect 11156 17116 11157 17156
rect 11115 17107 11157 17116
rect 11307 17156 11349 17165
rect 11307 17116 11308 17156
rect 11348 17116 11349 17156
rect 11307 17107 11349 17116
rect 11116 17072 11156 17107
rect 11116 17021 11156 17032
rect 11884 16997 11924 18544
rect 12940 18584 12980 18593
rect 12980 18544 13364 18584
rect 12940 18535 12980 18544
rect 13324 17996 13364 18544
rect 13324 17947 13364 17956
rect 12172 17744 12212 17755
rect 12172 17669 12212 17704
rect 11979 17660 12021 17669
rect 11979 17620 11980 17660
rect 12020 17620 12021 17660
rect 11979 17611 12021 17620
rect 12171 17660 12213 17669
rect 12171 17620 12172 17660
rect 12212 17620 12213 17660
rect 12171 17611 12213 17620
rect 12939 17660 12981 17669
rect 12939 17620 12940 17660
rect 12980 17620 12981 17660
rect 12939 17611 12981 17620
rect 11980 17072 12020 17611
rect 11980 17023 12020 17032
rect 11883 16988 11925 16997
rect 11883 16948 11884 16988
rect 11924 16948 11925 16988
rect 11883 16939 11925 16948
rect 11884 16484 11924 16939
rect 12363 16820 12405 16829
rect 12363 16780 12364 16820
rect 12404 16780 12405 16820
rect 12363 16771 12405 16780
rect 11692 16444 11924 16484
rect 11692 16400 11732 16444
rect 11692 16351 11732 16360
rect 11020 16267 11060 16276
rect 9483 16232 9525 16241
rect 9483 16192 9484 16232
rect 9524 16192 9525 16232
rect 9483 16183 9525 16192
rect 12364 16232 12404 16771
rect 12940 16400 12980 17611
rect 13131 16820 13173 16829
rect 13131 16780 13132 16820
rect 13172 16780 13173 16820
rect 13131 16771 13173 16780
rect 13132 16686 13172 16771
rect 12940 16351 12980 16360
rect 12364 16183 12404 16192
rect 12651 16232 12693 16241
rect 12651 16192 12652 16232
rect 12692 16192 12693 16232
rect 12651 16183 12693 16192
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 555 15728 597 15737
rect 555 15688 556 15728
rect 596 15688 597 15728
rect 555 15679 597 15688
rect 652 15728 692 15737
rect 652 14897 692 15688
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 9484 14972 9524 16183
rect 12652 16098 12692 16183
rect 13516 16148 13556 16157
rect 9484 14923 9524 14932
rect 651 14888 693 14897
rect 651 14848 652 14888
rect 692 14848 693 14888
rect 651 14839 693 14848
rect 9771 14720 9813 14729
rect 9771 14680 9772 14720
rect 9812 14680 9813 14720
rect 9771 14671 9813 14680
rect 652 14552 692 14561
rect 652 14057 692 14512
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 651 14048 693 14057
rect 651 14008 652 14048
rect 692 14008 693 14048
rect 651 13999 693 14008
rect 4204 14048 4244 14057
rect 4244 14008 4532 14048
rect 4204 13999 4244 14008
rect 3532 13796 3572 13805
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 651 13208 693 13217
rect 651 13168 652 13208
rect 692 13168 693 13208
rect 651 13159 693 13168
rect 2475 13208 2517 13217
rect 2475 13168 2476 13208
rect 2516 13168 2517 13208
rect 2475 13159 2517 13168
rect 2955 13208 2997 13217
rect 2955 13168 2956 13208
rect 2996 13168 2997 13208
rect 2955 13159 2997 13168
rect 3340 13208 3380 13217
rect 652 13040 692 13159
rect 652 12991 692 13000
rect 2092 13124 2132 13133
rect 652 12704 692 12713
rect 2092 12704 2132 13084
rect 2476 13074 2516 13159
rect 2188 12704 2228 12713
rect 2092 12664 2188 12704
rect 652 12377 692 12664
rect 2188 12655 2228 12664
rect 2572 12536 2612 12545
rect 2956 12536 2996 13159
rect 3340 12545 3380 13168
rect 2612 12496 2900 12536
rect 2572 12487 2612 12496
rect 2379 12452 2421 12461
rect 2379 12412 2380 12452
rect 2420 12412 2421 12452
rect 2379 12403 2421 12412
rect 651 12368 693 12377
rect 651 12328 652 12368
rect 692 12328 693 12368
rect 651 12319 693 12328
rect 2380 12318 2420 12403
rect 2860 11948 2900 12496
rect 2956 12377 2996 12496
rect 3339 12536 3381 12545
rect 3339 12496 3340 12536
rect 3380 12496 3381 12536
rect 3339 12487 3381 12496
rect 3532 12461 3572 13756
rect 4492 13460 4532 14008
rect 4492 13411 4532 13420
rect 9772 13217 9812 14671
rect 12172 14048 12212 14057
rect 11884 14008 12172 14048
rect 8043 13208 8085 13217
rect 8043 13168 8044 13208
rect 8084 13168 8085 13208
rect 8043 13159 8085 13168
rect 9196 13208 9236 13217
rect 7180 13124 7220 13133
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 3627 12536 3669 12545
rect 3627 12496 3628 12536
rect 3668 12496 3669 12536
rect 3627 12487 3669 12496
rect 3819 12536 3861 12545
rect 6220 12536 6260 12545
rect 3819 12496 3820 12536
rect 3860 12496 3861 12536
rect 3819 12487 3861 12496
rect 5644 12496 6220 12536
rect 3531 12452 3573 12461
rect 3531 12412 3532 12452
rect 3572 12412 3573 12452
rect 3531 12403 3573 12412
rect 2955 12368 2997 12377
rect 2955 12328 2956 12368
rect 2996 12328 2997 12368
rect 2955 12319 2997 12328
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 3244 11948 3284 11957
rect 2860 11908 3244 11948
rect 3244 11899 3284 11908
rect 3532 11789 3572 12403
rect 3436 11780 3476 11789
rect 3436 11537 3476 11740
rect 3531 11780 3573 11789
rect 3531 11740 3532 11780
rect 3572 11740 3573 11780
rect 3531 11731 3573 11740
rect 651 11528 693 11537
rect 651 11488 652 11528
rect 692 11488 693 11528
rect 651 11479 693 11488
rect 3435 11528 3477 11537
rect 3435 11488 3436 11528
rect 3476 11488 3477 11528
rect 3435 11479 3477 11488
rect 652 11394 692 11479
rect 652 11192 692 11201
rect 652 10697 692 11152
rect 651 10688 693 10697
rect 651 10648 652 10688
rect 692 10648 693 10688
rect 651 10639 693 10648
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 3628 10436 3668 12487
rect 3820 12402 3860 12487
rect 3723 12368 3765 12377
rect 3723 12328 3724 12368
rect 3764 12328 3765 12368
rect 3723 12319 3765 12328
rect 939 10100 981 10109
rect 939 10060 940 10100
rect 980 10060 981 10100
rect 939 10051 981 10060
rect 652 10016 692 10025
rect 652 9857 692 9976
rect 651 9848 693 9857
rect 651 9808 652 9848
rect 692 9808 693 9848
rect 651 9799 693 9808
rect 652 9680 692 9689
rect 652 9017 692 9640
rect 843 9176 885 9185
rect 843 9136 844 9176
rect 884 9136 885 9176
rect 843 9127 885 9136
rect 651 9008 693 9017
rect 651 8968 652 9008
rect 692 8968 693 9008
rect 651 8959 693 8968
rect 652 8504 692 8513
rect 556 8464 652 8504
rect 556 8177 596 8464
rect 652 8455 692 8464
rect 555 8168 597 8177
rect 555 8128 556 8168
rect 596 8128 597 8168
rect 555 8119 597 8128
rect 652 8168 692 8177
rect 652 7337 692 8128
rect 651 7328 693 7337
rect 651 7288 652 7328
rect 692 7288 693 7328
rect 651 7279 693 7288
rect 652 6992 692 7001
rect 652 6497 692 6952
rect 651 6488 693 6497
rect 651 6448 652 6488
rect 692 6448 693 6488
rect 651 6439 693 6448
rect 651 5648 693 5657
rect 651 5608 652 5648
rect 692 5608 693 5648
rect 651 5599 693 5608
rect 652 5480 692 5599
rect 652 5431 692 5440
rect 844 4892 884 9127
rect 844 4843 884 4852
rect 651 4808 693 4817
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 652 4674 692 4759
rect 844 4220 884 4229
rect 940 4220 980 10051
rect 2955 9680 2997 9689
rect 2955 9640 2956 9680
rect 2996 9640 2997 9680
rect 2955 9631 2997 9640
rect 3339 9680 3381 9689
rect 3339 9640 3340 9680
rect 3380 9640 3381 9680
rect 3339 9631 3381 9640
rect 2475 9512 2517 9521
rect 2475 9472 2476 9512
rect 2516 9472 2517 9512
rect 2475 9463 2517 9472
rect 2379 8756 2421 8765
rect 2379 8716 2380 8756
rect 2420 8716 2421 8756
rect 2379 8707 2421 8716
rect 2380 8672 2420 8707
rect 2380 8621 2420 8632
rect 1996 8588 2036 8597
rect 2036 8548 2324 8588
rect 1996 8539 2036 8548
rect 2284 8168 2324 8548
rect 2284 8119 2324 8128
rect 2476 7916 2516 9463
rect 2956 9428 2996 9631
rect 3243 9596 3285 9605
rect 3243 9556 3244 9596
rect 3284 9556 3285 9596
rect 3243 9547 3285 9556
rect 3147 9512 3189 9521
rect 3147 9472 3148 9512
rect 3188 9472 3189 9512
rect 3147 9463 3189 9472
rect 2956 9379 2996 9388
rect 3148 9378 3188 9463
rect 3244 9462 3284 9547
rect 3340 9512 3380 9631
rect 3340 9463 3380 9472
rect 3531 9512 3573 9521
rect 3531 9472 3532 9512
rect 3572 9472 3573 9512
rect 3531 9463 3573 9472
rect 3532 9378 3572 9463
rect 2764 9260 2804 9269
rect 2668 8084 2708 8093
rect 2764 8084 2804 9220
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 3051 8756 3093 8765
rect 3051 8716 3052 8756
rect 3092 8716 3093 8756
rect 3051 8707 3093 8716
rect 2708 8044 2804 8084
rect 2668 8035 2708 8044
rect 3052 8000 3092 8707
rect 3628 8681 3668 10396
rect 3724 8765 3764 12319
rect 4972 12284 5012 12293
rect 3915 11780 3957 11789
rect 3915 11740 3916 11780
rect 3956 11740 3957 11780
rect 3915 11731 3957 11740
rect 3916 11696 3956 11731
rect 3916 11645 3956 11656
rect 4011 11696 4053 11705
rect 4011 11656 4012 11696
rect 4052 11656 4053 11696
rect 4011 11647 4053 11656
rect 4108 11696 4148 11705
rect 4012 11562 4052 11647
rect 4108 11537 4148 11656
rect 4972 11696 5012 12244
rect 4972 11647 5012 11656
rect 5163 11696 5205 11705
rect 5163 11656 5164 11696
rect 5204 11656 5205 11696
rect 5163 11647 5205 11656
rect 5452 11696 5492 11705
rect 4300 11537 4340 11622
rect 5164 11562 5204 11647
rect 4107 11528 4149 11537
rect 4107 11488 4108 11528
rect 4148 11488 4149 11528
rect 4107 11479 4149 11488
rect 4299 11528 4341 11537
rect 4299 11488 4300 11528
rect 4340 11488 4341 11528
rect 4299 11479 4341 11488
rect 5355 11528 5397 11537
rect 5355 11488 5356 11528
rect 5396 11488 5397 11528
rect 5355 11479 5397 11488
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 4203 11276 4245 11285
rect 4203 11236 4204 11276
rect 4244 11236 4245 11276
rect 4203 11227 4245 11236
rect 4204 10184 4244 11227
rect 4204 10135 4244 10144
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 4395 9680 4437 9689
rect 4395 9640 4396 9680
rect 4436 9640 4437 9680
rect 4395 9631 4437 9640
rect 5259 9680 5301 9689
rect 5259 9640 5260 9680
rect 5300 9640 5301 9680
rect 5259 9631 5301 9640
rect 4396 9546 4436 9631
rect 5260 9546 5300 9631
rect 4204 9512 4244 9521
rect 5068 9512 5108 9521
rect 4244 9472 4340 9512
rect 4204 9463 4244 9472
rect 4300 8924 4340 9472
rect 4779 9260 4821 9269
rect 4779 9220 4780 9260
rect 4820 9220 4821 9260
rect 4779 9211 4821 9220
rect 4396 8924 4436 8933
rect 4300 8884 4396 8924
rect 4396 8875 4436 8884
rect 3723 8756 3765 8765
rect 3723 8716 3724 8756
rect 3764 8716 3765 8756
rect 3723 8707 3765 8716
rect 3243 8672 3285 8681
rect 3243 8632 3244 8672
rect 3284 8632 3285 8672
rect 3243 8623 3285 8632
rect 3627 8672 3669 8681
rect 3627 8632 3628 8672
rect 3668 8632 3669 8672
rect 3627 8623 3669 8632
rect 3915 8672 3957 8681
rect 3915 8632 3916 8672
rect 3956 8632 3957 8672
rect 3915 8623 3957 8632
rect 4780 8672 4820 9211
rect 4780 8623 4820 8632
rect 3244 8538 3284 8623
rect 3052 7951 3092 7960
rect 3916 8000 3956 8623
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 5068 8168 5108 9472
rect 5356 9512 5396 11479
rect 5452 9605 5492 11656
rect 5644 11612 5684 12496
rect 6220 12487 6260 12496
rect 6604 12536 6644 12547
rect 6604 12461 6644 12496
rect 6603 12452 6645 12461
rect 6603 12412 6604 12452
rect 6644 12412 6645 12452
rect 6603 12403 6645 12412
rect 5644 11563 5684 11572
rect 7180 11369 7220 13084
rect 8044 13074 8084 13159
rect 9196 12629 9236 13168
rect 9771 13208 9813 13217
rect 9771 13168 9772 13208
rect 9812 13168 9813 13208
rect 9771 13159 9813 13168
rect 11691 13208 11733 13217
rect 11691 13168 11692 13208
rect 11732 13168 11733 13208
rect 11691 13159 11733 13168
rect 9868 13040 9908 13049
rect 9484 13000 9868 13040
rect 8619 12620 8661 12629
rect 8619 12580 8620 12620
rect 8660 12580 8661 12620
rect 8619 12571 8661 12580
rect 9195 12620 9237 12629
rect 9195 12580 9196 12620
rect 9236 12580 9237 12620
rect 9195 12571 9237 12580
rect 9484 12620 9524 13000
rect 9868 12991 9908 13000
rect 11212 13040 11252 13049
rect 9484 12571 9524 12580
rect 9867 12620 9909 12629
rect 9867 12580 9868 12620
rect 9908 12580 9909 12620
rect 9867 12571 9909 12580
rect 7468 12536 7508 12545
rect 7179 11360 7221 11369
rect 7179 11320 7180 11360
rect 7220 11320 7221 11360
rect 7179 11311 7221 11320
rect 5451 9596 5493 9605
rect 5451 9556 5452 9596
rect 5492 9556 5493 9596
rect 5451 9547 5493 9556
rect 5356 9463 5396 9472
rect 5547 9260 5589 9269
rect 5547 9220 5548 9260
rect 5588 9220 5589 9260
rect 5547 9211 5589 9220
rect 7372 9260 7412 9269
rect 5548 9126 5588 9211
rect 7179 8840 7221 8849
rect 7179 8800 7180 8840
rect 7220 8800 7221 8840
rect 7179 8791 7221 8800
rect 5163 8756 5205 8765
rect 5163 8716 5164 8756
rect 5204 8716 5205 8756
rect 5163 8707 5205 8716
rect 5164 8672 5204 8707
rect 7180 8706 7220 8791
rect 5164 8621 5204 8632
rect 6027 8672 6069 8681
rect 6027 8632 6028 8672
rect 6068 8632 6069 8672
rect 6027 8623 6069 8632
rect 7372 8672 7412 9220
rect 7468 8681 7508 12496
rect 8620 12452 8660 12571
rect 9868 12536 9908 12571
rect 9868 12485 9908 12496
rect 10731 12536 10773 12545
rect 10731 12496 10732 12536
rect 10772 12496 10773 12536
rect 10731 12487 10773 12496
rect 8620 12403 8660 12412
rect 10732 12402 10772 12487
rect 11212 12461 11252 13000
rect 11692 12629 11732 13159
rect 11691 12620 11733 12629
rect 11691 12580 11692 12620
rect 11732 12580 11733 12620
rect 11691 12571 11733 12580
rect 11211 12452 11253 12461
rect 11211 12412 11212 12452
rect 11252 12412 11253 12452
rect 11211 12403 11253 12412
rect 8715 11360 8757 11369
rect 8715 11320 8716 11360
rect 8756 11320 8757 11360
rect 8715 11311 8757 11320
rect 8044 9512 8084 9521
rect 8044 8849 8084 9472
rect 8043 8840 8085 8849
rect 8043 8800 8044 8840
rect 8084 8800 8085 8840
rect 8043 8791 8085 8800
rect 7755 8756 7797 8765
rect 7755 8716 7756 8756
rect 7796 8716 7797 8756
rect 7755 8707 7797 8716
rect 7372 8623 7412 8632
rect 7467 8672 7509 8681
rect 7467 8632 7468 8672
rect 7508 8632 7509 8672
rect 7467 8623 7509 8632
rect 7756 8672 7796 8707
rect 6028 8538 6068 8623
rect 7756 8621 7796 8632
rect 8331 8672 8373 8681
rect 8331 8632 8332 8672
rect 8372 8632 8373 8672
rect 8331 8623 8373 8632
rect 8619 8672 8661 8681
rect 8619 8632 8620 8672
rect 8660 8632 8661 8672
rect 8619 8623 8661 8632
rect 5068 8119 5108 8128
rect 3916 7951 3956 7960
rect 2476 7867 2516 7876
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 884 4180 980 4220
rect 844 4171 884 4180
rect 651 3968 693 3977
rect 651 3928 652 3968
rect 692 3928 693 3968
rect 651 3919 693 3928
rect 652 3834 692 3919
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 843 3548 885 3557
rect 843 3508 844 3548
rect 884 3508 885 3548
rect 843 3499 885 3508
rect 844 3380 884 3499
rect 844 3331 884 3340
rect 7084 3464 7124 3473
rect 651 3212 693 3221
rect 651 3172 652 3212
rect 692 3172 693 3212
rect 651 3163 693 3172
rect 652 3078 692 3163
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 843 2708 885 2717
rect 843 2668 844 2708
rect 884 2668 885 2708
rect 843 2659 885 2668
rect 844 2574 884 2659
rect 7084 2465 7124 3424
rect 7468 3464 7508 3473
rect 7468 2801 7508 3424
rect 8332 3464 8372 8623
rect 8620 8538 8660 8623
rect 8716 8000 8756 11311
rect 11212 9521 11252 12403
rect 10059 9512 10101 9521
rect 10059 9472 10060 9512
rect 10100 9472 10101 9512
rect 10059 9463 10101 9472
rect 10636 9512 10676 9521
rect 9964 9260 10004 9269
rect 9771 8840 9813 8849
rect 9771 8800 9772 8840
rect 9812 8800 9813 8840
rect 9771 8791 9813 8800
rect 9772 8706 9812 8791
rect 9099 8672 9141 8681
rect 9099 8632 9100 8672
rect 9140 8632 9141 8672
rect 9099 8623 9141 8632
rect 9964 8672 10004 9220
rect 10060 8765 10100 9463
rect 10636 8849 10676 9472
rect 11211 9512 11253 9521
rect 11211 9472 11212 9512
rect 11252 9472 11253 9512
rect 11211 9463 11253 9472
rect 10635 8840 10677 8849
rect 10635 8800 10636 8840
rect 10676 8800 10677 8840
rect 10635 8791 10677 8800
rect 11692 8765 11732 12571
rect 11884 12452 11924 14008
rect 12172 13999 12212 14008
rect 13132 14048 13172 14057
rect 12267 13880 12309 13889
rect 12267 13840 12268 13880
rect 12308 13840 12309 13880
rect 12267 13831 12309 13840
rect 12843 13880 12885 13889
rect 12843 13840 12844 13880
rect 12884 13840 12885 13880
rect 12843 13831 12885 13840
rect 12268 13208 12308 13831
rect 12844 13746 12884 13831
rect 13132 13217 13172 14008
rect 12268 13159 12308 13168
rect 12651 13208 12693 13217
rect 12651 13168 12652 13208
rect 12692 13168 12693 13208
rect 12651 13159 12693 13168
rect 13131 13208 13173 13217
rect 13131 13168 13132 13208
rect 13172 13168 13173 13208
rect 13131 13159 13173 13168
rect 13516 13208 13556 16108
rect 13996 14048 14036 20719
rect 14572 20634 14612 20719
rect 14188 20600 14228 20609
rect 14188 20189 14228 20560
rect 14187 20180 14229 20189
rect 14187 20140 14188 20180
rect 14228 20140 14229 20180
rect 14187 20131 14229 20140
rect 14284 20096 14324 20105
rect 14284 17669 14324 20056
rect 15436 20012 15476 21568
rect 15916 21559 15956 21568
rect 21676 21608 21716 22828
rect 21676 21559 21716 21568
rect 21964 21692 22004 21701
rect 19947 21440 19989 21449
rect 19947 21400 19948 21440
rect 19988 21400 19989 21440
rect 19947 21391 19989 21400
rect 21003 21440 21045 21449
rect 21003 21400 21004 21440
rect 21044 21400 21045 21440
rect 21003 21391 21045 21400
rect 18232 21188 18600 21197
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18232 21139 18600 21148
rect 19472 20432 19840 20441
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19472 20383 19840 20392
rect 15436 19963 15476 19972
rect 18232 19676 18600 19685
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18232 19627 18600 19636
rect 19472 18920 19840 18929
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19472 18871 19840 18880
rect 19948 18752 19988 21391
rect 21004 21306 21044 21391
rect 21964 20861 22004 21652
rect 22060 21608 22100 25264
rect 22251 25264 22252 25304
rect 22292 25264 22293 25304
rect 22251 25255 22293 25264
rect 22827 25304 22869 25313
rect 22827 25264 22828 25304
rect 22868 25264 22869 25304
rect 22827 25255 22869 25264
rect 22828 25170 22868 25255
rect 22540 25136 22580 25145
rect 22540 23960 22580 25096
rect 22924 23960 22964 27616
rect 23020 24968 23060 29119
rect 23212 27749 23252 30640
rect 23308 29177 23348 31312
rect 25324 31352 25364 31361
rect 25324 30689 25364 31312
rect 25900 30848 25940 35176
rect 26284 34376 26324 35680
rect 27628 35671 27668 35680
rect 26284 33713 26324 34336
rect 26092 33704 26132 33713
rect 26092 31529 26132 33664
rect 26283 33704 26325 33713
rect 26283 33664 26284 33704
rect 26324 33664 26325 33704
rect 26283 33655 26325 33664
rect 26955 33704 26997 33713
rect 26955 33664 26956 33704
rect 26996 33664 26997 33704
rect 26955 33655 26997 33664
rect 26956 33570 26996 33655
rect 28108 33452 28148 33461
rect 27244 32873 27284 32958
rect 28108 32873 28148 33412
rect 27243 32864 27285 32873
rect 27243 32824 27244 32864
rect 27284 32824 27285 32864
rect 27243 32815 27285 32824
rect 27436 32864 27476 32873
rect 26572 32780 26612 32789
rect 27436 32780 27476 32824
rect 28107 32864 28149 32873
rect 28107 32824 28108 32864
rect 28148 32824 28149 32864
rect 28107 32815 28149 32824
rect 26476 32740 26572 32780
rect 26187 32192 26229 32201
rect 26187 32152 26188 32192
rect 26228 32152 26229 32192
rect 26187 32143 26229 32152
rect 26284 32192 26324 32201
rect 26188 32058 26228 32143
rect 26284 31604 26324 32152
rect 26284 31555 26324 31564
rect 26091 31520 26133 31529
rect 26091 31480 26092 31520
rect 26132 31480 26133 31520
rect 26091 31471 26133 31480
rect 25995 31352 26037 31361
rect 25995 31312 25996 31352
rect 26036 31312 26037 31352
rect 25995 31303 26037 31312
rect 25996 31218 26036 31303
rect 25996 30848 26036 30857
rect 25900 30808 25996 30848
rect 25996 30799 26036 30808
rect 25803 30764 25845 30773
rect 25803 30724 25804 30764
rect 25844 30724 25845 30764
rect 25803 30715 25845 30724
rect 24363 30680 24405 30689
rect 24363 30640 24364 30680
rect 24404 30640 24405 30680
rect 24363 30631 24405 30640
rect 25323 30680 25365 30689
rect 25323 30640 25324 30680
rect 25364 30640 25365 30680
rect 25323 30631 25365 30640
rect 25804 30680 25844 30715
rect 24364 30596 24404 30631
rect 25804 30629 25844 30640
rect 24364 30545 24404 30556
rect 25131 30428 25173 30437
rect 25131 30388 25132 30428
rect 25172 30388 25173 30428
rect 25131 30379 25173 30388
rect 25707 30428 25749 30437
rect 25707 30388 25708 30428
rect 25748 30388 25749 30428
rect 25707 30379 25749 30388
rect 25996 30428 26036 30437
rect 25132 30294 25172 30379
rect 25708 29840 25748 30379
rect 25708 29791 25748 29800
rect 23307 29168 23349 29177
rect 23307 29128 23308 29168
rect 23348 29128 23349 29168
rect 23307 29119 23349 29128
rect 25132 28328 25172 28337
rect 25132 27749 25172 28288
rect 23211 27740 23253 27749
rect 23211 27700 23212 27740
rect 23252 27700 23253 27740
rect 23211 27691 23253 27700
rect 23403 27740 23445 27749
rect 23403 27700 23404 27740
rect 23444 27700 23445 27740
rect 23403 27691 23445 27700
rect 25131 27740 25173 27749
rect 25131 27700 25132 27740
rect 25172 27700 25173 27740
rect 25131 27691 25173 27700
rect 23308 27656 23348 27665
rect 23308 27497 23348 27616
rect 23404 27581 23444 27691
rect 24843 27656 24885 27665
rect 24843 27616 24844 27656
rect 24884 27616 24885 27656
rect 24843 27607 24885 27616
rect 23403 27572 23445 27581
rect 23403 27532 23404 27572
rect 23444 27532 23445 27572
rect 23403 27523 23445 27532
rect 23307 27488 23349 27497
rect 23307 27448 23308 27488
rect 23348 27448 23349 27488
rect 23307 27439 23349 27448
rect 23787 26060 23829 26069
rect 23787 26020 23788 26060
rect 23828 26020 23829 26060
rect 23787 26011 23829 26020
rect 23788 25926 23828 26011
rect 23596 25892 23636 25901
rect 23211 25304 23253 25313
rect 23211 25264 23212 25304
rect 23252 25264 23253 25304
rect 23211 25255 23253 25264
rect 23596 25304 23636 25852
rect 23596 25255 23636 25264
rect 23980 25304 24020 25313
rect 23212 25170 23252 25255
rect 23308 25145 23348 25230
rect 23307 25136 23349 25145
rect 23307 25096 23308 25136
rect 23348 25096 23349 25136
rect 23307 25087 23349 25096
rect 23020 24928 23348 24968
rect 22540 23920 22676 23960
rect 22924 23920 23156 23960
rect 22348 23120 22388 23129
rect 22156 22532 22196 22541
rect 22348 22532 22388 23080
rect 22196 22492 22388 22532
rect 22156 22483 22196 22492
rect 22443 22364 22485 22373
rect 22443 22324 22444 22364
rect 22484 22324 22485 22364
rect 22443 22315 22485 22324
rect 22444 22230 22484 22315
rect 22060 21559 22100 21568
rect 22443 21608 22485 21617
rect 22443 21568 22444 21608
rect 22484 21568 22485 21608
rect 22443 21559 22485 21568
rect 22636 21608 22676 23920
rect 22731 23120 22773 23129
rect 22731 23080 22732 23120
rect 22772 23080 22773 23120
rect 22731 23071 22773 23080
rect 22732 21692 22772 23071
rect 23020 22868 23060 22877
rect 22732 21643 22772 21652
rect 22828 22828 23020 22868
rect 22828 21617 22868 22828
rect 23020 22819 23060 22828
rect 23020 22532 23060 22541
rect 23116 22532 23156 23920
rect 23060 22492 23156 22532
rect 23020 22483 23060 22492
rect 22923 22280 22965 22289
rect 22923 22240 22924 22280
rect 22964 22240 22965 22280
rect 22923 22231 22965 22240
rect 23211 22280 23253 22289
rect 23211 22240 23212 22280
rect 23252 22240 23253 22280
rect 23211 22231 23253 22240
rect 22636 21559 22676 21568
rect 22827 21608 22869 21617
rect 22827 21568 22828 21608
rect 22868 21568 22869 21608
rect 22827 21559 22869 21568
rect 22444 21474 22484 21559
rect 22828 21474 22868 21559
rect 21099 20852 21141 20861
rect 21099 20812 21100 20852
rect 21140 20812 21141 20852
rect 21099 20803 21141 20812
rect 21963 20852 22005 20861
rect 21963 20812 21964 20852
rect 22004 20812 22005 20852
rect 21963 20803 22005 20812
rect 21100 20096 21140 20803
rect 22924 20777 22964 22231
rect 23212 22146 23252 22231
rect 22923 20768 22965 20777
rect 22923 20728 22924 20768
rect 22964 20728 22965 20768
rect 22923 20719 22965 20728
rect 21100 20047 21140 20056
rect 19756 18712 19988 18752
rect 20428 19844 20468 19853
rect 19756 18668 19796 18712
rect 19756 18619 19796 18628
rect 18508 18584 18548 18593
rect 19372 18584 19412 18593
rect 18548 18544 18740 18584
rect 18508 18535 18548 18544
rect 17356 18332 17396 18341
rect 14283 17660 14325 17669
rect 14283 17620 14284 17660
rect 14324 17620 14325 17660
rect 14283 17611 14325 17620
rect 17259 17072 17301 17081
rect 17259 17032 17260 17072
rect 17300 17032 17301 17072
rect 17259 17023 17301 17032
rect 16492 16820 16532 16829
rect 16492 14720 16532 16780
rect 16492 14671 16532 14680
rect 17164 14552 17204 14561
rect 13996 13999 14036 14008
rect 14667 14048 14709 14057
rect 14667 14008 14668 14048
rect 14708 14008 14709 14048
rect 14667 13999 14709 14008
rect 15147 14048 15189 14057
rect 15147 14008 15148 14048
rect 15188 14008 15189 14048
rect 15147 13999 15189 14008
rect 15820 14048 15860 14057
rect 16012 14048 16052 14057
rect 15860 14008 16012 14048
rect 15820 13999 15860 14008
rect 16012 13999 16052 14008
rect 16395 14048 16437 14057
rect 16395 14008 16396 14048
rect 16436 14008 16437 14048
rect 16395 13999 16437 14008
rect 14668 13460 14708 13999
rect 15148 13914 15188 13999
rect 16396 13914 16436 13999
rect 14668 13411 14708 13420
rect 12652 13074 12692 13159
rect 13516 12545 13556 13168
rect 13515 12536 13557 12545
rect 13515 12496 13516 12536
rect 13556 12496 13557 12536
rect 13515 12487 13557 12496
rect 11884 12403 11924 12412
rect 17164 11705 17204 14512
rect 17260 14048 17300 17023
rect 17260 13999 17300 14008
rect 17356 13889 17396 18292
rect 18232 18164 18600 18173
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18232 18115 18600 18124
rect 18700 17753 18740 18544
rect 19276 18544 19372 18584
rect 17643 17744 17685 17753
rect 17643 17704 17644 17744
rect 17684 17704 17685 17744
rect 17643 17695 17685 17704
rect 18699 17744 18741 17753
rect 18699 17704 18700 17744
rect 18740 17704 18741 17744
rect 18699 17695 18741 17704
rect 18987 17744 19029 17753
rect 18987 17704 18988 17744
rect 19028 17704 19029 17744
rect 18987 17695 19029 17704
rect 17644 17081 17684 17695
rect 18891 17660 18933 17669
rect 18891 17620 18892 17660
rect 18932 17620 18933 17660
rect 18891 17611 18933 17620
rect 18507 17492 18549 17501
rect 18507 17452 18508 17492
rect 18548 17452 18549 17492
rect 18507 17443 18549 17452
rect 18508 17081 18548 17443
rect 18892 17156 18932 17611
rect 18988 17610 19028 17695
rect 19276 17501 19316 18544
rect 19372 18535 19412 18544
rect 19371 17744 19413 17753
rect 19371 17704 19372 17744
rect 19412 17704 19413 17744
rect 19371 17695 19413 17704
rect 19275 17492 19317 17501
rect 19275 17452 19276 17492
rect 19316 17452 19317 17492
rect 19275 17443 19317 17452
rect 18892 17107 18932 17116
rect 17643 17072 17685 17081
rect 17643 17032 17644 17072
rect 17684 17032 17685 17072
rect 17643 17023 17685 17032
rect 18123 17072 18165 17081
rect 18123 17032 18124 17072
rect 18164 17032 18165 17072
rect 18123 17023 18165 17032
rect 18507 17072 18549 17081
rect 18507 17032 18508 17072
rect 18548 17032 18549 17072
rect 18507 17023 18549 17032
rect 19180 17072 19220 17081
rect 17644 16938 17684 17023
rect 18124 14057 18164 17023
rect 18508 16938 18548 17023
rect 18232 16652 18600 16661
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18232 16603 18600 16612
rect 18232 15140 18600 15149
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18232 15091 18600 15100
rect 18891 14720 18933 14729
rect 18891 14680 18892 14720
rect 18932 14680 18933 14720
rect 18891 14671 18933 14680
rect 18123 14048 18165 14057
rect 18123 14008 18124 14048
rect 18164 14008 18165 14048
rect 18123 13999 18165 14008
rect 18603 14048 18645 14057
rect 18796 14048 18836 14057
rect 18603 14008 18604 14048
rect 18644 14008 18645 14048
rect 18603 13999 18645 14008
rect 18700 14008 18796 14048
rect 18411 13964 18453 13973
rect 18411 13924 18412 13964
rect 18452 13924 18453 13964
rect 18411 13915 18453 13924
rect 17355 13880 17397 13889
rect 17355 13840 17356 13880
rect 17396 13840 17397 13880
rect 17355 13831 17397 13840
rect 18412 13830 18452 13915
rect 18604 13914 18644 13999
rect 18700 13889 18740 14008
rect 18796 13999 18836 14008
rect 18699 13880 18741 13889
rect 18699 13840 18700 13880
rect 18740 13840 18741 13880
rect 18699 13831 18741 13840
rect 18232 13628 18600 13637
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18232 13579 18600 13588
rect 18700 13385 18740 13831
rect 18796 13796 18836 13805
rect 18699 13376 18741 13385
rect 18699 13336 18700 13376
rect 18740 13336 18741 13376
rect 18699 13327 18741 13336
rect 18700 13208 18740 13327
rect 18700 13159 18740 13168
rect 18604 13040 18644 13049
rect 17259 12536 17301 12545
rect 17259 12496 17260 12536
rect 17300 12496 17301 12536
rect 17259 12487 17301 12496
rect 18507 12536 18549 12545
rect 18507 12496 18508 12536
rect 18548 12496 18549 12536
rect 18507 12487 18549 12496
rect 18604 12536 18644 13000
rect 18796 12629 18836 13756
rect 18795 12620 18837 12629
rect 18795 12580 18796 12620
rect 18836 12580 18837 12620
rect 18795 12571 18837 12580
rect 18604 12487 18644 12496
rect 17260 11948 17300 12487
rect 18508 12402 18548 12487
rect 18795 12452 18837 12461
rect 18795 12412 18796 12452
rect 18836 12412 18837 12452
rect 18795 12403 18837 12412
rect 18796 12318 18836 12403
rect 18232 12116 18600 12125
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18232 12067 18600 12076
rect 17260 11899 17300 11908
rect 16299 11696 16341 11705
rect 16684 11696 16724 11705
rect 16299 11656 16300 11696
rect 16340 11656 16341 11696
rect 16299 11647 16341 11656
rect 16492 11656 16684 11696
rect 16012 11528 16052 11537
rect 15820 11488 16012 11528
rect 12940 10184 12980 10193
rect 12268 10016 12308 10025
rect 11884 9976 12268 10016
rect 11884 9596 11924 9976
rect 12268 9967 12308 9976
rect 11884 9547 11924 9556
rect 12267 9512 12309 9521
rect 12267 9472 12268 9512
rect 12308 9472 12309 9512
rect 12267 9463 12309 9472
rect 12268 9378 12308 9463
rect 12940 8849 12980 10144
rect 14283 10184 14325 10193
rect 14283 10144 14284 10184
rect 14324 10144 14325 10184
rect 14283 10135 14325 10144
rect 14284 9680 14324 10135
rect 14284 9631 14324 9640
rect 15820 9596 15860 11488
rect 16012 11479 16052 11488
rect 15916 11024 15956 11033
rect 15916 10184 15956 10984
rect 16011 10184 16053 10193
rect 15916 10144 16012 10184
rect 16052 10144 16053 10184
rect 16011 10135 16053 10144
rect 16300 10184 16340 11647
rect 16300 10135 16340 10144
rect 16012 10050 16052 10135
rect 16492 10100 16532 11656
rect 16684 11647 16724 11656
rect 17163 11696 17205 11705
rect 17163 11656 17164 11696
rect 17204 11656 17205 11696
rect 17163 11647 17205 11656
rect 17356 11696 17396 11705
rect 17164 11562 17204 11647
rect 17356 11276 17396 11656
rect 16588 11236 17396 11276
rect 18892 11696 18932 14671
rect 18988 14048 19028 14059
rect 18988 13973 19028 14008
rect 19083 14048 19125 14057
rect 19083 14008 19084 14048
rect 19124 14008 19125 14048
rect 19083 13999 19125 14008
rect 18987 13964 19029 13973
rect 18987 13924 18988 13964
rect 19028 13924 19029 13964
rect 18987 13915 19029 13924
rect 19084 13301 19124 13999
rect 19083 13292 19125 13301
rect 19083 13252 19084 13292
rect 19124 13252 19125 13292
rect 19083 13243 19125 13252
rect 19084 13208 19124 13243
rect 19084 13158 19124 13168
rect 16588 11192 16628 11236
rect 16588 11143 16628 11152
rect 18232 10604 18600 10613
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18232 10555 18600 10564
rect 16492 10051 16532 10060
rect 18892 9605 18932 11656
rect 18988 12284 19028 12293
rect 18988 10184 19028 12244
rect 19180 11948 19220 17032
rect 19372 16904 19412 17695
rect 20428 17669 20468 19804
rect 21963 18332 22005 18341
rect 21963 18292 21964 18332
rect 22004 18292 22005 18332
rect 21963 18283 22005 18292
rect 22827 18332 22869 18341
rect 22827 18292 22828 18332
rect 22868 18292 22869 18332
rect 22827 18283 22869 18292
rect 21388 17744 21428 17753
rect 20427 17660 20469 17669
rect 20427 17620 20428 17660
rect 20468 17620 20469 17660
rect 20427 17611 20469 17620
rect 21003 17660 21045 17669
rect 21003 17620 21004 17660
rect 21044 17620 21045 17660
rect 21003 17611 21045 17620
rect 21004 17526 21044 17611
rect 19472 17408 19840 17417
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19472 17359 19840 17368
rect 21388 17081 21428 17704
rect 21771 17660 21813 17669
rect 21771 17620 21772 17660
rect 21812 17620 21813 17660
rect 21771 17611 21813 17620
rect 21772 17240 21812 17611
rect 21867 17492 21909 17501
rect 21867 17452 21868 17492
rect 21908 17452 21909 17492
rect 21867 17443 21909 17452
rect 21772 17191 21812 17200
rect 21387 17072 21429 17081
rect 21387 17032 21388 17072
rect 21428 17032 21429 17072
rect 21387 17023 21429 17032
rect 19468 16904 19508 16913
rect 19372 16864 19468 16904
rect 19468 16855 19508 16864
rect 19472 15896 19840 15905
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19472 15847 19840 15856
rect 21868 14972 21908 17443
rect 21964 16988 22004 18283
rect 22828 18198 22868 18283
rect 22251 17744 22293 17753
rect 22251 17704 22252 17744
rect 22292 17704 22293 17744
rect 22251 17695 22293 17704
rect 22252 17610 22292 17695
rect 22731 17156 22773 17165
rect 22731 17116 22732 17156
rect 22772 17116 22773 17156
rect 22731 17107 22773 17116
rect 22732 17022 22772 17107
rect 21964 16939 22004 16948
rect 21868 14923 21908 14932
rect 21675 14888 21717 14897
rect 21675 14848 21676 14888
rect 21716 14848 21717 14888
rect 21675 14839 21717 14848
rect 21676 14720 21716 14839
rect 21676 14671 21716 14680
rect 22924 14720 22964 20719
rect 23308 19853 23348 24928
rect 23980 23129 24020 25264
rect 24844 25304 24884 27607
rect 25996 26069 26036 30388
rect 26092 30269 26132 31471
rect 26187 31352 26229 31361
rect 26187 31312 26188 31352
rect 26228 31312 26229 31352
rect 26187 31303 26229 31312
rect 26379 31352 26421 31361
rect 26476 31352 26516 32740
rect 26572 32731 26612 32740
rect 27340 32740 27476 32780
rect 28204 32780 28244 35848
rect 29068 35888 29108 35897
rect 29068 33713 29108 35848
rect 33196 35888 33236 36511
rect 34156 36426 34196 36511
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 35116 35981 35156 36511
rect 35596 36140 35636 36688
rect 35788 36679 35828 36688
rect 37132 36728 37172 36737
rect 37132 36140 37172 36688
rect 37515 36728 37557 36737
rect 37515 36688 37516 36728
rect 37556 36688 37557 36728
rect 37515 36679 37557 36688
rect 38379 36728 38421 36737
rect 38379 36688 38380 36728
rect 38420 36688 38421 36728
rect 38379 36679 38421 36688
rect 37516 36594 37556 36679
rect 38380 36594 38420 36679
rect 37420 36140 37460 36149
rect 37132 36100 37420 36140
rect 35596 36091 35636 36100
rect 37420 36091 37460 36100
rect 35115 35972 35157 35981
rect 35115 35932 35116 35972
rect 35156 35932 35157 35972
rect 35115 35923 35157 35932
rect 37131 35972 37173 35981
rect 37131 35932 37132 35972
rect 37172 35932 37173 35972
rect 37131 35923 37173 35932
rect 37612 35972 37652 35981
rect 33196 35839 33236 35848
rect 33580 35888 33620 35897
rect 33580 35225 33620 35848
rect 34444 35888 34484 35897
rect 33196 35216 33236 35225
rect 33196 34637 33236 35176
rect 33579 35216 33621 35225
rect 33579 35176 33580 35216
rect 33620 35176 33621 35216
rect 33579 35167 33621 35176
rect 34251 35216 34293 35225
rect 34251 35176 34252 35216
rect 34292 35176 34293 35216
rect 34251 35167 34293 35176
rect 34444 35216 34484 35848
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 36939 35384 36981 35393
rect 36939 35344 36940 35384
rect 36980 35344 36981 35384
rect 36939 35335 36981 35344
rect 36940 35250 36980 35335
rect 33580 35082 33620 35167
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 33195 34628 33237 34637
rect 33195 34588 33196 34628
rect 33236 34588 33237 34628
rect 33195 34579 33237 34588
rect 34155 34628 34197 34637
rect 34155 34588 34156 34628
rect 34196 34588 34197 34628
rect 34155 34579 34197 34588
rect 34156 34494 34196 34579
rect 29067 33704 29109 33713
rect 29067 33664 29068 33704
rect 29108 33664 29109 33704
rect 29067 33655 29109 33664
rect 29355 33704 29397 33713
rect 29355 33664 29356 33704
rect 29396 33664 29397 33704
rect 29355 33655 29397 33664
rect 28204 32740 28532 32780
rect 27340 32444 27380 32740
rect 26572 32404 27380 32444
rect 28108 32696 28148 32705
rect 26572 32360 26612 32404
rect 26572 32311 26612 32320
rect 28108 32276 28148 32656
rect 28108 32227 28148 32236
rect 28492 32192 28532 32740
rect 26379 31312 26380 31352
rect 26420 31312 26516 31352
rect 27051 31352 27093 31361
rect 27051 31312 27052 31352
rect 27092 31312 27093 31352
rect 26379 31303 26421 31312
rect 27051 31303 27093 31312
rect 26188 31218 26228 31303
rect 26380 31218 26420 31303
rect 26955 30764 26997 30773
rect 26955 30724 26956 30764
rect 26996 30724 26997 30764
rect 26955 30715 26997 30724
rect 26668 30680 26708 30689
rect 26091 30260 26133 30269
rect 26091 30220 26092 30260
rect 26132 30220 26133 30260
rect 26091 30211 26133 30220
rect 26092 29840 26132 30211
rect 26092 29791 26132 29800
rect 26091 29672 26133 29681
rect 26091 29632 26092 29672
rect 26132 29632 26133 29672
rect 26091 29623 26133 29632
rect 26092 28328 26132 29623
rect 26092 27665 26132 28288
rect 26284 28160 26324 28169
rect 26091 27656 26133 27665
rect 26091 27616 26092 27656
rect 26132 27616 26133 27656
rect 26091 27607 26133 27616
rect 26092 26825 26132 27607
rect 26284 27497 26324 28120
rect 26283 27488 26325 27497
rect 26283 27448 26284 27488
rect 26324 27448 26325 27488
rect 26283 27439 26325 27448
rect 26091 26816 26133 26825
rect 26091 26776 26092 26816
rect 26132 26776 26133 26816
rect 26091 26767 26133 26776
rect 25995 26060 26037 26069
rect 25995 26020 25996 26060
rect 26036 26020 26037 26060
rect 25995 26011 26037 26020
rect 26668 25565 26708 30640
rect 26956 30630 26996 30715
rect 27052 30680 27092 31303
rect 27052 30631 27092 30640
rect 27435 30680 27477 30689
rect 27435 30640 27436 30680
rect 27476 30640 27477 30680
rect 27435 30631 27477 30640
rect 27436 30546 27476 30631
rect 28492 30269 28532 32152
rect 29356 32192 29396 33655
rect 33352 33284 33720 33293
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33352 33235 33720 33244
rect 34252 32780 34292 35167
rect 34347 34460 34389 34469
rect 34347 34420 34348 34460
rect 34388 34420 34389 34460
rect 34347 34411 34389 34420
rect 34348 34326 34388 34411
rect 34252 32740 34388 32780
rect 29356 32143 29396 32152
rect 34348 32117 34388 32740
rect 34444 32201 34484 35176
rect 35788 35216 35828 35225
rect 35596 35132 35636 35141
rect 35788 35132 35828 35176
rect 36459 35216 36501 35225
rect 36459 35176 36460 35216
rect 36500 35176 36501 35216
rect 36459 35167 36501 35176
rect 36843 35216 36885 35225
rect 36843 35176 36844 35216
rect 36884 35176 36885 35216
rect 36843 35167 36885 35176
rect 37132 35216 37172 35923
rect 37612 35897 37652 35932
rect 38668 35897 38708 37192
rect 39532 36896 39572 37360
rect 39532 36847 39572 36856
rect 39628 37232 39668 37241
rect 39628 36812 39668 37192
rect 39820 37232 39860 37444
rect 40684 37400 40724 37409
rect 40012 37232 40052 37241
rect 39820 37192 40012 37232
rect 39724 36812 39764 36821
rect 39628 36772 39724 36812
rect 39724 36763 39764 36772
rect 37611 35888 37653 35897
rect 37611 35848 37612 35888
rect 37652 35848 37653 35888
rect 37611 35839 37653 35848
rect 38667 35888 38709 35897
rect 38667 35848 38668 35888
rect 38708 35848 38709 35888
rect 38667 35839 38709 35848
rect 39627 35888 39669 35897
rect 39627 35848 39628 35888
rect 39668 35848 39669 35888
rect 39627 35839 39669 35848
rect 39820 35888 39860 37192
rect 40012 37183 40052 37192
rect 40684 36905 40724 37360
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 95072 37064 95440 37073
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95072 37015 95440 37024
rect 40683 36896 40725 36905
rect 40683 36856 40684 36896
rect 40724 36856 40725 36896
rect 40683 36847 40725 36856
rect 42123 36896 42165 36905
rect 42123 36856 42124 36896
rect 42164 36856 42165 36896
rect 42123 36847 42165 36856
rect 42124 36762 42164 36847
rect 40108 36728 40148 36739
rect 40108 36653 40148 36688
rect 40971 36728 41013 36737
rect 40971 36688 40972 36728
rect 41012 36688 41013 36728
rect 40971 36679 41013 36688
rect 41547 36728 41589 36737
rect 41547 36688 41548 36728
rect 41588 36688 41589 36728
rect 41547 36679 41589 36688
rect 40107 36644 40149 36653
rect 40107 36604 40108 36644
rect 40148 36604 40149 36644
rect 40107 36595 40149 36604
rect 40683 36644 40725 36653
rect 40683 36604 40684 36644
rect 40724 36604 40725 36644
rect 40683 36595 40725 36604
rect 39820 35839 39860 35848
rect 37612 35393 37652 35839
rect 39628 35754 39668 35839
rect 39724 35804 39764 35813
rect 39724 35468 39764 35764
rect 39436 35428 39764 35468
rect 37611 35384 37653 35393
rect 37611 35344 37612 35384
rect 37652 35344 37653 35384
rect 37611 35335 37653 35344
rect 37323 35300 37365 35309
rect 37323 35260 37324 35300
rect 37364 35260 37365 35300
rect 37323 35251 37365 35260
rect 37132 35167 37172 35176
rect 37227 35216 37269 35225
rect 37227 35176 37228 35216
rect 37268 35176 37269 35216
rect 37227 35167 37269 35176
rect 37324 35216 37364 35251
rect 35636 35092 35828 35132
rect 35596 35083 35636 35092
rect 36460 34964 36500 35167
rect 36844 35082 36884 35167
rect 37228 35082 37268 35167
rect 37324 35165 37364 35176
rect 39051 35216 39093 35225
rect 39051 35176 39052 35216
rect 39092 35176 39093 35216
rect 39051 35167 39093 35176
rect 39436 35216 39476 35428
rect 39532 35300 39572 35309
rect 39572 35260 40340 35300
rect 39532 35251 39572 35260
rect 39436 35167 39476 35176
rect 39052 35082 39092 35167
rect 36460 34469 36500 34924
rect 36652 34964 36692 34973
rect 36459 34460 36501 34469
rect 36459 34420 36460 34460
rect 36500 34420 36501 34460
rect 36459 34411 36501 34420
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 36652 33209 36692 34924
rect 40300 33788 40340 35260
rect 40300 33739 40340 33748
rect 40684 33704 40724 36595
rect 40972 36594 41012 36679
rect 35499 33200 35541 33209
rect 35499 33160 35500 33200
rect 35540 33160 35541 33200
rect 35499 33151 35541 33160
rect 36651 33200 36693 33209
rect 36651 33160 36652 33200
rect 36692 33160 36693 33200
rect 36651 33151 36693 33160
rect 34592 32528 34960 32537
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34592 32479 34960 32488
rect 35500 32276 35540 33151
rect 35500 32227 35540 32236
rect 34443 32192 34485 32201
rect 34443 32152 34444 32192
rect 34484 32152 34485 32192
rect 34443 32143 34485 32152
rect 35019 32192 35061 32201
rect 35019 32152 35020 32192
rect 35060 32152 35061 32192
rect 35019 32143 35061 32152
rect 35884 32192 35924 32203
rect 34347 32108 34389 32117
rect 34347 32068 34348 32108
rect 34388 32068 34389 32108
rect 34347 32059 34389 32068
rect 30508 31940 30548 31949
rect 28875 30764 28917 30773
rect 28875 30724 28876 30764
rect 28916 30724 28917 30764
rect 28875 30715 28917 30724
rect 28491 30260 28533 30269
rect 28491 30220 28492 30260
rect 28532 30220 28533 30260
rect 28491 30211 28533 30220
rect 26956 29840 26996 29849
rect 26956 29681 26996 29800
rect 28396 29840 28436 29849
rect 26955 29672 26997 29681
rect 26955 29632 26956 29672
rect 26996 29632 26997 29672
rect 26955 29623 26997 29632
rect 28108 29672 28148 29681
rect 28396 29672 28436 29800
rect 28148 29632 28436 29672
rect 28011 29252 28053 29261
rect 28011 29212 28012 29252
rect 28052 29212 28053 29252
rect 28011 29203 28053 29212
rect 26956 28328 26996 28337
rect 28012 28328 28052 29203
rect 26996 28288 27668 28328
rect 26956 28279 26996 28288
rect 27628 28244 27668 28288
rect 28108 28328 28148 29632
rect 28491 29252 28533 29261
rect 28491 29212 28492 29252
rect 28532 29212 28533 29252
rect 28491 29203 28533 29212
rect 28492 29168 28532 29203
rect 28492 29117 28532 29128
rect 28683 29168 28725 29177
rect 28683 29128 28684 29168
rect 28724 29128 28725 29168
rect 28683 29119 28725 29128
rect 28684 29034 28724 29119
rect 28588 28916 28628 28925
rect 28628 28876 28820 28916
rect 28588 28867 28628 28876
rect 28300 28328 28340 28337
rect 28108 28288 28300 28328
rect 28012 28279 28052 28288
rect 28300 28279 28340 28288
rect 28780 28328 28820 28876
rect 28780 28279 28820 28288
rect 28876 28328 28916 30715
rect 30508 30680 30548 31900
rect 33352 31772 33720 31781
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33352 31723 33720 31732
rect 33484 31352 33524 31361
rect 32332 31184 32372 31193
rect 31083 30764 31125 30773
rect 31083 30724 31084 30764
rect 31124 30724 31125 30764
rect 31083 30715 31125 30724
rect 30604 30680 30644 30689
rect 30508 30640 30604 30680
rect 30604 30631 30644 30640
rect 30987 30680 31029 30689
rect 30987 30640 30988 30680
rect 31028 30640 31029 30680
rect 30987 30631 31029 30640
rect 30988 30546 31028 30631
rect 31084 30630 31124 30715
rect 32332 30689 32372 31144
rect 33484 30689 33524 31312
rect 34348 31352 34388 32059
rect 34348 31303 34388 31312
rect 34732 31277 34772 31362
rect 34731 31268 34773 31277
rect 34731 31228 34732 31268
rect 34772 31228 34773 31268
rect 34731 31219 34773 31228
rect 34592 31016 34960 31025
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34592 30967 34960 30976
rect 35020 30848 35060 32143
rect 35884 32117 35924 32152
rect 36747 32192 36789 32201
rect 36747 32152 36748 32192
rect 36788 32152 36789 32192
rect 36747 32143 36789 32152
rect 38380 32192 38420 32201
rect 35883 32108 35925 32117
rect 35883 32068 35884 32108
rect 35924 32068 35925 32108
rect 35883 32059 35925 32068
rect 36748 32058 36788 32143
rect 36939 31940 36981 31949
rect 36939 31900 36940 31940
rect 36980 31900 36981 31940
rect 36939 31891 36981 31900
rect 37900 31940 37940 31949
rect 36940 31352 36980 31891
rect 36940 31303 36980 31312
rect 37132 31352 37172 31361
rect 37900 31352 37940 31900
rect 38187 31940 38229 31949
rect 38187 31900 38188 31940
rect 38228 31900 38229 31940
rect 38187 31891 38229 31900
rect 38188 31806 38228 31891
rect 37996 31352 38036 31361
rect 36267 31268 36309 31277
rect 36267 31228 36268 31268
rect 36308 31228 36309 31268
rect 36267 31219 36309 31228
rect 36268 31134 36308 31219
rect 35020 30689 35060 30808
rect 37036 30848 37076 30857
rect 37132 30848 37172 31312
rect 37076 30808 37172 30848
rect 37708 31312 37996 31352
rect 37036 30799 37076 30808
rect 32331 30680 32373 30689
rect 32331 30640 32332 30680
rect 32372 30640 32373 30680
rect 32331 30631 32373 30640
rect 33483 30680 33525 30689
rect 33483 30640 33484 30680
rect 33524 30640 33525 30680
rect 33483 30631 33525 30640
rect 34155 30680 34197 30689
rect 34540 30680 34580 30689
rect 34155 30640 34156 30680
rect 34196 30640 34197 30680
rect 34155 30631 34197 30640
rect 34348 30640 34540 30680
rect 34156 30546 34196 30631
rect 29163 30260 29205 30269
rect 29163 30220 29164 30260
rect 29204 30220 29205 30260
rect 29163 30211 29205 30220
rect 33352 30260 33720 30269
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33352 30211 33720 30220
rect 29068 29672 29108 29681
rect 29068 29177 29108 29632
rect 29067 29168 29109 29177
rect 29067 29128 29068 29168
rect 29108 29128 29109 29168
rect 29067 29119 29109 29128
rect 29164 29168 29204 30211
rect 30411 29252 30453 29261
rect 30411 29212 30412 29252
rect 30452 29212 30453 29252
rect 30411 29203 30453 29212
rect 29164 29119 29204 29128
rect 30124 29168 30164 29177
rect 28876 28279 28916 28288
rect 27820 28244 27860 28253
rect 27628 28204 27820 28244
rect 27820 28195 27860 28204
rect 29068 28160 29108 28169
rect 29108 28120 29780 28160
rect 29068 28111 29108 28120
rect 29740 27656 29780 28120
rect 29740 27607 29780 27616
rect 28971 26816 29013 26825
rect 28971 26776 28972 26816
rect 29012 26776 29013 26816
rect 28971 26767 29013 26776
rect 29836 26816 29876 26825
rect 28972 26682 29012 26767
rect 27820 26648 27860 26657
rect 25995 25556 26037 25565
rect 25995 25516 25996 25556
rect 26036 25516 26037 25556
rect 25995 25507 26037 25516
rect 26667 25556 26709 25565
rect 26667 25516 26668 25556
rect 26708 25516 26709 25556
rect 26667 25507 26709 25516
rect 25996 25422 26036 25507
rect 27820 25313 27860 26608
rect 29836 26489 29876 26776
rect 29835 26480 29877 26489
rect 29835 26440 29836 26480
rect 29876 26440 29877 26480
rect 29835 26431 29877 26440
rect 30124 26237 30164 29128
rect 30412 29118 30452 29203
rect 31084 29168 31124 29179
rect 33292 29168 33332 29177
rect 31084 29093 31124 29128
rect 33196 29128 33292 29168
rect 31083 29084 31125 29093
rect 31083 29044 31084 29084
rect 31124 29044 31125 29084
rect 31083 29035 31125 29044
rect 32139 29084 32181 29093
rect 32139 29044 32140 29084
rect 32180 29044 32181 29084
rect 32139 29035 32181 29044
rect 32140 28950 32180 29035
rect 30412 27404 30452 27413
rect 30220 27364 30412 27404
rect 30220 26816 30260 27364
rect 30412 27355 30452 27364
rect 30220 26767 30260 26776
rect 32139 26816 32181 26825
rect 32139 26776 32140 26816
rect 32180 26776 32181 26816
rect 32139 26767 32181 26776
rect 32140 26682 32180 26767
rect 31467 26648 31509 26657
rect 31467 26608 31468 26648
rect 31508 26608 31509 26648
rect 31467 26599 31509 26608
rect 32043 26648 32085 26657
rect 32043 26608 32044 26648
rect 32084 26608 32085 26648
rect 32043 26599 32085 26608
rect 31468 26514 31508 26599
rect 30219 26480 30261 26489
rect 30219 26440 30220 26480
rect 30260 26440 30261 26480
rect 30219 26431 30261 26440
rect 30220 26312 30260 26431
rect 30220 26263 30260 26272
rect 29835 26228 29877 26237
rect 29835 26188 29836 26228
rect 29876 26188 29877 26228
rect 29835 26179 29877 26188
rect 30123 26228 30165 26237
rect 30123 26188 30124 26228
rect 30164 26188 30165 26228
rect 30123 26179 30165 26188
rect 29836 26144 29876 26179
rect 29836 26093 29876 26104
rect 30699 26144 30741 26153
rect 30699 26104 30700 26144
rect 30740 26104 30741 26144
rect 30699 26095 30741 26104
rect 30892 26144 30932 26153
rect 30700 26010 30740 26095
rect 30892 25565 30932 26104
rect 31275 26144 31317 26153
rect 31275 26104 31276 26144
rect 31316 26104 31317 26144
rect 31275 26095 31317 26104
rect 30891 25556 30933 25565
rect 30891 25516 30892 25556
rect 30932 25516 30933 25556
rect 30891 25507 30933 25516
rect 24844 25255 24884 25264
rect 27819 25304 27861 25313
rect 27819 25264 27820 25304
rect 27860 25264 27861 25304
rect 27819 25255 27861 25264
rect 25707 23288 25749 23297
rect 25707 23248 25708 23288
rect 25748 23248 25749 23288
rect 25707 23239 25749 23248
rect 26187 23288 26229 23297
rect 26187 23248 26188 23288
rect 26228 23248 26229 23288
rect 26187 23239 26229 23248
rect 23979 23120 24021 23129
rect 23979 23080 23980 23120
rect 24020 23080 24021 23120
rect 23979 23071 24021 23080
rect 24843 23120 24885 23129
rect 24843 23080 24844 23120
rect 24884 23080 24885 23120
rect 24843 23071 24885 23080
rect 25708 23120 25748 23239
rect 25708 23071 25748 23080
rect 26188 23120 26228 23239
rect 26188 23071 26228 23080
rect 27148 23120 27188 23129
rect 28780 23120 28820 23129
rect 23980 22289 24020 23071
rect 24844 22986 24884 23071
rect 23979 22280 24021 22289
rect 23979 22240 23980 22280
rect 24020 22240 24021 22280
rect 23979 22231 24021 22240
rect 26091 20852 26133 20861
rect 26091 20812 26092 20852
rect 26132 20812 26133 20852
rect 26091 20803 26133 20812
rect 26571 20852 26613 20861
rect 26571 20812 26572 20852
rect 26612 20812 26613 20852
rect 26571 20803 26613 20812
rect 26859 20852 26901 20861
rect 26859 20812 26860 20852
rect 26900 20812 26901 20852
rect 26859 20803 26901 20812
rect 26092 20718 26132 20803
rect 25900 20600 25940 20609
rect 25900 20189 25940 20560
rect 24939 20180 24981 20189
rect 24939 20140 24940 20180
rect 24980 20140 24981 20180
rect 24939 20131 24981 20140
rect 25899 20180 25941 20189
rect 25899 20140 25900 20180
rect 25940 20140 25941 20180
rect 25899 20131 25941 20140
rect 24940 20046 24980 20131
rect 25324 20096 25364 20105
rect 23307 19844 23349 19853
rect 23307 19804 23308 19844
rect 23348 19804 23349 19844
rect 23307 19795 23349 19804
rect 23115 17072 23157 17081
rect 23115 17032 23116 17072
rect 23156 17032 23157 17072
rect 23115 17023 23157 17032
rect 23116 14897 23156 17023
rect 23115 14888 23157 14897
rect 23115 14848 23116 14888
rect 23156 14848 23157 14888
rect 23115 14839 23157 14848
rect 23116 14754 23156 14839
rect 23308 14729 23348 19795
rect 23500 18584 23540 18593
rect 23404 17996 23444 18005
rect 23500 17996 23540 18544
rect 25132 18584 25172 18593
rect 25324 18584 25364 20056
rect 26187 20096 26229 20105
rect 26187 20056 26188 20096
rect 26228 20056 26229 20096
rect 26187 20047 26229 20056
rect 25516 18584 25556 18593
rect 25324 18544 25516 18584
rect 26188 18584 26228 20047
rect 26572 19256 26612 20803
rect 26860 20718 26900 20803
rect 26572 19207 26612 19216
rect 26764 19256 26804 19265
rect 26668 19172 26708 19181
rect 26380 18584 26420 18593
rect 26188 18544 26380 18584
rect 25132 18005 25172 18544
rect 25516 18173 25556 18544
rect 25515 18164 25557 18173
rect 25515 18124 25516 18164
rect 25556 18124 25557 18164
rect 25515 18115 25557 18124
rect 23444 17956 23540 17996
rect 25131 17996 25173 18005
rect 25131 17956 25132 17996
rect 25172 17956 25173 17996
rect 23404 17947 23444 17956
rect 25131 17947 25173 17956
rect 23979 17912 24021 17921
rect 23979 17872 23980 17912
rect 24020 17872 24021 17912
rect 23979 17863 24021 17872
rect 24651 17912 24693 17921
rect 24651 17872 24652 17912
rect 24692 17872 24693 17912
rect 24651 17863 24693 17872
rect 23980 17828 24020 17863
rect 23980 17777 24020 17788
rect 24652 17778 24692 17863
rect 25324 17744 25364 17753
rect 25132 17704 25324 17744
rect 23979 17660 24021 17669
rect 23979 17620 23980 17660
rect 24020 17620 24021 17660
rect 23979 17611 24021 17620
rect 23788 17576 23828 17585
rect 23788 17165 23828 17536
rect 23787 17156 23829 17165
rect 23787 17116 23788 17156
rect 23828 17116 23829 17156
rect 23787 17107 23829 17116
rect 23980 17072 24020 17611
rect 25132 17240 25172 17704
rect 25324 17695 25364 17704
rect 25516 17501 25556 18115
rect 25899 17996 25941 18005
rect 25899 17956 25900 17996
rect 25940 17956 25941 17996
rect 25899 17947 25941 17956
rect 25900 17862 25940 17947
rect 26091 17828 26133 17837
rect 26091 17788 26092 17828
rect 26132 17788 26133 17828
rect 26091 17779 26133 17788
rect 26092 17694 26132 17779
rect 26380 17669 26420 18544
rect 26668 18005 26708 19132
rect 26764 18593 26804 19216
rect 26956 19088 26996 19097
rect 26996 19048 27092 19088
rect 26956 19039 26996 19048
rect 26763 18584 26805 18593
rect 26763 18544 26764 18584
rect 26804 18544 26805 18584
rect 26763 18535 26805 18544
rect 27052 18080 27092 19048
rect 27148 18500 27188 23080
rect 28204 23080 28780 23120
rect 28204 22532 28244 23080
rect 28780 23071 28820 23080
rect 29451 23120 29493 23129
rect 29451 23080 29452 23120
rect 29492 23080 29493 23120
rect 29451 23071 29493 23080
rect 29643 23120 29685 23129
rect 29643 23080 29644 23120
rect 29684 23080 29685 23120
rect 29643 23071 29685 23080
rect 29452 22986 29492 23071
rect 29644 23036 29684 23071
rect 29644 22985 29684 22996
rect 29835 22868 29877 22877
rect 29835 22828 29836 22868
rect 29876 22828 29877 22868
rect 29835 22819 29877 22828
rect 30603 22868 30645 22877
rect 30603 22828 30604 22868
rect 30644 22828 30645 22868
rect 30603 22819 30645 22828
rect 29836 22734 29876 22819
rect 28204 22483 28244 22492
rect 29356 22280 29396 22289
rect 27532 20768 27572 20777
rect 27340 20728 27532 20768
rect 27340 20264 27380 20728
rect 27532 20719 27572 20728
rect 27340 20215 27380 20224
rect 29356 20105 29396 22240
rect 30219 22280 30261 22289
rect 30219 22240 30220 22280
rect 30260 22240 30261 22280
rect 30219 22231 30261 22240
rect 30604 22280 30644 22819
rect 30604 22231 30644 22240
rect 31084 22364 31124 22373
rect 30220 21617 30260 22231
rect 30892 22112 30932 22121
rect 30700 22072 30892 22112
rect 31084 22112 31124 22324
rect 31276 22289 31316 26095
rect 31851 25556 31893 25565
rect 31851 25516 31852 25556
rect 31892 25516 31893 25556
rect 31851 25507 31893 25516
rect 31852 25422 31892 25507
rect 32044 25388 32084 26599
rect 33196 26153 33236 29128
rect 33292 29119 33332 29128
rect 34156 29168 34196 29177
rect 33352 28748 33720 28757
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33352 28699 33720 28708
rect 33352 27236 33720 27245
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33352 27187 33720 27196
rect 33291 26816 33333 26825
rect 33291 26776 33292 26816
rect 33332 26776 33333 26816
rect 33291 26767 33333 26776
rect 33292 26312 33332 26767
rect 33292 26263 33332 26272
rect 34156 26237 34196 29128
rect 34155 26228 34197 26237
rect 34155 26188 34156 26228
rect 34196 26188 34197 26228
rect 34155 26179 34197 26188
rect 32139 26144 32181 26153
rect 33195 26144 33237 26153
rect 32139 26104 32140 26144
rect 32180 26104 32181 26144
rect 32139 26095 32181 26104
rect 33100 26104 33196 26144
rect 33236 26104 33237 26144
rect 32140 26010 32180 26095
rect 32044 24884 32084 25348
rect 32811 25388 32853 25397
rect 32811 25348 32812 25388
rect 32852 25348 32853 25388
rect 32811 25339 32853 25348
rect 31852 24844 32084 24884
rect 31755 24632 31797 24641
rect 31755 24592 31756 24632
rect 31796 24592 31797 24632
rect 31755 24583 31797 24592
rect 31852 24632 31892 24844
rect 32716 24800 32756 24828
rect 32812 24800 32852 25339
rect 31948 24760 32372 24800
rect 31948 24716 31988 24760
rect 31948 24667 31988 24676
rect 31852 24583 31892 24592
rect 32044 24632 32084 24641
rect 31756 23204 31796 24583
rect 31756 23155 31796 23164
rect 31659 23120 31701 23129
rect 31659 23080 31660 23120
rect 31700 23080 31701 23120
rect 31659 23071 31701 23080
rect 31852 23120 31892 23129
rect 31660 22986 31700 23071
rect 31275 22280 31317 22289
rect 31275 22240 31276 22280
rect 31316 22240 31317 22280
rect 31275 22231 31317 22240
rect 31563 22280 31605 22289
rect 31563 22240 31564 22280
rect 31604 22240 31605 22280
rect 31563 22231 31605 22240
rect 31276 22112 31316 22121
rect 31084 22072 31276 22112
rect 30700 21860 30740 22072
rect 30892 22063 30932 22072
rect 30316 21820 30740 21860
rect 30316 21692 30356 21820
rect 31276 21785 31316 22072
rect 31275 21776 31317 21785
rect 31275 21736 31276 21776
rect 31316 21736 31317 21776
rect 31275 21727 31317 21736
rect 30316 21643 30356 21652
rect 30219 21608 30261 21617
rect 30219 21568 30220 21608
rect 30260 21568 30261 21608
rect 30219 21559 30261 21568
rect 30699 21608 30741 21617
rect 30699 21568 30700 21608
rect 30740 21568 30741 21608
rect 30699 21559 30741 21568
rect 31564 21608 31604 22231
rect 31852 21785 31892 23080
rect 32044 23045 32084 24592
rect 32235 24632 32277 24641
rect 32235 24592 32236 24632
rect 32276 24592 32277 24632
rect 32332 24632 32372 24760
rect 32756 24760 32852 24800
rect 32716 24751 32756 24760
rect 33100 24716 33140 26104
rect 33195 26095 33237 26104
rect 33352 25724 33720 25733
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33352 25675 33720 25684
rect 34348 25556 34388 30640
rect 34540 30631 34580 30640
rect 35019 30680 35061 30689
rect 35019 30640 35020 30680
rect 35060 30640 35061 30680
rect 35019 30631 35061 30640
rect 36652 30680 36692 30689
rect 36692 30640 37268 30680
rect 36652 30631 36692 30640
rect 34443 30428 34485 30437
rect 34443 30388 34444 30428
rect 34484 30388 34485 30428
rect 34443 30379 34485 30388
rect 35979 30428 36021 30437
rect 35979 30388 35980 30428
rect 36020 30388 36021 30428
rect 35979 30379 36021 30388
rect 34444 29252 34484 30379
rect 35980 30294 36020 30379
rect 37228 29756 37268 30640
rect 37419 29840 37461 29849
rect 37419 29800 37420 29840
rect 37460 29800 37461 29840
rect 37419 29791 37461 29800
rect 37708 29840 37748 31312
rect 37996 31303 38036 31312
rect 37804 31184 37844 31193
rect 37804 29849 37844 31144
rect 38187 31184 38229 31193
rect 38187 31144 38188 31184
rect 38228 31144 38229 31184
rect 38187 31135 38229 31144
rect 37995 30848 38037 30857
rect 37995 30808 37996 30848
rect 38036 30808 38037 30848
rect 37995 30799 38037 30808
rect 37996 30092 38036 30799
rect 38188 30680 38228 31135
rect 38380 30857 38420 32152
rect 38475 32192 38517 32201
rect 38475 32152 38476 32192
rect 38516 32152 38517 32192
rect 38475 32143 38517 32152
rect 38476 32058 38516 32143
rect 39051 32108 39093 32117
rect 39051 32068 39052 32108
rect 39092 32068 39093 32108
rect 39051 32059 39093 32068
rect 38668 31184 38708 31193
rect 38379 30848 38421 30857
rect 38379 30808 38380 30848
rect 38420 30808 38421 30848
rect 38379 30799 38421 30808
rect 38228 30640 38420 30680
rect 38188 30631 38228 30640
rect 37996 30043 38036 30052
rect 37708 29791 37748 29800
rect 37803 29840 37845 29849
rect 37900 29840 37940 29849
rect 37803 29800 37804 29840
rect 37844 29800 37900 29840
rect 37803 29791 37845 29800
rect 37900 29791 37940 29800
rect 38091 29840 38133 29849
rect 38091 29800 38092 29840
rect 38132 29800 38133 29840
rect 38091 29791 38133 29800
rect 37228 29707 37268 29716
rect 37420 29706 37460 29791
rect 37804 29706 37844 29791
rect 38092 29706 38132 29791
rect 34592 29504 34960 29513
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34592 29455 34960 29464
rect 34540 29252 34580 29261
rect 34444 29212 34540 29252
rect 34540 29203 34580 29212
rect 34592 27992 34960 28001
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34592 27943 34960 27952
rect 37516 26816 37556 26825
rect 37131 26732 37173 26741
rect 37131 26692 37132 26732
rect 37172 26692 37173 26732
rect 37131 26683 37173 26692
rect 37132 26598 37172 26683
rect 34592 26480 34960 26489
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34592 26431 34960 26440
rect 34923 26228 34965 26237
rect 34923 26188 34924 26228
rect 34964 26188 34965 26228
rect 34923 26179 34965 26188
rect 34348 25507 34388 25516
rect 34540 26144 34580 26153
rect 34540 25397 34580 26104
rect 34924 26144 34964 26179
rect 34924 26093 34964 26104
rect 35787 26144 35829 26153
rect 35787 26104 35788 26144
rect 35828 26104 35829 26144
rect 35787 26095 35829 26104
rect 35788 26010 35828 26095
rect 37516 26069 37556 26776
rect 38380 26816 38420 30640
rect 38668 29849 38708 31144
rect 39052 30773 39092 32059
rect 40684 30773 40724 33664
rect 41548 33704 41588 36679
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 93832 36308 94200 36317
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 93832 36259 94200 36268
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 95072 35552 95440 35561
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95072 35503 95440 35512
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 93832 34796 94200 34805
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 93832 34747 94200 34756
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 95072 34040 95440 34049
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95072 33991 95440 34000
rect 41548 31436 41588 33664
rect 42699 33452 42741 33461
rect 42699 33412 42700 33452
rect 42740 33412 42741 33452
rect 42699 33403 42741 33412
rect 43371 33452 43413 33461
rect 43371 33412 43372 33452
rect 43412 33412 43413 33452
rect 43371 33403 43413 33412
rect 42700 33318 42740 33403
rect 42795 32276 42837 32285
rect 42892 32276 42932 32285
rect 42795 32236 42796 32276
rect 42836 32236 42892 32276
rect 42795 32227 42837 32236
rect 42892 32227 42932 32236
rect 42988 32192 43028 32201
rect 42988 31529 43028 32152
rect 43372 32192 43412 33403
rect 48472 33284 48840 33293
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48472 33235 48840 33244
rect 63592 33284 63960 33293
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63592 33235 63960 33244
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 93832 33284 94200 33293
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 93832 33235 94200 33244
rect 49712 32528 50080 32537
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 49712 32479 50080 32488
rect 64832 32528 65200 32537
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 64832 32479 65200 32488
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 95072 32528 95440 32537
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95072 32479 95440 32488
rect 43372 32143 43412 32152
rect 48940 32192 48980 32201
rect 48268 31940 48308 31949
rect 42315 31520 42357 31529
rect 42315 31480 42316 31520
rect 42356 31480 42357 31520
rect 42315 31471 42357 31480
rect 42987 31520 43029 31529
rect 42987 31480 42988 31520
rect 43028 31480 43029 31520
rect 48268 31520 48308 31900
rect 48472 31772 48840 31781
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48472 31723 48840 31732
rect 48940 31529 48980 32152
rect 63592 31772 63960 31781
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63592 31723 63960 31732
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 93832 31772 94200 31781
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 93832 31723 94200 31732
rect 48939 31520 48981 31529
rect 48268 31480 48500 31520
rect 42987 31471 43029 31480
rect 41548 31387 41588 31396
rect 41931 31184 41973 31193
rect 41931 31144 41932 31184
rect 41972 31144 41973 31184
rect 41931 31135 41973 31144
rect 41932 31050 41972 31135
rect 42316 30848 42356 31471
rect 46732 31436 46772 31445
rect 46636 31396 46732 31436
rect 42316 30799 42356 30808
rect 42412 31352 42452 31361
rect 39051 30764 39093 30773
rect 39051 30724 39052 30764
rect 39092 30724 39093 30764
rect 39051 30715 39093 30724
rect 40683 30764 40725 30773
rect 40683 30724 40684 30764
rect 40724 30724 40725 30764
rect 40683 30715 40725 30724
rect 41163 30764 41205 30773
rect 41163 30724 41164 30764
rect 41204 30724 41205 30764
rect 41163 30715 41205 30724
rect 39052 30680 39092 30715
rect 39052 30629 39092 30640
rect 39435 30680 39477 30689
rect 39435 30640 39436 30680
rect 39476 30640 39477 30680
rect 39435 30631 39477 30640
rect 39436 30546 39476 30631
rect 41164 30630 41204 30715
rect 42028 30680 42068 30689
rect 42028 30521 42068 30640
rect 42027 30512 42069 30521
rect 42027 30472 42028 30512
rect 42068 30472 42069 30512
rect 42027 30463 42069 30472
rect 42412 29849 42452 31312
rect 42699 30680 42741 30689
rect 42699 30640 42700 30680
rect 42740 30640 42741 30680
rect 42699 30631 42741 30640
rect 43467 30680 43509 30689
rect 43467 30640 43468 30680
rect 43508 30640 43509 30680
rect 43467 30631 43509 30640
rect 44332 30680 44372 30689
rect 38667 29840 38709 29849
rect 38667 29800 38668 29840
rect 38708 29800 38709 29840
rect 38667 29791 38709 29800
rect 42411 29840 42453 29849
rect 42411 29800 42412 29840
rect 42452 29800 42453 29840
rect 42411 29791 42453 29800
rect 41740 28328 41780 28337
rect 39531 26900 39573 26909
rect 39531 26860 39532 26900
rect 39572 26860 39573 26900
rect 39531 26851 39573 26860
rect 40395 26900 40437 26909
rect 40395 26860 40396 26900
rect 40436 26860 40437 26900
rect 40395 26851 40437 26860
rect 38380 26767 38420 26776
rect 39532 26766 39572 26851
rect 40396 26816 40436 26851
rect 40396 26765 40436 26776
rect 38187 26732 38229 26741
rect 38187 26692 38188 26732
rect 38228 26692 38229 26732
rect 38187 26683 38229 26692
rect 38188 26312 38228 26683
rect 38188 26263 38228 26272
rect 39724 26648 39764 26657
rect 39724 26069 39764 26608
rect 41740 26237 41780 28288
rect 42412 27656 42452 29791
rect 42603 29000 42645 29009
rect 42603 28960 42604 29000
rect 42644 28960 42645 29000
rect 42603 28951 42645 28960
rect 42604 28328 42644 28951
rect 42604 28279 42644 28288
rect 42508 27656 42548 27665
rect 42412 27616 42508 27656
rect 42508 27607 42548 27616
rect 41739 26228 41781 26237
rect 41739 26188 41740 26228
rect 41780 26188 41781 26228
rect 41739 26179 41781 26188
rect 41356 26144 41396 26153
rect 37515 26060 37557 26069
rect 37515 26020 37516 26060
rect 37556 26020 37557 26060
rect 37515 26011 37557 26020
rect 38379 26060 38421 26069
rect 38379 26020 38380 26060
rect 38420 26020 38421 26060
rect 38379 26011 38421 26020
rect 39723 26060 39765 26069
rect 39723 26020 39724 26060
rect 39764 26020 39765 26060
rect 39723 26011 39765 26020
rect 36939 25892 36981 25901
rect 36939 25852 36940 25892
rect 36980 25852 36981 25892
rect 36939 25843 36981 25852
rect 36940 25758 36980 25843
rect 34539 25388 34581 25397
rect 34539 25348 34540 25388
rect 34580 25348 34581 25388
rect 34539 25339 34581 25348
rect 34060 25304 34100 25313
rect 32524 24632 32564 24641
rect 32332 24592 32524 24632
rect 32235 24583 32277 24592
rect 32524 24583 32564 24592
rect 32236 24498 32276 24583
rect 32043 23036 32085 23045
rect 32043 22996 32044 23036
rect 32084 22996 32085 23036
rect 32043 22987 32085 22996
rect 32523 23036 32565 23045
rect 32523 22996 32524 23036
rect 32564 22996 32565 23036
rect 32523 22987 32565 22996
rect 32524 22902 32564 22987
rect 32332 22868 32372 22877
rect 32140 22828 32332 22868
rect 31948 22280 31988 22289
rect 32140 22280 32180 22828
rect 32332 22819 32372 22828
rect 32523 22364 32565 22373
rect 32523 22324 32524 22364
rect 32564 22324 32565 22364
rect 32523 22315 32565 22324
rect 31988 22240 32084 22280
rect 31948 22231 31988 22240
rect 31851 21776 31893 21785
rect 31851 21736 31852 21776
rect 31892 21736 31893 21776
rect 32044 21776 32084 22240
rect 32140 22231 32180 22240
rect 32524 22280 32564 22315
rect 33100 22289 33140 24676
rect 33964 25264 34060 25304
rect 33964 24632 34004 25264
rect 34060 25255 34100 25264
rect 35019 25304 35061 25313
rect 35019 25264 35020 25304
rect 35060 25264 35061 25304
rect 35019 25255 35061 25264
rect 34592 24968 34960 24977
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34592 24919 34960 24928
rect 33964 24583 34004 24592
rect 33352 24212 33720 24221
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33352 24163 33720 24172
rect 34592 23456 34960 23465
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34592 23407 34960 23416
rect 35020 23129 35060 25255
rect 36843 24380 36885 24389
rect 36843 24340 36844 24380
rect 36884 24340 36885 24380
rect 36843 24331 36885 24340
rect 36844 23792 36884 24331
rect 37516 23801 37556 26011
rect 38380 25926 38420 26011
rect 39627 25388 39669 25397
rect 39627 25348 39628 25388
rect 39668 25348 39669 25388
rect 39627 25339 39669 25348
rect 39532 25304 39572 25313
rect 39532 24809 39572 25264
rect 39628 25254 39668 25339
rect 39724 25304 39764 26011
rect 40299 25892 40341 25901
rect 40299 25852 40300 25892
rect 40340 25852 40341 25892
rect 40299 25843 40341 25852
rect 40683 25892 40725 25901
rect 40683 25852 40684 25892
rect 40724 25852 40725 25892
rect 40683 25843 40725 25852
rect 39724 25255 39764 25264
rect 40300 25304 40340 25843
rect 40300 25255 40340 25264
rect 40684 25304 40724 25843
rect 41259 25388 41301 25397
rect 41259 25348 41260 25388
rect 41300 25348 41301 25388
rect 41259 25339 41301 25348
rect 40684 25255 40724 25264
rect 41260 25304 41300 25339
rect 41260 25253 41300 25264
rect 41356 25229 41396 26104
rect 41740 26144 41780 26179
rect 41740 26094 41780 26104
rect 42604 26144 42644 26153
rect 42700 26144 42740 30631
rect 43468 30546 43508 30631
rect 43083 30512 43125 30521
rect 43083 30472 43084 30512
rect 43124 30472 43125 30512
rect 43083 30463 43125 30472
rect 43084 30092 43124 30463
rect 43084 30043 43124 30052
rect 42796 29840 42836 29849
rect 42796 29009 42836 29800
rect 43276 29672 43316 29681
rect 43180 29632 43276 29672
rect 43180 29093 43220 29632
rect 43276 29623 43316 29632
rect 43179 29084 43221 29093
rect 43179 29044 43180 29084
rect 43220 29044 43221 29084
rect 43179 29035 43221 29044
rect 42795 29000 42837 29009
rect 42795 28960 42796 29000
rect 42836 28960 42837 29000
rect 42795 28951 42837 28960
rect 42644 26104 42740 26144
rect 42604 26095 42644 26104
rect 41644 25304 41684 25313
rect 41355 25220 41397 25229
rect 41355 25180 41356 25220
rect 41396 25180 41397 25220
rect 41355 25171 41397 25180
rect 40780 25136 40820 25145
rect 37899 24800 37941 24809
rect 37899 24760 37900 24800
rect 37940 24760 37941 24800
rect 37899 24751 37941 24760
rect 38667 24800 38709 24809
rect 38667 24760 38668 24800
rect 38708 24760 38709 24800
rect 38667 24751 38709 24760
rect 38955 24800 38997 24809
rect 38955 24760 38956 24800
rect 38996 24760 38997 24800
rect 38955 24751 38997 24760
rect 39531 24800 39573 24809
rect 39531 24760 39532 24800
rect 39572 24760 39573 24800
rect 39531 24751 39573 24760
rect 37900 24548 37940 24751
rect 38668 24666 38708 24751
rect 37900 24499 37940 24508
rect 37707 24380 37749 24389
rect 37707 24340 37708 24380
rect 37748 24340 37749 24380
rect 37707 24331 37749 24340
rect 37708 24246 37748 24331
rect 36844 23743 36884 23752
rect 37227 23792 37269 23801
rect 37227 23752 37228 23792
rect 37268 23752 37269 23792
rect 37227 23743 37269 23752
rect 37515 23792 37557 23801
rect 37515 23752 37516 23792
rect 37556 23752 37557 23792
rect 37515 23743 37557 23752
rect 37803 23792 37845 23801
rect 37803 23752 37804 23792
rect 37844 23752 37845 23792
rect 37803 23743 37845 23752
rect 38091 23792 38133 23801
rect 38091 23752 38092 23792
rect 38132 23752 38133 23792
rect 38091 23743 38133 23752
rect 37228 23658 37268 23743
rect 33676 23120 33716 23129
rect 33771 23120 33813 23129
rect 33716 23080 33772 23120
rect 33812 23080 33813 23120
rect 33676 23071 33716 23080
rect 33771 23071 33813 23080
rect 34636 23120 34676 23129
rect 33196 22868 33236 22877
rect 32524 22229 32564 22240
rect 33099 22280 33141 22289
rect 33099 22240 33100 22280
rect 33140 22240 33141 22280
rect 33099 22231 33141 22240
rect 32716 21776 32756 21785
rect 32044 21736 32716 21776
rect 31851 21727 31893 21736
rect 32716 21727 32756 21736
rect 31564 21559 31604 21568
rect 30700 21474 30740 21559
rect 33196 20189 33236 22828
rect 33352 22700 33720 22709
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33352 22651 33720 22660
rect 33772 22532 33812 23071
rect 33963 23036 34005 23045
rect 33963 22996 33964 23036
rect 34004 22996 34005 23036
rect 33963 22987 34005 22996
rect 33964 22784 34004 22987
rect 33676 22492 33812 22532
rect 33868 22744 34004 22784
rect 33387 22280 33429 22289
rect 33387 22240 33388 22280
rect 33428 22240 33429 22280
rect 33387 22231 33429 22240
rect 33388 22146 33428 22231
rect 33676 21356 33716 22492
rect 33771 21776 33813 21785
rect 33771 21736 33772 21776
rect 33812 21736 33813 21776
rect 33771 21727 33813 21736
rect 33772 21642 33812 21727
rect 33868 21608 33908 22744
rect 34540 22532 34580 22541
rect 34636 22532 34676 23080
rect 35019 23120 35061 23129
rect 35019 23080 35020 23120
rect 35060 23080 35061 23120
rect 35019 23071 35061 23080
rect 37419 22868 37461 22877
rect 37419 22828 37420 22868
rect 37460 22828 37461 22868
rect 37419 22819 37461 22828
rect 34580 22492 34676 22532
rect 34540 22483 34580 22492
rect 34592 21944 34960 21953
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34592 21895 34960 21904
rect 37420 21692 37460 22819
rect 37420 21643 37460 21652
rect 33868 21559 33908 21568
rect 37804 21608 37844 23743
rect 38092 23658 38132 23743
rect 38956 23120 38996 24751
rect 39340 24632 39380 24641
rect 39244 24044 39284 24053
rect 39340 24044 39380 24592
rect 39284 24004 39380 24044
rect 39244 23995 39284 24004
rect 40780 23960 40820 25096
rect 40684 23920 40820 23960
rect 39051 23288 39093 23297
rect 39051 23248 39052 23288
rect 39092 23248 39093 23288
rect 39051 23239 39093 23248
rect 39052 23154 39092 23239
rect 38956 23071 38996 23080
rect 38763 22868 38805 22877
rect 38763 22828 38764 22868
rect 38804 22828 38805 22868
rect 38763 22819 38805 22828
rect 38764 22734 38804 22819
rect 37804 21559 37844 21568
rect 38668 21608 38708 21617
rect 34060 21356 34100 21365
rect 33676 21316 33812 21356
rect 33352 21188 33720 21197
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33352 21139 33720 21148
rect 33195 20180 33237 20189
rect 33195 20140 33196 20180
rect 33236 20140 33237 20180
rect 33195 20131 33237 20140
rect 29163 20096 29205 20105
rect 29163 20056 29164 20096
rect 29204 20056 29205 20096
rect 29163 20047 29205 20056
rect 29355 20096 29397 20105
rect 29355 20056 29356 20096
rect 29396 20056 29397 20096
rect 29355 20047 29397 20056
rect 30123 20096 30165 20105
rect 30123 20056 30124 20096
rect 30164 20056 30165 20096
rect 30123 20047 30165 20056
rect 30508 20096 30548 20105
rect 29164 19962 29204 20047
rect 30124 19962 30164 20047
rect 30411 20012 30453 20021
rect 30508 20012 30548 20056
rect 30411 19972 30412 20012
rect 30452 19972 30548 20012
rect 31468 20096 31508 20105
rect 30411 19963 30453 19972
rect 29836 19844 29876 19853
rect 27628 19256 27668 19265
rect 27532 18752 27572 18761
rect 27628 18752 27668 19216
rect 29836 18929 29876 19804
rect 30795 19844 30837 19853
rect 30795 19804 30796 19844
rect 30836 19804 30837 19844
rect 30795 19795 30837 19804
rect 30796 19710 30836 19795
rect 31468 19517 31508 20056
rect 33352 19676 33720 19685
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33352 19627 33720 19636
rect 33772 19517 33812 21316
rect 34060 20105 34100 21316
rect 34592 20432 34960 20441
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34592 20383 34960 20392
rect 34923 20180 34965 20189
rect 34923 20140 34924 20180
rect 34964 20140 34965 20180
rect 34923 20131 34965 20140
rect 34059 20096 34101 20105
rect 34059 20056 34060 20096
rect 34100 20056 34101 20096
rect 34059 20047 34101 20056
rect 31467 19508 31509 19517
rect 31467 19468 31468 19508
rect 31508 19468 31509 19508
rect 31467 19459 31509 19468
rect 33771 19508 33813 19517
rect 33771 19468 33772 19508
rect 33812 19468 33813 19508
rect 33771 19459 33813 19468
rect 34924 19256 34964 20131
rect 38668 20105 38708 21568
rect 39819 21440 39861 21449
rect 39819 21400 39820 21440
rect 39860 21400 39861 21440
rect 39819 21391 39861 21400
rect 40491 21440 40533 21449
rect 40491 21400 40492 21440
rect 40532 21400 40533 21440
rect 40491 21391 40533 21400
rect 39820 21306 39860 21391
rect 38956 20768 38996 20777
rect 36075 20096 36117 20105
rect 36075 20056 36076 20096
rect 36116 20056 36117 20096
rect 36075 20047 36117 20056
rect 36460 20096 36500 20105
rect 36076 19962 36116 20047
rect 34924 19207 34964 19216
rect 32235 19088 32277 19097
rect 32235 19048 32236 19088
rect 32276 19048 32277 19088
rect 32235 19039 32277 19048
rect 35403 19088 35445 19097
rect 35403 19048 35404 19088
rect 35444 19048 35445 19088
rect 35403 19039 35445 19048
rect 29835 18920 29877 18929
rect 29835 18880 29836 18920
rect 29876 18880 29877 18920
rect 29835 18871 29877 18880
rect 31179 18920 31221 18929
rect 31179 18880 31180 18920
rect 31220 18880 31221 18920
rect 31179 18871 31221 18880
rect 27572 18712 27668 18752
rect 27532 18703 27572 18712
rect 27148 18460 27668 18500
rect 27243 18248 27285 18257
rect 27243 18208 27244 18248
rect 27284 18208 27285 18248
rect 27243 18199 27285 18208
rect 26764 18040 27188 18080
rect 26667 17996 26709 18005
rect 26667 17956 26668 17996
rect 26708 17956 26709 17996
rect 26667 17947 26709 17956
rect 26475 17912 26517 17921
rect 26475 17872 26476 17912
rect 26516 17872 26517 17912
rect 26475 17863 26517 17872
rect 26476 17744 26516 17863
rect 26667 17828 26709 17837
rect 26764 17828 26804 18040
rect 26667 17788 26668 17828
rect 26708 17788 26804 17828
rect 27148 17828 27188 18040
rect 27148 17788 27191 17828
rect 26667 17779 26719 17788
rect 26679 17759 26719 17779
rect 26476 17695 26516 17704
rect 26571 17744 26613 17753
rect 26571 17704 26572 17744
rect 26612 17704 26613 17744
rect 26571 17695 26613 17704
rect 26379 17660 26421 17669
rect 26379 17620 26380 17660
rect 26420 17620 26421 17660
rect 26379 17611 26421 17620
rect 26572 17610 26612 17695
rect 26679 17675 26719 17719
rect 27151 17744 27191 17788
rect 27151 17695 27191 17704
rect 27052 17576 27092 17585
rect 27244 17576 27284 18199
rect 27531 17996 27573 18005
rect 27531 17956 27532 17996
rect 27572 17956 27573 17996
rect 27531 17947 27573 17956
rect 27532 17744 27572 17947
rect 27532 17695 27572 17704
rect 27092 17536 27284 17576
rect 27340 17576 27380 17585
rect 27052 17527 27092 17536
rect 25515 17492 25557 17501
rect 25515 17452 25516 17492
rect 25556 17452 25557 17492
rect 25515 17443 25557 17452
rect 25132 17191 25172 17200
rect 27340 17165 27380 17536
rect 27339 17156 27381 17165
rect 27339 17116 27340 17156
rect 27380 17116 27381 17156
rect 27339 17107 27381 17116
rect 23980 17023 24020 17032
rect 27628 15485 27668 18460
rect 30315 18164 30357 18173
rect 30315 18124 30316 18164
rect 30356 18124 30357 18164
rect 30315 18115 30357 18124
rect 30316 17753 30356 18115
rect 27819 17744 27861 17753
rect 27819 17704 27820 17744
rect 27860 17704 27861 17744
rect 27819 17695 27861 17704
rect 30315 17744 30357 17753
rect 30315 17704 30316 17744
rect 30356 17704 30357 17744
rect 30315 17695 30357 17704
rect 31180 17744 31220 18871
rect 31180 17695 31220 17704
rect 31371 17744 31413 17753
rect 31371 17704 31372 17744
rect 31412 17704 31413 17744
rect 31371 17695 31413 17704
rect 27820 17610 27860 17695
rect 28011 17660 28053 17669
rect 28011 17620 28012 17660
rect 28052 17620 28053 17660
rect 28011 17611 28053 17620
rect 29931 17660 29973 17669
rect 29931 17620 29932 17660
rect 29972 17620 29973 17660
rect 29931 17611 29973 17620
rect 28012 17526 28052 17611
rect 29932 17526 29972 17611
rect 30316 17610 30356 17695
rect 30987 17156 31029 17165
rect 30987 17116 30988 17156
rect 31028 17116 31029 17156
rect 30987 17107 31029 17116
rect 30988 17022 31028 17107
rect 31372 17072 31412 17695
rect 32236 17072 32276 19039
rect 35404 18954 35444 19039
rect 36460 18929 36500 20056
rect 37323 20096 37365 20105
rect 37323 20056 37324 20096
rect 37364 20056 37365 20096
rect 37323 20047 37365 20056
rect 38667 20096 38709 20105
rect 38667 20056 38668 20096
rect 38708 20056 38709 20096
rect 38667 20047 38709 20056
rect 36939 19508 36981 19517
rect 36939 19468 36940 19508
rect 36980 19468 36981 19508
rect 36939 19459 36981 19468
rect 34592 18920 34960 18929
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34592 18871 34960 18880
rect 36459 18920 36501 18929
rect 36459 18880 36460 18920
rect 36500 18880 36501 18920
rect 36459 18871 36501 18880
rect 33352 18164 33720 18173
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33352 18115 33720 18124
rect 32331 17828 32373 17837
rect 32331 17788 32332 17828
rect 32372 17788 32373 17828
rect 32331 17779 32373 17788
rect 32332 17694 32372 17779
rect 33867 17744 33909 17753
rect 33867 17704 33868 17744
rect 33908 17704 33909 17744
rect 33867 17695 33909 17704
rect 33580 17072 33620 17081
rect 30604 15560 30644 15569
rect 27627 15476 27669 15485
rect 27627 15436 27628 15476
rect 27668 15436 27669 15476
rect 27627 15427 27669 15436
rect 30604 15140 30644 15520
rect 30988 15560 31028 15569
rect 31372 15560 31412 17032
rect 31028 15520 31412 15560
rect 31852 17032 32236 17072
rect 31852 15560 31892 17032
rect 32236 17023 32276 17032
rect 33004 17032 33580 17072
rect 33004 15728 33044 17032
rect 33580 17023 33620 17032
rect 33868 17072 33908 17695
rect 34592 17408 34960 17417
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34592 17359 34960 17368
rect 34059 17156 34101 17165
rect 34059 17116 34060 17156
rect 34100 17116 34101 17156
rect 34059 17107 34101 17116
rect 36171 17156 36213 17165
rect 36171 17116 36172 17156
rect 36212 17116 36213 17156
rect 36171 17107 36213 17116
rect 33868 17023 33908 17032
rect 34060 17022 34100 17107
rect 33388 16829 33428 16914
rect 33387 16820 33429 16829
rect 33387 16780 33388 16820
rect 33428 16780 33429 16820
rect 33387 16771 33429 16780
rect 34923 16820 34965 16829
rect 34923 16780 34924 16820
rect 34964 16780 34965 16820
rect 34923 16771 34965 16780
rect 33352 16652 33720 16661
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33352 16603 33720 16612
rect 34924 16232 34964 16771
rect 36076 16232 36116 16241
rect 34924 16183 34964 16192
rect 35788 16192 36076 16232
rect 35596 16064 35636 16073
rect 35636 16024 35732 16064
rect 35596 16015 35636 16024
rect 34592 15896 34960 15905
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34592 15847 34960 15856
rect 33004 15679 33044 15688
rect 35692 15569 35732 16024
rect 35788 15644 35828 16192
rect 36076 16183 36116 16192
rect 36172 16232 36212 17107
rect 36364 17072 36404 17081
rect 36364 16316 36404 17032
rect 36364 16267 36404 16276
rect 36172 16183 36212 16192
rect 35788 15595 35828 15604
rect 30988 15511 31028 15520
rect 31852 15511 31892 15520
rect 35691 15560 35733 15569
rect 35691 15520 35692 15560
rect 35732 15520 35733 15560
rect 35691 15511 35733 15520
rect 35884 15560 35924 15569
rect 36076 15560 36116 15569
rect 35924 15520 36076 15560
rect 35884 15511 35924 15520
rect 36076 15511 36116 15520
rect 36267 15560 36309 15569
rect 36267 15520 36268 15560
rect 36308 15520 36309 15560
rect 36267 15511 36309 15520
rect 36748 15560 36788 15569
rect 34059 15476 34101 15485
rect 34059 15436 34060 15476
rect 34100 15436 34101 15476
rect 34059 15427 34101 15436
rect 30412 15100 30644 15140
rect 33352 15140 33720 15149
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 23500 14888 23540 14897
rect 22924 14671 22964 14680
rect 23307 14720 23349 14729
rect 23307 14680 23308 14720
rect 23348 14680 23349 14720
rect 23307 14671 23349 14680
rect 19472 14384 19840 14393
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19472 14335 19840 14344
rect 19659 14048 19701 14057
rect 19659 14008 19660 14048
rect 19700 14008 19701 14048
rect 19659 13999 19701 14008
rect 19660 13914 19700 13999
rect 20427 13376 20469 13385
rect 20427 13336 20428 13376
rect 20468 13336 20469 13376
rect 20427 13327 20469 13336
rect 23308 13376 23348 13385
rect 20235 13292 20277 13301
rect 20235 13252 20236 13292
rect 20276 13252 20277 13292
rect 20235 13243 20277 13252
rect 19371 13208 19413 13217
rect 19371 13168 19372 13208
rect 19412 13168 19413 13208
rect 19371 13159 19413 13168
rect 20236 13208 20276 13243
rect 19372 13074 19412 13159
rect 20236 13157 20276 13168
rect 20331 13208 20373 13217
rect 20331 13168 20332 13208
rect 20372 13168 20373 13208
rect 20331 13159 20373 13168
rect 20428 13208 20468 13327
rect 20428 13159 20468 13168
rect 20332 13074 20372 13159
rect 23308 13133 23348 13336
rect 23500 13217 23540 14848
rect 26572 14048 26612 14057
rect 26284 14008 26572 14048
rect 25324 13964 25364 13975
rect 25324 13889 25364 13924
rect 23883 13880 23925 13889
rect 23883 13840 23884 13880
rect 23924 13840 23925 13880
rect 23883 13831 23925 13840
rect 25131 13880 25173 13889
rect 25131 13840 25132 13880
rect 25172 13840 25173 13880
rect 25131 13831 25173 13840
rect 25323 13880 25365 13889
rect 25323 13840 25324 13880
rect 25364 13840 25365 13880
rect 25323 13831 25365 13840
rect 25899 13880 25941 13889
rect 25899 13840 25900 13880
rect 25940 13840 25941 13880
rect 25899 13831 25941 13840
rect 23499 13208 23541 13217
rect 23499 13168 23500 13208
rect 23540 13168 23541 13208
rect 23499 13159 23541 13168
rect 23884 13208 23924 13831
rect 25132 13746 25172 13831
rect 25900 13746 25940 13831
rect 26284 13460 26324 14008
rect 26572 13999 26612 14008
rect 28875 13880 28917 13889
rect 28875 13840 28876 13880
rect 28916 13840 28917 13880
rect 28875 13831 28917 13840
rect 26284 13411 26324 13420
rect 28588 13292 28628 13301
rect 23884 13159 23924 13168
rect 24267 13208 24309 13217
rect 24267 13168 24268 13208
rect 24308 13168 24309 13208
rect 24267 13159 24309 13168
rect 25132 13208 25172 13217
rect 23307 13124 23349 13133
rect 23307 13084 23308 13124
rect 23348 13084 23349 13124
rect 23307 13075 23349 13084
rect 23500 13074 23540 13159
rect 24268 13074 24308 13159
rect 20044 13040 20084 13049
rect 19472 12872 19840 12881
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19472 12823 19840 12832
rect 19947 12620 19989 12629
rect 19947 12580 19948 12620
rect 19988 12580 19989 12620
rect 19947 12571 19989 12580
rect 19660 12536 19700 12547
rect 19660 12461 19700 12496
rect 19851 12536 19893 12545
rect 19851 12496 19852 12536
rect 19892 12496 19893 12536
rect 19851 12487 19893 12496
rect 19948 12536 19988 12571
rect 19659 12452 19701 12461
rect 19659 12412 19660 12452
rect 19700 12412 19701 12452
rect 19659 12403 19701 12412
rect 19852 12402 19892 12487
rect 19948 12485 19988 12496
rect 20044 12536 20084 13000
rect 25132 12629 25172 13168
rect 28011 13124 28053 13133
rect 28011 13084 28012 13124
rect 28052 13084 28053 13124
rect 28011 13075 28053 13084
rect 27627 13040 27669 13049
rect 27627 13000 27628 13040
rect 27668 13000 27669 13040
rect 27627 12991 27669 13000
rect 25131 12620 25173 12629
rect 25131 12580 25132 12620
rect 25172 12580 25173 12620
rect 25131 12571 25173 12580
rect 27628 12620 27668 12991
rect 27628 12571 27668 12580
rect 20044 12487 20084 12496
rect 20139 12536 20181 12545
rect 20139 12496 20140 12536
rect 20180 12496 20181 12536
rect 20139 12487 20181 12496
rect 21291 12536 21333 12545
rect 21291 12496 21292 12536
rect 21332 12496 21333 12536
rect 21291 12487 21333 12496
rect 28012 12536 28052 13075
rect 28588 13049 28628 13252
rect 28876 13208 28916 13831
rect 28876 13159 28916 13168
rect 28971 13208 29013 13217
rect 28971 13168 28972 13208
rect 29012 13168 29013 13208
rect 28971 13159 29013 13168
rect 29068 13208 29108 13217
rect 28972 13074 29012 13159
rect 29068 13049 29108 13168
rect 30124 13208 30164 13217
rect 28395 13040 28437 13049
rect 28395 13000 28396 13040
rect 28436 13000 28437 13040
rect 28395 12991 28437 13000
rect 28587 13040 28629 13049
rect 28587 13000 28588 13040
rect 28628 13000 28629 13040
rect 28587 12991 28629 13000
rect 29067 13040 29109 13049
rect 29067 13000 29068 13040
rect 29108 13000 29109 13040
rect 29067 12991 29109 13000
rect 29451 13040 29493 13049
rect 29451 13000 29452 13040
rect 29492 13000 29493 13040
rect 29451 12991 29493 13000
rect 28396 12906 28436 12991
rect 29452 12906 29492 12991
rect 30028 12704 30068 12713
rect 30124 12704 30164 13168
rect 30412 13124 30452 15100
rect 33352 15091 33720 15100
rect 32523 14048 32565 14057
rect 32523 14008 32524 14048
rect 32564 14008 32565 14048
rect 32523 13999 32565 14008
rect 33675 14048 33717 14057
rect 33675 14008 33676 14048
rect 33716 14008 33717 14048
rect 33675 13999 33717 14008
rect 34060 14048 34100 15427
rect 35692 15426 35732 15511
rect 35979 15308 36021 15317
rect 35979 15268 35980 15308
rect 36020 15268 36021 15308
rect 35979 15259 36021 15268
rect 35980 14720 36020 15259
rect 36268 14720 36308 15511
rect 36748 15317 36788 15520
rect 36747 15308 36789 15317
rect 36747 15268 36748 15308
rect 36788 15268 36789 15308
rect 36747 15259 36789 15268
rect 36940 15140 36980 19459
rect 37324 19097 37364 20047
rect 38956 19853 38996 20728
rect 39628 20768 39668 20777
rect 40492 20768 40532 21391
rect 39668 20728 39956 20768
rect 39628 20719 39668 20728
rect 39820 20600 39860 20609
rect 39820 20348 39860 20560
rect 39724 20308 39860 20348
rect 39724 20096 39764 20308
rect 38475 19844 38517 19853
rect 38475 19804 38476 19844
rect 38516 19804 38517 19844
rect 38475 19795 38517 19804
rect 38955 19844 38997 19853
rect 38955 19804 38956 19844
rect 38996 19804 38997 19844
rect 38955 19795 38997 19804
rect 39339 19844 39381 19853
rect 39339 19804 39340 19844
rect 39380 19804 39381 19844
rect 39339 19795 39381 19804
rect 38476 19710 38516 19795
rect 39340 19256 39380 19795
rect 39340 19207 39380 19216
rect 39724 19256 39764 20056
rect 39819 20096 39861 20105
rect 39819 20056 39820 20096
rect 39860 20056 39861 20096
rect 39819 20047 39861 20056
rect 39916 20096 39956 20728
rect 40492 20719 40532 20728
rect 40587 20180 40629 20189
rect 40587 20140 40588 20180
rect 40628 20140 40629 20180
rect 40587 20131 40629 20140
rect 39916 20047 39956 20056
rect 40588 20096 40628 20131
rect 39820 19962 39860 20047
rect 40588 20045 40628 20056
rect 40684 20096 40724 23920
rect 41644 23885 41684 25264
rect 41739 25220 41781 25229
rect 41739 25180 41740 25220
rect 41780 25180 41781 25220
rect 41739 25171 41781 25180
rect 41740 25086 41780 25171
rect 42316 24632 42356 24641
rect 41643 23876 41685 23885
rect 41643 23836 41644 23876
rect 41684 23836 41685 23876
rect 41643 23827 41685 23836
rect 42316 23801 42356 24592
rect 43180 24464 43220 29035
rect 44332 29009 44372 30640
rect 44716 30680 44756 30689
rect 44716 29765 44756 30640
rect 46155 30680 46197 30689
rect 46155 30640 46156 30680
rect 46196 30640 46197 30680
rect 46155 30631 46197 30640
rect 45675 30596 45717 30605
rect 45675 30556 45676 30596
rect 45716 30556 45717 30596
rect 45675 30547 45717 30556
rect 45676 30092 45716 30547
rect 46156 30546 46196 30631
rect 46636 30269 46676 31396
rect 46732 31387 46772 31396
rect 47500 31352 47540 31361
rect 48364 31352 48404 31361
rect 47116 31268 47156 31277
rect 46924 31228 47116 31268
rect 46924 31184 46964 31228
rect 47116 31219 47156 31228
rect 46924 31135 46964 31144
rect 47500 30773 47540 31312
rect 48268 31312 48364 31352
rect 47499 30764 47541 30773
rect 47499 30724 47500 30764
rect 47540 30724 47541 30764
rect 47499 30715 47541 30724
rect 46731 30680 46773 30689
rect 46731 30640 46732 30680
rect 46772 30640 46773 30680
rect 46731 30631 46773 30640
rect 46635 30260 46677 30269
rect 46635 30220 46636 30260
rect 46676 30220 46677 30260
rect 46635 30211 46677 30220
rect 45676 30043 45716 30052
rect 45868 29840 45908 29849
rect 44715 29756 44757 29765
rect 44715 29716 44716 29756
rect 44756 29716 44757 29756
rect 44715 29707 44757 29716
rect 45868 29177 45908 29800
rect 46251 29840 46293 29849
rect 46251 29800 46252 29840
rect 46292 29800 46293 29840
rect 46251 29791 46293 29800
rect 46252 29706 46292 29791
rect 46636 29681 46676 30211
rect 46732 30092 46772 30631
rect 46732 30043 46772 30052
rect 47404 29840 47444 29849
rect 46924 29800 47404 29840
rect 45963 29672 46005 29681
rect 45963 29632 45964 29672
rect 46004 29632 46005 29672
rect 45963 29623 46005 29632
rect 46635 29672 46677 29681
rect 46635 29632 46636 29672
rect 46676 29632 46677 29672
rect 46635 29623 46677 29632
rect 45964 29538 46004 29623
rect 46924 29252 46964 29800
rect 47404 29791 47444 29800
rect 46924 29203 46964 29212
rect 45867 29168 45909 29177
rect 45867 29128 45868 29168
rect 45908 29128 45909 29168
rect 45867 29119 45909 29128
rect 46827 29168 46869 29177
rect 46827 29128 46828 29168
rect 46868 29128 46869 29168
rect 46827 29119 46869 29128
rect 47020 29168 47060 29177
rect 44139 29000 44181 29009
rect 44139 28960 44140 29000
rect 44180 28960 44181 29000
rect 44139 28951 44181 28960
rect 44331 29000 44373 29009
rect 44331 28960 44332 29000
rect 44372 28960 44373 29000
rect 44331 28951 44373 28960
rect 43755 27740 43797 27749
rect 43755 27700 43756 27740
rect 43796 27700 43797 27740
rect 43755 27691 43797 27700
rect 43372 27656 43412 27665
rect 43372 26153 43412 27616
rect 43756 27606 43796 27691
rect 44140 27656 44180 28951
rect 45868 28421 45908 29119
rect 46828 29034 46868 29119
rect 44907 28412 44949 28421
rect 44907 28372 44908 28412
rect 44948 28372 44949 28412
rect 44907 28363 44949 28372
rect 45675 28412 45717 28421
rect 45675 28372 45676 28412
rect 45716 28372 45717 28412
rect 45675 28363 45717 28372
rect 45867 28412 45909 28421
rect 45867 28372 45868 28412
rect 45908 28372 45909 28412
rect 45867 28363 45909 28372
rect 44908 28278 44948 28363
rect 45676 28278 45716 28363
rect 46348 28328 46388 28337
rect 46156 28288 46348 28328
rect 44716 28160 44756 28169
rect 44716 27749 44756 28120
rect 46156 27824 46196 28288
rect 46348 28279 46388 28288
rect 46156 27775 46196 27784
rect 44715 27740 44757 27749
rect 44715 27700 44716 27740
rect 44756 27700 44757 27740
rect 44715 27691 44757 27700
rect 47020 27740 47060 29128
rect 47403 29084 47445 29093
rect 47500 29084 47540 30715
rect 48268 30689 48308 31312
rect 48364 31303 48404 31312
rect 48267 30680 48309 30689
rect 48267 30640 48268 30680
rect 48308 30640 48309 30680
rect 48267 30631 48309 30640
rect 48364 30680 48404 30689
rect 48460 30680 48500 31480
rect 48939 31480 48940 31520
rect 48980 31480 48981 31520
rect 48939 31471 48981 31480
rect 49515 31520 49557 31529
rect 49515 31480 49516 31520
rect 49556 31480 49557 31520
rect 49515 31471 49557 31480
rect 49516 31386 49556 31471
rect 50956 31352 50996 31361
rect 50996 31312 51572 31352
rect 50956 31303 50996 31312
rect 50284 31184 50324 31193
rect 49712 31016 50080 31025
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 49712 30967 50080 30976
rect 48940 30848 48980 30857
rect 48980 30808 49172 30848
rect 48940 30799 48980 30808
rect 49132 30764 49172 30808
rect 49132 30715 49172 30724
rect 49515 30764 49557 30773
rect 49515 30724 49516 30764
rect 49556 30724 49557 30764
rect 49515 30715 49557 30724
rect 48404 30640 48500 30680
rect 48556 30680 48596 30691
rect 47787 30428 47829 30437
rect 47787 30388 47788 30428
rect 47828 30388 47829 30428
rect 47787 30379 47829 30388
rect 47788 29840 47828 30379
rect 48364 30269 48404 30640
rect 48556 30605 48596 30640
rect 49516 30680 49556 30715
rect 49516 30629 49556 30640
rect 50284 30605 50324 31144
rect 51532 30848 51572 31312
rect 64832 31016 65200 31025
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 64832 30967 65200 30976
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 95072 31016 95440 31025
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95072 30967 95440 30976
rect 51532 30799 51572 30808
rect 50379 30680 50421 30689
rect 50379 30640 50380 30680
rect 50420 30640 50421 30680
rect 50379 30631 50421 30640
rect 48555 30596 48597 30605
rect 48555 30556 48556 30596
rect 48596 30556 48597 30596
rect 48555 30547 48597 30556
rect 48747 30596 48789 30605
rect 48747 30556 48748 30596
rect 48788 30556 48789 30596
rect 48747 30547 48789 30556
rect 50283 30596 50325 30605
rect 50283 30556 50284 30596
rect 50324 30556 50325 30596
rect 50283 30547 50325 30556
rect 48460 30437 48500 30522
rect 48748 30462 48788 30547
rect 50380 30546 50420 30631
rect 48459 30428 48501 30437
rect 48459 30388 48460 30428
rect 48500 30388 48501 30428
rect 48459 30379 48501 30388
rect 48363 30260 48405 30269
rect 48363 30220 48364 30260
rect 48404 30220 48405 30260
rect 48363 30211 48405 30220
rect 48472 30260 48840 30269
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48472 30211 48840 30220
rect 63592 30260 63960 30269
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63592 30211 63960 30220
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 93832 30260 94200 30269
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 93832 30211 94200 30220
rect 47788 29791 47828 29800
rect 47883 29756 47925 29765
rect 47883 29716 47884 29756
rect 47924 29716 47925 29756
rect 47883 29707 47925 29716
rect 47884 29622 47924 29707
rect 49712 29504 50080 29513
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 49712 29455 50080 29464
rect 64832 29504 65200 29513
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 64832 29455 65200 29464
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 95072 29504 95440 29513
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95072 29455 95440 29464
rect 47403 29044 47404 29084
rect 47444 29044 47540 29084
rect 47403 29035 47445 29044
rect 47212 27740 47252 27749
rect 47020 27700 47212 27740
rect 44044 27068 44084 27077
rect 44140 27068 44180 27616
rect 44084 27028 44180 27068
rect 45004 27656 45044 27665
rect 44044 27019 44084 27028
rect 44428 26816 44468 26825
rect 43371 26144 43413 26153
rect 43371 26104 43372 26144
rect 43412 26104 43413 26144
rect 43371 26095 43413 26104
rect 43372 25313 43412 26095
rect 43755 25892 43797 25901
rect 43755 25852 43756 25892
rect 43796 25852 43797 25892
rect 43755 25843 43797 25852
rect 43756 25758 43796 25843
rect 43371 25304 43413 25313
rect 43371 25264 43372 25304
rect 43412 25264 43413 25304
rect 43371 25255 43413 25264
rect 43275 25220 43317 25229
rect 43275 25180 43276 25220
rect 43316 25180 43317 25220
rect 43275 25171 43317 25180
rect 43276 24632 43316 25171
rect 43276 24583 43316 24592
rect 43180 24424 43316 24464
rect 42891 23876 42933 23885
rect 42891 23836 42892 23876
rect 42932 23836 42933 23876
rect 42891 23827 42933 23836
rect 43180 23876 43220 23885
rect 42315 23792 42357 23801
rect 42315 23752 42316 23792
rect 42356 23752 42357 23792
rect 42315 23743 42357 23752
rect 42795 23792 42837 23801
rect 42795 23752 42796 23792
rect 42836 23752 42837 23792
rect 42795 23743 42837 23752
rect 42219 23456 42261 23465
rect 42219 23416 42220 23456
rect 42260 23416 42261 23456
rect 42219 23407 42261 23416
rect 42220 22364 42260 23407
rect 42316 23129 42356 23743
rect 42796 23465 42836 23743
rect 42892 23742 42932 23827
rect 42988 23792 43028 23801
rect 43180 23792 43220 23836
rect 43028 23752 43220 23792
rect 42795 23456 42837 23465
rect 42795 23416 42796 23456
rect 42836 23416 42837 23456
rect 42795 23407 42837 23416
rect 42700 23288 42740 23297
rect 42988 23288 43028 23752
rect 42740 23248 43028 23288
rect 42700 23239 42740 23248
rect 42315 23120 42357 23129
rect 42315 23080 42316 23120
rect 42356 23080 42357 23120
rect 42315 23071 42357 23080
rect 43276 23045 43316 24424
rect 44428 23960 44468 26776
rect 45004 23960 45044 27616
rect 47020 27572 47060 27700
rect 47212 27691 47252 27700
rect 47020 27523 47060 27532
rect 46828 27404 46868 27413
rect 46868 27364 47060 27404
rect 46828 27355 46868 27364
rect 47020 26816 47060 27364
rect 47020 26767 47060 26776
rect 47404 26816 47444 29035
rect 48472 28748 48840 28757
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48472 28699 48840 28708
rect 63592 28748 63960 28757
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63592 28699 63960 28708
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 93832 28748 94200 28757
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 93832 28699 94200 28708
rect 49712 27992 50080 28001
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 49712 27943 50080 27952
rect 64832 27992 65200 28001
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 64832 27943 65200 27952
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 95072 27992 95440 28001
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95072 27943 95440 27952
rect 47884 27656 47924 27665
rect 47884 27077 47924 27616
rect 48472 27236 48840 27245
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48472 27187 48840 27196
rect 63592 27236 63960 27245
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63592 27187 63960 27196
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 93832 27236 94200 27245
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 93832 27187 94200 27196
rect 47883 27068 47925 27077
rect 47883 27028 47884 27068
rect 47924 27028 47925 27068
rect 47883 27019 47925 27028
rect 49419 27068 49461 27077
rect 49419 27028 49420 27068
rect 49460 27028 49461 27068
rect 49419 27019 49461 27028
rect 49420 26934 49460 27019
rect 47404 26767 47444 26776
rect 48268 26816 48308 26825
rect 46635 26144 46677 26153
rect 46635 26104 46636 26144
rect 46676 26104 46677 26144
rect 46635 26095 46677 26104
rect 46636 26010 46676 26095
rect 46348 25892 46388 25901
rect 46348 25229 46388 25852
rect 46347 25220 46389 25229
rect 46347 25180 46348 25220
rect 46388 25180 46389 25220
rect 46347 25171 46389 25180
rect 47307 25220 47349 25229
rect 47307 25180 47308 25220
rect 47348 25180 47349 25220
rect 47307 25171 47349 25180
rect 44332 23920 44468 23960
rect 44716 23920 45044 23960
rect 43755 23792 43797 23801
rect 43755 23752 43756 23792
rect 43796 23752 43797 23792
rect 43755 23743 43797 23752
rect 43756 23658 43796 23743
rect 43371 23624 43413 23633
rect 43371 23584 43372 23624
rect 43412 23584 43413 23624
rect 43371 23575 43413 23584
rect 43372 23490 43412 23575
rect 43372 23120 43412 23129
rect 42987 23036 43029 23045
rect 42987 22996 42988 23036
rect 43028 22996 43029 23036
rect 42987 22987 43029 22996
rect 43275 23036 43317 23045
rect 43275 22996 43276 23036
rect 43316 22996 43317 23036
rect 43372 23036 43412 23080
rect 43851 23120 43893 23129
rect 43851 23080 43852 23120
rect 43892 23080 43893 23120
rect 43851 23071 43893 23080
rect 43564 23036 43604 23045
rect 43372 22996 43564 23036
rect 43275 22987 43317 22996
rect 43564 22987 43604 22996
rect 42220 22315 42260 22324
rect 42988 22280 43028 22987
rect 42988 22231 43028 22240
rect 43852 22280 43892 23071
rect 43852 22231 43892 22240
rect 42604 22196 42644 22205
rect 42412 22112 42452 22121
rect 42604 22112 42644 22156
rect 42452 22072 42644 22112
rect 42412 22063 42452 22072
rect 40684 20047 40724 20056
rect 41739 20096 41781 20105
rect 41739 20056 41740 20096
rect 41780 20056 41781 20096
rect 41739 20047 41781 20056
rect 40875 20012 40917 20021
rect 40875 19972 40876 20012
rect 40916 19972 40917 20012
rect 40875 19963 40917 19972
rect 40876 19878 40916 19963
rect 41740 19962 41780 20047
rect 39724 19207 39764 19216
rect 41068 19844 41108 19853
rect 37323 19088 37365 19097
rect 37323 19048 37324 19088
rect 37364 19048 37365 19088
rect 37323 19039 37365 19048
rect 38475 19088 38517 19097
rect 38475 19048 38476 19088
rect 38516 19048 38517 19088
rect 38475 19039 38517 19048
rect 39819 19088 39861 19097
rect 39819 19048 39820 19088
rect 39860 19048 39861 19088
rect 39819 19039 39861 19048
rect 40683 19088 40725 19097
rect 40683 19048 40684 19088
rect 40724 19048 40725 19088
rect 40683 19039 40725 19048
rect 37611 18920 37653 18929
rect 37611 18880 37612 18920
rect 37652 18880 37653 18920
rect 37611 18871 37653 18880
rect 37612 17081 37652 18871
rect 37036 17072 37076 17081
rect 37228 17072 37268 17081
rect 37076 17032 37228 17072
rect 37036 17023 37076 17032
rect 37228 17023 37268 17032
rect 37611 17072 37653 17081
rect 37611 17032 37612 17072
rect 37652 17032 37653 17072
rect 37611 17023 37653 17032
rect 38476 17072 38516 19039
rect 39820 18954 39860 19039
rect 40684 18584 40724 19039
rect 41068 18668 41108 19804
rect 41068 18619 41108 18628
rect 41452 18584 41492 18593
rect 40684 18535 40724 18544
rect 41356 18544 41452 18584
rect 40012 18332 40052 18341
rect 39627 17744 39669 17753
rect 39627 17704 39628 17744
rect 39668 17704 39669 17744
rect 39627 17695 39669 17704
rect 39628 17240 39668 17695
rect 39628 17191 39668 17200
rect 40012 17156 40052 18292
rect 41356 17165 41396 18544
rect 41452 18535 41492 18544
rect 42316 18584 42356 18593
rect 41547 17828 41589 17837
rect 41547 17788 41548 17828
rect 41588 17788 41589 17828
rect 41547 17779 41589 17788
rect 41931 17828 41973 17837
rect 41931 17788 41932 17828
rect 41972 17788 41973 17828
rect 41931 17779 41973 17788
rect 41451 17744 41493 17753
rect 41451 17704 41452 17744
rect 41492 17704 41493 17744
rect 41451 17695 41493 17704
rect 41452 17610 41492 17695
rect 40012 17107 40052 17116
rect 41355 17156 41397 17165
rect 41355 17116 41356 17156
rect 41396 17116 41397 17156
rect 41355 17107 41397 17116
rect 38476 17023 38516 17032
rect 40395 17072 40437 17081
rect 40395 17032 40396 17072
rect 40436 17032 40437 17072
rect 40395 17023 40437 17032
rect 41259 17072 41301 17081
rect 41259 17032 41260 17072
rect 41300 17032 41301 17072
rect 41259 17023 41301 17032
rect 37612 15140 37652 17023
rect 40396 16938 40436 17023
rect 41260 16938 41300 17023
rect 41356 16997 41396 17107
rect 41355 16988 41397 16997
rect 41548 16988 41588 17779
rect 41835 17744 41877 17753
rect 41835 17704 41836 17744
rect 41876 17704 41877 17744
rect 41835 17695 41877 17704
rect 41836 17610 41876 17695
rect 41932 17660 41972 17779
rect 41932 17611 41972 17620
rect 42316 17081 42356 18544
rect 43468 18332 43508 18341
rect 43468 17753 43508 18292
rect 43467 17744 43509 17753
rect 43467 17704 43468 17744
rect 43508 17704 43509 17744
rect 43467 17695 43509 17704
rect 42315 17072 42357 17081
rect 42315 17032 42316 17072
rect 42356 17032 42357 17072
rect 42315 17023 42357 17032
rect 42699 17072 42741 17081
rect 42699 17032 42700 17072
rect 42740 17032 42741 17072
rect 42699 17023 42741 17032
rect 41355 16948 41356 16988
rect 41396 16948 41397 16988
rect 41355 16939 41397 16948
rect 41452 16948 41588 16988
rect 41739 16988 41781 16997
rect 41739 16948 41740 16988
rect 41780 16948 41781 16988
rect 40876 15308 40916 15317
rect 40876 15140 40916 15268
rect 36940 15100 37076 15140
rect 37612 15100 37748 15140
rect 36020 14680 36116 14720
rect 35980 14671 36020 14680
rect 34592 14384 34960 14393
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34592 14335 34960 14344
rect 36076 14216 36116 14680
rect 36268 14671 36308 14680
rect 36460 14552 36500 14561
rect 36500 14512 36980 14552
rect 36460 14503 36500 14512
rect 36076 14167 36116 14176
rect 34060 13999 34100 14008
rect 34924 14048 34964 14057
rect 36940 14048 36980 14512
rect 34964 14008 35060 14048
rect 34924 13999 34964 14008
rect 32524 13460 32564 13999
rect 33676 13914 33716 13999
rect 33352 13628 33720 13637
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33352 13579 33720 13588
rect 32524 13411 32564 13420
rect 30507 13208 30549 13217
rect 30507 13168 30508 13208
rect 30548 13168 30549 13208
rect 30507 13159 30549 13168
rect 30892 13208 30932 13217
rect 32332 13208 32372 13217
rect 30932 13168 31316 13208
rect 30892 13159 30932 13168
rect 30412 13075 30452 13084
rect 30508 13074 30548 13159
rect 30068 12664 30164 12704
rect 30028 12655 30068 12664
rect 28875 12620 28917 12629
rect 28875 12580 28876 12620
rect 28916 12580 28917 12620
rect 28875 12571 28917 12580
rect 20140 12402 20180 12487
rect 21292 12402 21332 12487
rect 21963 12284 22005 12293
rect 21963 12244 21964 12284
rect 22004 12244 22005 12284
rect 21963 12235 22005 12244
rect 23019 12284 23061 12293
rect 23019 12244 23020 12284
rect 23060 12244 23061 12284
rect 23019 12235 23061 12244
rect 21964 12150 22004 12235
rect 19180 11899 19220 11908
rect 19372 11528 19412 11537
rect 18988 10135 19028 10144
rect 19276 11488 19372 11528
rect 15916 9596 15956 9605
rect 15820 9556 15916 9596
rect 15916 9547 15956 9556
rect 18891 9596 18933 9605
rect 18891 9556 18892 9596
rect 18932 9556 18933 9596
rect 18891 9547 18933 9556
rect 13131 9512 13173 9521
rect 13131 9472 13132 9512
rect 13172 9472 13173 9512
rect 13131 9463 13173 9472
rect 16300 9512 16340 9521
rect 13132 9378 13172 9463
rect 12363 8840 12405 8849
rect 12363 8800 12364 8840
rect 12404 8800 12405 8840
rect 12363 8791 12405 8800
rect 12939 8840 12981 8849
rect 12939 8800 12940 8840
rect 12980 8800 12981 8840
rect 12939 8791 12981 8800
rect 10059 8756 10101 8765
rect 10059 8716 10060 8756
rect 10100 8716 10101 8756
rect 10059 8707 10101 8716
rect 10347 8756 10389 8765
rect 10347 8716 10348 8756
rect 10388 8716 10389 8756
rect 10347 8707 10389 8716
rect 11691 8756 11733 8765
rect 11691 8716 11692 8756
rect 11732 8716 11828 8756
rect 11691 8707 11733 8716
rect 9964 8623 10004 8632
rect 10348 8672 10388 8707
rect 9100 8168 9140 8623
rect 10348 8621 10388 8632
rect 11211 8672 11253 8681
rect 11211 8632 11212 8672
rect 11252 8632 11253 8672
rect 11211 8623 11253 8632
rect 11212 8538 11252 8623
rect 9100 8119 9140 8128
rect 8716 7951 8756 7960
rect 10924 7160 10964 7169
rect 10924 6320 10964 7120
rect 11788 7160 11828 8716
rect 12364 8706 12404 8791
rect 16300 7253 16340 9472
rect 17163 9512 17205 9521
rect 17163 9472 17164 9512
rect 17204 9472 17205 9512
rect 17163 9463 17205 9472
rect 17164 8849 17204 9463
rect 18892 9428 18932 9437
rect 18316 9260 18356 9269
rect 18356 9220 18836 9260
rect 18316 9211 18356 9220
rect 18232 9092 18600 9101
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18232 9043 18600 9052
rect 17163 8840 17205 8849
rect 17163 8800 17164 8840
rect 17204 8800 17205 8840
rect 17163 8791 17205 8800
rect 17451 8840 17493 8849
rect 17451 8800 17452 8840
rect 17492 8800 17493 8840
rect 17451 8791 17493 8800
rect 16107 7244 16149 7253
rect 16107 7204 16108 7244
rect 16148 7204 16149 7244
rect 16107 7195 16149 7204
rect 16299 7244 16341 7253
rect 16299 7204 16300 7244
rect 16340 7204 16341 7244
rect 16299 7195 16341 7204
rect 16587 7244 16629 7253
rect 16587 7204 16588 7244
rect 16628 7204 16629 7244
rect 16587 7195 16629 7204
rect 11788 7111 11828 7120
rect 10732 6280 10964 6320
rect 8372 3424 8564 3464
rect 8332 3415 8372 3424
rect 7467 2792 7509 2801
rect 7467 2752 7468 2792
rect 7508 2752 7509 2792
rect 7467 2743 7509 2752
rect 7659 2792 7701 2801
rect 7659 2752 7660 2792
rect 7700 2752 7701 2792
rect 7659 2743 7701 2752
rect 7660 2624 7700 2743
rect 7660 2575 7700 2584
rect 8524 2624 8564 3424
rect 9484 3212 9524 3221
rect 9524 3172 9620 3212
rect 9484 3163 9524 3172
rect 8524 2575 8564 2584
rect 7276 2540 7316 2549
rect 652 2456 692 2465
rect 652 2297 692 2416
rect 7083 2456 7125 2465
rect 7083 2416 7084 2456
rect 7124 2416 7125 2456
rect 7083 2407 7125 2416
rect 651 2288 693 2297
rect 651 2248 652 2288
rect 692 2248 693 2288
rect 651 2239 693 2248
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 7276 2129 7316 2500
rect 8427 2540 8469 2549
rect 8427 2500 8428 2540
rect 8468 2500 8469 2540
rect 8427 2491 8469 2500
rect 7851 2456 7893 2465
rect 7851 2416 7852 2456
rect 7892 2416 7893 2456
rect 7851 2407 7893 2416
rect 7275 2120 7317 2129
rect 7275 2080 7276 2120
rect 7316 2080 7317 2120
rect 7275 2071 7317 2080
rect 7852 2120 7892 2407
rect 7852 2071 7892 2080
rect 8235 2120 8277 2129
rect 8235 2080 8236 2120
rect 8276 2080 8277 2120
rect 8235 2071 8277 2080
rect 8043 2036 8085 2045
rect 8043 1996 8044 2036
rect 8084 1996 8085 2036
rect 8043 1987 8085 1996
rect 8044 1868 8084 1987
rect 8236 1986 8276 2071
rect 8044 1819 8084 1828
rect 8428 1868 8468 2491
rect 8907 2120 8949 2129
rect 8907 2080 8908 2120
rect 8948 2080 8949 2120
rect 8907 2071 8949 2080
rect 8908 1986 8948 2071
rect 9580 1952 9620 3172
rect 10732 2801 10772 6280
rect 13036 5648 13076 5657
rect 15148 5648 15188 5657
rect 13076 5608 13652 5648
rect 13036 5599 13076 5608
rect 12364 5480 12404 5489
rect 11500 4976 11540 4985
rect 11883 4976 11925 4985
rect 11540 4936 11828 4976
rect 11500 4927 11540 4936
rect 10828 4220 10868 4229
rect 10828 3473 10868 4180
rect 11595 4136 11637 4145
rect 11595 4096 11596 4136
rect 11636 4096 11637 4136
rect 11595 4087 11637 4096
rect 11212 4052 11252 4061
rect 11020 4012 11212 4052
rect 11020 3968 11060 4012
rect 11212 4003 11252 4012
rect 11596 4002 11636 4087
rect 11020 3919 11060 3928
rect 11788 3632 11828 4936
rect 11883 4936 11884 4976
rect 11924 4936 11925 4976
rect 11883 4927 11925 4936
rect 11884 4145 11924 4927
rect 11883 4136 11925 4145
rect 11883 4096 11884 4136
rect 11924 4096 11925 4136
rect 11883 4087 11925 4096
rect 11788 3583 11828 3592
rect 12364 3632 12404 5440
rect 12748 4976 12788 4985
rect 12460 4136 12500 4145
rect 12748 4136 12788 4936
rect 13612 4388 13652 5608
rect 13900 4724 13940 4733
rect 13612 4339 13652 4348
rect 13708 4684 13900 4724
rect 12500 4096 12788 4136
rect 12460 4087 12500 4096
rect 12556 3632 12596 3641
rect 12364 3592 12556 3632
rect 11499 3548 11541 3557
rect 11499 3508 11500 3548
rect 11540 3508 11541 3548
rect 11499 3499 11541 3508
rect 11979 3548 12021 3557
rect 11979 3508 11980 3548
rect 12020 3508 12021 3548
rect 11979 3499 12021 3508
rect 10827 3464 10869 3473
rect 10827 3424 10828 3464
rect 10868 3424 10869 3464
rect 10827 3415 10869 3424
rect 10924 3464 10964 3473
rect 10731 2792 10773 2801
rect 10731 2752 10732 2792
rect 10772 2752 10773 2792
rect 10731 2743 10773 2752
rect 9676 2708 9716 2717
rect 9716 2668 9908 2708
rect 9676 2659 9716 2668
rect 9868 2624 9908 2668
rect 9868 2575 9908 2584
rect 10924 2549 10964 3424
rect 11115 3464 11157 3473
rect 11115 3424 11116 3464
rect 11156 3424 11157 3464
rect 11115 3415 11157 3424
rect 11308 3464 11348 3473
rect 11116 3330 11156 3415
rect 11020 3212 11060 3221
rect 11020 2633 11060 3172
rect 11019 2624 11061 2633
rect 11019 2584 11020 2624
rect 11060 2584 11061 2624
rect 11019 2575 11061 2584
rect 10539 2540 10581 2549
rect 10539 2500 10540 2540
rect 10580 2500 10581 2540
rect 10539 2491 10581 2500
rect 10923 2540 10965 2549
rect 10923 2500 10924 2540
rect 10964 2500 10965 2540
rect 10923 2491 10965 2500
rect 10540 2406 10580 2491
rect 11308 2129 11348 3424
rect 11500 3464 11540 3499
rect 11500 3413 11540 3424
rect 11980 3380 12020 3499
rect 12364 3473 12404 3592
rect 12556 3583 12596 3592
rect 12651 3548 12693 3557
rect 12651 3508 12652 3548
rect 12692 3508 12693 3548
rect 12651 3499 12693 3508
rect 12363 3464 12405 3473
rect 12363 3424 12364 3464
rect 12404 3424 12405 3464
rect 12363 3415 12405 3424
rect 12652 3464 12692 3499
rect 12748 3473 12788 4096
rect 13035 3548 13077 3557
rect 13035 3508 13036 3548
rect 13076 3508 13077 3548
rect 13035 3499 13077 3508
rect 12652 3413 12692 3424
rect 12747 3464 12789 3473
rect 12747 3424 12748 3464
rect 12788 3424 12789 3464
rect 12747 3415 12789 3424
rect 13036 3414 13076 3499
rect 13708 3464 13748 4684
rect 13900 4675 13940 4684
rect 13708 3415 13748 3424
rect 11980 3331 12020 3340
rect 11404 3212 11444 3221
rect 12844 3212 12884 3221
rect 11444 3172 11732 3212
rect 11404 3163 11444 3172
rect 11692 2876 11732 3172
rect 11692 2836 12020 2876
rect 11691 2624 11733 2633
rect 11691 2584 11692 2624
rect 11732 2584 11733 2624
rect 11691 2575 11733 2584
rect 11980 2624 12020 2836
rect 12844 2633 12884 3172
rect 15148 2801 15188 5608
rect 16108 5648 16148 7195
rect 16203 7160 16245 7169
rect 16203 7120 16204 7160
rect 16244 7120 16245 7160
rect 16203 7111 16245 7120
rect 16588 7160 16628 7195
rect 16204 7026 16244 7111
rect 16588 7109 16628 7120
rect 17452 7160 17492 8791
rect 18796 8681 18836 9220
rect 18795 8672 18837 8681
rect 18795 8632 18796 8672
rect 18836 8632 18837 8672
rect 18795 8623 18837 8632
rect 18700 8084 18740 8093
rect 17452 7111 17492 7120
rect 17932 8044 18700 8084
rect 16108 5599 16148 5608
rect 17260 5564 17300 5573
rect 15628 5480 15668 5489
rect 15628 4985 15668 5440
rect 15627 4976 15669 4985
rect 15627 4936 15628 4976
rect 15668 4936 15669 4976
rect 15627 4927 15669 4936
rect 17260 3473 17300 5524
rect 15339 3464 15381 3473
rect 15339 3424 15340 3464
rect 15380 3424 15381 3464
rect 15339 3415 15381 3424
rect 17259 3464 17301 3473
rect 17259 3424 17260 3464
rect 17300 3424 17301 3464
rect 17259 3415 17301 3424
rect 17644 3464 17684 3473
rect 14475 2792 14517 2801
rect 14475 2752 14476 2792
rect 14516 2752 14517 2792
rect 14475 2743 14517 2752
rect 15147 2792 15189 2801
rect 15147 2752 15148 2792
rect 15188 2752 15189 2792
rect 15147 2743 15189 2752
rect 11980 2575 12020 2584
rect 12843 2624 12885 2633
rect 12843 2584 12844 2624
rect 12884 2584 12885 2624
rect 12843 2575 12885 2584
rect 14091 2624 14133 2633
rect 14091 2584 14092 2624
rect 14132 2584 14133 2624
rect 14091 2575 14133 2584
rect 14476 2624 14516 2743
rect 14476 2575 14516 2584
rect 15340 2624 15380 3415
rect 17644 2717 17684 3424
rect 17835 2876 17877 2885
rect 17835 2836 17836 2876
rect 17876 2836 17877 2876
rect 17835 2827 17877 2836
rect 17643 2708 17685 2717
rect 17643 2668 17644 2708
rect 17684 2668 17685 2708
rect 17643 2659 17685 2668
rect 15340 2575 15380 2584
rect 17836 2624 17876 2827
rect 17932 2801 17972 8044
rect 18700 8035 18740 8044
rect 18796 8000 18836 8623
rect 18796 7951 18836 7960
rect 18699 7916 18741 7925
rect 18699 7876 18700 7916
rect 18740 7876 18741 7916
rect 18699 7867 18741 7876
rect 18232 7580 18600 7589
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18232 7531 18600 7540
rect 18604 7412 18644 7421
rect 18700 7412 18740 7867
rect 18644 7372 18740 7412
rect 18604 7363 18644 7372
rect 18892 6245 18932 9388
rect 19179 8840 19221 8849
rect 19179 8800 19180 8840
rect 19220 8800 19221 8840
rect 19179 8791 19221 8800
rect 19180 8706 19220 8791
rect 19276 8672 19316 11488
rect 19372 11479 19412 11488
rect 19472 11360 19840 11369
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19472 11311 19840 11320
rect 23020 11108 23060 12235
rect 28012 11705 28052 12496
rect 28876 12536 28916 12571
rect 28876 12485 28916 12496
rect 31179 12452 31221 12461
rect 31179 12412 31180 12452
rect 31220 12412 31221 12452
rect 31179 12403 31221 12412
rect 28011 11696 28053 11705
rect 28011 11656 28012 11696
rect 28052 11656 28053 11696
rect 28011 11647 28053 11656
rect 28299 11696 28341 11705
rect 28299 11656 28300 11696
rect 28340 11656 28341 11696
rect 28299 11647 28341 11656
rect 31180 11696 31220 12403
rect 31276 11948 31316 13168
rect 32332 13049 32372 13168
rect 32236 13040 32276 13049
rect 32236 12461 32276 13000
rect 32331 13040 32373 13049
rect 32331 13000 32332 13040
rect 32372 13000 32373 13040
rect 32331 12991 32373 13000
rect 34592 12872 34960 12881
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34592 12823 34960 12832
rect 35020 12629 35060 14008
rect 36940 13999 36980 14008
rect 32619 12620 32661 12629
rect 32619 12580 32620 12620
rect 32660 12580 32661 12620
rect 32619 12571 32661 12580
rect 35019 12620 35061 12629
rect 35019 12580 35020 12620
rect 35060 12580 35061 12620
rect 35019 12571 35061 12580
rect 32620 12486 32660 12571
rect 33483 12536 33525 12545
rect 33483 12496 33484 12536
rect 33524 12496 33525 12536
rect 33483 12487 33525 12496
rect 34444 12536 34484 12545
rect 32235 12452 32277 12461
rect 32235 12412 32236 12452
rect 32276 12412 32277 12452
rect 32235 12403 32277 12412
rect 32236 12318 32276 12403
rect 33484 12402 33524 12487
rect 33771 12452 33813 12461
rect 33771 12412 33772 12452
rect 33812 12412 33813 12452
rect 33771 12403 33813 12412
rect 33772 12318 33812 12403
rect 32044 12284 32084 12293
rect 31276 11899 31316 11908
rect 31564 12244 32044 12284
rect 31180 11647 31220 11656
rect 31372 11696 31412 11705
rect 23020 11059 23060 11068
rect 19371 11024 19413 11033
rect 19371 10984 19372 11024
rect 19412 10984 19413 11024
rect 19371 10975 19413 10984
rect 23403 11024 23445 11033
rect 23403 10984 23404 11024
rect 23444 10984 23445 11024
rect 23403 10975 23445 10984
rect 24268 11024 24308 11033
rect 19372 10184 19412 10975
rect 19372 10135 19412 10144
rect 20235 10184 20277 10193
rect 20235 10144 20236 10184
rect 20276 10144 20277 10184
rect 20235 10135 20277 10144
rect 19472 9848 19840 9857
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19472 9799 19840 9808
rect 19659 9596 19701 9605
rect 19659 9556 19660 9596
rect 19700 9556 19701 9596
rect 19659 9547 19701 9556
rect 19660 9512 19700 9547
rect 19660 9461 19700 9472
rect 20236 8849 20276 10135
rect 21388 10016 21428 10025
rect 21100 9976 21388 10016
rect 20235 8840 20277 8849
rect 20235 8800 20236 8840
rect 20276 8800 20277 8840
rect 20235 8791 20277 8800
rect 19372 8672 19412 8681
rect 19276 8632 19372 8672
rect 19372 8623 19412 8632
rect 19755 8672 19797 8681
rect 19755 8632 19756 8672
rect 19796 8632 19797 8672
rect 19755 8623 19797 8632
rect 19756 8538 19796 8623
rect 19852 8597 19892 8682
rect 21100 8681 21140 9976
rect 21388 9967 21428 9976
rect 22251 8756 22293 8765
rect 22251 8716 22252 8756
rect 22292 8716 22293 8756
rect 22251 8707 22293 8716
rect 19948 8672 19988 8681
rect 19851 8588 19893 8597
rect 19851 8548 19852 8588
rect 19892 8548 19893 8588
rect 19851 8539 19893 8548
rect 19472 8336 19840 8345
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19472 8287 19840 8296
rect 19180 8000 19220 8011
rect 19180 7925 19220 7960
rect 19948 7925 19988 8632
rect 20331 8672 20373 8681
rect 20331 8632 20332 8672
rect 20372 8632 20373 8672
rect 20331 8623 20373 8632
rect 20907 8672 20949 8681
rect 20907 8632 20908 8672
rect 20948 8632 20949 8672
rect 20907 8623 20949 8632
rect 21099 8672 21141 8681
rect 21099 8632 21100 8672
rect 21140 8632 21141 8672
rect 21099 8623 21141 8632
rect 21580 8672 21620 8683
rect 19179 7916 19221 7925
rect 19179 7876 19180 7916
rect 19220 7876 19221 7916
rect 19179 7867 19221 7876
rect 19947 7916 19989 7925
rect 19947 7876 19948 7916
rect 19988 7876 19989 7916
rect 19947 7867 19989 7876
rect 20332 7412 20372 8623
rect 20908 8538 20948 8623
rect 21100 8538 21140 8623
rect 21580 8597 21620 8632
rect 21676 8672 21716 8681
rect 22059 8672 22101 8681
rect 21716 8632 21908 8672
rect 21676 8623 21716 8632
rect 21579 8588 21621 8597
rect 21579 8548 21580 8588
rect 21620 8548 21621 8588
rect 21579 8539 21621 8548
rect 21003 8504 21045 8513
rect 21292 8504 21332 8513
rect 21003 8464 21004 8504
rect 21044 8464 21045 8504
rect 21003 8455 21045 8464
rect 21196 8464 21292 8504
rect 21004 8370 21044 8455
rect 20332 7363 20372 7372
rect 19472 6824 19840 6833
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19472 6775 19840 6784
rect 18123 6236 18165 6245
rect 18123 6196 18124 6236
rect 18164 6196 18165 6236
rect 18123 6187 18165 6196
rect 18891 6236 18933 6245
rect 18891 6196 18892 6236
rect 18932 6196 18933 6236
rect 18891 6187 18933 6196
rect 18124 5648 18164 6187
rect 18232 6068 18600 6077
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18232 6019 18600 6028
rect 18124 5599 18164 5608
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 21196 4220 21236 8464
rect 21292 8455 21332 8464
rect 21868 8168 21908 8632
rect 22059 8632 22060 8672
rect 22100 8632 22101 8672
rect 22059 8623 22101 8632
rect 22252 8672 22292 8707
rect 21868 8119 21908 8128
rect 22060 8000 22100 8623
rect 22156 8588 22196 8597
rect 22156 8009 22196 8548
rect 22060 7951 22100 7960
rect 22155 8000 22197 8009
rect 22155 7960 22156 8000
rect 22196 7960 22197 8000
rect 22252 8000 22292 8632
rect 22923 8588 22965 8597
rect 22923 8548 22924 8588
rect 22964 8548 22965 8588
rect 22923 8539 22965 8548
rect 22348 8000 22388 8009
rect 22252 7960 22348 8000
rect 22155 7951 22197 7960
rect 22348 7951 22388 7960
rect 22924 8000 22964 8539
rect 23019 8504 23061 8513
rect 23019 8464 23020 8504
rect 23060 8464 23061 8504
rect 23019 8455 23061 8464
rect 22924 7951 22964 7960
rect 23020 8000 23060 8455
rect 23211 8168 23253 8177
rect 23211 8128 23212 8168
rect 23252 8128 23253 8168
rect 23211 8119 23253 8128
rect 23212 8034 23252 8119
rect 23020 7951 23060 7960
rect 23115 8000 23157 8009
rect 23115 7960 23116 8000
rect 23156 7960 23157 8000
rect 23115 7951 23157 7960
rect 23116 7866 23156 7951
rect 23404 7337 23444 10975
rect 24268 10193 24308 10984
rect 25420 10772 25460 10781
rect 25460 10732 25556 10772
rect 25420 10723 25460 10732
rect 25420 10268 25460 10277
rect 24267 10184 24309 10193
rect 24267 10144 24268 10184
rect 24308 10144 24309 10184
rect 24267 10135 24309 10144
rect 25420 10109 25460 10228
rect 25419 10100 25461 10109
rect 25419 10060 25420 10100
rect 25460 10060 25461 10100
rect 25419 10051 25461 10060
rect 25516 9521 25556 10732
rect 25612 10184 25652 10193
rect 25515 9512 25557 9521
rect 25515 9472 25516 9512
rect 25556 9472 25557 9512
rect 25515 9463 25557 9472
rect 25515 9260 25557 9269
rect 25515 9220 25516 9260
rect 25556 9220 25557 9260
rect 25515 9211 25557 9220
rect 25516 9126 25556 9211
rect 25612 8933 25652 10144
rect 25708 10184 25748 10193
rect 25708 9596 25748 10144
rect 26476 9680 26516 9689
rect 26516 9640 26900 9680
rect 25708 9556 25940 9596
rect 25611 8924 25653 8933
rect 25611 8884 25612 8924
rect 25652 8884 25653 8924
rect 25611 8875 25653 8884
rect 24939 8840 24981 8849
rect 24939 8800 24940 8840
rect 24980 8800 24981 8840
rect 24939 8791 24981 8800
rect 24940 8168 24980 8791
rect 25708 8177 25748 9556
rect 25900 9507 25940 9556
rect 25804 9470 25844 9479
rect 25900 9458 25940 9467
rect 25996 9512 26036 9523
rect 25996 9437 26036 9472
rect 26379 9512 26421 9521
rect 26379 9472 26380 9512
rect 26420 9472 26421 9512
rect 26379 9463 26421 9472
rect 25804 9353 25844 9430
rect 25995 9428 26037 9437
rect 25995 9388 25996 9428
rect 26036 9388 26037 9428
rect 25995 9379 26037 9388
rect 26380 9378 26420 9463
rect 25803 9344 25845 9353
rect 25803 9304 25804 9344
rect 25844 9304 25845 9344
rect 25803 9295 25845 9304
rect 26187 9344 26229 9353
rect 26187 9304 26188 9344
rect 26228 9304 26229 9344
rect 26187 9295 26229 9304
rect 25803 8924 25845 8933
rect 25803 8884 25804 8924
rect 25844 8884 25845 8924
rect 25803 8875 25845 8884
rect 25804 8504 25844 8875
rect 25995 8672 26037 8681
rect 25995 8632 25996 8672
rect 26036 8632 26037 8672
rect 25995 8623 26037 8632
rect 26092 8672 26132 8681
rect 26188 8672 26228 9295
rect 26476 8849 26516 9640
rect 26763 9512 26805 9521
rect 26763 9472 26764 9512
rect 26804 9472 26805 9512
rect 26763 9463 26805 9472
rect 26860 9512 26900 9640
rect 26860 9463 26900 9472
rect 26764 9344 26804 9463
rect 26860 9344 26900 9353
rect 26764 9304 26860 9344
rect 26860 9295 26900 9304
rect 26667 9260 26709 9269
rect 26667 9220 26668 9260
rect 26708 9220 26709 9260
rect 26667 9211 26709 9220
rect 26668 9126 26708 9211
rect 26475 8840 26517 8849
rect 26475 8800 26476 8840
rect 26516 8800 26517 8840
rect 26475 8791 26517 8800
rect 26132 8632 26228 8672
rect 26092 8623 26132 8632
rect 25996 8538 26036 8623
rect 25804 8455 25844 8464
rect 24940 8119 24980 8128
rect 25707 8168 25749 8177
rect 25707 8128 25708 8168
rect 25748 8128 25749 8168
rect 25707 8119 25749 8128
rect 27339 8084 27381 8093
rect 27339 8044 27340 8084
rect 27380 8044 27381 8084
rect 27339 8035 27381 8044
rect 26092 8000 26132 8009
rect 22347 7328 22389 7337
rect 22347 7288 22348 7328
rect 22388 7288 22389 7328
rect 22347 7279 22389 7288
rect 23403 7328 23445 7337
rect 23403 7288 23404 7328
rect 23444 7288 23445 7328
rect 23403 7279 23445 7288
rect 21484 7160 21524 7169
rect 22348 7160 22388 7279
rect 21524 7120 21716 7160
rect 21484 7111 21524 7120
rect 21580 6488 21620 6497
rect 21580 6245 21620 6448
rect 21676 6320 21716 7120
rect 22348 7111 22388 7120
rect 22923 7160 22965 7169
rect 22923 7120 22924 7160
rect 22964 7120 22965 7160
rect 22923 7111 22965 7120
rect 23596 7160 23636 7169
rect 22731 7076 22773 7085
rect 22731 7036 22732 7076
rect 22772 7036 22773 7076
rect 22731 7027 22773 7036
rect 22732 6942 22772 7027
rect 22924 7026 22964 7111
rect 23596 7001 23636 7120
rect 25995 7076 26037 7085
rect 25995 7036 25996 7076
rect 26036 7036 26037 7076
rect 25995 7027 26037 7036
rect 23595 6992 23637 7001
rect 23595 6952 23596 6992
rect 23636 6952 23637 6992
rect 23595 6943 23637 6952
rect 25996 6942 26036 7027
rect 22540 6488 22580 6497
rect 22580 6448 22676 6488
rect 22540 6439 22580 6448
rect 21868 6320 21908 6329
rect 21676 6280 21868 6320
rect 21868 6271 21908 6280
rect 21579 6236 21621 6245
rect 21579 6196 21580 6236
rect 21620 6196 21621 6236
rect 21579 6187 21621 6196
rect 21100 4180 21236 4220
rect 20043 4136 20085 4145
rect 20043 4096 20044 4136
rect 20084 4096 20085 4136
rect 20043 4087 20085 4096
rect 20523 4136 20565 4145
rect 20523 4096 20524 4136
rect 20564 4096 20565 4136
rect 20523 4087 20565 4096
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 20044 3632 20084 4087
rect 20524 4002 20564 4087
rect 21100 3641 21140 4180
rect 21772 4136 21812 4145
rect 21196 4052 21236 4061
rect 21388 4052 21428 4061
rect 21236 4012 21388 4052
rect 21196 4003 21236 4012
rect 21388 4003 21428 4012
rect 21772 3641 21812 4096
rect 22636 4136 22676 6448
rect 24555 4976 24597 4985
rect 24555 4936 24556 4976
rect 24596 4936 24597 4976
rect 24555 4927 24597 4936
rect 25611 4976 25653 4985
rect 25611 4936 25612 4976
rect 25652 4936 25653 4976
rect 25611 4927 25653 4936
rect 23787 4220 23829 4229
rect 23787 4180 23788 4220
rect 23828 4180 23829 4220
rect 23787 4171 23829 4180
rect 24363 4220 24405 4229
rect 24363 4180 24364 4220
rect 24404 4180 24405 4220
rect 24363 4171 24405 4180
rect 20044 3583 20084 3592
rect 21099 3632 21141 3641
rect 21099 3592 21100 3632
rect 21140 3592 21141 3632
rect 21099 3583 21141 3592
rect 21771 3632 21813 3641
rect 21771 3592 21772 3632
rect 21812 3592 21813 3632
rect 21771 3583 21813 3592
rect 22539 3548 22581 3557
rect 22539 3508 22540 3548
rect 22580 3508 22581 3548
rect 22539 3499 22581 3508
rect 18028 3464 18068 3473
rect 18028 2885 18068 3424
rect 18699 3464 18741 3473
rect 18699 3424 18700 3464
rect 18740 3424 18741 3464
rect 18699 3415 18741 3424
rect 18891 3464 18933 3473
rect 18891 3424 18892 3464
rect 18932 3424 18933 3464
rect 18891 3415 18933 3424
rect 21100 3464 21140 3473
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 18027 2876 18069 2885
rect 18027 2836 18028 2876
rect 18068 2836 18069 2876
rect 18027 2827 18069 2836
rect 17931 2792 17973 2801
rect 17931 2752 17932 2792
rect 17972 2752 17973 2792
rect 17931 2743 17973 2752
rect 17836 2575 17876 2584
rect 18700 2624 18740 3415
rect 18892 3330 18932 3415
rect 21100 2885 21140 3424
rect 21772 3464 21812 3473
rect 22156 3464 22196 3473
rect 21812 3424 22156 3464
rect 21772 3415 21812 3424
rect 22156 3415 22196 3424
rect 22540 3464 22580 3499
rect 22636 3473 22676 4096
rect 23788 4086 23828 4171
rect 24364 4136 24404 4171
rect 24364 4085 24404 4096
rect 24556 3632 24596 4927
rect 25612 4842 25652 4927
rect 25036 3968 25076 3977
rect 24556 3583 24596 3592
rect 24748 3928 25036 3968
rect 24748 3548 24788 3928
rect 25036 3919 25076 3928
rect 24748 3499 24788 3508
rect 25131 3548 25173 3557
rect 25131 3508 25132 3548
rect 25172 3508 25173 3548
rect 25131 3499 25173 3508
rect 22540 3413 22580 3424
rect 22635 3464 22677 3473
rect 22635 3424 22636 3464
rect 22676 3424 22677 3464
rect 22635 3415 22677 3424
rect 23403 3464 23445 3473
rect 23403 3424 23404 3464
rect 23444 3424 23445 3464
rect 23403 3415 23445 3424
rect 25132 3464 25172 3499
rect 23404 3330 23444 3415
rect 25132 3413 25172 3424
rect 25995 3464 26037 3473
rect 26092 3464 26132 7960
rect 26956 8000 26996 8009
rect 26956 7337 26996 7960
rect 27340 7950 27380 8035
rect 26955 7328 26997 7337
rect 26955 7288 26956 7328
rect 26996 7288 26997 7328
rect 26955 7279 26997 7288
rect 26667 7160 26709 7169
rect 26667 7120 26668 7160
rect 26708 7120 26709 7160
rect 26667 7111 26709 7120
rect 26668 7026 26708 7111
rect 28300 4985 28340 11647
rect 31372 11369 31412 11656
rect 31467 11696 31509 11705
rect 31467 11656 31468 11696
rect 31508 11656 31509 11696
rect 31467 11647 31509 11656
rect 31564 11696 31604 12244
rect 32044 12235 32084 12244
rect 32812 12284 32852 12293
rect 32812 11705 32852 12244
rect 33352 12116 33720 12125
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33352 12067 33720 12076
rect 34444 11957 34484 12496
rect 36171 12536 36213 12545
rect 36171 12496 36172 12536
rect 36212 12496 36213 12536
rect 36171 12487 36213 12496
rect 33963 11948 34005 11957
rect 33963 11908 33964 11948
rect 34004 11908 34005 11948
rect 33963 11899 34005 11908
rect 34443 11948 34485 11957
rect 34443 11908 34444 11948
rect 34484 11908 34485 11948
rect 34443 11899 34485 11908
rect 33964 11814 34004 11899
rect 31564 11647 31604 11656
rect 31947 11696 31989 11705
rect 31947 11656 31948 11696
rect 31988 11656 31989 11696
rect 31947 11647 31989 11656
rect 32331 11696 32373 11705
rect 32331 11656 32332 11696
rect 32372 11656 32373 11696
rect 32331 11647 32373 11656
rect 32811 11696 32853 11705
rect 32811 11656 32812 11696
rect 32852 11656 32853 11696
rect 32811 11647 32853 11656
rect 31371 11360 31413 11369
rect 31371 11320 31372 11360
rect 31412 11320 31413 11360
rect 31371 11311 31413 11320
rect 31083 10184 31125 10193
rect 31083 10144 31084 10184
rect 31124 10144 31125 10184
rect 31083 10135 31125 10144
rect 31468 10184 31508 11647
rect 31948 11562 31988 11647
rect 31851 11360 31893 11369
rect 31851 11320 31852 11360
rect 31892 11320 31893 11360
rect 31851 11311 31893 11320
rect 31852 10940 31892 11311
rect 31852 10891 31892 10900
rect 31660 10772 31700 10781
rect 31660 10193 31700 10732
rect 31468 10135 31508 10144
rect 31659 10184 31701 10193
rect 31659 10144 31660 10184
rect 31700 10144 31701 10184
rect 31659 10135 31701 10144
rect 32332 10184 32372 11647
rect 32812 11562 32852 11647
rect 36172 11369 36212 12487
rect 32811 11360 32853 11369
rect 32811 11320 32812 11360
rect 32852 11320 32853 11360
rect 32811 11311 32853 11320
rect 34592 11360 34960 11369
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34592 11311 34960 11320
rect 36171 11360 36213 11369
rect 36171 11320 36172 11360
rect 36212 11320 36213 11360
rect 36171 11311 36213 11320
rect 32812 11192 32852 11311
rect 32812 11143 32852 11152
rect 36172 11108 36212 11311
rect 36172 11059 36212 11068
rect 33484 11024 33524 11033
rect 37036 11024 37076 15100
rect 37612 13796 37652 13805
rect 37228 13756 37612 13796
rect 37228 13208 37268 13756
rect 37612 13747 37652 13756
rect 37228 13159 37268 13168
rect 37612 13208 37652 13217
rect 37708 13208 37748 15100
rect 40780 15100 40916 15140
rect 40780 14720 40820 15100
rect 40780 14645 40820 14680
rect 40875 14720 40917 14729
rect 40875 14680 40876 14720
rect 40916 14680 40917 14720
rect 40875 14671 40917 14680
rect 40972 14720 41012 14729
rect 40203 14636 40245 14645
rect 40203 14596 40204 14636
rect 40244 14596 40245 14636
rect 40203 14587 40245 14596
rect 40779 14636 40821 14645
rect 40779 14596 40780 14636
rect 40820 14596 40821 14636
rect 40779 14587 40821 14596
rect 38956 14048 38996 14057
rect 38475 13208 38517 13217
rect 37652 13168 37844 13208
rect 37612 13159 37652 13168
rect 33524 10984 33812 11024
rect 33484 10975 33524 10984
rect 33352 10604 33720 10613
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33352 10555 33720 10564
rect 33484 10436 33524 10445
rect 33772 10436 33812 10984
rect 33524 10396 33812 10436
rect 33484 10387 33524 10396
rect 32332 10135 32372 10144
rect 31084 10050 31124 10135
rect 34592 9848 34960 9857
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34592 9799 34960 9808
rect 33352 9092 33720 9101
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33352 9043 33720 9052
rect 30028 8840 30068 8849
rect 29740 8800 30028 8840
rect 29356 8672 29396 8681
rect 28684 8504 28724 8513
rect 28684 8093 28724 8464
rect 29356 8168 29396 8632
rect 29548 8168 29588 8177
rect 29356 8128 29548 8168
rect 29548 8119 29588 8128
rect 28683 8084 28725 8093
rect 28683 8044 28684 8084
rect 28724 8044 28725 8084
rect 28683 8035 28725 8044
rect 29643 8000 29685 8009
rect 29643 7960 29644 8000
rect 29684 7960 29685 8000
rect 29643 7951 29685 7960
rect 29740 8000 29780 8800
rect 30028 8791 30068 8800
rect 30028 8672 30068 8681
rect 29740 7951 29780 7960
rect 29836 8000 29876 8009
rect 29644 7866 29684 7951
rect 29836 7328 29876 7960
rect 29356 7288 29876 7328
rect 29067 7244 29109 7253
rect 29067 7204 29068 7244
rect 29108 7204 29109 7244
rect 29067 7195 29109 7204
rect 28588 7160 28628 7169
rect 28395 6992 28437 7001
rect 28395 6952 28396 6992
rect 28436 6952 28437 6992
rect 28395 6943 28437 6952
rect 28396 6858 28436 6943
rect 28588 6665 28628 7120
rect 28875 7160 28917 7169
rect 28875 7120 28876 7160
rect 28916 7120 28917 7160
rect 28875 7111 28917 7120
rect 28876 7026 28916 7111
rect 29068 7110 29108 7195
rect 29356 7160 29396 7288
rect 29356 7111 29396 7120
rect 29452 7160 29492 7169
rect 29452 7001 29492 7120
rect 29451 6992 29493 7001
rect 29451 6952 29452 6992
rect 29492 6952 29493 6992
rect 29451 6943 29493 6952
rect 28587 6656 28629 6665
rect 28587 6616 28588 6656
rect 28628 6616 28629 6656
rect 28587 6607 28629 6616
rect 29451 6656 29493 6665
rect 29451 6616 29452 6656
rect 29492 6616 29493 6656
rect 29451 6607 29493 6616
rect 29643 6656 29685 6665
rect 29643 6616 29644 6656
rect 29684 6616 29685 6656
rect 29643 6607 29685 6616
rect 29452 6522 29492 6607
rect 28780 6488 28820 6497
rect 29644 6488 29684 6607
rect 29740 6572 29780 7288
rect 30028 7169 30068 8632
rect 30220 8672 30260 8681
rect 30260 8632 30452 8672
rect 30220 8623 30260 8632
rect 30315 8000 30357 8009
rect 30315 7960 30316 8000
rect 30356 7960 30357 8000
rect 30315 7951 30357 7960
rect 30316 7866 30356 7951
rect 30027 7160 30069 7169
rect 30027 7120 30028 7160
rect 30068 7120 30069 7160
rect 30027 7111 30069 7120
rect 30219 7160 30261 7169
rect 30219 7120 30220 7160
rect 30260 7120 30261 7160
rect 30219 7111 30261 7120
rect 30412 7160 30452 8632
rect 35979 8504 36021 8513
rect 35979 8464 35980 8504
rect 36020 8464 36021 8504
rect 35979 8455 36021 8464
rect 34592 8336 34960 8345
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34592 8287 34960 8296
rect 30988 8000 31028 8009
rect 30700 7412 30740 7421
rect 30988 7412 31028 7960
rect 32908 8000 32948 8009
rect 33484 8000 33524 8009
rect 32948 7960 33484 8000
rect 32908 7951 32948 7960
rect 33484 7951 33524 7960
rect 34732 8000 34772 8009
rect 31083 7748 31125 7757
rect 31083 7708 31084 7748
rect 31124 7708 31125 7748
rect 31083 7699 31125 7708
rect 32235 7748 32277 7757
rect 32235 7708 32236 7748
rect 32276 7708 32277 7748
rect 32235 7699 32277 7708
rect 30740 7372 31028 7412
rect 30700 7363 30740 7372
rect 30604 7169 30644 7254
rect 30028 7026 30068 7111
rect 29931 6992 29973 7001
rect 29931 6952 29932 6992
rect 29972 6952 29973 6992
rect 29931 6943 29973 6952
rect 29932 6858 29972 6943
rect 29740 6523 29780 6532
rect 28820 6448 28916 6488
rect 28780 6439 28820 6448
rect 26284 4976 26324 4985
rect 26476 4976 26516 4985
rect 26324 4936 26476 4976
rect 26284 4927 26324 4936
rect 26476 4927 26516 4936
rect 26859 4976 26901 4985
rect 26859 4936 26860 4976
rect 26900 4936 26901 4976
rect 26859 4927 26901 4936
rect 27724 4976 27764 4985
rect 26860 3557 26900 4927
rect 27724 4145 27764 4936
rect 28299 4976 28341 4985
rect 28299 4936 28300 4976
rect 28340 4936 28341 4976
rect 28299 4927 28341 4936
rect 27052 4136 27092 4145
rect 27052 3632 27092 4096
rect 27723 4136 27765 4145
rect 27723 4096 27724 4136
rect 27764 4096 27765 4136
rect 27723 4087 27765 4096
rect 28300 4136 28340 4927
rect 28876 4892 28916 6448
rect 29644 6439 29684 6448
rect 29835 6488 29877 6497
rect 29835 6448 29836 6488
rect 29876 6448 29877 6488
rect 29835 6439 29877 6448
rect 29836 6354 29876 6439
rect 28876 4843 28916 4852
rect 30220 4388 30260 7111
rect 30412 6992 30452 7120
rect 30603 7160 30645 7169
rect 30603 7120 30604 7160
rect 30644 7120 30645 7160
rect 30603 7111 30645 7120
rect 30796 7160 30836 7169
rect 31084 7160 31124 7699
rect 32236 7614 32276 7699
rect 33352 7580 33720 7589
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33352 7531 33720 7540
rect 30836 7120 31124 7160
rect 32332 7160 32372 7171
rect 34636 7160 34676 7169
rect 34732 7160 34772 7960
rect 35596 8000 35636 8009
rect 35596 7841 35636 7960
rect 35980 8000 36020 8455
rect 37036 8009 37076 10984
rect 35980 7951 36020 7960
rect 37035 8000 37077 8009
rect 37035 7960 37036 8000
rect 37076 7960 37077 8000
rect 37035 7951 37077 7960
rect 37227 8000 37269 8009
rect 37227 7960 37228 8000
rect 37268 7960 37269 8000
rect 37804 8000 37844 13168
rect 38475 13168 38476 13208
rect 38516 13168 38517 13208
rect 38475 13159 38517 13168
rect 38476 13074 38516 13159
rect 38956 11369 38996 14008
rect 39627 14048 39669 14057
rect 39627 14008 39628 14048
rect 39668 14008 39669 14048
rect 39627 13999 39669 14008
rect 39916 14048 39956 14057
rect 39244 13796 39284 13805
rect 39244 13217 39284 13756
rect 39628 13460 39668 13999
rect 39916 13889 39956 14008
rect 39915 13880 39957 13889
rect 39915 13840 39916 13880
rect 39956 13840 39957 13880
rect 39915 13831 39957 13840
rect 39668 13420 39860 13460
rect 39628 13411 39668 13420
rect 39243 13208 39285 13217
rect 39243 13168 39244 13208
rect 39284 13168 39285 13208
rect 39243 13159 39285 13168
rect 39531 13208 39573 13217
rect 39531 13168 39532 13208
rect 39572 13168 39573 13208
rect 39531 13159 39573 13168
rect 39820 13208 39860 13420
rect 39820 13159 39860 13168
rect 40204 13208 40244 14587
rect 40876 14586 40916 14671
rect 40972 14216 41012 14680
rect 41452 14720 41492 16948
rect 41739 16939 41781 16948
rect 41547 16820 41589 16829
rect 41547 16780 41548 16820
rect 41588 16780 41589 16820
rect 41547 16771 41589 16780
rect 41548 15560 41588 16771
rect 41548 15511 41588 15520
rect 41740 15560 41780 16939
rect 42411 16820 42453 16829
rect 42411 16780 42412 16820
rect 42452 16780 42453 16820
rect 42411 16771 42453 16780
rect 42412 16686 42452 16771
rect 42603 15728 42645 15737
rect 42603 15688 42604 15728
rect 42644 15688 42645 15728
rect 42603 15679 42645 15688
rect 41740 15140 41780 15520
rect 42604 15560 42644 15679
rect 42604 15485 42644 15520
rect 42603 15476 42645 15485
rect 42603 15436 42604 15476
rect 42644 15436 42645 15476
rect 42603 15427 42645 15436
rect 42604 15396 42644 15427
rect 41740 15100 41876 15140
rect 41452 14671 41492 14680
rect 41547 14720 41589 14729
rect 41547 14680 41548 14720
rect 41588 14680 41589 14720
rect 41547 14671 41589 14680
rect 41548 14586 41588 14671
rect 40972 14167 41012 14176
rect 41260 14552 41300 14561
rect 41260 14057 41300 14512
rect 40299 14048 40341 14057
rect 40299 14008 40300 14048
rect 40340 14008 40341 14048
rect 40299 13999 40341 14008
rect 41259 14048 41301 14057
rect 41259 14008 41260 14048
rect 41300 14008 41301 14048
rect 41259 13999 41301 14008
rect 40300 13914 40340 13999
rect 40204 13159 40244 13168
rect 41452 13796 41492 13805
rect 41452 13208 41492 13756
rect 41452 13159 41492 13168
rect 41836 13208 41876 15100
rect 42123 14048 42165 14057
rect 42123 14008 42124 14048
rect 42164 14008 42165 14048
rect 42123 13999 42165 14008
rect 42124 13914 42164 13999
rect 42700 13889 42740 17023
rect 44332 15737 44372 23920
rect 44428 23792 44468 23801
rect 44468 23752 44660 23792
rect 44428 23743 44468 23752
rect 44620 22532 44660 23752
rect 44716 23129 44756 23920
rect 45963 23624 46005 23633
rect 45963 23584 45964 23624
rect 46004 23584 46005 23624
rect 45963 23575 46005 23584
rect 45964 23204 46004 23575
rect 45964 23155 46004 23164
rect 44715 23120 44757 23129
rect 44715 23080 44716 23120
rect 44756 23080 44757 23120
rect 44715 23071 44757 23080
rect 45580 23120 45620 23131
rect 44716 22986 44756 23071
rect 45580 23045 45620 23080
rect 45579 23036 45621 23045
rect 45579 22996 45580 23036
rect 45620 22996 45621 23036
rect 45579 22987 45621 22996
rect 45004 22532 45044 22541
rect 44620 22492 45004 22532
rect 45004 22483 45044 22492
rect 47308 22280 47348 25171
rect 48268 23960 48308 26776
rect 49712 26480 50080 26489
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 49712 26431 50080 26440
rect 64832 26480 65200 26489
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 64832 26431 65200 26440
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 95072 26480 95440 26489
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95072 26431 95440 26440
rect 48472 25724 48840 25733
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48472 25675 48840 25684
rect 63592 25724 63960 25733
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63592 25675 63960 25684
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 93832 25724 94200 25733
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 93832 25675 94200 25684
rect 49712 24968 50080 24977
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 49712 24919 50080 24928
rect 64832 24968 65200 24977
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 64832 24919 65200 24928
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 95072 24968 95440 24977
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95072 24919 95440 24928
rect 48472 24212 48840 24221
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48472 24163 48840 24172
rect 63592 24212 63960 24221
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63592 24163 63960 24172
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 93832 24212 94200 24221
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 93832 24163 94200 24172
rect 47980 23920 48308 23960
rect 47308 22231 47348 22240
rect 47884 23120 47924 23129
rect 47884 21785 47924 23080
rect 47980 22448 48020 23920
rect 49712 23456 50080 23465
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 49712 23407 50080 23416
rect 64832 23456 65200 23465
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 64832 23407 65200 23416
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 95072 23456 95440 23465
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95072 23407 95440 23416
rect 48268 23120 48308 23131
rect 48268 23045 48308 23080
rect 49131 23120 49173 23129
rect 49131 23080 49132 23120
rect 49172 23080 49173 23120
rect 49131 23071 49173 23080
rect 48267 23036 48309 23045
rect 48267 22996 48268 23036
rect 48308 22996 48309 23036
rect 48267 22987 48309 22996
rect 48939 23036 48981 23045
rect 48939 22996 48940 23036
rect 48980 22996 48981 23036
rect 48939 22987 48981 22996
rect 48472 22700 48840 22709
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48472 22651 48840 22660
rect 47980 22289 48020 22408
rect 47979 22280 48021 22289
rect 47979 22240 47980 22280
rect 48020 22240 48021 22280
rect 47979 22231 48021 22240
rect 48844 22280 48884 22289
rect 48940 22280 48980 22987
rect 49132 22986 49172 23071
rect 50284 22868 50324 22877
rect 50188 22828 50284 22868
rect 48884 22240 48980 22280
rect 49707 22280 49749 22289
rect 49707 22240 49708 22280
rect 49748 22240 49749 22280
rect 48844 22231 48884 22240
rect 49707 22231 49749 22240
rect 47883 21776 47925 21785
rect 47883 21736 47884 21776
rect 47924 21736 47925 21776
rect 47883 21727 47925 21736
rect 47980 19265 48020 22231
rect 48460 22196 48500 22205
rect 48500 22156 48788 22196
rect 48460 22147 48500 22156
rect 48075 21776 48117 21785
rect 48075 21736 48076 21776
rect 48116 21736 48117 21776
rect 48748 21776 48788 22156
rect 49708 22146 49748 22231
rect 49712 21944 50080 21953
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 49712 21895 50080 21904
rect 49036 21776 49076 21785
rect 48748 21736 49036 21776
rect 48075 21727 48117 21736
rect 49036 21727 49076 21736
rect 48076 21642 48116 21727
rect 50092 21608 50132 21617
rect 50188 21608 50228 22828
rect 50284 22819 50324 22828
rect 63592 22700 63960 22709
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63592 22651 63960 22660
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 93832 22700 94200 22709
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 93832 22651 94200 22660
rect 50132 21568 50228 21608
rect 50860 22112 50900 22121
rect 50860 21608 50900 22072
rect 64832 21944 65200 21953
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 64832 21895 65200 21904
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 95072 21944 95440 21953
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95072 21895 95440 21904
rect 50956 21608 50996 21617
rect 50860 21568 50956 21608
rect 50092 21559 50132 21568
rect 50956 21559 50996 21568
rect 48268 21524 48308 21535
rect 48268 21449 48308 21484
rect 49227 21524 49269 21533
rect 50283 21524 50325 21533
rect 49227 21484 49228 21524
rect 49268 21484 49269 21524
rect 49227 21475 49269 21484
rect 50188 21484 50284 21524
rect 50324 21484 50325 21524
rect 48267 21440 48309 21449
rect 48267 21400 48268 21440
rect 48308 21400 48309 21440
rect 48267 21391 48309 21400
rect 49228 21390 49268 21475
rect 49419 21440 49461 21449
rect 49419 21400 49420 21440
rect 49460 21400 49556 21440
rect 49419 21391 49461 21400
rect 49420 21306 49460 21391
rect 48472 21188 48840 21197
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48472 21139 48840 21148
rect 48171 20096 48213 20105
rect 48076 20056 48172 20096
rect 48212 20056 48213 20096
rect 46732 19256 46772 19265
rect 47595 19256 47637 19265
rect 46772 19216 46868 19256
rect 46732 19207 46772 19216
rect 46347 19172 46389 19181
rect 46347 19132 46348 19172
rect 46388 19132 46389 19172
rect 46347 19123 46389 19132
rect 46348 19038 46388 19123
rect 46732 18584 46772 18593
rect 46732 18005 46772 18544
rect 46828 18509 46868 19216
rect 47595 19216 47596 19256
rect 47636 19216 47637 19256
rect 47595 19207 47637 19216
rect 47979 19256 48021 19265
rect 47979 19216 47980 19256
rect 48020 19216 48021 19256
rect 47979 19207 48021 19216
rect 47211 19172 47253 19181
rect 47211 19132 47212 19172
rect 47252 19132 47253 19172
rect 47211 19123 47253 19132
rect 47116 18584 47156 18595
rect 47116 18509 47156 18544
rect 46827 18500 46869 18509
rect 46827 18460 46828 18500
rect 46868 18460 46869 18500
rect 46827 18451 46869 18460
rect 47115 18500 47157 18509
rect 47115 18460 47116 18500
rect 47156 18460 47157 18500
rect 47115 18451 47157 18460
rect 46731 17996 46773 18005
rect 46731 17956 46732 17996
rect 46772 17956 46773 17996
rect 46731 17947 46773 17956
rect 44331 15728 44373 15737
rect 44331 15688 44332 15728
rect 44372 15688 44373 15728
rect 44331 15679 44373 15688
rect 45099 15728 45141 15737
rect 45099 15688 45100 15728
rect 45140 15688 45141 15728
rect 45099 15679 45141 15688
rect 45100 14720 45140 15679
rect 47116 14972 47156 18451
rect 47212 17996 47252 19123
rect 47596 19122 47636 19207
rect 47980 18593 48020 19207
rect 47979 18584 48021 18593
rect 47979 18544 47980 18584
rect 48020 18544 48021 18584
rect 47979 18535 48021 18544
rect 47980 18450 48020 18535
rect 47212 17947 47252 17956
rect 47595 17996 47637 18005
rect 47595 17956 47596 17996
rect 47636 17956 47637 17996
rect 47595 17947 47637 17956
rect 47787 17996 47829 18005
rect 47787 17956 47788 17996
rect 47828 17956 47829 17996
rect 47787 17947 47829 17956
rect 47596 17862 47636 17947
rect 47403 17828 47445 17837
rect 47403 17788 47404 17828
rect 47444 17788 47445 17828
rect 47403 17779 47445 17788
rect 47788 17828 47828 17947
rect 48076 17837 48116 20056
rect 48171 20047 48213 20056
rect 48844 20096 48884 20105
rect 49323 20096 49365 20105
rect 48884 20056 48980 20096
rect 48844 20047 48884 20056
rect 48172 19962 48212 20047
rect 48472 19676 48840 19685
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48472 19627 48840 19636
rect 48748 19508 48788 19517
rect 48940 19508 48980 20056
rect 49323 20056 49324 20096
rect 49364 20056 49365 20096
rect 49323 20047 49365 20056
rect 49516 20096 49556 21400
rect 49712 20432 50080 20441
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 49712 20383 50080 20392
rect 49803 20180 49845 20189
rect 49803 20140 49804 20180
rect 49844 20140 49845 20180
rect 49803 20131 49845 20140
rect 49516 20047 49556 20056
rect 49708 20096 49748 20105
rect 49324 19962 49364 20047
rect 48788 19468 48980 19508
rect 49420 19844 49460 19853
rect 48748 19459 48788 19468
rect 49420 19265 49460 19804
rect 49419 19256 49461 19265
rect 49419 19216 49420 19256
rect 49460 19216 49461 19256
rect 49419 19207 49461 19216
rect 49708 19088 49748 20056
rect 49804 20046 49844 20131
rect 49900 20096 49940 20105
rect 50188 20096 50228 21484
rect 50283 21475 50325 21484
rect 50284 21390 50324 21475
rect 63592 21188 63960 21197
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63592 21139 63960 21148
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 93832 21188 94200 21197
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 93832 21139 94200 21148
rect 64832 20432 65200 20441
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 64832 20383 65200 20392
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 95072 20432 95440 20441
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95072 20383 95440 20392
rect 50475 20180 50517 20189
rect 50475 20140 50476 20180
rect 50516 20140 50517 20180
rect 50475 20131 50517 20140
rect 49940 20056 50228 20096
rect 49900 20047 49940 20056
rect 50187 19256 50229 19265
rect 50187 19216 50188 19256
rect 50228 19216 50229 19256
rect 50187 19207 50229 19216
rect 50476 19256 50516 20131
rect 63592 19676 63960 19685
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63592 19627 63960 19636
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 93832 19676 94200 19685
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 93832 19627 94200 19636
rect 50476 19207 50516 19216
rect 50188 19122 50228 19207
rect 49612 19048 49748 19088
rect 50667 19088 50709 19097
rect 50667 19048 50668 19088
rect 50708 19048 50709 19088
rect 49132 18332 49172 18341
rect 49172 18292 49268 18332
rect 49132 18283 49172 18292
rect 48472 18164 48840 18173
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48472 18115 48840 18124
rect 48171 17996 48213 18005
rect 48171 17956 48172 17996
rect 48212 17956 48213 17996
rect 48171 17947 48213 17956
rect 48555 17996 48597 18005
rect 48555 17956 48556 17996
rect 48596 17956 48597 17996
rect 48555 17947 48597 17956
rect 47788 17779 47828 17788
rect 48075 17828 48117 17837
rect 48075 17788 48076 17828
rect 48116 17788 48117 17828
rect 48075 17779 48117 17788
rect 47404 17694 47444 17779
rect 48076 17576 48116 17779
rect 48172 17744 48212 17947
rect 48556 17862 48596 17947
rect 48172 17695 48212 17704
rect 49228 17744 49268 18292
rect 49612 18005 49652 19048
rect 50667 19039 50709 19048
rect 52011 19088 52053 19097
rect 52011 19048 52012 19088
rect 52052 19048 52053 19088
rect 52011 19039 52053 19048
rect 50668 18954 50708 19039
rect 49712 18920 50080 18929
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 49712 18871 50080 18880
rect 52012 18668 52052 19039
rect 64832 18920 65200 18929
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 64832 18871 65200 18880
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 95072 18920 95440 18929
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95072 18871 95440 18880
rect 52012 18619 52052 18628
rect 52396 18584 52436 18593
rect 52299 18500 52341 18509
rect 52396 18500 52436 18544
rect 53259 18584 53301 18593
rect 53259 18544 53260 18584
rect 53300 18544 53301 18584
rect 53259 18535 53301 18544
rect 52299 18460 52300 18500
rect 52340 18460 52436 18500
rect 52299 18451 52341 18460
rect 53260 18450 53300 18535
rect 54412 18332 54452 18341
rect 49611 17996 49653 18005
rect 49611 17956 49612 17996
rect 49652 17956 49653 17996
rect 49611 17947 49653 17956
rect 49228 17695 49268 17704
rect 48076 17527 48116 17536
rect 48364 17576 48404 17585
rect 48364 15653 48404 17536
rect 49712 17408 50080 17417
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 49712 17359 50080 17368
rect 54412 17072 54452 18292
rect 63592 18164 63960 18173
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63592 18115 63960 18124
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 93832 18164 94200 18173
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 93832 18115 94200 18124
rect 64832 17408 65200 17417
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 64832 17359 65200 17368
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 95072 17408 95440 17417
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95072 17359 95440 17368
rect 54988 17240 55028 17249
rect 54796 17200 54988 17240
rect 54508 17072 54548 17081
rect 54412 17032 54508 17072
rect 54508 17023 54548 17032
rect 48472 16652 48840 16661
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48472 16603 48840 16612
rect 49712 15896 50080 15905
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 49712 15847 50080 15856
rect 48363 15644 48405 15653
rect 48363 15604 48364 15644
rect 48404 15604 48405 15644
rect 48363 15595 48405 15604
rect 49227 15644 49269 15653
rect 49227 15604 49228 15644
rect 49268 15604 49269 15644
rect 49227 15595 49269 15604
rect 49228 15510 49268 15595
rect 49612 15560 49652 15569
rect 48472 15140 48840 15149
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48472 15091 48840 15100
rect 47116 14923 47156 14932
rect 49612 14729 49652 15520
rect 50476 15560 50516 15569
rect 45100 14671 45140 14680
rect 46059 14720 46101 14729
rect 46059 14680 46060 14720
rect 46100 14680 46101 14720
rect 46059 14671 46101 14680
rect 46635 14720 46677 14729
rect 46635 14680 46636 14720
rect 46676 14680 46677 14720
rect 46635 14671 46677 14680
rect 47596 14720 47636 14729
rect 49611 14720 49653 14729
rect 47636 14680 47924 14720
rect 47596 14671 47636 14680
rect 46060 14586 46100 14671
rect 46636 14586 46676 14671
rect 47884 14057 47924 14680
rect 49611 14680 49612 14720
rect 49652 14680 49653 14720
rect 49611 14671 49653 14680
rect 50379 14552 50421 14561
rect 50379 14512 50380 14552
rect 50420 14512 50421 14552
rect 50379 14503 50421 14512
rect 49712 14384 50080 14393
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 49712 14335 50080 14344
rect 50380 14132 50420 14503
rect 50380 14083 50420 14092
rect 47883 14048 47925 14057
rect 47883 14008 47884 14048
rect 47924 14008 47925 14048
rect 47883 13999 47925 14008
rect 49132 14048 49172 14057
rect 42699 13880 42741 13889
rect 42699 13840 42700 13880
rect 42740 13840 42741 13880
rect 42699 13831 42741 13840
rect 41836 13159 41876 13168
rect 42700 13208 42740 13831
rect 42700 13159 42740 13168
rect 45291 13208 45333 13217
rect 45291 13168 45292 13208
rect 45332 13168 45333 13208
rect 45291 13159 45333 13168
rect 47115 13208 47157 13217
rect 47115 13168 47116 13208
rect 47156 13168 47157 13208
rect 47884 13208 47924 13999
rect 47979 13880 48021 13889
rect 47979 13840 47980 13880
rect 48020 13840 48021 13880
rect 47979 13831 48021 13840
rect 47980 13746 48020 13831
rect 48363 13796 48405 13805
rect 48363 13756 48364 13796
rect 48404 13756 48405 13796
rect 48363 13747 48405 13756
rect 47980 13208 48020 13217
rect 47884 13168 47980 13208
rect 47115 13159 47157 13168
rect 47980 13159 48020 13168
rect 48364 13208 48404 13747
rect 48472 13628 48840 13637
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48472 13579 48840 13588
rect 49132 13217 49172 14008
rect 49995 14048 50037 14057
rect 49995 14008 49996 14048
rect 50036 14008 50037 14048
rect 49995 13999 50037 14008
rect 49996 13914 50036 13999
rect 49611 13880 49653 13889
rect 49611 13840 49612 13880
rect 49652 13840 49653 13880
rect 49611 13831 49653 13840
rect 48364 13159 48404 13168
rect 49131 13208 49173 13217
rect 49131 13168 49132 13208
rect 49172 13168 49173 13208
rect 49131 13159 49173 13168
rect 49323 13208 49365 13217
rect 49323 13168 49324 13208
rect 49364 13168 49365 13208
rect 49323 13159 49365 13168
rect 38955 11360 38997 11369
rect 38955 11320 38956 11360
rect 38996 11320 38997 11360
rect 38955 11311 38997 11320
rect 38379 11024 38421 11033
rect 38379 10984 38380 11024
rect 38420 10984 38421 11024
rect 38379 10975 38421 10984
rect 38380 10436 38420 10975
rect 38380 10387 38420 10396
rect 39532 10184 39572 13159
rect 40300 13040 40340 13049
rect 43852 13040 43892 13049
rect 40340 13000 40724 13040
rect 40300 12991 40340 13000
rect 40684 11696 40724 13000
rect 43892 13000 44084 13040
rect 43852 12991 43892 13000
rect 40684 11647 40724 11656
rect 41356 11528 41396 11537
rect 40780 11488 41356 11528
rect 39915 11024 39957 11033
rect 39915 10984 39916 11024
rect 39956 10984 39957 11024
rect 39915 10975 39957 10984
rect 40299 11024 40341 11033
rect 40299 10984 40300 11024
rect 40340 10984 40341 11024
rect 40299 10975 40341 10984
rect 39916 10890 39956 10975
rect 39532 10135 39572 10144
rect 39916 9512 39956 9521
rect 39820 9472 39916 9512
rect 38763 9260 38805 9269
rect 38763 9220 38764 9260
rect 38804 9220 38805 9260
rect 38763 9211 38805 9220
rect 39531 9260 39573 9269
rect 39531 9220 39532 9260
rect 39572 9220 39573 9260
rect 39531 9211 39573 9220
rect 38764 9126 38804 9211
rect 38763 8840 38805 8849
rect 38763 8800 38764 8840
rect 38804 8800 38805 8840
rect 38763 8791 38805 8800
rect 38379 8504 38421 8513
rect 38379 8464 38380 8504
rect 38420 8464 38421 8504
rect 38379 8455 38421 8464
rect 38380 8370 38420 8455
rect 38667 8084 38709 8093
rect 38667 8044 38668 8084
rect 38708 8044 38709 8084
rect 38667 8035 38709 8044
rect 37900 8000 37940 8009
rect 37804 7960 37900 8000
rect 37227 7951 37269 7960
rect 37228 7866 37268 7951
rect 35595 7832 35637 7841
rect 35595 7792 35596 7832
rect 35636 7792 35637 7832
rect 35595 7783 35637 7792
rect 30796 6992 30836 7120
rect 32332 7085 32372 7120
rect 34444 7120 34636 7160
rect 34676 7120 34772 7160
rect 35500 7160 35540 7169
rect 35596 7160 35636 7783
rect 35540 7120 35636 7160
rect 36556 7748 36596 7757
rect 32331 7076 32373 7085
rect 32331 7036 32332 7076
rect 32372 7036 32373 7076
rect 32331 7027 32373 7036
rect 30412 6952 30836 6992
rect 31660 6992 31700 7001
rect 31660 6497 31700 6952
rect 33483 6992 33525 7001
rect 33483 6952 33484 6992
rect 33524 6952 33525 6992
rect 33483 6943 33525 6952
rect 33484 6858 33524 6943
rect 31659 6488 31701 6497
rect 31659 6448 31660 6488
rect 31700 6448 31701 6488
rect 31659 6439 31701 6448
rect 34444 6320 34484 7120
rect 34636 7111 34676 7120
rect 34592 6824 34960 6833
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34592 6775 34960 6784
rect 34348 6280 34484 6320
rect 33352 6068 33720 6077
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33352 6019 33720 6028
rect 33867 5648 33909 5657
rect 33867 5608 33868 5648
rect 33908 5608 33909 5648
rect 33867 5599 33909 5608
rect 33868 5514 33908 5599
rect 33388 5480 33428 5489
rect 33388 5069 33428 5440
rect 34348 5069 34388 6280
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 33387 5060 33429 5069
rect 33387 5020 33388 5060
rect 33428 5020 33429 5060
rect 33387 5011 33429 5020
rect 34347 5060 34389 5069
rect 34347 5020 34348 5060
rect 34388 5020 34389 5060
rect 34347 5011 34389 5020
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 30316 4388 30356 4397
rect 30220 4348 30316 4388
rect 30316 4339 30356 4348
rect 34348 4145 34388 5011
rect 34443 4220 34485 4229
rect 34443 4180 34444 4220
rect 34484 4180 34485 4220
rect 34443 4171 34485 4180
rect 28300 4087 28340 4096
rect 29163 4136 29205 4145
rect 29163 4096 29164 4136
rect 29204 4096 29205 4136
rect 29163 4087 29205 4096
rect 34347 4136 34389 4145
rect 34347 4096 34348 4136
rect 34388 4096 34389 4136
rect 34347 4087 34389 4096
rect 27916 4052 27956 4061
rect 27724 3968 27764 3977
rect 27916 3968 27956 4012
rect 29164 4002 29204 4087
rect 27764 3928 27956 3968
rect 33387 3968 33429 3977
rect 33387 3928 33388 3968
rect 33428 3928 33429 3968
rect 27724 3919 27764 3928
rect 33387 3919 33429 3928
rect 34251 3968 34293 3977
rect 34251 3928 34252 3968
rect 34292 3928 34293 3968
rect 34251 3919 34293 3928
rect 27148 3632 27188 3641
rect 27052 3592 27148 3632
rect 27148 3583 27188 3592
rect 26859 3548 26901 3557
rect 26859 3508 26860 3548
rect 26900 3508 26901 3548
rect 26859 3499 26901 3508
rect 33388 3548 33428 3919
rect 34252 3834 34292 3919
rect 33388 3499 33428 3508
rect 25995 3424 25996 3464
rect 26036 3424 26132 3464
rect 33772 3464 33812 3473
rect 34348 3464 34388 4087
rect 34444 4086 34484 4171
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 34636 3464 34676 3473
rect 34348 3424 34636 3464
rect 25995 3415 26037 3424
rect 25996 3330 26036 3415
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 19851 2876 19893 2885
rect 19851 2836 19852 2876
rect 19892 2836 19893 2876
rect 19851 2827 19893 2836
rect 21099 2876 21141 2885
rect 21099 2836 21100 2876
rect 21140 2836 21141 2876
rect 21099 2827 21141 2836
rect 19852 2742 19892 2827
rect 33772 2717 33812 3424
rect 34636 3415 34676 3424
rect 35500 2717 35540 7120
rect 35883 7076 35925 7085
rect 35883 7036 35884 7076
rect 35924 7036 35925 7076
rect 35883 7027 35925 7036
rect 35884 6942 35924 7027
rect 36556 6497 36596 7708
rect 36555 6488 36597 6497
rect 36555 6448 36556 6488
rect 36596 6448 36597 6488
rect 36555 6439 36597 6448
rect 36556 5657 36596 6439
rect 37900 6320 37940 7960
rect 38091 7832 38133 7841
rect 38091 7792 38092 7832
rect 38132 7792 38133 7832
rect 38091 7783 38133 7792
rect 38092 7698 38132 7783
rect 38668 7160 38708 8035
rect 38764 8000 38804 8791
rect 39051 8756 39093 8765
rect 39051 8716 39052 8756
rect 39092 8716 39093 8756
rect 39051 8707 39093 8716
rect 39052 8672 39092 8707
rect 39052 8621 39092 8632
rect 39532 8672 39572 9211
rect 39532 8623 39572 8632
rect 38764 7951 38804 7960
rect 38668 7111 38708 7120
rect 37995 7076 38037 7085
rect 37995 7036 37996 7076
rect 38036 7036 38037 7076
rect 37995 7027 38037 7036
rect 37996 6942 38036 7027
rect 38763 6992 38805 7001
rect 38763 6952 38764 6992
rect 38804 6952 38805 6992
rect 38763 6943 38805 6952
rect 39531 6992 39573 7001
rect 39531 6952 39532 6992
rect 39572 6952 39573 6992
rect 39531 6943 39573 6952
rect 38572 6329 38612 6414
rect 38764 6404 38804 6943
rect 39532 6858 39572 6943
rect 39820 6656 39860 9472
rect 39916 9463 39956 9472
rect 40203 9512 40245 9521
rect 40203 9472 40204 9512
rect 40244 9472 40245 9512
rect 40203 9463 40245 9472
rect 40204 8840 40244 9463
rect 39915 8084 39957 8093
rect 39915 8044 39916 8084
rect 39956 8044 39957 8084
rect 39915 8035 39957 8044
rect 39916 7950 39956 8035
rect 40108 8000 40148 8009
rect 40204 8000 40244 8800
rect 40148 7960 40244 8000
rect 40300 8000 40340 10975
rect 40588 10772 40628 10781
rect 40396 10184 40436 10193
rect 40396 9512 40436 10144
rect 40588 9689 40628 10732
rect 40780 10184 40820 11488
rect 41356 11479 41396 11488
rect 40875 11108 40917 11117
rect 40875 11068 40876 11108
rect 40916 11068 40917 11108
rect 40875 11059 40917 11068
rect 43659 11108 43701 11117
rect 43659 11068 43660 11108
rect 43700 11068 43701 11108
rect 43659 11059 43701 11068
rect 40780 10135 40820 10144
rect 40587 9680 40629 9689
rect 40587 9640 40588 9680
rect 40628 9640 40629 9680
rect 40587 9631 40629 9640
rect 40780 9512 40820 9521
rect 40396 9472 40780 9512
rect 40684 8849 40724 9472
rect 40780 9463 40820 9472
rect 40876 9344 40916 11059
rect 43660 10974 43700 11059
rect 43852 11024 43892 11033
rect 44044 11024 44084 13000
rect 44140 11024 44180 11033
rect 43892 10984 43988 11024
rect 44044 10984 44140 11024
rect 43852 10975 43892 10984
rect 41163 10772 41205 10781
rect 41163 10732 41164 10772
rect 41204 10732 41205 10772
rect 41163 10723 41205 10732
rect 41164 9596 41204 10723
rect 43948 10436 43988 10984
rect 44140 10975 44180 10984
rect 45004 11024 45044 11033
rect 44331 10772 44373 10781
rect 44331 10732 44332 10772
rect 44372 10732 44373 10772
rect 44331 10723 44373 10732
rect 44332 10638 44372 10723
rect 44140 10436 44180 10445
rect 43948 10396 44140 10436
rect 44140 10387 44180 10396
rect 45004 9689 45044 10984
rect 45292 10184 45332 13159
rect 47116 13074 47156 13159
rect 49324 13074 49364 13159
rect 45963 13040 46005 13049
rect 45963 13000 45964 13040
rect 46004 13000 46005 13040
rect 45963 12991 46005 13000
rect 46827 13040 46869 13049
rect 46827 13000 46828 13040
rect 46868 13000 46869 13040
rect 46827 12991 46869 13000
rect 45964 12906 46004 12991
rect 46828 11696 46868 12991
rect 48472 12116 48840 12125
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48472 12067 48840 12076
rect 46828 11647 46868 11656
rect 47500 11528 47540 11537
rect 46924 11488 47500 11528
rect 46156 10184 46196 10193
rect 45292 10135 45332 10144
rect 45868 10144 46156 10184
rect 41355 9680 41397 9689
rect 41355 9640 41356 9680
rect 41396 9640 41397 9680
rect 41355 9631 41397 9640
rect 45003 9680 45045 9689
rect 45003 9640 45004 9680
rect 45044 9640 45045 9680
rect 45003 9631 45045 9640
rect 41164 9547 41204 9556
rect 41356 9512 41396 9631
rect 41356 9463 41396 9472
rect 41547 9512 41589 9521
rect 41547 9472 41548 9512
rect 41588 9472 41589 9512
rect 41547 9463 41589 9472
rect 41548 9378 41588 9463
rect 40780 9304 40916 9344
rect 40683 8840 40725 8849
rect 40683 8800 40684 8840
rect 40724 8800 40725 8840
rect 40683 8791 40725 8800
rect 40587 8756 40629 8765
rect 40587 8716 40588 8756
rect 40628 8716 40629 8756
rect 40587 8707 40629 8716
rect 40588 8622 40628 8707
rect 40780 8672 40820 9304
rect 41452 9260 41492 9269
rect 40780 8623 40820 8632
rect 40876 9220 41452 9260
rect 40876 8672 40916 9220
rect 41452 9211 41492 9220
rect 41547 8840 41589 8849
rect 41547 8800 41548 8840
rect 41588 8800 41589 8840
rect 41547 8791 41589 8800
rect 40876 8623 40916 8632
rect 40396 8000 40436 8009
rect 40300 7960 40396 8000
rect 40108 7951 40148 7960
rect 40396 7951 40436 7960
rect 40204 7160 40244 7169
rect 40011 6992 40053 7001
rect 40011 6952 40012 6992
rect 40052 6952 40053 6992
rect 40011 6943 40053 6952
rect 39820 6607 39860 6616
rect 39339 6488 39381 6497
rect 39339 6448 39340 6488
rect 39380 6448 39381 6488
rect 39339 6439 39381 6448
rect 38764 6355 38804 6364
rect 39340 6354 39380 6439
rect 38571 6320 38613 6329
rect 37900 6280 38132 6320
rect 37707 6236 37749 6245
rect 37707 6196 37708 6236
rect 37748 6196 37749 6236
rect 37707 6187 37749 6196
rect 36555 5648 36597 5657
rect 36555 5608 36556 5648
rect 36596 5608 36597 5648
rect 36555 5599 36597 5608
rect 37708 5648 37748 6187
rect 37708 5599 37748 5608
rect 38092 5648 38132 6280
rect 38571 6280 38572 6320
rect 38612 6280 38613 6320
rect 38571 6271 38613 6280
rect 39628 6320 39668 6329
rect 38092 5599 38132 5608
rect 38956 5648 38996 5657
rect 38956 4892 38996 5608
rect 39628 4901 39668 6280
rect 39243 4892 39285 4901
rect 38956 4852 39244 4892
rect 39284 4852 39285 4892
rect 39243 4843 39285 4852
rect 39627 4892 39669 4901
rect 39627 4852 39628 4892
rect 39668 4852 39669 4892
rect 39627 4843 39669 4852
rect 38955 4220 38997 4229
rect 38955 4180 38956 4220
rect 38996 4180 38997 4220
rect 38955 4171 38997 4180
rect 38284 4136 38324 4145
rect 37995 3800 38037 3809
rect 37995 3760 37996 3800
rect 38036 3760 38037 3800
rect 37995 3751 38037 3760
rect 35787 3632 35829 3641
rect 35787 3592 35788 3632
rect 35828 3592 35829 3632
rect 35787 3583 35829 3592
rect 35788 3498 35828 3583
rect 33771 2708 33813 2717
rect 33771 2668 33772 2708
rect 33812 2668 33813 2708
rect 33771 2659 33813 2668
rect 35499 2708 35541 2717
rect 35499 2668 35500 2708
rect 35540 2668 35541 2708
rect 35499 2659 35541 2668
rect 37131 2708 37173 2717
rect 37131 2668 37132 2708
rect 37172 2668 37173 2708
rect 37131 2659 37173 2668
rect 18700 2575 18740 2584
rect 36747 2624 36789 2633
rect 36747 2584 36748 2624
rect 36788 2584 36789 2624
rect 36747 2575 36789 2584
rect 37132 2624 37172 2659
rect 11692 2490 11732 2575
rect 12171 2540 12213 2549
rect 12171 2500 12172 2540
rect 12212 2500 12213 2540
rect 12171 2491 12213 2500
rect 12172 2406 12212 2491
rect 14092 2490 14132 2575
rect 17452 2540 17492 2549
rect 17492 2500 17780 2540
rect 17452 2491 17492 2500
rect 16492 2456 16532 2465
rect 16532 2416 17108 2456
rect 16492 2407 16532 2416
rect 11307 2120 11349 2129
rect 11307 2080 11308 2120
rect 11348 2080 11349 2120
rect 11307 2071 11349 2080
rect 9580 1903 9620 1912
rect 17068 1952 17108 2416
rect 17740 2120 17780 2500
rect 36748 2490 36788 2575
rect 37132 2573 37172 2584
rect 37996 2624 38036 3751
rect 38284 3641 38324 4096
rect 38956 4086 38996 4171
rect 39244 3809 39284 4843
rect 40012 4136 40052 6943
rect 40108 5900 40148 5909
rect 40204 5900 40244 7120
rect 40148 5860 40244 5900
rect 40108 5851 40148 5860
rect 41548 5060 41588 8791
rect 45868 8681 45908 10144
rect 46156 10135 46196 10144
rect 46924 10184 46964 11488
rect 47500 11479 47540 11488
rect 49612 11192 49652 13831
rect 50476 13469 50516 15520
rect 52780 15560 52820 15571
rect 52780 15485 52820 15520
rect 51627 15476 51669 15485
rect 51627 15436 51628 15476
rect 51668 15436 51669 15476
rect 51627 15427 51669 15436
rect 52779 15476 52821 15485
rect 52779 15436 52780 15476
rect 52820 15436 52821 15476
rect 52779 15427 52821 15436
rect 53451 15476 53493 15485
rect 53451 15436 53452 15476
rect 53492 15436 53493 15476
rect 53451 15427 53493 15436
rect 51628 15342 51668 15427
rect 51435 15308 51477 15317
rect 51435 15268 51436 15308
rect 51476 15268 51477 15308
rect 51435 15259 51477 15268
rect 52107 15308 52149 15317
rect 52107 15268 52108 15308
rect 52148 15268 52149 15308
rect 52107 15259 52149 15268
rect 51244 14720 51284 14729
rect 51244 14309 51284 14680
rect 51436 14720 51476 15259
rect 52108 15174 52148 15259
rect 52588 14804 52628 14813
rect 52300 14764 52588 14804
rect 51436 14671 51476 14680
rect 52203 14720 52245 14729
rect 52203 14680 52204 14720
rect 52244 14680 52245 14720
rect 52203 14671 52245 14680
rect 52300 14720 52340 14764
rect 52588 14755 52628 14764
rect 52300 14671 52340 14680
rect 52779 14720 52821 14729
rect 52779 14680 52780 14720
rect 52820 14680 52821 14720
rect 52779 14671 52821 14680
rect 52876 14720 52916 14731
rect 51339 14636 51381 14645
rect 51339 14596 51340 14636
rect 51380 14596 51381 14636
rect 51339 14587 51381 14596
rect 51340 14502 51380 14587
rect 51627 14552 51669 14561
rect 51627 14512 51628 14552
rect 51668 14512 51669 14552
rect 51627 14503 51669 14512
rect 51628 14418 51668 14503
rect 51243 14300 51285 14309
rect 51243 14260 51244 14300
rect 51284 14260 51285 14300
rect 51243 14251 51285 14260
rect 51243 14132 51285 14141
rect 51243 14092 51244 14132
rect 51284 14092 51285 14132
rect 51243 14083 51285 14092
rect 51244 14048 51284 14083
rect 52012 14048 52052 14057
rect 51244 13997 51284 14008
rect 51820 14008 52012 14048
rect 50571 13796 50613 13805
rect 50571 13756 50572 13796
rect 50612 13756 50613 13796
rect 50571 13747 50613 13756
rect 50572 13662 50612 13747
rect 49995 13460 50037 13469
rect 49995 13420 49996 13460
rect 50036 13420 50037 13460
rect 49995 13411 50037 13420
rect 50475 13460 50517 13469
rect 50475 13420 50476 13460
rect 50516 13420 50517 13460
rect 50475 13411 50517 13420
rect 51820 13460 51860 14008
rect 52012 13999 52052 14008
rect 51820 13411 51860 13420
rect 49996 13326 50036 13411
rect 52204 13301 52244 14671
rect 52780 14586 52820 14671
rect 52876 14645 52916 14680
rect 52875 14636 52917 14645
rect 52875 14596 52876 14636
rect 52916 14596 52917 14636
rect 52875 14587 52917 14596
rect 52683 14300 52725 14309
rect 52683 14260 52684 14300
rect 52724 14260 52725 14300
rect 52683 14251 52725 14260
rect 53067 14300 53109 14309
rect 53067 14260 53068 14300
rect 53108 14260 53109 14300
rect 53067 14251 53109 14260
rect 52684 14216 52724 14251
rect 52684 14165 52724 14176
rect 52875 14132 52917 14141
rect 52972 14132 53012 14141
rect 52875 14092 52876 14132
rect 52916 14092 52972 14132
rect 52875 14083 52917 14092
rect 52972 14083 53012 14092
rect 53068 14048 53108 14251
rect 53068 13999 53108 14008
rect 53452 14048 53492 15427
rect 54796 14729 54836 17200
rect 54988 17191 55028 17200
rect 54892 17072 54932 17081
rect 54892 16988 54932 17032
rect 56428 17072 56468 17081
rect 55276 16988 55316 16997
rect 54892 16948 55276 16988
rect 55276 16939 55316 16948
rect 55947 15812 55989 15821
rect 55947 15772 55948 15812
rect 55988 15772 55989 15812
rect 55947 15763 55989 15772
rect 54795 14720 54837 14729
rect 54795 14680 54796 14720
rect 54836 14680 54837 14720
rect 54795 14671 54837 14680
rect 55948 14216 55988 15763
rect 55948 14167 55988 14176
rect 56331 14132 56373 14141
rect 56331 14092 56332 14132
rect 56372 14092 56373 14132
rect 56331 14083 56373 14092
rect 53452 13999 53492 14008
rect 54604 14048 54644 14057
rect 52971 13460 53013 13469
rect 52971 13420 52972 13460
rect 53012 13420 53013 13460
rect 54604 13460 54644 14008
rect 55468 14048 55508 14057
rect 54892 13460 54932 13469
rect 54604 13420 54892 13460
rect 52971 13411 53013 13420
rect 54892 13411 54932 13420
rect 52203 13292 52245 13301
rect 52203 13252 52204 13292
rect 52244 13252 52245 13292
rect 52203 13243 52245 13252
rect 52875 13292 52917 13301
rect 52875 13252 52876 13292
rect 52916 13252 52917 13292
rect 52875 13243 52917 13252
rect 50283 13208 50325 13217
rect 50283 13168 50284 13208
rect 50324 13168 50325 13208
rect 50283 13159 50325 13168
rect 52299 13208 52341 13217
rect 52299 13168 52300 13208
rect 52340 13168 52341 13208
rect 52299 13159 52341 13168
rect 50284 13074 50324 13159
rect 49712 12872 50080 12881
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 49712 12823 50080 12832
rect 49712 11360 50080 11369
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 49712 11311 50080 11320
rect 49612 11152 49940 11192
rect 48472 10604 48840 10613
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48472 10555 48840 10564
rect 47019 10268 47061 10277
rect 48172 10268 48212 10277
rect 47019 10228 47020 10268
rect 47060 10228 47061 10268
rect 47019 10219 47061 10228
rect 47980 10228 48172 10268
rect 46539 10100 46581 10109
rect 46539 10060 46540 10100
rect 46580 10060 46581 10100
rect 46539 10051 46581 10060
rect 46540 9966 46580 10051
rect 46924 9848 46964 10144
rect 47020 10134 47060 10219
rect 47115 10184 47157 10193
rect 47115 10144 47116 10184
rect 47156 10144 47157 10184
rect 47115 10135 47157 10144
rect 47883 10184 47925 10193
rect 47883 10144 47884 10184
rect 47924 10144 47925 10184
rect 47883 10135 47925 10144
rect 47980 10184 48020 10228
rect 48172 10219 48212 10228
rect 48459 10268 48501 10277
rect 48459 10228 48460 10268
rect 48500 10228 48501 10268
rect 48459 10219 48501 10228
rect 47980 10135 48020 10144
rect 48460 10184 48500 10219
rect 47116 10050 47156 10135
rect 47307 10100 47349 10109
rect 47307 10060 47308 10100
rect 47348 10060 47349 10100
rect 47307 10051 47349 10060
rect 47308 9966 47348 10051
rect 46924 9808 47348 9848
rect 47211 9680 47253 9689
rect 47211 9640 47212 9680
rect 47252 9640 47253 9680
rect 47211 9631 47253 9640
rect 47212 9546 47252 9631
rect 47308 9512 47348 9808
rect 47884 9680 47924 10135
rect 48460 10133 48500 10144
rect 48555 10184 48597 10193
rect 48555 10144 48556 10184
rect 48596 10144 48597 10184
rect 48555 10135 48597 10144
rect 49803 10184 49845 10193
rect 49803 10144 49804 10184
rect 49844 10144 49845 10184
rect 49803 10135 49845 10144
rect 49900 10184 49940 11152
rect 52300 10436 52340 13159
rect 52779 10772 52821 10781
rect 52779 10732 52780 10772
rect 52820 10732 52821 10772
rect 52779 10723 52821 10732
rect 52300 10387 52340 10396
rect 49900 10135 49940 10144
rect 50283 10184 50325 10193
rect 50283 10144 50284 10184
rect 50324 10144 50325 10184
rect 50283 10135 50325 10144
rect 50763 10184 50805 10193
rect 50763 10144 50764 10184
rect 50804 10144 50805 10184
rect 50763 10135 50805 10144
rect 51724 10184 51764 10193
rect 48556 10050 48596 10135
rect 49804 10100 49844 10135
rect 49804 10049 49844 10060
rect 50284 10050 50324 10135
rect 49712 9848 50080 9857
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 49712 9799 50080 9808
rect 47884 9631 47924 9640
rect 47308 9463 47348 9472
rect 47691 9512 47733 9521
rect 48555 9512 48597 9521
rect 47691 9472 47692 9512
rect 47732 9472 47828 9512
rect 47691 9463 47733 9472
rect 47692 9378 47732 9463
rect 47788 8924 47828 9472
rect 48555 9472 48556 9512
rect 48596 9472 48597 9512
rect 48555 9463 48597 9472
rect 48556 9378 48596 9463
rect 48472 9092 48840 9101
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48472 9043 48840 9052
rect 47884 8924 47924 8933
rect 47788 8884 47884 8924
rect 47884 8875 47924 8884
rect 45867 8672 45909 8681
rect 45867 8632 45868 8672
rect 45908 8632 45909 8672
rect 45867 8623 45909 8632
rect 46732 8672 46772 8681
rect 45484 8588 45524 8597
rect 45484 8168 45524 8548
rect 45868 8538 45908 8623
rect 45580 8168 45620 8177
rect 45484 8128 45580 8168
rect 45580 8119 45620 8128
rect 46252 8000 46292 8009
rect 45388 7960 46252 8000
rect 45292 6656 45332 6665
rect 45388 6656 45428 7960
rect 46252 7951 46292 7960
rect 45332 6616 45428 6656
rect 45292 6607 45332 6616
rect 44812 6488 44852 6497
rect 44812 5657 44852 6448
rect 45195 6488 45237 6497
rect 45195 6448 45196 6488
rect 45236 6448 45237 6488
rect 45195 6439 45237 6448
rect 45580 6488 45620 6497
rect 45196 6354 45236 6439
rect 45580 6320 45620 6448
rect 46251 6488 46293 6497
rect 46251 6448 46252 6488
rect 46292 6448 46293 6488
rect 46251 6439 46293 6448
rect 46443 6488 46485 6497
rect 46443 6448 46444 6488
rect 46484 6448 46485 6488
rect 46443 6439 46485 6448
rect 46252 6354 46292 6439
rect 45388 6280 45620 6320
rect 43659 5648 43701 5657
rect 43659 5608 43660 5648
rect 43700 5608 43701 5648
rect 43659 5599 43701 5608
rect 44811 5648 44853 5657
rect 44811 5608 44812 5648
rect 44852 5608 44853 5648
rect 44811 5599 44853 5608
rect 45291 5648 45333 5657
rect 45291 5608 45292 5648
rect 45332 5608 45333 5648
rect 45291 5599 45333 5608
rect 43660 5144 43700 5599
rect 45292 5514 45332 5599
rect 43660 5095 43700 5104
rect 45388 5060 45428 6280
rect 46444 5648 46484 6439
rect 46444 5599 46484 5608
rect 46539 5648 46581 5657
rect 46539 5608 46540 5648
rect 46580 5608 46581 5648
rect 46539 5599 46581 5608
rect 46636 5648 46676 5659
rect 45963 5564 46005 5573
rect 45963 5524 45964 5564
rect 46004 5524 46005 5564
rect 45963 5515 46005 5524
rect 45964 5430 46004 5515
rect 46540 5514 46580 5599
rect 46636 5573 46676 5608
rect 46635 5564 46677 5573
rect 46635 5524 46636 5564
rect 46676 5524 46677 5564
rect 46635 5515 46677 5524
rect 41548 5020 41684 5060
rect 41260 4976 41300 4985
rect 40684 4936 41260 4976
rect 40684 4388 40724 4936
rect 41260 4927 41300 4936
rect 41644 4976 41684 5020
rect 45292 5020 45428 5060
rect 41644 4927 41684 4936
rect 42507 4976 42549 4985
rect 42507 4936 42508 4976
rect 42548 4936 42549 4976
rect 42507 4927 42549 4936
rect 42508 4842 42548 4927
rect 45292 4892 45332 5020
rect 45292 4843 45332 4852
rect 46444 4976 46484 4985
rect 46732 4976 46772 8632
rect 47115 8672 47157 8681
rect 47115 8632 47116 8672
rect 47156 8632 47157 8672
rect 47115 8623 47157 8632
rect 47116 7169 47156 8623
rect 49712 8336 50080 8345
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 49712 8287 50080 8296
rect 48472 7580 48840 7589
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48472 7531 48840 7540
rect 50764 7412 50804 10135
rect 51724 8009 51764 10144
rect 52780 10184 52820 10723
rect 52780 10135 52820 10144
rect 51819 9680 51861 9689
rect 51819 9640 51820 9680
rect 51860 9640 51861 9680
rect 51819 9631 51861 9640
rect 51820 9546 51860 9631
rect 52300 9512 52340 9521
rect 52876 9512 52916 13243
rect 52972 13208 53012 13411
rect 53835 13292 53877 13301
rect 53835 13252 53836 13292
rect 53876 13252 53877 13292
rect 53835 13243 53877 13252
rect 52972 13159 53012 13168
rect 53836 13208 53876 13243
rect 53836 13157 53876 13168
rect 54603 13208 54645 13217
rect 54603 13168 54604 13208
rect 54644 13168 54645 13208
rect 54603 13159 54645 13168
rect 54220 13124 54260 13133
rect 54260 13084 54548 13124
rect 54220 13075 54260 13084
rect 54508 12704 54548 13084
rect 54604 13074 54644 13159
rect 55083 13040 55125 13049
rect 55083 13000 55084 13040
rect 55124 13000 55125 13040
rect 55083 12991 55125 13000
rect 55084 12906 55124 12991
rect 54892 12704 54932 12713
rect 54508 12664 54892 12704
rect 54892 12655 54932 12664
rect 55179 12704 55221 12713
rect 55179 12664 55180 12704
rect 55220 12664 55221 12704
rect 55179 12655 55221 12664
rect 55180 12570 55220 12655
rect 55468 12629 55508 14008
rect 55852 14048 55892 14057
rect 55467 12620 55509 12629
rect 55467 12580 55468 12620
rect 55508 12580 55509 12620
rect 55467 12571 55509 12580
rect 55084 12536 55124 12545
rect 55084 11201 55124 12496
rect 54027 11192 54069 11201
rect 54027 11152 54028 11192
rect 54068 11152 54069 11192
rect 54027 11143 54069 11152
rect 54699 11192 54741 11201
rect 54699 11152 54700 11192
rect 54740 11152 54741 11192
rect 54699 11143 54741 11152
rect 55083 11192 55125 11201
rect 55083 11152 55084 11192
rect 55124 11152 55125 11192
rect 55083 11143 55125 11152
rect 55755 11192 55797 11201
rect 55755 11152 55756 11192
rect 55796 11152 55797 11192
rect 55755 11143 55797 11152
rect 54028 10940 54068 11143
rect 54700 11058 54740 11143
rect 55372 11024 55412 11033
rect 54028 10891 54068 10900
rect 55180 10984 55372 11024
rect 53835 10772 53877 10781
rect 53835 10732 53836 10772
rect 53876 10732 53877 10772
rect 53835 10723 53877 10732
rect 53836 10638 53876 10723
rect 55180 10436 55220 10984
rect 55372 10975 55412 10984
rect 55756 11024 55796 11143
rect 55852 11108 55892 14008
rect 56332 13998 56372 14083
rect 56236 13124 56276 13133
rect 56139 13040 56181 13049
rect 56139 13000 56140 13040
rect 56180 13000 56181 13040
rect 56139 12991 56181 13000
rect 55852 11059 55892 11068
rect 55756 10975 55796 10984
rect 55948 11024 55988 11033
rect 55180 10387 55220 10396
rect 54891 10352 54933 10361
rect 54891 10312 54892 10352
rect 54932 10312 54933 10352
rect 54891 10303 54933 10312
rect 55563 10352 55605 10361
rect 55563 10312 55564 10352
rect 55604 10312 55605 10352
rect 55563 10303 55605 10312
rect 53164 10184 53204 10193
rect 54028 10184 54068 10193
rect 53164 9689 53204 10144
rect 53836 10144 54028 10184
rect 53163 9680 53205 9689
rect 53163 9640 53164 9680
rect 53204 9640 53205 9680
rect 53163 9631 53205 9640
rect 53067 9512 53109 9521
rect 52340 9472 52876 9512
rect 52300 9463 52340 9472
rect 52876 9463 52916 9472
rect 52972 9472 53068 9512
rect 53108 9472 53109 9512
rect 51820 9260 51860 9269
rect 50955 8000 50997 8009
rect 50955 7960 50956 8000
rect 50996 7960 50997 8000
rect 50955 7951 50997 7960
rect 51723 8000 51765 8009
rect 51723 7960 51724 8000
rect 51764 7960 51765 8000
rect 51723 7951 51765 7960
rect 50956 7866 50996 7951
rect 50764 7363 50804 7372
rect 51148 7748 51188 7757
rect 47115 7160 47157 7169
rect 47115 7120 47116 7160
rect 47156 7120 47157 7160
rect 47115 7111 47157 7120
rect 48747 7160 48789 7169
rect 48747 7120 48748 7160
rect 48788 7120 48789 7160
rect 48747 7111 48789 7120
rect 49612 7160 49652 7169
rect 46484 4936 46772 4976
rect 47116 4976 47156 7111
rect 48364 7076 48404 7085
rect 48404 7036 48692 7076
rect 48364 7027 48404 7036
rect 48652 6656 48692 7036
rect 48748 7026 48788 7111
rect 48652 6607 48692 6616
rect 47403 6488 47445 6497
rect 47403 6448 47404 6488
rect 47444 6448 47445 6488
rect 47403 6439 47445 6448
rect 47979 6488 48021 6497
rect 47979 6448 47980 6488
rect 48020 6448 48021 6488
rect 47979 6439 48021 6448
rect 47404 5900 47444 6439
rect 47980 6354 48020 6439
rect 48472 6068 48840 6077
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48472 6019 48840 6028
rect 49612 5909 49652 7120
rect 49712 6824 50080 6833
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 49712 6775 50080 6784
rect 51148 6497 51188 7708
rect 51820 7169 51860 9220
rect 51819 7160 51861 7169
rect 51819 7120 51820 7160
rect 51860 7120 51861 7160
rect 51819 7111 51861 7120
rect 51147 6488 51189 6497
rect 51147 6448 51148 6488
rect 51188 6448 51189 6488
rect 51147 6439 51189 6448
rect 47404 5851 47444 5860
rect 48363 5900 48405 5909
rect 48363 5860 48364 5900
rect 48404 5860 48405 5900
rect 48363 5851 48405 5860
rect 49611 5900 49653 5909
rect 49611 5860 49612 5900
rect 49652 5860 49653 5900
rect 49611 5851 49653 5860
rect 48364 5766 48404 5851
rect 51148 5657 51188 6439
rect 52204 5732 52244 5741
rect 52108 5692 52204 5732
rect 47211 5648 47253 5657
rect 47211 5608 47212 5648
rect 47252 5608 47253 5648
rect 47211 5599 47253 5608
rect 47308 5648 47348 5657
rect 48651 5648 48693 5657
rect 47348 5608 47636 5648
rect 47308 5599 47348 5608
rect 47212 5514 47252 5599
rect 47308 4976 47348 4985
rect 47116 4936 47308 4976
rect 40684 4339 40724 4348
rect 40203 4220 40245 4229
rect 40203 4180 40204 4220
rect 40244 4180 40245 4220
rect 40203 4171 40245 4180
rect 40491 4220 40533 4229
rect 40491 4180 40492 4220
rect 40532 4180 40533 4220
rect 40491 4171 40533 4180
rect 40012 4087 40052 4096
rect 40107 4136 40149 4145
rect 40107 4096 40108 4136
rect 40148 4096 40149 4136
rect 40107 4087 40149 4096
rect 40204 4136 40244 4171
rect 40108 4002 40148 4087
rect 40204 4085 40244 4096
rect 40492 4136 40532 4171
rect 40492 4085 40532 4096
rect 41068 4136 41108 4145
rect 40396 3968 40436 3977
rect 39243 3800 39285 3809
rect 39243 3760 39244 3800
rect 39284 3760 39285 3800
rect 39243 3751 39285 3760
rect 38283 3632 38325 3641
rect 38283 3592 38284 3632
rect 38324 3592 38325 3632
rect 38283 3583 38325 3592
rect 40299 3548 40341 3557
rect 40299 3508 40300 3548
rect 40340 3508 40341 3548
rect 40299 3499 40341 3508
rect 38860 3464 38900 3473
rect 38379 3380 38421 3389
rect 38379 3340 38380 3380
rect 38420 3340 38421 3380
rect 38379 3331 38421 3340
rect 38380 3246 38420 3331
rect 38188 3212 38228 3221
rect 38188 2633 38228 3172
rect 38860 2876 38900 3424
rect 40011 3464 40053 3473
rect 40011 3424 40012 3464
rect 40052 3424 40053 3464
rect 40011 3415 40053 3424
rect 40204 3464 40244 3475
rect 39531 3380 39573 3389
rect 39531 3340 39532 3380
rect 39572 3340 39573 3380
rect 39531 3331 39573 3340
rect 40012 3380 40052 3415
rect 40204 3389 40244 3424
rect 40300 3414 40340 3499
rect 40396 3473 40436 3928
rect 40587 3800 40629 3809
rect 40587 3760 40588 3800
rect 40628 3760 40629 3800
rect 40587 3751 40629 3760
rect 40395 3464 40437 3473
rect 40395 3424 40396 3464
rect 40436 3424 40437 3464
rect 40395 3415 40437 3424
rect 39532 3246 39572 3331
rect 40012 3329 40052 3340
rect 40203 3380 40245 3389
rect 40203 3340 40204 3380
rect 40244 3340 40245 3380
rect 40203 3331 40245 3340
rect 40396 3330 40436 3415
rect 39820 3212 39860 3221
rect 39628 3172 39820 3212
rect 39148 2876 39188 2885
rect 38860 2836 39148 2876
rect 39148 2827 39188 2836
rect 37996 2575 38036 2584
rect 38187 2624 38229 2633
rect 38187 2584 38188 2624
rect 38228 2584 38229 2624
rect 38187 2575 38229 2584
rect 39340 2624 39380 2633
rect 39628 2624 39668 3172
rect 39820 3163 39860 3172
rect 39380 2584 39668 2624
rect 39723 2624 39765 2633
rect 39723 2584 39724 2624
rect 39764 2584 39765 2624
rect 39340 2575 39380 2584
rect 39723 2575 39765 2584
rect 40588 2624 40628 3751
rect 41068 3557 41108 4096
rect 41355 4136 41397 4145
rect 41355 4096 41356 4136
rect 41396 4096 41397 4136
rect 41355 4087 41397 4096
rect 41356 4002 41396 4087
rect 41548 3968 41588 3977
rect 41643 3968 41685 3977
rect 41588 3928 41644 3968
rect 41684 3928 41685 3968
rect 41548 3919 41588 3928
rect 41643 3919 41685 3928
rect 44043 3968 44085 3977
rect 44043 3928 44044 3968
rect 44084 3928 44085 3968
rect 44043 3919 44085 3928
rect 41067 3548 41109 3557
rect 41067 3508 41068 3548
rect 41108 3508 41109 3548
rect 41067 3499 41109 3508
rect 40971 3464 41013 3473
rect 40971 3424 40972 3464
rect 41012 3424 41013 3464
rect 40971 3415 41013 3424
rect 41644 3464 41684 3473
rect 40972 3330 41012 3415
rect 41644 2876 41684 3424
rect 41740 2876 41780 2885
rect 41644 2836 41740 2876
rect 41740 2827 41780 2836
rect 40588 2575 40628 2584
rect 44044 2624 44084 3919
rect 46444 3809 46484 4936
rect 45291 3800 45333 3809
rect 45291 3760 45292 3800
rect 45332 3760 45333 3800
rect 45291 3751 45333 3760
rect 46443 3800 46485 3809
rect 46443 3760 46444 3800
rect 46484 3760 46485 3800
rect 46443 3751 46485 3760
rect 44044 2575 44084 2584
rect 44427 2624 44469 2633
rect 44427 2584 44428 2624
rect 44468 2584 44469 2624
rect 44427 2575 44469 2584
rect 45292 2624 45332 3751
rect 47115 3464 47157 3473
rect 47115 3424 47116 3464
rect 47156 3424 47157 3464
rect 47115 3415 47157 3424
rect 46443 2876 46485 2885
rect 46443 2836 46444 2876
rect 46484 2836 46485 2876
rect 46443 2827 46485 2836
rect 47116 2876 47156 3415
rect 47116 2827 47156 2836
rect 46444 2742 46484 2827
rect 47308 2633 47348 4936
rect 47596 3632 47636 5608
rect 48651 5608 48652 5648
rect 48692 5608 48693 5648
rect 48651 5599 48693 5608
rect 51147 5648 51189 5657
rect 51147 5608 51148 5648
rect 51188 5608 51189 5648
rect 51147 5599 51189 5608
rect 48652 5514 48692 5599
rect 48172 5480 48212 5489
rect 48212 5440 48308 5480
rect 48172 5431 48212 5440
rect 47691 5060 47733 5069
rect 47691 5020 47692 5060
rect 47732 5020 47733 5060
rect 47691 5011 47733 5020
rect 47692 4926 47732 5011
rect 48268 3809 48308 5440
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 51915 5060 51957 5069
rect 51915 5020 51916 5060
rect 51956 5020 51957 5060
rect 51915 5011 51957 5020
rect 51916 4926 51956 5011
rect 52108 4985 52148 5692
rect 52204 5683 52244 5692
rect 52972 5648 53012 9472
rect 53067 9463 53109 9472
rect 53068 9378 53108 9463
rect 53739 6656 53781 6665
rect 53739 6616 53740 6656
rect 53780 6616 53781 6656
rect 53739 6607 53781 6616
rect 53740 6488 53780 6607
rect 53740 6439 53780 6448
rect 52588 5564 52628 5573
rect 52396 5480 52436 5489
rect 52588 5480 52628 5524
rect 52436 5440 52628 5480
rect 52396 5431 52436 5440
rect 52204 5144 52244 5153
rect 52107 4976 52149 4985
rect 52107 4936 52108 4976
rect 52148 4936 52149 4976
rect 52107 4927 52149 4936
rect 52108 4842 52148 4927
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 48267 3800 48309 3809
rect 48267 3760 48268 3800
rect 48308 3760 48309 3800
rect 48267 3751 48309 3760
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 47596 3583 47636 3592
rect 47691 3464 47733 3473
rect 47691 3424 47692 3464
rect 47732 3424 47733 3464
rect 47691 3415 47733 3424
rect 48076 3464 48116 3473
rect 47692 3330 47732 3415
rect 48076 2885 48116 3424
rect 48075 2876 48117 2885
rect 48075 2836 48076 2876
rect 48116 2836 48117 2876
rect 48075 2827 48117 2836
rect 45292 2575 45332 2584
rect 47307 2624 47349 2633
rect 47307 2584 47308 2624
rect 47348 2584 47349 2624
rect 47307 2575 47349 2584
rect 48268 2624 48308 3751
rect 52204 3716 52244 5104
rect 52972 4649 53012 5608
rect 53068 6320 53108 6329
rect 53068 4985 53108 6280
rect 53836 6236 53876 10144
rect 54028 10135 54068 10144
rect 54892 9596 54932 10303
rect 55564 10218 55604 10303
rect 55948 10277 55988 10984
rect 55755 10268 55797 10277
rect 55755 10228 55756 10268
rect 55796 10228 55797 10268
rect 55755 10219 55797 10228
rect 55947 10268 55989 10277
rect 55947 10228 55948 10268
rect 55988 10228 55989 10268
rect 55947 10219 55989 10228
rect 55756 10134 55796 10219
rect 54892 9547 54932 9556
rect 55275 9512 55317 9521
rect 55275 9472 55276 9512
rect 55316 9472 55317 9512
rect 55275 9463 55317 9472
rect 56140 9512 56180 12991
rect 56236 12704 56276 13084
rect 56428 13049 56468 17032
rect 57292 17072 57332 17081
rect 57004 14804 57044 14813
rect 57004 14561 57044 14764
rect 56812 14552 56852 14561
rect 56812 14141 56852 14512
rect 57003 14552 57045 14561
rect 57003 14512 57004 14552
rect 57044 14512 57045 14552
rect 57003 14503 57045 14512
rect 56811 14132 56853 14141
rect 56811 14092 56812 14132
rect 56852 14092 56853 14132
rect 56811 14083 56853 14092
rect 56716 14048 56756 14059
rect 56716 13973 56756 14008
rect 56715 13964 56757 13973
rect 56620 13924 56716 13964
rect 56756 13924 56757 13964
rect 56620 13208 56660 13924
rect 56715 13915 56757 13924
rect 56620 13159 56660 13168
rect 56427 13040 56469 13049
rect 56427 13000 56428 13040
rect 56468 13000 56469 13040
rect 56427 12991 56469 13000
rect 56236 12655 56276 12664
rect 56427 12704 56469 12713
rect 56427 12664 56428 12704
rect 56468 12664 56469 12704
rect 56427 12655 56469 12664
rect 56428 12536 56468 12655
rect 56715 12620 56757 12629
rect 56715 12580 56716 12620
rect 56756 12580 56757 12620
rect 56715 12571 56757 12580
rect 56620 12536 56660 12545
rect 56428 12496 56620 12536
rect 56428 12452 56468 12496
rect 56620 12487 56660 12496
rect 56716 12486 56756 12571
rect 56812 12536 56852 12545
rect 57004 12536 57044 14503
rect 57292 13973 57332 17032
rect 57676 17072 57716 17081
rect 57676 15821 57716 17032
rect 63592 16652 63960 16661
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63592 16603 63960 16612
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 93832 16652 94200 16661
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 93832 16603 94200 16612
rect 64832 15896 65200 15905
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 64832 15847 65200 15856
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 95072 15896 95440 15905
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95072 15847 95440 15856
rect 57675 15812 57717 15821
rect 57675 15772 57676 15812
rect 57716 15772 57717 15812
rect 57675 15763 57717 15772
rect 63592 15140 63960 15149
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63592 15091 63960 15100
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 93832 15140 94200 15149
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 93832 15091 94200 15100
rect 58636 14720 58676 14729
rect 57963 14552 58005 14561
rect 57963 14512 57964 14552
rect 58004 14512 58005 14552
rect 57963 14503 58005 14512
rect 57964 14418 58004 14503
rect 58636 14216 58676 14680
rect 64832 14384 65200 14393
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 64832 14335 65200 14344
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 95072 14384 95440 14393
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95072 14335 95440 14344
rect 58732 14216 58772 14225
rect 58636 14176 58732 14216
rect 58732 14167 58772 14176
rect 57580 14048 57620 14057
rect 57484 14008 57580 14048
rect 57291 13964 57333 13973
rect 57291 13924 57292 13964
rect 57332 13924 57333 13964
rect 57291 13915 57333 13924
rect 57484 13208 57524 14008
rect 57580 13999 57620 14008
rect 63592 13628 63960 13637
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63592 13579 63960 13588
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 93832 13628 94200 13637
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 93832 13579 94200 13588
rect 57484 13049 57524 13168
rect 57483 13040 57525 13049
rect 58636 13040 58676 13049
rect 57483 13000 57484 13040
rect 57524 13000 57525 13040
rect 57483 12991 57525 13000
rect 58348 13000 58636 13040
rect 57675 12704 57717 12713
rect 57675 12664 57676 12704
rect 57716 12664 57717 12704
rect 57675 12655 57717 12664
rect 57676 12620 57716 12655
rect 57676 12569 57716 12580
rect 56852 12496 57044 12536
rect 58348 12536 58388 13000
rect 58636 12991 58676 13000
rect 64832 12872 65200 12881
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 64832 12823 65200 12832
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 95072 12872 95440 12881
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95072 12823 95440 12832
rect 56812 12487 56852 12496
rect 58348 12487 58388 12496
rect 56428 12403 56468 12412
rect 63592 12116 63960 12125
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63592 12067 63960 12076
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 93832 12116 94200 12125
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 93832 12067 94200 12076
rect 64832 11360 65200 11369
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 64832 11311 65200 11320
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 95072 11360 95440 11369
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95072 11311 95440 11320
rect 63592 10604 63960 10613
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63592 10555 63960 10564
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 93832 10604 94200 10613
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 93832 10555 94200 10564
rect 56619 10268 56661 10277
rect 56619 10228 56620 10268
rect 56660 10228 56661 10268
rect 56619 10219 56661 10228
rect 56620 10134 56660 10219
rect 57292 10184 57332 10193
rect 57292 9680 57332 10144
rect 64832 9848 65200 9857
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 64832 9799 65200 9808
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 95072 9848 95440 9857
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95072 9799 95440 9808
rect 57292 9631 57332 9640
rect 56140 9463 56180 9472
rect 55276 9378 55316 9463
rect 63592 9092 63960 9101
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63592 9043 63960 9052
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 93832 9092 94200 9101
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 93832 9043 94200 9052
rect 64832 8336 65200 8345
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 64832 8287 65200 8296
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 95072 8336 95440 8345
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95072 8287 95440 8296
rect 63592 7580 63960 7589
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63592 7531 63960 7540
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 93832 7580 94200 7589
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 93832 7531 94200 7540
rect 64832 6824 65200 6833
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 64832 6775 65200 6784
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 95072 6824 95440 6833
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95072 6775 95440 6784
rect 54987 6656 55029 6665
rect 54987 6616 54988 6656
rect 55028 6616 55029 6656
rect 54987 6607 55029 6616
rect 54027 6488 54069 6497
rect 54027 6448 54028 6488
rect 54068 6448 54069 6488
rect 54027 6439 54069 6448
rect 54028 6354 54068 6439
rect 54316 6320 54356 6329
rect 54124 6280 54316 6320
rect 54124 6236 54164 6280
rect 54316 6271 54356 6280
rect 53836 6196 54164 6236
rect 53836 5648 53876 6196
rect 54988 5900 55028 6607
rect 63592 6068 63960 6077
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63592 6019 63960 6028
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 93832 6068 94200 6077
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 93832 6019 94200 6028
rect 54988 5851 55028 5860
rect 53067 4976 53109 4985
rect 53067 4936 53068 4976
rect 53108 4936 53109 4976
rect 53067 4927 53109 4936
rect 52971 4640 53013 4649
rect 52971 4600 52972 4640
rect 53012 4600 53013 4640
rect 52971 4591 53013 4600
rect 51916 3676 52244 3716
rect 51723 3464 51765 3473
rect 51723 3424 51724 3464
rect 51764 3424 51765 3464
rect 51723 3415 51765 3424
rect 51916 3464 51956 3676
rect 52204 3632 52244 3676
rect 52300 3632 52340 3641
rect 53644 3632 53684 3641
rect 52204 3592 52300 3632
rect 52300 3583 52340 3592
rect 53452 3592 53644 3632
rect 52011 3548 52053 3557
rect 52011 3508 52012 3548
rect 52052 3508 52053 3548
rect 52011 3499 52053 3508
rect 53163 3548 53205 3557
rect 53163 3508 53164 3548
rect 53204 3508 53205 3548
rect 53163 3499 53205 3508
rect 51435 3380 51477 3389
rect 51435 3340 51436 3380
rect 51476 3340 51477 3380
rect 51435 3331 51477 3340
rect 51436 3246 51476 3331
rect 51244 3212 51284 3221
rect 50476 3172 51244 3212
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 49515 2708 49557 2717
rect 49515 2668 49516 2708
rect 49556 2668 49557 2708
rect 49515 2659 49557 2668
rect 48268 2575 48308 2584
rect 49131 2624 49173 2633
rect 49131 2584 49132 2624
rect 49172 2584 49173 2624
rect 49131 2575 49173 2584
rect 49516 2624 49556 2659
rect 39724 2490 39764 2575
rect 44428 2490 44468 2575
rect 49132 2490 49172 2575
rect 49516 2573 49556 2584
rect 50476 2624 50516 3172
rect 51244 3163 51284 3172
rect 50476 2575 50516 2584
rect 50859 2624 50901 2633
rect 50859 2584 50860 2624
rect 50900 2584 50901 2624
rect 50859 2575 50901 2584
rect 51724 2624 51764 3415
rect 51916 3389 51956 3424
rect 52012 3414 52052 3499
rect 52108 3464 52148 3473
rect 51915 3380 51957 3389
rect 51915 3340 51916 3380
rect 51956 3340 51957 3380
rect 51915 3331 51957 3340
rect 51916 3300 51956 3331
rect 52108 2801 52148 3424
rect 52972 3464 53012 3473
rect 52876 2876 52916 2885
rect 52972 2876 53012 3424
rect 53164 3464 53204 3499
rect 53164 3413 53204 3424
rect 52916 2836 53012 2876
rect 52876 2827 52916 2836
rect 52107 2792 52149 2801
rect 52107 2752 52108 2792
rect 52148 2752 52149 2792
rect 52107 2743 52149 2752
rect 53452 2717 53492 3592
rect 53644 3583 53684 3592
rect 53836 3473 53876 5608
rect 56619 5648 56661 5657
rect 56619 5608 56620 5648
rect 56660 5608 56661 5648
rect 56619 5599 56661 5608
rect 57195 5648 57237 5657
rect 57195 5608 57196 5648
rect 57236 5608 57237 5648
rect 57195 5599 57237 5608
rect 56620 5514 56660 5599
rect 54411 5480 54453 5489
rect 54411 5440 54412 5480
rect 54452 5440 54453 5480
rect 54411 5431 54453 5440
rect 55947 5480 55989 5489
rect 55947 5440 55948 5480
rect 55988 5440 55989 5480
rect 55947 5431 55989 5440
rect 54027 4976 54069 4985
rect 54027 4936 54028 4976
rect 54068 4936 54069 4976
rect 54027 4927 54069 4936
rect 54028 4136 54068 4927
rect 54412 4892 54452 5431
rect 55948 5346 55988 5431
rect 54028 4087 54068 4096
rect 54220 4852 54412 4892
rect 54220 4136 54260 4852
rect 54412 4843 54452 4852
rect 54796 4976 54836 4985
rect 54604 4808 54644 4817
rect 54796 4808 54836 4936
rect 54644 4768 54836 4808
rect 55180 4976 55220 4985
rect 54604 4759 54644 4768
rect 55180 4649 55220 4936
rect 56044 4976 56084 4985
rect 54795 4640 54837 4649
rect 54795 4600 54796 4640
rect 54836 4600 54837 4640
rect 54795 4591 54837 4600
rect 55179 4640 55221 4649
rect 55179 4600 55180 4640
rect 55220 4600 55221 4640
rect 55179 4591 55221 4600
rect 54220 4087 54260 4096
rect 54124 4052 54164 4061
rect 53548 3464 53588 3473
rect 53548 3296 53588 3424
rect 53835 3464 53877 3473
rect 53835 3424 53836 3464
rect 53876 3424 53877 3464
rect 53835 3415 53877 3424
rect 54124 3296 54164 4012
rect 53548 3256 54164 3296
rect 54412 3464 54452 3473
rect 54412 2876 54452 3424
rect 54796 3464 54836 4591
rect 55852 3968 55892 3977
rect 54796 3415 54836 3424
rect 55659 3464 55701 3473
rect 55659 3424 55660 3464
rect 55700 3424 55701 3464
rect 55659 3415 55701 3424
rect 55660 3330 55700 3415
rect 54508 2876 54548 2885
rect 54412 2836 54508 2876
rect 54508 2827 54548 2836
rect 55852 2717 55892 3928
rect 56044 3473 56084 4936
rect 57196 4892 57236 5599
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 95072 5312 95440 5321
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95072 5263 95440 5272
rect 57196 4843 57236 4852
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 93832 4556 94200 4565
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 93832 4507 94200 4516
rect 56524 4136 56564 4145
rect 56564 4096 56852 4136
rect 56524 4087 56564 4096
rect 56812 3632 56852 4096
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 95072 3800 95440 3809
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95072 3751 95440 3760
rect 56812 3583 56852 3592
rect 56043 3464 56085 3473
rect 56043 3424 56044 3464
rect 56084 3424 56085 3464
rect 56043 3415 56085 3424
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 93832 3044 94200 3053
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 93832 2995 94200 3004
rect 53451 2708 53493 2717
rect 53451 2668 53452 2708
rect 53492 2668 53493 2708
rect 53451 2659 53493 2668
rect 54699 2708 54741 2717
rect 54699 2668 54700 2708
rect 54740 2668 54741 2708
rect 54699 2659 54741 2668
rect 55851 2708 55893 2717
rect 55851 2668 55852 2708
rect 55892 2668 55893 2708
rect 55851 2659 55893 2668
rect 51724 2575 51764 2584
rect 50860 2490 50900 2575
rect 54700 2574 54740 2659
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 95072 2288 95440 2297
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95072 2239 95440 2248
rect 17740 2071 17780 2080
rect 17068 1903 17108 1912
rect 8428 1819 8468 1828
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 93832 1532 94200 1541
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 93832 1483 94200 1492
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
rect 95072 776 95440 785
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95072 727 95440 736
<< via2 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 268 37528 308 37568
rect 76 36688 116 36728
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 6124 35848 6164 35888
rect 6700 35848 6740 35888
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 6124 35092 6164 35132
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 6700 35176 6740 35216
rect 10540 36604 10580 36644
rect 9676 35764 9716 35804
rect 7276 35092 7316 35132
rect 8812 35176 8852 35216
rect 6700 35008 6740 35048
rect 6988 35008 7028 35048
rect 7564 35008 7604 35048
rect 6316 34588 6356 34628
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 8908 35092 8948 35132
rect 7180 34588 7220 34628
rect 7372 34168 7412 34208
rect 8140 34168 8180 34208
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 3148 32152 3188 32192
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 7180 33580 7220 33620
rect 3820 32152 3860 32192
rect 6316 32152 6356 32192
rect 2380 31396 2420 31436
rect 3532 31396 3572 31436
rect 2284 31312 2324 31352
rect 2956 31312 2996 31352
rect 4012 31396 4052 31436
rect 2668 31060 2708 31100
rect 3532 30640 3572 30680
rect 7660 31312 7700 31352
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 4204 30640 4244 30680
rect 5644 30640 5684 30680
rect 7276 30640 7316 30680
rect 4108 30388 4148 30428
rect 5164 30388 5204 30428
rect 4492 30304 4532 30344
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 6508 30304 6548 30344
rect 3532 28960 3572 29000
rect 4204 28960 4244 29000
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 5068 28960 5108 29000
rect 2668 27616 2708 27656
rect 2284 27448 2324 27488
rect 2380 25852 2420 25892
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 5836 28540 5876 28580
rect 6124 28288 6164 28328
rect 8524 28540 8564 28580
rect 8812 28288 8852 28328
rect 5260 28120 5300 28160
rect 6412 28120 6452 28160
rect 3628 27700 3668 27740
rect 5164 27700 5204 27740
rect 3244 27448 3284 27488
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 3436 26020 3476 26060
rect 3244 25852 3284 25892
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 4300 27616 4340 27656
rect 6700 27700 6740 27740
rect 8620 27700 8660 27740
rect 4684 27028 4724 27068
rect 5260 27028 5300 27068
rect 5644 27028 5684 27068
rect 10540 35764 10580 35804
rect 9100 34168 9140 34208
rect 10444 34168 10484 34208
rect 10060 33580 10100 33620
rect 9004 31312 9044 31352
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 25708 37444 25748 37484
rect 26188 37444 26228 37484
rect 26764 37444 26804 37484
rect 18124 37192 18164 37232
rect 18796 37192 18836 37232
rect 21772 37192 21812 37232
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 16780 36772 16820 36812
rect 17932 36772 17972 36812
rect 12076 36604 12116 36644
rect 11884 36520 11924 36560
rect 13324 36520 13364 36560
rect 16204 36520 16244 36560
rect 17164 36520 17204 36560
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 18220 35932 18260 35972
rect 19084 35932 19124 35972
rect 15820 35764 15860 35804
rect 11884 34336 11924 34376
rect 12268 34336 12308 34376
rect 12460 34336 12500 34376
rect 12172 33580 12212 33620
rect 11404 32656 11444 32696
rect 9676 31312 9716 31352
rect 9676 30388 9716 30428
rect 10540 32152 10580 32192
rect 13132 34000 13172 34040
rect 15628 34000 15668 34040
rect 14476 32824 14516 32864
rect 15532 32824 15572 32864
rect 15724 33580 15764 33620
rect 17068 35848 17108 35888
rect 18028 35848 18068 35888
rect 16876 35764 16916 35804
rect 21868 36772 21908 36812
rect 22252 36688 22292 36728
rect 25132 37192 25172 37232
rect 25516 37192 25556 37232
rect 22636 36772 22676 36812
rect 22540 36604 22580 36644
rect 21964 35848 22004 35888
rect 18028 35176 18068 35216
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 18796 35176 18836 35216
rect 20524 35176 20564 35216
rect 17068 35092 17108 35132
rect 18124 35092 18164 35132
rect 18412 35092 18452 35132
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 16396 33580 16436 33620
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 18124 32908 18164 32948
rect 16396 32824 16436 32864
rect 18028 32824 18068 32864
rect 14860 32656 14900 32696
rect 16204 32656 16244 32696
rect 11116 30388 11156 30428
rect 9772 29128 9812 29168
rect 10444 29128 10484 29168
rect 9484 28960 9524 29000
rect 11404 28960 11444 29000
rect 12460 28960 12500 29000
rect 13036 28960 13076 29000
rect 8908 26776 8948 26816
rect 9484 26776 9524 26816
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 4108 26020 4148 26060
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 268 23248 308 23288
rect 3628 23584 3668 23624
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 4300 23584 4340 23624
rect 4492 23584 4532 23624
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 8812 23752 8852 23792
rect 11020 27532 11060 27572
rect 10060 26776 10100 26816
rect 9868 26272 9908 26312
rect 10060 26272 10100 26312
rect 15916 30136 15956 30176
rect 17452 31900 17492 31940
rect 18028 31900 18068 31940
rect 17548 30220 17588 30260
rect 17932 30220 17972 30260
rect 18028 30136 18068 30176
rect 18220 31900 18260 31940
rect 18700 31900 18740 31940
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 21196 34504 21236 34544
rect 25516 36688 25556 36728
rect 22156 34504 22196 34544
rect 23116 34504 23156 34544
rect 19180 34252 19220 34292
rect 20908 34252 20948 34292
rect 21484 34336 21524 34376
rect 23308 34420 23348 34460
rect 24076 34420 24116 34460
rect 23116 34336 23156 34376
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 21292 34000 21332 34040
rect 22348 34000 22388 34040
rect 18988 32908 19028 32948
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 19180 31900 19220 31940
rect 20140 31900 20180 31940
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 26284 36604 26324 36644
rect 28204 36688 28244 36728
rect 29644 36688 29684 36728
rect 30220 36688 30260 36728
rect 25708 35848 25748 35888
rect 26380 35848 26420 35888
rect 27436 35932 27476 35972
rect 33196 36520 33236 36560
rect 34156 36520 34196 36560
rect 34348 36520 34388 36560
rect 35116 36520 35156 36560
rect 28972 35932 29012 35972
rect 25324 34336 25364 34376
rect 25324 33664 25364 33704
rect 24652 32152 24692 32192
rect 22348 31480 22388 31520
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 13132 28288 13172 28328
rect 14092 28288 14132 28328
rect 12076 27532 12116 27572
rect 13708 27532 13748 27572
rect 13132 26776 13172 26816
rect 18124 30052 18164 30092
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 19180 30052 19220 30092
rect 20332 30724 20372 30764
rect 21964 30724 22004 30764
rect 20140 30136 20180 30176
rect 20044 30052 20084 30092
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 15724 26776 15764 26816
rect 16108 26776 16148 26816
rect 16588 26776 16628 26816
rect 18796 26776 18836 26816
rect 19372 26776 19412 26816
rect 19564 26776 19604 26816
rect 15148 26608 15188 26648
rect 17068 26608 17108 26648
rect 11788 26272 11828 26312
rect 13996 26272 14036 26312
rect 13996 25180 14036 25220
rect 15628 25180 15668 25220
rect 6316 23668 6356 23708
rect 6124 23584 6164 23624
rect 5740 23164 5780 23204
rect 4204 23080 4244 23120
rect 5260 23080 5300 23120
rect 3052 22996 3092 23036
rect 2668 21652 2708 21692
rect 652 21568 692 21608
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 4204 22660 4244 22700
rect 5548 22660 5588 22700
rect 3628 22492 3668 22532
rect 7564 23164 7604 23204
rect 9100 23668 9140 23708
rect 7948 22996 7988 23036
rect 4300 22492 4340 22532
rect 4492 22492 4532 22532
rect 6028 22492 6068 22532
rect 3436 21652 3476 21692
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 652 20728 692 20768
rect 2860 20140 2900 20180
rect 3628 20140 3668 20180
rect 76 20056 116 20096
rect 652 19888 692 19928
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 652 19048 692 19088
rect 1708 19048 1748 19088
rect 2668 19048 2708 19088
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 10060 23752 10100 23792
rect 10348 23752 10388 23792
rect 11500 23584 11540 23624
rect 12844 23584 12884 23624
rect 14764 23752 14804 23792
rect 17260 25264 17300 25304
rect 17836 25264 17876 25304
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 19372 26104 19412 26144
rect 22060 27700 22100 27740
rect 23020 29128 23060 29168
rect 22156 27532 22196 27572
rect 20908 27364 20948 27404
rect 21868 27364 21908 27404
rect 20524 26776 20564 26816
rect 18124 25516 18164 25556
rect 18988 25516 19028 25556
rect 18604 24592 18644 24632
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 19084 24592 19124 24632
rect 16492 23752 16532 23792
rect 18604 23752 18644 23792
rect 12844 23080 12884 23120
rect 10156 22996 10196 23036
rect 9964 22828 10004 22868
rect 11116 22828 11156 22868
rect 13516 22828 13556 22868
rect 13900 22828 13940 22868
rect 11596 22408 11636 22448
rect 4108 20140 4148 20180
rect 9100 20140 9140 20180
rect 9484 20140 9524 20180
rect 9868 20140 9908 20180
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 7468 18712 7508 18752
rect 9964 18712 10004 18752
rect 652 18208 692 18248
rect 2956 18544 2996 18584
rect 3916 18544 3956 18584
rect 5356 18544 5396 18584
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 6796 18460 6836 18500
rect 5644 18292 5684 18332
rect 6604 18292 6644 18332
rect 2092 17704 2132 17744
rect 4492 17704 4532 17744
rect 5356 17704 5396 17744
rect 4108 17620 4148 17660
rect 5260 17620 5300 17660
rect 652 17368 692 17408
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 6028 17788 6068 17828
rect 7948 18544 7988 18584
rect 7660 18460 7700 18500
rect 7660 17956 7700 17996
rect 6988 17704 7028 17744
rect 8044 17704 8084 17744
rect 6028 17116 6068 17156
rect 8812 17956 8852 17996
rect 8332 17704 8372 17744
rect 9484 18544 9524 18584
rect 9004 17704 9044 17744
rect 5452 16948 5492 16988
rect 7372 16948 7412 16988
rect 8236 16948 8276 16988
rect 8428 16948 8468 16988
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 652 16528 692 16568
rect 14476 23080 14516 23120
rect 14092 22408 14132 22448
rect 14092 22240 14132 22280
rect 19372 23752 19412 23792
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 19756 22828 19796 22868
rect 16492 22324 16532 22364
rect 14860 22240 14900 22280
rect 17356 22240 17396 22280
rect 20332 26104 20372 26144
rect 21100 26104 21140 26144
rect 20236 22828 20276 22868
rect 20140 22324 20180 22364
rect 22156 26776 22196 26816
rect 21964 25096 22004 25136
rect 21868 23080 21908 23120
rect 20332 22240 20372 22280
rect 21004 22240 21044 22280
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 14860 21736 14900 21776
rect 15244 21736 15284 21776
rect 13996 20728 14036 20768
rect 14572 20728 14612 20768
rect 13420 20140 13460 20180
rect 12076 18964 12116 19004
rect 13036 18964 13076 19004
rect 11020 18712 11060 18752
rect 11788 18712 11828 18752
rect 12268 18712 12308 18752
rect 11020 17704 11060 17744
rect 10156 17116 10196 17156
rect 10348 16948 10388 16988
rect 11116 17116 11156 17156
rect 11308 17116 11348 17156
rect 11980 17620 12020 17660
rect 12172 17620 12212 17660
rect 12940 17620 12980 17660
rect 11884 16948 11924 16988
rect 12364 16780 12404 16820
rect 9484 16192 9524 16232
rect 13132 16780 13172 16820
rect 12652 16192 12692 16232
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 556 15688 596 15728
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 652 14848 692 14888
rect 9772 14680 9812 14720
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 652 14008 692 14048
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 652 13168 692 13208
rect 2476 13168 2516 13208
rect 2956 13168 2996 13208
rect 2380 12412 2420 12452
rect 652 12328 692 12368
rect 3340 12496 3380 12536
rect 8044 13168 8084 13208
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 3628 12496 3668 12536
rect 3820 12496 3860 12536
rect 3532 12412 3572 12452
rect 2956 12328 2996 12368
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 3532 11740 3572 11780
rect 652 11488 692 11528
rect 3436 11488 3476 11528
rect 652 10648 692 10688
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 3724 12328 3764 12368
rect 940 10060 980 10100
rect 652 9808 692 9848
rect 844 9136 884 9176
rect 652 8968 692 9008
rect 556 8128 596 8168
rect 652 7288 692 7328
rect 652 6448 692 6488
rect 652 5608 692 5648
rect 652 4768 692 4808
rect 2956 9640 2996 9680
rect 3340 9640 3380 9680
rect 2476 9472 2516 9512
rect 2380 8716 2420 8756
rect 3244 9556 3284 9596
rect 3148 9472 3188 9512
rect 3532 9472 3572 9512
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 3052 8716 3092 8756
rect 3916 11740 3956 11780
rect 4012 11656 4052 11696
rect 5164 11656 5204 11696
rect 4108 11488 4148 11528
rect 4300 11488 4340 11528
rect 5356 11488 5396 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 4204 11236 4244 11276
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 4396 9640 4436 9680
rect 5260 9640 5300 9680
rect 4780 9220 4820 9260
rect 3724 8716 3764 8756
rect 3244 8632 3284 8672
rect 3628 8632 3668 8672
rect 3916 8632 3956 8672
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 6604 12412 6644 12452
rect 9772 13168 9812 13208
rect 11692 13168 11732 13208
rect 8620 12580 8660 12620
rect 9196 12580 9236 12620
rect 9868 12580 9908 12620
rect 7180 11320 7220 11360
rect 5452 9556 5492 9596
rect 5548 9220 5588 9260
rect 7180 8800 7220 8840
rect 5164 8716 5204 8756
rect 6028 8632 6068 8672
rect 10732 12496 10772 12536
rect 11692 12580 11732 12620
rect 11212 12412 11252 12452
rect 8716 11320 8756 11360
rect 8044 8800 8084 8840
rect 7756 8716 7796 8756
rect 7468 8632 7508 8672
rect 8332 8632 8372 8672
rect 8620 8632 8660 8672
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 652 3928 692 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 844 3508 884 3548
rect 652 3172 692 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 844 2668 884 2708
rect 10060 9472 10100 9512
rect 9772 8800 9812 8840
rect 9100 8632 9140 8672
rect 11212 9472 11252 9512
rect 10636 8800 10676 8840
rect 12268 13840 12308 13880
rect 12844 13840 12884 13880
rect 12652 13168 12692 13208
rect 13132 13168 13172 13208
rect 14188 20140 14228 20180
rect 19948 21400 19988 21440
rect 21004 21400 21044 21440
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 22252 25264 22292 25304
rect 22828 25264 22868 25304
rect 26284 33664 26324 33704
rect 26956 33664 26996 33704
rect 27244 32824 27284 32864
rect 28108 32824 28148 32864
rect 26188 32152 26228 32192
rect 26092 31480 26132 31520
rect 25996 31312 26036 31352
rect 25804 30724 25844 30764
rect 24364 30640 24404 30680
rect 25324 30640 25364 30680
rect 25132 30388 25172 30428
rect 25708 30388 25748 30428
rect 23308 29128 23348 29168
rect 23212 27700 23252 27740
rect 23404 27700 23444 27740
rect 25132 27700 25172 27740
rect 24844 27616 24884 27656
rect 23404 27532 23444 27572
rect 23308 27448 23348 27488
rect 23788 26020 23828 26060
rect 23212 25264 23252 25304
rect 23308 25096 23348 25136
rect 22444 22324 22484 22364
rect 22444 21568 22484 21608
rect 22732 23080 22772 23120
rect 22924 22240 22964 22280
rect 23212 22240 23252 22280
rect 22828 21568 22868 21608
rect 21100 20812 21140 20852
rect 21964 20812 22004 20852
rect 22924 20728 22964 20768
rect 14284 17620 14324 17660
rect 17260 17032 17300 17072
rect 14668 14008 14708 14048
rect 15148 14008 15188 14048
rect 16396 14008 16436 14048
rect 13516 12496 13556 12536
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 17644 17704 17684 17744
rect 18700 17704 18740 17744
rect 18988 17704 19028 17744
rect 18892 17620 18932 17660
rect 18508 17452 18548 17492
rect 19372 17704 19412 17744
rect 19276 17452 19316 17492
rect 17644 17032 17684 17072
rect 18124 17032 18164 17072
rect 18508 17032 18548 17072
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 18892 14680 18932 14720
rect 18124 14008 18164 14048
rect 18604 14008 18644 14048
rect 18412 13924 18452 13964
rect 17356 13840 17396 13880
rect 18700 13840 18740 13880
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 18700 13336 18740 13376
rect 17260 12496 17300 12536
rect 18508 12496 18548 12536
rect 18796 12580 18836 12620
rect 18796 12412 18836 12452
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 16300 11656 16340 11696
rect 12268 9472 12308 9512
rect 14284 10144 14324 10184
rect 16012 10144 16052 10184
rect 17164 11656 17204 11696
rect 19084 14008 19124 14048
rect 18988 13924 19028 13964
rect 19084 13252 19124 13292
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 21964 18292 22004 18332
rect 22828 18292 22868 18332
rect 20428 17620 20468 17660
rect 21004 17620 21044 17660
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 21772 17620 21812 17660
rect 21868 17452 21908 17492
rect 21388 17032 21428 17072
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 22252 17704 22292 17744
rect 22732 17116 22772 17156
rect 21676 14848 21716 14888
rect 26188 31312 26228 31352
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 37516 36688 37556 36728
rect 38380 36688 38420 36728
rect 35116 35932 35156 35972
rect 37132 35932 37172 35972
rect 33580 35176 33620 35216
rect 34252 35176 34292 35216
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 36940 35344 36980 35384
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 33196 34588 33236 34628
rect 34156 34588 34196 34628
rect 29068 33664 29108 33704
rect 29356 33664 29396 33704
rect 26380 31312 26420 31352
rect 27052 31312 27092 31352
rect 26956 30724 26996 30764
rect 26092 30220 26132 30260
rect 26092 29632 26132 29672
rect 26092 27616 26132 27656
rect 26284 27448 26324 27488
rect 26092 26776 26132 26816
rect 25996 26020 26036 26060
rect 27436 30640 27476 30680
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 34348 34420 34388 34460
rect 36460 35176 36500 35216
rect 36844 35176 36884 35216
rect 37612 35848 37652 35888
rect 38668 35848 38708 35888
rect 39628 35848 39668 35888
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 40684 36856 40724 36896
rect 42124 36856 42164 36896
rect 40972 36688 41012 36728
rect 41548 36688 41588 36728
rect 40108 36604 40148 36644
rect 40684 36604 40724 36644
rect 37612 35344 37652 35384
rect 37324 35260 37364 35300
rect 37228 35176 37268 35216
rect 39052 35176 39092 35216
rect 36460 34420 36500 34460
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 35500 33160 35540 33200
rect 36652 33160 36692 33200
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 34444 32152 34484 32192
rect 35020 32152 35060 32192
rect 34348 32068 34388 32108
rect 28876 30724 28916 30764
rect 28492 30220 28532 30260
rect 26956 29632 26996 29672
rect 28012 29212 28052 29252
rect 28492 29212 28532 29252
rect 28684 29128 28724 29168
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 31084 30724 31124 30764
rect 30988 30640 31028 30680
rect 34732 31228 34772 31268
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 36748 32152 36788 32192
rect 35884 32068 35924 32108
rect 36940 31900 36980 31940
rect 38188 31900 38228 31940
rect 36268 31228 36308 31268
rect 32332 30640 32372 30680
rect 33484 30640 33524 30680
rect 34156 30640 34196 30680
rect 29164 30220 29204 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 29068 29128 29108 29168
rect 30412 29212 30452 29252
rect 28972 26776 29012 26816
rect 25996 25516 26036 25556
rect 26668 25516 26708 25556
rect 29836 26440 29876 26480
rect 31084 29044 31124 29084
rect 32140 29044 32180 29084
rect 32140 26776 32180 26816
rect 31468 26608 31508 26648
rect 32044 26608 32084 26648
rect 30220 26440 30260 26480
rect 29836 26188 29876 26228
rect 30124 26188 30164 26228
rect 30700 26104 30740 26144
rect 31276 26104 31316 26144
rect 30892 25516 30932 25556
rect 27820 25264 27860 25304
rect 25708 23248 25748 23288
rect 26188 23248 26228 23288
rect 23980 23080 24020 23120
rect 24844 23080 24884 23120
rect 23980 22240 24020 22280
rect 26092 20812 26132 20852
rect 26572 20812 26612 20852
rect 26860 20812 26900 20852
rect 24940 20140 24980 20180
rect 25900 20140 25940 20180
rect 23308 19804 23348 19844
rect 23116 17032 23156 17072
rect 23116 14848 23156 14888
rect 26188 20056 26228 20096
rect 25516 18124 25556 18164
rect 25132 17956 25172 17996
rect 23980 17872 24020 17912
rect 24652 17872 24692 17912
rect 23980 17620 24020 17660
rect 23788 17116 23828 17156
rect 25900 17956 25940 17996
rect 26092 17788 26132 17828
rect 26764 18544 26804 18584
rect 29452 23080 29492 23120
rect 29644 23080 29684 23120
rect 29836 22828 29876 22868
rect 30604 22828 30644 22868
rect 30220 22240 30260 22280
rect 31852 25516 31892 25556
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 33292 26776 33332 26816
rect 34156 26188 34196 26228
rect 32140 26104 32180 26144
rect 33196 26104 33236 26144
rect 32812 25348 32852 25388
rect 31756 24592 31796 24632
rect 31660 23080 31700 23120
rect 31276 22240 31316 22280
rect 31564 22240 31604 22280
rect 31276 21736 31316 21776
rect 30220 21568 30260 21608
rect 30700 21568 30740 21608
rect 32236 24592 32276 24632
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 35020 30640 35060 30680
rect 34444 30388 34484 30428
rect 35980 30388 36020 30428
rect 37420 29800 37460 29840
rect 38188 31144 38228 31184
rect 37996 30808 38036 30848
rect 38476 32152 38516 32192
rect 39052 32068 39092 32108
rect 38380 30808 38420 30848
rect 37804 29800 37844 29840
rect 38092 29800 38132 29840
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 37132 26692 37172 26732
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 34924 26188 34964 26228
rect 35788 26104 35828 26144
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 42700 33412 42740 33452
rect 43372 33412 43412 33452
rect 42796 32236 42836 32276
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 42316 31480 42356 31520
rect 42988 31480 43028 31520
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 41932 31144 41972 31184
rect 39052 30724 39092 30764
rect 40684 30724 40724 30764
rect 41164 30724 41204 30764
rect 39436 30640 39476 30680
rect 42028 30472 42068 30512
rect 42700 30640 42740 30680
rect 43468 30640 43508 30680
rect 38668 29800 38708 29840
rect 42412 29800 42452 29840
rect 39532 26860 39572 26900
rect 40396 26860 40436 26900
rect 38188 26692 38228 26732
rect 42604 28960 42644 29000
rect 41740 26188 41780 26228
rect 37516 26020 37556 26060
rect 38380 26020 38420 26060
rect 39724 26020 39764 26060
rect 36940 25852 36980 25892
rect 34540 25348 34580 25388
rect 32044 22996 32084 23036
rect 32524 22996 32564 23036
rect 32524 22324 32564 22364
rect 31852 21736 31892 21776
rect 35020 25264 35060 25304
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 36844 24340 36884 24380
rect 39628 25348 39668 25388
rect 40300 25852 40340 25892
rect 40684 25852 40724 25892
rect 41260 25348 41300 25388
rect 43084 30472 43124 30512
rect 43180 29044 43220 29084
rect 42796 28960 42836 29000
rect 41356 25180 41396 25220
rect 37900 24760 37940 24800
rect 38668 24760 38708 24800
rect 38956 24760 38996 24800
rect 39532 24760 39572 24800
rect 37708 24340 37748 24380
rect 37228 23752 37268 23792
rect 37516 23752 37556 23792
rect 37804 23752 37844 23792
rect 38092 23752 38132 23792
rect 33772 23080 33812 23120
rect 33100 22240 33140 22280
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 33964 22996 34004 23036
rect 33388 22240 33428 22280
rect 33772 21736 33812 21776
rect 35020 23080 35060 23120
rect 37420 22828 37460 22868
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 39052 23248 39092 23288
rect 38764 22828 38804 22868
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 33196 20140 33236 20180
rect 29164 20056 29204 20096
rect 29356 20056 29396 20096
rect 30124 20056 30164 20096
rect 30412 19972 30452 20012
rect 30796 19804 30836 19844
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 34924 20140 34964 20180
rect 34060 20056 34100 20096
rect 31468 19468 31508 19508
rect 33772 19468 33812 19508
rect 39820 21400 39860 21440
rect 40492 21400 40532 21440
rect 36076 20056 36116 20096
rect 32236 19048 32276 19088
rect 35404 19048 35444 19088
rect 29836 18880 29876 18920
rect 31180 18880 31220 18920
rect 27244 18208 27284 18248
rect 26668 17956 26708 17996
rect 26476 17872 26516 17912
rect 26668 17788 26708 17828
rect 26572 17704 26612 17744
rect 26380 17620 26420 17660
rect 27532 17956 27572 17996
rect 25516 17452 25556 17492
rect 27340 17116 27380 17156
rect 30316 18124 30356 18164
rect 27820 17704 27860 17744
rect 30316 17704 30356 17744
rect 31372 17704 31412 17744
rect 28012 17620 28052 17660
rect 29932 17620 29972 17660
rect 30988 17116 31028 17156
rect 37324 20056 37364 20096
rect 38668 20056 38708 20096
rect 36940 19468 36980 19508
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 36460 18880 36500 18920
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 32332 17788 32372 17828
rect 33868 17704 33908 17744
rect 27628 15436 27668 15476
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 34060 17116 34100 17156
rect 36172 17116 36212 17156
rect 33388 16780 33428 16820
rect 34924 16780 34964 16820
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 35692 15520 35732 15560
rect 36268 15520 36308 15560
rect 34060 15436 34100 15476
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 23308 14680 23348 14720
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 19660 14008 19700 14048
rect 20428 13336 20468 13376
rect 20236 13252 20276 13292
rect 19372 13168 19412 13208
rect 20332 13168 20372 13208
rect 23884 13840 23924 13880
rect 25132 13840 25172 13880
rect 25324 13840 25364 13880
rect 25900 13840 25940 13880
rect 23500 13168 23540 13208
rect 28876 13840 28916 13880
rect 24268 13168 24308 13208
rect 23308 13084 23348 13124
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 19948 12580 19988 12620
rect 19852 12496 19892 12536
rect 19660 12412 19700 12452
rect 28012 13084 28052 13124
rect 27628 13000 27668 13040
rect 25132 12580 25172 12620
rect 20140 12496 20180 12536
rect 21292 12496 21332 12536
rect 28972 13168 29012 13208
rect 28396 13000 28436 13040
rect 28588 13000 28628 13040
rect 29068 13000 29108 13040
rect 29452 13000 29492 13040
rect 32524 14008 32564 14048
rect 33676 14008 33716 14048
rect 35980 15268 36020 15308
rect 36748 15268 36788 15308
rect 38476 19804 38516 19844
rect 38956 19804 38996 19844
rect 39340 19804 39380 19844
rect 39820 20056 39860 20096
rect 40588 20140 40628 20180
rect 41740 25180 41780 25220
rect 41644 23836 41684 23876
rect 46156 30640 46196 30680
rect 45676 30556 45716 30596
rect 47500 30724 47540 30764
rect 46732 30640 46772 30680
rect 46636 30220 46676 30260
rect 44716 29716 44756 29756
rect 46252 29800 46292 29840
rect 45964 29632 46004 29672
rect 46636 29632 46676 29672
rect 45868 29128 45908 29168
rect 46828 29128 46868 29168
rect 44140 28960 44180 29000
rect 44332 28960 44372 29000
rect 43756 27700 43796 27740
rect 44908 28372 44948 28412
rect 45676 28372 45716 28412
rect 45868 28372 45908 28412
rect 44716 27700 44756 27740
rect 48268 30640 48308 30680
rect 48940 31480 48980 31520
rect 49516 31480 49556 31520
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 49516 30724 49556 30764
rect 47788 30388 47828 30428
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 50380 30640 50420 30680
rect 48556 30556 48596 30596
rect 48748 30556 48788 30596
rect 50284 30556 50324 30596
rect 48460 30388 48500 30428
rect 48364 30220 48404 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 47884 29716 47924 29756
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 47404 29044 47444 29084
rect 43372 26104 43412 26144
rect 43756 25852 43796 25892
rect 43372 25264 43412 25304
rect 43276 25180 43316 25220
rect 42892 23836 42932 23876
rect 42316 23752 42356 23792
rect 42796 23752 42836 23792
rect 42220 23416 42260 23456
rect 42796 23416 42836 23456
rect 42316 23080 42356 23120
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 47884 27028 47924 27068
rect 49420 27028 49460 27068
rect 46636 26104 46676 26144
rect 46348 25180 46388 25220
rect 47308 25180 47348 25220
rect 43756 23752 43796 23792
rect 43372 23584 43412 23624
rect 42988 22996 43028 23036
rect 43276 22996 43316 23036
rect 43852 23080 43892 23120
rect 41740 20056 41780 20096
rect 40876 19972 40916 20012
rect 37324 19048 37364 19088
rect 38476 19048 38516 19088
rect 39820 19048 39860 19088
rect 40684 19048 40724 19088
rect 37612 18880 37652 18920
rect 37612 17032 37652 17072
rect 39628 17704 39668 17744
rect 41548 17788 41588 17828
rect 41932 17788 41972 17828
rect 41452 17704 41492 17744
rect 41356 17116 41396 17156
rect 40396 17032 40436 17072
rect 41260 17032 41300 17072
rect 41836 17704 41876 17744
rect 43468 17704 43508 17744
rect 42316 17032 42356 17072
rect 42700 17032 42740 17072
rect 41356 16948 41396 16988
rect 41740 16948 41780 16988
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 30508 13168 30548 13208
rect 28876 12580 28916 12620
rect 21964 12244 22004 12284
rect 23020 12244 23060 12284
rect 18892 9556 18932 9596
rect 13132 9472 13172 9512
rect 12364 8800 12404 8840
rect 12940 8800 12980 8840
rect 10060 8716 10100 8756
rect 10348 8716 10388 8756
rect 11692 8716 11732 8756
rect 11212 8632 11252 8672
rect 17164 9472 17204 9512
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 17164 8800 17204 8840
rect 17452 8800 17492 8840
rect 16108 7204 16148 7244
rect 16300 7204 16340 7244
rect 16588 7204 16628 7244
rect 7468 2752 7508 2792
rect 7660 2752 7700 2792
rect 7084 2416 7124 2456
rect 652 2248 692 2288
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 8428 2500 8468 2540
rect 7852 2416 7892 2456
rect 7276 2080 7316 2120
rect 8236 2080 8276 2120
rect 8044 1996 8084 2036
rect 8908 2080 8948 2120
rect 11596 4096 11636 4136
rect 11884 4936 11924 4976
rect 11884 4096 11924 4136
rect 11500 3508 11540 3548
rect 11980 3508 12020 3548
rect 10828 3424 10868 3464
rect 10732 2752 10772 2792
rect 11116 3424 11156 3464
rect 11020 2584 11060 2624
rect 10540 2500 10580 2540
rect 10924 2500 10964 2540
rect 12652 3508 12692 3548
rect 12364 3424 12404 3464
rect 13036 3508 13076 3548
rect 12748 3424 12788 3464
rect 11692 2584 11732 2624
rect 16204 7120 16244 7160
rect 18796 8632 18836 8672
rect 15628 4936 15668 4976
rect 15340 3424 15380 3464
rect 17260 3424 17300 3464
rect 14476 2752 14516 2792
rect 15148 2752 15188 2792
rect 12844 2584 12884 2624
rect 14092 2584 14132 2624
rect 17836 2836 17876 2876
rect 17644 2668 17684 2708
rect 18700 7876 18740 7916
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 19180 8800 19220 8840
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 31180 12412 31220 12452
rect 28012 11656 28052 11696
rect 28300 11656 28340 11696
rect 32332 13000 32372 13040
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 32620 12580 32660 12620
rect 35020 12580 35060 12620
rect 33484 12496 33524 12536
rect 32236 12412 32276 12452
rect 33772 12412 33812 12452
rect 19372 10984 19412 11024
rect 23404 10984 23444 11024
rect 20236 10144 20276 10184
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 19660 9556 19700 9596
rect 20236 8800 20276 8840
rect 19756 8632 19796 8672
rect 22252 8716 22292 8756
rect 19852 8548 19892 8588
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 20332 8632 20372 8672
rect 20908 8632 20948 8672
rect 21100 8632 21140 8672
rect 19180 7876 19220 7916
rect 19948 7876 19988 7916
rect 21580 8548 21620 8588
rect 21004 8464 21044 8504
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 18124 6196 18164 6236
rect 18892 6196 18932 6236
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 22060 8632 22100 8672
rect 22156 7960 22196 8000
rect 22924 8548 22964 8588
rect 23020 8464 23060 8504
rect 23212 8128 23252 8168
rect 23116 7960 23156 8000
rect 24268 10144 24308 10184
rect 25420 10060 25460 10100
rect 25516 9472 25556 9512
rect 25516 9220 25556 9260
rect 25612 8884 25652 8924
rect 24940 8800 24980 8840
rect 26380 9472 26420 9512
rect 25996 9388 26036 9428
rect 25804 9304 25844 9344
rect 26188 9304 26228 9344
rect 25804 8884 25844 8924
rect 25996 8632 26036 8672
rect 26764 9472 26804 9512
rect 26668 9220 26708 9260
rect 26476 8800 26516 8840
rect 25708 8128 25748 8168
rect 27340 8044 27380 8084
rect 22348 7288 22388 7328
rect 23404 7288 23444 7328
rect 22924 7120 22964 7160
rect 22732 7036 22772 7076
rect 25996 7036 26036 7076
rect 23596 6952 23636 6992
rect 21580 6196 21620 6236
rect 20044 4096 20084 4136
rect 20524 4096 20564 4136
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 24556 4936 24596 4976
rect 25612 4936 25652 4976
rect 23788 4180 23828 4220
rect 24364 4180 24404 4220
rect 21100 3592 21140 3632
rect 21772 3592 21812 3632
rect 22540 3508 22580 3548
rect 18700 3424 18740 3464
rect 18892 3424 18932 3464
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 18028 2836 18068 2876
rect 17932 2752 17972 2792
rect 25132 3508 25172 3548
rect 22636 3424 22676 3464
rect 23404 3424 23444 3464
rect 26956 7288 26996 7328
rect 26668 7120 26708 7160
rect 31468 11656 31508 11696
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 36172 12496 36212 12536
rect 33964 11908 34004 11948
rect 34444 11908 34484 11948
rect 31948 11656 31988 11696
rect 32332 11656 32372 11696
rect 32812 11656 32852 11696
rect 31372 11320 31412 11360
rect 31084 10144 31124 10184
rect 31852 11320 31892 11360
rect 31660 10144 31700 10184
rect 32812 11320 32852 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 36172 11320 36212 11360
rect 40876 14680 40916 14720
rect 40204 14596 40244 14636
rect 40780 14596 40820 14636
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 28684 8044 28724 8084
rect 29644 7960 29684 8000
rect 29068 7204 29108 7244
rect 28396 6952 28436 6992
rect 28876 7120 28916 7160
rect 29452 6952 29492 6992
rect 28588 6616 28628 6656
rect 29452 6616 29492 6656
rect 29644 6616 29684 6656
rect 30316 7960 30356 8000
rect 30028 7120 30068 7160
rect 30220 7120 30260 7160
rect 35980 8464 36020 8504
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 31084 7708 31124 7748
rect 32236 7708 32276 7748
rect 29932 6952 29972 6992
rect 26860 4936 26900 4976
rect 28300 4936 28340 4976
rect 27724 4096 27764 4136
rect 29836 6448 29876 6488
rect 30604 7120 30644 7160
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 37036 7960 37076 8000
rect 37228 7960 37268 8000
rect 38476 13168 38516 13208
rect 39628 14008 39668 14048
rect 39916 13840 39956 13880
rect 39244 13168 39284 13208
rect 39532 13168 39572 13208
rect 41548 16780 41588 16820
rect 42412 16780 42452 16820
rect 42604 15688 42644 15728
rect 42604 15436 42644 15476
rect 41548 14680 41588 14720
rect 40300 14008 40340 14048
rect 41260 14008 41300 14048
rect 42124 14008 42164 14048
rect 45964 23584 46004 23624
rect 44716 23080 44756 23120
rect 45580 22996 45620 23036
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 49132 23080 49172 23120
rect 48268 22996 48308 23036
rect 48940 22996 48980 23036
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 47980 22240 48020 22280
rect 49708 22240 49748 22280
rect 47884 21736 47924 21776
rect 48076 21736 48116 21776
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 49228 21484 49268 21524
rect 50284 21484 50324 21524
rect 48268 21400 48308 21440
rect 49420 21400 49460 21440
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 48172 20056 48212 20096
rect 46348 19132 46388 19172
rect 47596 19216 47636 19256
rect 47980 19216 48020 19256
rect 47212 19132 47252 19172
rect 46828 18460 46868 18500
rect 47116 18460 47156 18500
rect 46732 17956 46772 17996
rect 44332 15688 44372 15728
rect 45100 15688 45140 15728
rect 47980 18544 48020 18584
rect 47596 17956 47636 17996
rect 47788 17956 47828 17996
rect 47404 17788 47444 17828
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 49324 20056 49364 20096
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 49804 20140 49844 20180
rect 49420 19216 49460 19256
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 50476 20140 50516 20180
rect 50188 19216 50228 19256
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 50668 19048 50708 19088
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 48172 17956 48212 17996
rect 48556 17956 48596 17996
rect 48076 17788 48116 17828
rect 52012 19048 52052 19088
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 53260 18544 53300 18584
rect 52300 18460 52340 18500
rect 49612 17956 49652 17996
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 48364 15604 48404 15644
rect 49228 15604 49268 15644
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 46060 14680 46100 14720
rect 46636 14680 46676 14720
rect 49612 14680 49652 14720
rect 50380 14512 50420 14552
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 47884 14008 47924 14048
rect 42700 13840 42740 13880
rect 45292 13168 45332 13208
rect 47116 13168 47156 13208
rect 47980 13840 48020 13880
rect 48364 13756 48404 13796
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 49996 14008 50036 14048
rect 49612 13840 49652 13880
rect 49132 13168 49172 13208
rect 49324 13168 49364 13208
rect 38956 11320 38996 11360
rect 38380 10984 38420 11024
rect 39916 10984 39956 11024
rect 40300 10984 40340 11024
rect 38764 9220 38804 9260
rect 39532 9220 39572 9260
rect 38764 8800 38804 8840
rect 38380 8464 38420 8504
rect 38668 8044 38708 8084
rect 35596 7792 35636 7832
rect 32332 7036 32372 7076
rect 33484 6952 33524 6992
rect 31660 6448 31700 6488
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 33868 5608 33908 5648
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 33388 5020 33428 5060
rect 34348 5020 34388 5060
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 34444 4180 34484 4220
rect 29164 4096 29204 4136
rect 34348 4096 34388 4136
rect 33388 3928 33428 3968
rect 34252 3928 34292 3968
rect 26860 3508 26900 3548
rect 25996 3424 26036 3464
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 19852 2836 19892 2876
rect 21100 2836 21140 2876
rect 35884 7036 35924 7076
rect 36556 6448 36596 6488
rect 38092 7792 38132 7832
rect 39052 8716 39092 8756
rect 37996 7036 38036 7076
rect 38764 6952 38804 6992
rect 39532 6952 39572 6992
rect 40204 9472 40244 9512
rect 39916 8044 39956 8084
rect 40876 11068 40916 11108
rect 43660 11068 43700 11108
rect 40588 9640 40628 9680
rect 41164 10732 41204 10772
rect 44332 10732 44372 10772
rect 45964 13000 46004 13040
rect 46828 13000 46868 13040
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 41356 9640 41396 9680
rect 45004 9640 45044 9680
rect 41548 9472 41588 9512
rect 40684 8800 40724 8840
rect 40588 8716 40628 8756
rect 41548 8800 41588 8840
rect 40012 6952 40052 6992
rect 39340 6448 39380 6488
rect 37708 6196 37748 6236
rect 36556 5608 36596 5648
rect 38572 6280 38612 6320
rect 39244 4852 39284 4892
rect 39628 4852 39668 4892
rect 38956 4180 38996 4220
rect 37996 3760 38036 3800
rect 35788 3592 35828 3632
rect 33772 2668 33812 2708
rect 35500 2668 35540 2708
rect 37132 2668 37172 2708
rect 36748 2584 36788 2624
rect 12172 2500 12212 2540
rect 11308 2080 11348 2120
rect 51628 15436 51668 15476
rect 52780 15436 52820 15476
rect 53452 15436 53492 15476
rect 51436 15268 51476 15308
rect 52108 15268 52148 15308
rect 52204 14680 52244 14720
rect 52780 14680 52820 14720
rect 51340 14596 51380 14636
rect 51628 14512 51668 14552
rect 51244 14260 51284 14300
rect 51244 14092 51284 14132
rect 50572 13756 50612 13796
rect 49996 13420 50036 13460
rect 50476 13420 50516 13460
rect 52876 14596 52916 14636
rect 52684 14260 52724 14300
rect 53068 14260 53108 14300
rect 52876 14092 52916 14132
rect 55948 15772 55988 15812
rect 54796 14680 54836 14720
rect 56332 14092 56372 14132
rect 52972 13420 53012 13460
rect 52204 13252 52244 13292
rect 52876 13252 52916 13292
rect 50284 13168 50324 13208
rect 52300 13168 52340 13208
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 47020 10228 47060 10268
rect 46540 10060 46580 10100
rect 47116 10144 47156 10184
rect 47884 10144 47924 10184
rect 48460 10228 48500 10268
rect 47308 10060 47348 10100
rect 47212 9640 47252 9680
rect 48556 10144 48596 10184
rect 49804 10144 49844 10184
rect 52780 10732 52820 10772
rect 50284 10144 50324 10184
rect 50764 10144 50804 10184
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 47692 9472 47732 9512
rect 48556 9472 48596 9512
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 45868 8632 45908 8672
rect 45196 6448 45236 6488
rect 46252 6448 46292 6488
rect 46444 6448 46484 6488
rect 43660 5608 43700 5648
rect 44812 5608 44852 5648
rect 45292 5608 45332 5648
rect 46540 5608 46580 5648
rect 45964 5524 46004 5564
rect 46636 5524 46676 5564
rect 42508 4936 42548 4976
rect 47116 8632 47156 8672
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 51820 9640 51860 9680
rect 53836 13252 53876 13292
rect 54604 13168 54644 13208
rect 55084 13000 55124 13040
rect 55180 12664 55220 12704
rect 55468 12580 55508 12620
rect 54028 11152 54068 11192
rect 54700 11152 54740 11192
rect 55084 11152 55124 11192
rect 55756 11152 55796 11192
rect 53836 10732 53876 10772
rect 56140 13000 56180 13040
rect 54892 10312 54932 10352
rect 55564 10312 55604 10352
rect 53164 9640 53204 9680
rect 53068 9472 53108 9512
rect 50956 7960 50996 8000
rect 51724 7960 51764 8000
rect 47116 7120 47156 7160
rect 48748 7120 48788 7160
rect 47404 6448 47444 6488
rect 47980 6448 48020 6488
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 51820 7120 51860 7160
rect 51148 6448 51188 6488
rect 48364 5860 48404 5900
rect 49612 5860 49652 5900
rect 47212 5608 47252 5648
rect 40204 4180 40244 4220
rect 40492 4180 40532 4220
rect 40108 4096 40148 4136
rect 39244 3760 39284 3800
rect 38284 3592 38324 3632
rect 40300 3508 40340 3548
rect 38380 3340 38420 3380
rect 40012 3424 40052 3464
rect 39532 3340 39572 3380
rect 40588 3760 40628 3800
rect 40396 3424 40436 3464
rect 40204 3340 40244 3380
rect 38188 2584 38228 2624
rect 39724 2584 39764 2624
rect 41356 4096 41396 4136
rect 41644 3928 41684 3968
rect 44044 3928 44084 3968
rect 41068 3508 41108 3548
rect 40972 3424 41012 3464
rect 45292 3760 45332 3800
rect 46444 3760 46484 3800
rect 44428 2584 44468 2624
rect 47116 3424 47156 3464
rect 46444 2836 46484 2876
rect 48652 5608 48692 5648
rect 51148 5608 51188 5648
rect 47692 5020 47732 5060
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 51916 5020 51956 5060
rect 53740 6616 53780 6656
rect 52108 4936 52148 4976
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 48268 3760 48308 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 47692 3424 47732 3464
rect 48076 2836 48116 2876
rect 47308 2584 47348 2624
rect 55756 10228 55796 10268
rect 55948 10228 55988 10268
rect 55276 9472 55316 9512
rect 57004 14512 57044 14552
rect 56812 14092 56852 14132
rect 56716 13924 56756 13964
rect 56428 13000 56468 13040
rect 56428 12664 56468 12704
rect 56716 12580 56756 12620
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 57676 15772 57716 15812
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 57964 14512 58004 14552
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 57292 13924 57332 13964
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 57484 13000 57524 13040
rect 57676 12664 57716 12704
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 56620 10228 56660 10268
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 54988 6616 55028 6656
rect 54028 6448 54068 6488
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 53068 4936 53108 4976
rect 52972 4600 53012 4640
rect 51724 3424 51764 3464
rect 52012 3508 52052 3548
rect 53164 3508 53204 3548
rect 51436 3340 51476 3380
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 49516 2668 49556 2708
rect 49132 2584 49172 2624
rect 50860 2584 50900 2624
rect 51916 3340 51956 3380
rect 52108 2752 52148 2792
rect 56620 5608 56660 5648
rect 57196 5608 57236 5648
rect 54412 5440 54452 5480
rect 55948 5440 55988 5480
rect 54028 4936 54068 4976
rect 54796 4600 54836 4640
rect 55180 4600 55220 4640
rect 53836 3424 53876 3464
rect 55660 3424 55700 3464
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 56044 3424 56084 3464
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 53452 2668 53492 2708
rect 54700 2668 54740 2708
rect 55852 2668 55892 2708
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal3 >>
rect 4343 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 4729 38576
rect 19463 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 19849 38576
rect 34583 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 34969 38576
rect 49703 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 50089 38576
rect 64823 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 65209 38576
rect 79943 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 80329 38576
rect 95063 38536 95072 38576
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95440 38536 95449 38576
rect 3103 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 3489 37820
rect 18223 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 18609 37820
rect 33343 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 33729 37820
rect 48463 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 48849 37820
rect 63583 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 63969 37820
rect 78703 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 79089 37820
rect 93823 37780 93832 37820
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 94200 37780 94209 37820
rect 0 37568 80 37588
rect 0 37528 268 37568
rect 308 37528 317 37568
rect 0 37508 80 37528
rect 25699 37444 25708 37484
rect 25748 37444 26188 37484
rect 26228 37444 26764 37484
rect 26804 37444 26813 37484
rect 18115 37192 18124 37232
rect 18164 37192 18796 37232
rect 18836 37192 21772 37232
rect 21812 37192 21821 37232
rect 25123 37192 25132 37232
rect 25172 37192 25516 37232
rect 25556 37192 25565 37232
rect 4343 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 4729 37064
rect 19463 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 19849 37064
rect 34583 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 34969 37064
rect 49703 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 50089 37064
rect 64823 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 65209 37064
rect 79943 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 80329 37064
rect 95063 37024 95072 37064
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95440 37024 95449 37064
rect 40675 36856 40684 36896
rect 40724 36856 42124 36896
rect 42164 36856 42173 36896
rect 16771 36772 16780 36812
rect 16820 36772 17932 36812
rect 17972 36772 17981 36812
rect 21859 36772 21868 36812
rect 21908 36772 22636 36812
rect 22676 36772 22685 36812
rect 0 36728 80 36748
rect 0 36688 76 36728
rect 116 36688 125 36728
rect 22243 36688 22252 36728
rect 22292 36688 25516 36728
rect 25556 36688 28204 36728
rect 28244 36688 28253 36728
rect 29635 36688 29644 36728
rect 29684 36688 30220 36728
rect 30260 36688 30269 36728
rect 37507 36688 37516 36728
rect 37556 36688 37565 36728
rect 38371 36688 38380 36728
rect 38420 36688 40972 36728
rect 41012 36688 41548 36728
rect 41588 36688 41597 36728
rect 0 36668 80 36688
rect 37516 36644 37556 36688
rect 10531 36604 10540 36644
rect 10580 36604 12076 36644
rect 12116 36604 12125 36644
rect 22531 36604 22540 36644
rect 22580 36604 26284 36644
rect 26324 36604 26333 36644
rect 37516 36604 40108 36644
rect 40148 36604 40684 36644
rect 40724 36604 40733 36644
rect 11875 36520 11884 36560
rect 11924 36520 13324 36560
rect 13364 36520 13373 36560
rect 16195 36520 16204 36560
rect 16244 36520 17164 36560
rect 17204 36520 17213 36560
rect 33187 36520 33196 36560
rect 33236 36520 34156 36560
rect 34196 36520 34205 36560
rect 34339 36520 34348 36560
rect 34388 36520 35116 36560
rect 35156 36520 35165 36560
rect 3103 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 3489 36308
rect 18223 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 18609 36308
rect 33343 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 33729 36308
rect 48463 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 48849 36308
rect 63583 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 63969 36308
rect 78703 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 79089 36308
rect 93823 36268 93832 36308
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 94200 36268 94209 36308
rect 18211 35932 18220 35972
rect 18260 35932 19084 35972
rect 19124 35932 19133 35972
rect 26380 35932 27436 35972
rect 27476 35932 28972 35972
rect 29012 35932 29021 35972
rect 35107 35932 35116 35972
rect 35156 35932 37132 35972
rect 37172 35932 37181 35972
rect 0 35828 80 35908
rect 26380 35888 26420 35932
rect 6115 35848 6124 35888
rect 6164 35848 6700 35888
rect 6740 35848 6749 35888
rect 17059 35848 17068 35888
rect 17108 35848 18028 35888
rect 18068 35848 18077 35888
rect 21955 35848 21964 35888
rect 22004 35848 25708 35888
rect 25748 35848 25757 35888
rect 26371 35848 26380 35888
rect 26420 35848 26429 35888
rect 37603 35848 37612 35888
rect 37652 35848 38668 35888
rect 38708 35848 39628 35888
rect 39668 35848 39677 35888
rect 9667 35764 9676 35804
rect 9716 35764 10540 35804
rect 10580 35764 10589 35804
rect 15811 35764 15820 35804
rect 15860 35764 16876 35804
rect 16916 35764 16925 35804
rect 4343 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 4729 35552
rect 19463 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 19849 35552
rect 34583 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 34969 35552
rect 49703 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 50089 35552
rect 64823 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 65209 35552
rect 79943 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 80329 35552
rect 95063 35512 95072 35552
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95440 35512 95449 35552
rect 36931 35344 36940 35384
rect 36980 35344 37612 35384
rect 37652 35344 37661 35384
rect 36844 35260 37324 35300
rect 37364 35260 37373 35300
rect 36844 35216 36884 35260
rect 6691 35176 6700 35216
rect 6740 35176 8812 35216
rect 8852 35176 8861 35216
rect 18019 35176 18028 35216
rect 18068 35176 18796 35216
rect 18836 35176 20524 35216
rect 20564 35176 20573 35216
rect 33571 35176 33580 35216
rect 33620 35176 34252 35216
rect 34292 35176 34301 35216
rect 36451 35176 36460 35216
rect 36500 35176 36844 35216
rect 36884 35176 36893 35216
rect 37219 35176 37228 35216
rect 37268 35176 39052 35216
rect 39092 35176 39101 35216
rect 6115 35092 6124 35132
rect 6164 35092 7276 35132
rect 7316 35092 8908 35132
rect 8948 35092 8957 35132
rect 17059 35092 17068 35132
rect 17108 35092 18124 35132
rect 18164 35092 18412 35132
rect 18452 35092 18461 35132
rect 0 34988 80 35068
rect 6691 35008 6700 35048
rect 6740 35008 6988 35048
rect 7028 35008 7564 35048
rect 7604 35008 7613 35048
rect 3103 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 3489 34796
rect 18223 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 18609 34796
rect 33343 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 33729 34796
rect 48463 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 48849 34796
rect 63583 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 63969 34796
rect 78703 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 79089 34796
rect 93823 34756 93832 34796
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 94200 34756 94209 34796
rect 6307 34588 6316 34628
rect 6356 34588 7180 34628
rect 7220 34588 7229 34628
rect 33187 34588 33196 34628
rect 33236 34588 34156 34628
rect 34196 34588 34205 34628
rect 21187 34504 21196 34544
rect 21236 34504 22156 34544
rect 22196 34504 23116 34544
rect 23156 34504 23165 34544
rect 23299 34420 23308 34460
rect 23348 34420 24076 34460
rect 24116 34420 24125 34460
rect 34339 34420 34348 34460
rect 34388 34420 36460 34460
rect 36500 34420 36509 34460
rect 11875 34336 11884 34376
rect 11924 34336 12268 34376
rect 12308 34336 12460 34376
rect 12500 34336 12509 34376
rect 21475 34336 21484 34376
rect 21524 34336 23116 34376
rect 23156 34336 25324 34376
rect 25364 34336 25373 34376
rect 19171 34252 19180 34292
rect 19220 34252 20908 34292
rect 20948 34252 20957 34292
rect 0 34148 80 34228
rect 7363 34168 7372 34208
rect 7412 34168 8140 34208
rect 8180 34168 9100 34208
rect 9140 34168 10444 34208
rect 10484 34168 10493 34208
rect 4343 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 4729 34040
rect 13123 34000 13132 34040
rect 13172 34000 15628 34040
rect 15668 34000 15677 34040
rect 19463 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 19849 34040
rect 21283 34000 21292 34040
rect 21332 34000 22348 34040
rect 22388 34000 22397 34040
rect 34583 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 34969 34040
rect 49703 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 50089 34040
rect 64823 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 65209 34040
rect 79943 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 80329 34040
rect 95063 34000 95072 34040
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95440 34000 95449 34040
rect 25315 33664 25324 33704
rect 25364 33664 26284 33704
rect 26324 33664 26956 33704
rect 26996 33664 29068 33704
rect 29108 33664 29356 33704
rect 29396 33664 29405 33704
rect 7171 33580 7180 33620
rect 7220 33580 10060 33620
rect 10100 33580 12172 33620
rect 12212 33580 12221 33620
rect 15715 33580 15724 33620
rect 15764 33580 16396 33620
rect 16436 33580 16445 33620
rect 42691 33412 42700 33452
rect 42740 33412 43372 33452
rect 43412 33412 43421 33452
rect 0 33308 80 33388
rect 3103 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 3489 33284
rect 18223 33244 18232 33284
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18600 33244 18609 33284
rect 33343 33244 33352 33284
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33720 33244 33729 33284
rect 48463 33244 48472 33284
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48840 33244 48849 33284
rect 63583 33244 63592 33284
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63960 33244 63969 33284
rect 78703 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 79089 33284
rect 93823 33244 93832 33284
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 94200 33244 94209 33284
rect 35491 33160 35500 33200
rect 35540 33160 36652 33200
rect 36692 33160 36701 33200
rect 18115 32908 18124 32948
rect 18164 32908 18988 32948
rect 19028 32908 19037 32948
rect 14467 32824 14476 32864
rect 14516 32824 15532 32864
rect 15572 32824 15581 32864
rect 16387 32824 16396 32864
rect 16436 32824 18028 32864
rect 18068 32824 18077 32864
rect 27235 32824 27244 32864
rect 27284 32824 28108 32864
rect 28148 32824 28157 32864
rect 11395 32656 11404 32696
rect 11444 32656 14860 32696
rect 14900 32656 16204 32696
rect 16244 32656 16253 32696
rect 0 32468 80 32548
rect 4343 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 4729 32528
rect 19463 32488 19472 32528
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19840 32488 19849 32528
rect 34583 32488 34592 32528
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34960 32488 34969 32528
rect 49703 32488 49712 32528
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 50080 32488 50089 32528
rect 64823 32488 64832 32528
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 65200 32488 65209 32528
rect 79943 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 80329 32528
rect 95063 32488 95072 32528
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95440 32488 95449 32528
rect 42787 32236 42796 32276
rect 42836 32236 42845 32276
rect 42796 32192 42836 32236
rect 3139 32152 3148 32192
rect 3188 32152 3820 32192
rect 3860 32152 6316 32192
rect 6356 32152 10540 32192
rect 10580 32152 10589 32192
rect 24643 32152 24652 32192
rect 24692 32152 26188 32192
rect 26228 32152 26237 32192
rect 34435 32152 34444 32192
rect 34484 32152 35020 32192
rect 35060 32152 36748 32192
rect 36788 32152 36797 32192
rect 38467 32152 38476 32192
rect 38516 32152 42836 32192
rect 34339 32068 34348 32108
rect 34388 32068 35884 32108
rect 35924 32068 39052 32108
rect 39092 32068 39101 32108
rect 17443 31900 17452 31940
rect 17492 31900 18028 31940
rect 18068 31900 18077 31940
rect 18211 31900 18220 31940
rect 18260 31900 18700 31940
rect 18740 31900 19180 31940
rect 19220 31900 20140 31940
rect 20180 31900 20189 31940
rect 36931 31900 36940 31940
rect 36980 31900 38188 31940
rect 38228 31900 38237 31940
rect 3103 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 3489 31772
rect 18223 31732 18232 31772
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18600 31732 18609 31772
rect 33343 31732 33352 31772
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33720 31732 33729 31772
rect 48463 31732 48472 31772
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48840 31732 48849 31772
rect 63583 31732 63592 31772
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63960 31732 63969 31772
rect 78703 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 79089 31772
rect 93823 31732 93832 31772
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 94200 31732 94209 31772
rect 0 31628 80 31708
rect 22339 31480 22348 31520
rect 22388 31480 26092 31520
rect 26132 31480 26141 31520
rect 42307 31480 42316 31520
rect 42356 31480 42988 31520
rect 43028 31480 43037 31520
rect 48931 31480 48940 31520
rect 48980 31480 49516 31520
rect 49556 31480 49565 31520
rect 2371 31396 2380 31436
rect 2420 31396 3532 31436
rect 3572 31396 4012 31436
rect 4052 31396 4061 31436
rect 2275 31312 2284 31352
rect 2324 31312 2956 31352
rect 2996 31312 7660 31352
rect 7700 31312 9004 31352
rect 9044 31312 9676 31352
rect 9716 31312 9725 31352
rect 25987 31312 25996 31352
rect 26036 31312 26188 31352
rect 26228 31312 26237 31352
rect 26371 31312 26380 31352
rect 26420 31312 27052 31352
rect 27092 31312 27101 31352
rect 2668 31100 2708 31312
rect 34723 31228 34732 31268
rect 34772 31228 36268 31268
rect 36308 31228 36317 31268
rect 38179 31144 38188 31184
rect 38228 31144 41932 31184
rect 41972 31144 41981 31184
rect 2659 31060 2668 31100
rect 2708 31060 2717 31100
rect 4343 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 4729 31016
rect 19463 30976 19472 31016
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19840 30976 19849 31016
rect 34583 30976 34592 31016
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34960 30976 34969 31016
rect 49703 30976 49712 31016
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 50080 30976 50089 31016
rect 64823 30976 64832 31016
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 65200 30976 65209 31016
rect 79943 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 80329 31016
rect 95063 30976 95072 31016
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95440 30976 95449 31016
rect 0 30788 80 30868
rect 37987 30808 37996 30848
rect 38036 30808 38380 30848
rect 38420 30808 38429 30848
rect 20323 30724 20332 30764
rect 20372 30724 21964 30764
rect 22004 30724 22013 30764
rect 25795 30724 25804 30764
rect 25844 30724 26956 30764
rect 26996 30724 27005 30764
rect 28867 30724 28876 30764
rect 28916 30724 31084 30764
rect 31124 30724 31133 30764
rect 39043 30724 39052 30764
rect 39092 30724 40684 30764
rect 40724 30724 41164 30764
rect 41204 30724 41213 30764
rect 47491 30724 47500 30764
rect 47540 30724 49516 30764
rect 49556 30724 49565 30764
rect 3523 30640 3532 30680
rect 3572 30640 4204 30680
rect 4244 30640 4253 30680
rect 5635 30640 5644 30680
rect 5684 30640 7276 30680
rect 7316 30640 7325 30680
rect 24355 30640 24364 30680
rect 24404 30640 25324 30680
rect 25364 30640 27436 30680
rect 27476 30640 27485 30680
rect 30979 30640 30988 30680
rect 31028 30640 32332 30680
rect 32372 30640 32381 30680
rect 33475 30640 33484 30680
rect 33524 30640 34156 30680
rect 34196 30640 35020 30680
rect 35060 30640 35069 30680
rect 39427 30640 39436 30680
rect 39476 30640 41600 30680
rect 42691 30640 42700 30680
rect 42740 30640 43468 30680
rect 43508 30640 46156 30680
rect 46196 30640 46732 30680
rect 46772 30640 48268 30680
rect 48308 30640 50380 30680
rect 50420 30640 50429 30680
rect 41560 30596 41600 30640
rect 41560 30556 45676 30596
rect 45716 30556 45725 30596
rect 48547 30556 48556 30596
rect 48596 30556 48748 30596
rect 48788 30556 50284 30596
rect 50324 30556 50333 30596
rect 42019 30472 42028 30512
rect 42068 30472 43084 30512
rect 43124 30472 43133 30512
rect 4099 30388 4108 30428
rect 4148 30388 5164 30428
rect 5204 30388 5213 30428
rect 9667 30388 9676 30428
rect 9716 30388 11116 30428
rect 11156 30388 11165 30428
rect 25123 30388 25132 30428
rect 25172 30388 25708 30428
rect 25748 30388 25757 30428
rect 34435 30388 34444 30428
rect 34484 30388 35980 30428
rect 36020 30388 36029 30428
rect 47779 30388 47788 30428
rect 47828 30388 48460 30428
rect 48500 30388 48509 30428
rect 4483 30304 4492 30344
rect 4532 30304 6508 30344
rect 6548 30304 6557 30344
rect 3103 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 3489 30260
rect 17539 30220 17548 30260
rect 17588 30220 17932 30260
rect 17972 30220 17981 30260
rect 18223 30220 18232 30260
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18600 30220 18609 30260
rect 26083 30220 26092 30260
rect 26132 30220 28492 30260
rect 28532 30220 29164 30260
rect 29204 30220 29213 30260
rect 33343 30220 33352 30260
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33720 30220 33729 30260
rect 46627 30220 46636 30260
rect 46676 30220 48364 30260
rect 48404 30220 48413 30260
rect 48463 30220 48472 30260
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48840 30220 48849 30260
rect 63583 30220 63592 30260
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63960 30220 63969 30260
rect 78703 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 79089 30260
rect 93823 30220 93832 30260
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 94200 30220 94209 30260
rect 15907 30136 15916 30176
rect 15956 30136 18028 30176
rect 18068 30136 20140 30176
rect 20180 30136 20189 30176
rect 18115 30052 18124 30092
rect 18164 30052 19180 30092
rect 19220 30052 20044 30092
rect 20084 30052 20093 30092
rect 0 29948 80 30028
rect 37411 29800 37420 29840
rect 37460 29800 37804 29840
rect 37844 29800 37853 29840
rect 38083 29800 38092 29840
rect 38132 29800 38668 29840
rect 38708 29800 38717 29840
rect 42403 29800 42412 29840
rect 42452 29800 46252 29840
rect 46292 29800 46301 29840
rect 44707 29716 44716 29756
rect 44756 29716 47884 29756
rect 47924 29716 47933 29756
rect 26083 29632 26092 29672
rect 26132 29632 26956 29672
rect 26996 29632 27005 29672
rect 45955 29632 45964 29672
rect 46004 29632 46636 29672
rect 46676 29632 46685 29672
rect 4343 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 4729 29504
rect 19463 29464 19472 29504
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19840 29464 19849 29504
rect 34583 29464 34592 29504
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34960 29464 34969 29504
rect 49703 29464 49712 29504
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 50080 29464 50089 29504
rect 64823 29464 64832 29504
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 65200 29464 65209 29504
rect 79943 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 80329 29504
rect 95063 29464 95072 29504
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95440 29464 95449 29504
rect 28003 29212 28012 29252
rect 28052 29212 28492 29252
rect 28532 29212 30412 29252
rect 30452 29212 30461 29252
rect 0 29108 80 29188
rect 9763 29128 9772 29168
rect 9812 29128 10444 29168
rect 10484 29128 23020 29168
rect 23060 29128 23308 29168
rect 23348 29128 23357 29168
rect 28675 29128 28684 29168
rect 28724 29128 29068 29168
rect 29108 29128 29117 29168
rect 45859 29128 45868 29168
rect 45908 29128 46828 29168
rect 46868 29128 46877 29168
rect 31075 29044 31084 29084
rect 31124 29044 32140 29084
rect 32180 29044 32189 29084
rect 43171 29044 43180 29084
rect 43220 29044 47404 29084
rect 47444 29044 47453 29084
rect 3523 28960 3532 29000
rect 3572 28960 4204 29000
rect 4244 28960 5068 29000
rect 5108 28960 5117 29000
rect 9475 28960 9484 29000
rect 9524 28960 11404 29000
rect 11444 28960 11453 29000
rect 12451 28960 12460 29000
rect 12500 28960 13036 29000
rect 13076 28960 13085 29000
rect 42595 28960 42604 29000
rect 42644 28960 42796 29000
rect 42836 28960 44140 29000
rect 44180 28960 44332 29000
rect 44372 28960 44381 29000
rect 3103 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 3489 28748
rect 18223 28708 18232 28748
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18600 28708 18609 28748
rect 33343 28708 33352 28748
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33720 28708 33729 28748
rect 48463 28708 48472 28748
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48840 28708 48849 28748
rect 63583 28708 63592 28748
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63960 28708 63969 28748
rect 78703 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 79089 28748
rect 93823 28708 93832 28748
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 94200 28708 94209 28748
rect 5827 28540 5836 28580
rect 5876 28540 8524 28580
rect 8564 28540 8573 28580
rect 44899 28372 44908 28412
rect 44948 28372 45676 28412
rect 45716 28372 45868 28412
rect 45908 28372 45917 28412
rect 0 28268 80 28348
rect 6115 28288 6124 28328
rect 6164 28288 8812 28328
rect 8852 28288 8861 28328
rect 13123 28288 13132 28328
rect 13172 28288 14092 28328
rect 14132 28288 14141 28328
rect 5251 28120 5260 28160
rect 5300 28120 6412 28160
rect 6452 28120 6461 28160
rect 4343 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 4729 27992
rect 19463 27952 19472 27992
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19840 27952 19849 27992
rect 34583 27952 34592 27992
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34960 27952 34969 27992
rect 49703 27952 49712 27992
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 50080 27952 50089 27992
rect 64823 27952 64832 27992
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 65200 27952 65209 27992
rect 79943 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 80329 27992
rect 95063 27952 95072 27992
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95440 27952 95449 27992
rect 3619 27700 3628 27740
rect 3668 27700 5164 27740
rect 5204 27700 5213 27740
rect 6691 27700 6700 27740
rect 6740 27700 8620 27740
rect 8660 27700 8669 27740
rect 22051 27700 22060 27740
rect 22100 27700 23212 27740
rect 23252 27700 23261 27740
rect 23395 27700 23404 27740
rect 23444 27700 25132 27740
rect 25172 27700 25181 27740
rect 43747 27700 43756 27740
rect 43796 27700 44716 27740
rect 44756 27700 44765 27740
rect 23212 27656 23252 27700
rect 2659 27616 2668 27656
rect 2708 27616 4300 27656
rect 4340 27616 4349 27656
rect 23212 27616 24844 27656
rect 24884 27616 26092 27656
rect 26132 27616 26141 27656
rect 11011 27532 11020 27572
rect 11060 27532 12076 27572
rect 12116 27532 13708 27572
rect 13748 27532 13757 27572
rect 22147 27532 22156 27572
rect 22196 27532 23404 27572
rect 23444 27532 23453 27572
rect 0 27428 80 27508
rect 2275 27448 2284 27488
rect 2324 27448 3244 27488
rect 3284 27448 3293 27488
rect 23299 27448 23308 27488
rect 23348 27448 26284 27488
rect 26324 27448 26333 27488
rect 20899 27364 20908 27404
rect 20948 27364 21868 27404
rect 21908 27364 21917 27404
rect 3103 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 3489 27236
rect 18223 27196 18232 27236
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18600 27196 18609 27236
rect 33343 27196 33352 27236
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33720 27196 33729 27236
rect 48463 27196 48472 27236
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48840 27196 48849 27236
rect 63583 27196 63592 27236
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63960 27196 63969 27236
rect 78703 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 79089 27236
rect 93823 27196 93832 27236
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 94200 27196 94209 27236
rect 4675 27028 4684 27068
rect 4724 27028 5260 27068
rect 5300 27028 5644 27068
rect 5684 27028 5693 27068
rect 47875 27028 47884 27068
rect 47924 27028 49420 27068
rect 49460 27028 49469 27068
rect 39523 26860 39532 26900
rect 39572 26860 40396 26900
rect 40436 26860 40445 26900
rect 8899 26776 8908 26816
rect 8948 26776 9484 26816
rect 9524 26776 10060 26816
rect 10100 26776 10109 26816
rect 13123 26776 13132 26816
rect 13172 26776 15724 26816
rect 15764 26776 16108 26816
rect 16148 26776 16157 26816
rect 16579 26776 16588 26816
rect 16628 26776 18796 26816
rect 18836 26776 19372 26816
rect 19412 26776 19564 26816
rect 19604 26776 19613 26816
rect 20515 26776 20524 26816
rect 20564 26776 22156 26816
rect 22196 26776 22205 26816
rect 26083 26776 26092 26816
rect 26132 26776 28972 26816
rect 29012 26776 29021 26816
rect 32131 26776 32140 26816
rect 32180 26776 33292 26816
rect 33332 26776 33341 26816
rect 37123 26692 37132 26732
rect 37172 26692 38188 26732
rect 38228 26692 38237 26732
rect 0 26588 80 26668
rect 15139 26608 15148 26648
rect 15188 26608 17068 26648
rect 17108 26608 17117 26648
rect 31459 26608 31468 26648
rect 31508 26608 32044 26648
rect 32084 26608 32093 26648
rect 4343 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 4729 26480
rect 19463 26440 19472 26480
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19840 26440 19849 26480
rect 29827 26440 29836 26480
rect 29876 26440 30220 26480
rect 30260 26440 30269 26480
rect 34583 26440 34592 26480
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34960 26440 34969 26480
rect 49703 26440 49712 26480
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 50080 26440 50089 26480
rect 64823 26440 64832 26480
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 65200 26440 65209 26480
rect 79943 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 80329 26480
rect 95063 26440 95072 26480
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95440 26440 95449 26480
rect 9859 26272 9868 26312
rect 9908 26272 10060 26312
rect 10100 26272 11788 26312
rect 11828 26272 13996 26312
rect 14036 26272 14045 26312
rect 29827 26188 29836 26228
rect 29876 26188 30124 26228
rect 30164 26188 34156 26228
rect 34196 26188 34924 26228
rect 34964 26188 41740 26228
rect 41780 26188 41789 26228
rect 19363 26104 19372 26144
rect 19412 26104 20332 26144
rect 20372 26104 21100 26144
rect 21140 26104 21149 26144
rect 30691 26104 30700 26144
rect 30740 26104 31276 26144
rect 31316 26104 31325 26144
rect 32131 26104 32140 26144
rect 32180 26104 33196 26144
rect 33236 26104 35788 26144
rect 35828 26104 35837 26144
rect 43363 26104 43372 26144
rect 43412 26104 46636 26144
rect 46676 26104 46685 26144
rect 31276 26060 31316 26104
rect 3427 26020 3436 26060
rect 3476 26020 4108 26060
rect 4148 26020 4157 26060
rect 23779 26020 23788 26060
rect 23828 26020 25996 26060
rect 26036 26020 26045 26060
rect 31276 26020 37516 26060
rect 37556 26020 37565 26060
rect 38371 26020 38380 26060
rect 38420 26020 39724 26060
rect 39764 26020 39773 26060
rect 2371 25852 2380 25892
rect 2420 25852 3244 25892
rect 3284 25852 3293 25892
rect 36931 25852 36940 25892
rect 36980 25852 40300 25892
rect 40340 25852 40349 25892
rect 40675 25852 40684 25892
rect 40724 25852 43756 25892
rect 43796 25852 43805 25892
rect 0 25748 80 25828
rect 3103 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 3489 25724
rect 18223 25684 18232 25724
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18600 25684 18609 25724
rect 33343 25684 33352 25724
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33720 25684 33729 25724
rect 48463 25684 48472 25724
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48840 25684 48849 25724
rect 63583 25684 63592 25724
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63960 25684 63969 25724
rect 78703 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 79089 25724
rect 93823 25684 93832 25724
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 94200 25684 94209 25724
rect 18115 25516 18124 25556
rect 18164 25516 18988 25556
rect 19028 25516 19037 25556
rect 25987 25516 25996 25556
rect 26036 25516 26668 25556
rect 26708 25516 26717 25556
rect 30883 25516 30892 25556
rect 30932 25516 31852 25556
rect 31892 25516 31901 25556
rect 32803 25348 32812 25388
rect 32852 25348 34540 25388
rect 34580 25348 34589 25388
rect 39619 25348 39628 25388
rect 39668 25348 41260 25388
rect 41300 25348 41309 25388
rect 17251 25264 17260 25304
rect 17300 25264 17836 25304
rect 17876 25264 17885 25304
rect 22243 25264 22252 25304
rect 22292 25264 22828 25304
rect 22868 25264 22877 25304
rect 23203 25264 23212 25304
rect 23252 25264 27820 25304
rect 27860 25264 27869 25304
rect 35011 25264 35020 25304
rect 35060 25264 43372 25304
rect 43412 25264 43421 25304
rect 13987 25180 13996 25220
rect 14036 25180 15628 25220
rect 15668 25180 15677 25220
rect 41347 25180 41356 25220
rect 41396 25180 41740 25220
rect 41780 25180 41789 25220
rect 43267 25180 43276 25220
rect 43316 25180 46348 25220
rect 46388 25180 47308 25220
rect 47348 25180 47357 25220
rect 21955 25096 21964 25136
rect 22004 25096 23308 25136
rect 23348 25096 23357 25136
rect 0 24908 80 24988
rect 4343 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 4729 24968
rect 19463 24928 19472 24968
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19840 24928 19849 24968
rect 34583 24928 34592 24968
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34960 24928 34969 24968
rect 49703 24928 49712 24968
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 50080 24928 50089 24968
rect 64823 24928 64832 24968
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 65200 24928 65209 24968
rect 79943 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 80329 24968
rect 95063 24928 95072 24968
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95440 24928 95449 24968
rect 37891 24760 37900 24800
rect 37940 24760 38668 24800
rect 38708 24760 38956 24800
rect 38996 24760 39532 24800
rect 39572 24760 39581 24800
rect 18595 24592 18604 24632
rect 18644 24592 19084 24632
rect 19124 24592 19133 24632
rect 31747 24592 31756 24632
rect 31796 24592 32236 24632
rect 32276 24592 32285 24632
rect 36835 24340 36844 24380
rect 36884 24340 37708 24380
rect 37748 24340 37757 24380
rect 3103 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 3489 24212
rect 18223 24172 18232 24212
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18600 24172 18609 24212
rect 33343 24172 33352 24212
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33720 24172 33729 24212
rect 48463 24172 48472 24212
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48840 24172 48849 24212
rect 63583 24172 63592 24212
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63960 24172 63969 24212
rect 78703 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 79089 24212
rect 93823 24172 93832 24212
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 94200 24172 94209 24212
rect 0 24068 80 24148
rect 41635 23836 41644 23876
rect 41684 23836 42892 23876
rect 42932 23836 42941 23876
rect 8803 23752 8812 23792
rect 8852 23752 10060 23792
rect 10100 23752 10348 23792
rect 10388 23752 10397 23792
rect 14755 23752 14764 23792
rect 14804 23752 16492 23792
rect 16532 23752 16541 23792
rect 18595 23752 18604 23792
rect 18644 23752 19372 23792
rect 19412 23752 19421 23792
rect 37219 23752 37228 23792
rect 37268 23752 37516 23792
rect 37556 23752 37804 23792
rect 37844 23752 37853 23792
rect 38083 23752 38092 23792
rect 38132 23752 42316 23792
rect 42356 23752 42365 23792
rect 42787 23752 42796 23792
rect 42836 23752 43756 23792
rect 43796 23752 43805 23792
rect 6307 23668 6316 23708
rect 6356 23668 9100 23708
rect 9140 23668 9149 23708
rect 3619 23584 3628 23624
rect 3668 23584 4300 23624
rect 4340 23584 4492 23624
rect 4532 23584 6124 23624
rect 6164 23584 6173 23624
rect 11491 23584 11500 23624
rect 11540 23584 12844 23624
rect 12884 23584 12893 23624
rect 43363 23584 43372 23624
rect 43412 23584 45964 23624
rect 46004 23584 46013 23624
rect 4343 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 4729 23456
rect 19463 23416 19472 23456
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19840 23416 19849 23456
rect 34583 23416 34592 23456
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34960 23416 34969 23456
rect 41560 23416 42220 23456
rect 42260 23416 42796 23456
rect 42836 23416 42845 23456
rect 49703 23416 49712 23456
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 50080 23416 50089 23456
rect 64823 23416 64832 23456
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 65200 23416 65209 23456
rect 79943 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 80329 23456
rect 95063 23416 95072 23456
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95440 23416 95449 23456
rect 0 23228 80 23308
rect 41560 23288 41600 23416
rect 259 23248 268 23288
rect 308 23248 25708 23288
rect 25748 23248 26188 23288
rect 26228 23248 26237 23288
rect 39043 23248 39052 23288
rect 39092 23248 41600 23288
rect 5731 23164 5740 23204
rect 5780 23164 7564 23204
rect 7604 23164 7613 23204
rect 4195 23080 4204 23120
rect 4244 23080 5260 23120
rect 5300 23080 5309 23120
rect 12835 23080 12844 23120
rect 12884 23080 14476 23120
rect 14516 23080 14525 23120
rect 21859 23080 21868 23120
rect 21908 23080 22732 23120
rect 22772 23080 22781 23120
rect 23971 23080 23980 23120
rect 24020 23080 24844 23120
rect 24884 23080 24893 23120
rect 29443 23080 29452 23120
rect 29492 23080 29644 23120
rect 29684 23080 31660 23120
rect 31700 23080 31709 23120
rect 33763 23080 33772 23120
rect 33812 23080 35020 23120
rect 35060 23080 35069 23120
rect 42307 23080 42316 23120
rect 42356 23080 43852 23120
rect 43892 23080 44716 23120
rect 44756 23080 49132 23120
rect 49172 23080 49181 23120
rect 3043 22996 3052 23036
rect 3092 22996 7948 23036
rect 7988 22996 10156 23036
rect 10196 22996 10205 23036
rect 32035 22996 32044 23036
rect 32084 22996 32524 23036
rect 32564 22996 33964 23036
rect 34004 22996 34013 23036
rect 42979 22996 42988 23036
rect 43028 22996 43276 23036
rect 43316 22996 45580 23036
rect 45620 22996 48268 23036
rect 48308 22996 48940 23036
rect 48980 22996 48989 23036
rect 9955 22828 9964 22868
rect 10004 22828 11116 22868
rect 11156 22828 11165 22868
rect 13507 22828 13516 22868
rect 13556 22828 13900 22868
rect 13940 22828 13949 22868
rect 19747 22828 19756 22868
rect 19796 22828 20236 22868
rect 20276 22828 20285 22868
rect 29827 22828 29836 22868
rect 29876 22828 30604 22868
rect 30644 22828 30653 22868
rect 37411 22828 37420 22868
rect 37460 22828 38764 22868
rect 38804 22828 38813 22868
rect 3103 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 3489 22700
rect 4195 22660 4204 22700
rect 4244 22660 5548 22700
rect 5588 22660 5597 22700
rect 18223 22660 18232 22700
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18600 22660 18609 22700
rect 33343 22660 33352 22700
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33720 22660 33729 22700
rect 48463 22660 48472 22700
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48840 22660 48849 22700
rect 63583 22660 63592 22700
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63960 22660 63969 22700
rect 78703 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 79089 22700
rect 93823 22660 93832 22700
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 94200 22660 94209 22700
rect 3619 22492 3628 22532
rect 3668 22492 4300 22532
rect 4340 22492 4492 22532
rect 4532 22492 6028 22532
rect 6068 22492 6077 22532
rect 0 22388 80 22468
rect 11587 22408 11596 22448
rect 11636 22408 14092 22448
rect 14132 22408 14141 22448
rect 16483 22324 16492 22364
rect 16532 22324 20140 22364
rect 20180 22324 22444 22364
rect 22484 22324 22493 22364
rect 31276 22324 32524 22364
rect 32564 22324 32573 22364
rect 31276 22280 31316 22324
rect 14083 22240 14092 22280
rect 14132 22240 14860 22280
rect 14900 22240 14909 22280
rect 17347 22240 17356 22280
rect 17396 22240 20332 22280
rect 20372 22240 21004 22280
rect 21044 22240 21053 22280
rect 22915 22240 22924 22280
rect 22964 22240 23212 22280
rect 23252 22240 23980 22280
rect 24020 22240 24029 22280
rect 30211 22240 30220 22280
rect 30260 22240 31276 22280
rect 31316 22240 31325 22280
rect 31555 22240 31564 22280
rect 31604 22240 33100 22280
rect 33140 22240 33388 22280
rect 33428 22240 33437 22280
rect 47971 22240 47980 22280
rect 48020 22240 49708 22280
rect 49748 22240 49757 22280
rect 4343 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 4729 21944
rect 19463 21904 19472 21944
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19840 21904 19849 21944
rect 34583 21904 34592 21944
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34960 21904 34969 21944
rect 49703 21904 49712 21944
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 50080 21904 50089 21944
rect 64823 21904 64832 21944
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 65200 21904 65209 21944
rect 79943 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 80329 21944
rect 95063 21904 95072 21944
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95440 21904 95449 21944
rect 14851 21736 14860 21776
rect 14900 21736 15244 21776
rect 15284 21736 15293 21776
rect 31267 21736 31276 21776
rect 31316 21736 31852 21776
rect 31892 21736 33772 21776
rect 33812 21736 33821 21776
rect 47875 21736 47884 21776
rect 47924 21736 48076 21776
rect 48116 21736 48125 21776
rect 2659 21652 2668 21692
rect 2708 21652 3436 21692
rect 3476 21652 3485 21692
rect 0 21608 80 21628
rect 0 21568 652 21608
rect 692 21568 701 21608
rect 22435 21568 22444 21608
rect 22484 21568 22828 21608
rect 22868 21568 22877 21608
rect 30211 21568 30220 21608
rect 30260 21568 30700 21608
rect 30740 21568 30749 21608
rect 0 21548 80 21568
rect 49219 21484 49228 21524
rect 49268 21484 50284 21524
rect 50324 21484 50333 21524
rect 19939 21400 19948 21440
rect 19988 21400 21004 21440
rect 21044 21400 21053 21440
rect 39811 21400 39820 21440
rect 39860 21400 40492 21440
rect 40532 21400 40541 21440
rect 48259 21400 48268 21440
rect 48308 21400 49420 21440
rect 49460 21400 49469 21440
rect 3103 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 3489 21188
rect 18223 21148 18232 21188
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18600 21148 18609 21188
rect 33343 21148 33352 21188
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33720 21148 33729 21188
rect 48463 21148 48472 21188
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48840 21148 48849 21188
rect 63583 21148 63592 21188
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63960 21148 63969 21188
rect 78703 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 79089 21188
rect 93823 21148 93832 21188
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 94200 21148 94209 21188
rect 21091 20812 21100 20852
rect 21140 20812 21964 20852
rect 22004 20812 22013 20852
rect 26083 20812 26092 20852
rect 26132 20812 26572 20852
rect 26612 20812 26860 20852
rect 26900 20812 26909 20852
rect 0 20768 80 20788
rect 0 20728 652 20768
rect 692 20728 701 20768
rect 13987 20728 13996 20768
rect 14036 20728 14572 20768
rect 14612 20728 22924 20768
rect 22964 20728 22973 20768
rect 0 20708 80 20728
rect 4343 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 4729 20432
rect 19463 20392 19472 20432
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19840 20392 19849 20432
rect 34583 20392 34592 20432
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34960 20392 34969 20432
rect 49703 20392 49712 20432
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 50080 20392 50089 20432
rect 64823 20392 64832 20432
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 65200 20392 65209 20432
rect 79943 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 80329 20432
rect 95063 20392 95072 20432
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95440 20392 95449 20432
rect 2851 20140 2860 20180
rect 2900 20140 3628 20180
rect 3668 20140 4108 20180
rect 4148 20140 4157 20180
rect 9091 20140 9100 20180
rect 9140 20140 9484 20180
rect 9524 20140 9868 20180
rect 9908 20140 13420 20180
rect 13460 20140 14188 20180
rect 14228 20140 14237 20180
rect 24931 20140 24940 20180
rect 24980 20140 25900 20180
rect 25940 20140 25949 20180
rect 32740 20140 33196 20180
rect 33236 20140 34924 20180
rect 34964 20140 34973 20180
rect 39820 20140 40588 20180
rect 40628 20140 40637 20180
rect 49795 20140 49804 20180
rect 49844 20140 50476 20180
rect 50516 20140 50525 20180
rect 32740 20096 32780 20140
rect 39820 20096 39860 20140
rect 67 20056 76 20096
rect 116 20056 23960 20096
rect 26179 20056 26188 20096
rect 26228 20056 29164 20096
rect 29204 20056 29356 20096
rect 29396 20056 29405 20096
rect 30115 20056 30124 20096
rect 30164 20056 32780 20096
rect 34051 20056 34060 20096
rect 34100 20056 36076 20096
rect 36116 20056 36125 20096
rect 37315 20056 37324 20096
rect 37364 20056 38668 20096
rect 38708 20056 38717 20096
rect 39811 20056 39820 20096
rect 39860 20056 39869 20096
rect 41560 20056 41740 20096
rect 41780 20056 41789 20096
rect 48163 20056 48172 20096
rect 48212 20056 49324 20096
rect 49364 20056 49373 20096
rect 23920 20012 23960 20056
rect 41560 20012 41600 20056
rect 23920 19972 30412 20012
rect 30452 19972 30461 20012
rect 40867 19972 40876 20012
rect 40916 19972 41600 20012
rect 0 19928 80 19948
rect 0 19888 652 19928
rect 692 19888 701 19928
rect 0 19868 80 19888
rect 23299 19804 23308 19844
rect 23348 19804 30796 19844
rect 30836 19804 30845 19844
rect 38467 19804 38476 19844
rect 38516 19804 38956 19844
rect 38996 19804 39340 19844
rect 39380 19804 39389 19844
rect 3103 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 3489 19676
rect 18223 19636 18232 19676
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18600 19636 18609 19676
rect 33343 19636 33352 19676
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33720 19636 33729 19676
rect 48463 19636 48472 19676
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48840 19636 48849 19676
rect 63583 19636 63592 19676
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63960 19636 63969 19676
rect 78703 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 79089 19676
rect 93823 19636 93832 19676
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 94200 19636 94209 19676
rect 31459 19468 31468 19508
rect 31508 19468 33772 19508
rect 33812 19468 36940 19508
rect 36980 19468 36989 19508
rect 47587 19216 47596 19256
rect 47636 19216 47980 19256
rect 48020 19216 48029 19256
rect 49411 19216 49420 19256
rect 49460 19216 50188 19256
rect 50228 19216 50237 19256
rect 46339 19132 46348 19172
rect 46388 19132 47212 19172
rect 47252 19132 47261 19172
rect 0 19088 80 19108
rect 0 19048 652 19088
rect 692 19048 701 19088
rect 1699 19048 1708 19088
rect 1748 19048 2668 19088
rect 2708 19048 2717 19088
rect 32227 19048 32236 19088
rect 32276 19048 35404 19088
rect 35444 19048 37324 19088
rect 37364 19048 38476 19088
rect 38516 19048 38525 19088
rect 39811 19048 39820 19088
rect 39860 19048 40684 19088
rect 40724 19048 40733 19088
rect 50659 19048 50668 19088
rect 50708 19048 52012 19088
rect 52052 19048 52061 19088
rect 0 19028 80 19048
rect 12067 18964 12076 19004
rect 12116 18964 13036 19004
rect 13076 18964 13085 19004
rect 4343 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 4729 18920
rect 19463 18880 19472 18920
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19840 18880 19849 18920
rect 29827 18880 29836 18920
rect 29876 18880 31180 18920
rect 31220 18880 31229 18920
rect 34583 18880 34592 18920
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34960 18880 34969 18920
rect 36451 18880 36460 18920
rect 36500 18880 37612 18920
rect 37652 18880 37661 18920
rect 49703 18880 49712 18920
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 50080 18880 50089 18920
rect 64823 18880 64832 18920
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 65200 18880 65209 18920
rect 79943 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 80329 18920
rect 95063 18880 95072 18920
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95440 18880 95449 18920
rect 7459 18712 7468 18752
rect 7508 18712 9964 18752
rect 10004 18712 10013 18752
rect 11011 18712 11020 18752
rect 11060 18712 11788 18752
rect 11828 18712 12268 18752
rect 12308 18712 12317 18752
rect 2947 18544 2956 18584
rect 2996 18544 3916 18584
rect 3956 18544 5356 18584
rect 5396 18544 5405 18584
rect 7939 18544 7948 18584
rect 7988 18544 9484 18584
rect 9524 18544 9533 18584
rect 23920 18544 26764 18584
rect 26804 18544 27284 18584
rect 47971 18544 47980 18584
rect 48020 18544 53260 18584
rect 53300 18544 53309 18584
rect 6787 18460 6796 18500
rect 6836 18460 7660 18500
rect 7700 18460 7709 18500
rect 23920 18332 23960 18544
rect 5635 18292 5644 18332
rect 5684 18292 6604 18332
rect 6644 18292 6653 18332
rect 21955 18292 21964 18332
rect 22004 18292 22828 18332
rect 22868 18292 23960 18332
rect 0 18248 80 18268
rect 27244 18248 27284 18544
rect 46819 18460 46828 18500
rect 46868 18460 47116 18500
rect 47156 18460 52300 18500
rect 52340 18460 52349 18500
rect 0 18208 652 18248
rect 692 18208 701 18248
rect 27235 18208 27244 18248
rect 27284 18208 27293 18248
rect 0 18188 80 18208
rect 3103 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 3489 18164
rect 18223 18124 18232 18164
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18600 18124 18609 18164
rect 25507 18124 25516 18164
rect 25556 18124 30316 18164
rect 30356 18124 30365 18164
rect 33343 18124 33352 18164
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33720 18124 33729 18164
rect 48463 18124 48472 18164
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48840 18124 48849 18164
rect 63583 18124 63592 18164
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63960 18124 63969 18164
rect 78703 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 79089 18164
rect 93823 18124 93832 18164
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 94200 18124 94209 18164
rect 7651 17956 7660 17996
rect 7700 17956 8812 17996
rect 8852 17956 8861 17996
rect 25123 17956 25132 17996
rect 25172 17956 25900 17996
rect 25940 17956 25949 17996
rect 26659 17956 26668 17996
rect 26708 17956 27532 17996
rect 27572 17956 27581 17996
rect 46723 17956 46732 17996
rect 46772 17956 47596 17996
rect 47636 17956 47645 17996
rect 47779 17956 47788 17996
rect 47828 17956 48172 17996
rect 48212 17956 48556 17996
rect 48596 17956 49612 17996
rect 49652 17956 49661 17996
rect 23971 17872 23980 17912
rect 24020 17872 24652 17912
rect 24692 17872 26476 17912
rect 26516 17872 26525 17912
rect 4492 17788 6028 17828
rect 6068 17788 6077 17828
rect 26083 17788 26092 17828
rect 26132 17788 26668 17828
rect 26708 17788 26717 17828
rect 32323 17788 32332 17828
rect 32372 17788 32780 17828
rect 41539 17788 41548 17828
rect 41588 17788 41932 17828
rect 41972 17788 41981 17828
rect 47395 17788 47404 17828
rect 47444 17788 48076 17828
rect 48116 17788 48125 17828
rect 4492 17744 4532 17788
rect 32740 17744 32780 17788
rect 2083 17704 2092 17744
rect 2132 17704 4492 17744
rect 4532 17704 4541 17744
rect 5347 17704 5356 17744
rect 5396 17704 6988 17744
rect 7028 17704 7037 17744
rect 8035 17704 8044 17744
rect 8084 17704 8332 17744
rect 8372 17704 8381 17744
rect 8995 17704 9004 17744
rect 9044 17704 11020 17744
rect 11060 17704 11069 17744
rect 17635 17704 17644 17744
rect 17684 17704 18700 17744
rect 18740 17704 18988 17744
rect 19028 17704 19372 17744
rect 19412 17704 22252 17744
rect 22292 17704 22301 17744
rect 26563 17704 26572 17744
rect 26612 17704 27820 17744
rect 27860 17704 27869 17744
rect 30307 17704 30316 17744
rect 30356 17704 31372 17744
rect 31412 17704 31421 17744
rect 32740 17704 33868 17744
rect 33908 17704 33917 17744
rect 39619 17704 39628 17744
rect 39668 17704 41452 17744
rect 41492 17704 41501 17744
rect 41827 17704 41836 17744
rect 41876 17704 43468 17744
rect 43508 17704 43517 17744
rect 4099 17620 4108 17660
rect 4148 17620 5260 17660
rect 5300 17620 5309 17660
rect 11971 17620 11980 17660
rect 12020 17620 12172 17660
rect 12212 17620 12940 17660
rect 12980 17620 14284 17660
rect 14324 17620 14333 17660
rect 18883 17620 18892 17660
rect 18932 17620 20428 17660
rect 20468 17620 20477 17660
rect 20995 17620 21004 17660
rect 21044 17620 21772 17660
rect 21812 17620 21821 17660
rect 23971 17620 23980 17660
rect 24020 17620 26380 17660
rect 26420 17620 26429 17660
rect 28003 17620 28012 17660
rect 28052 17620 29932 17660
rect 29972 17620 29981 17660
rect 18499 17452 18508 17492
rect 18548 17452 19276 17492
rect 19316 17452 21868 17492
rect 21908 17452 25516 17492
rect 25556 17452 25565 17492
rect 0 17408 80 17428
rect 0 17368 652 17408
rect 692 17368 701 17408
rect 4343 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 4729 17408
rect 19463 17368 19472 17408
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19840 17368 19849 17408
rect 34583 17368 34592 17408
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34960 17368 34969 17408
rect 49703 17368 49712 17408
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 50080 17368 50089 17408
rect 64823 17368 64832 17408
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 65200 17368 65209 17408
rect 79943 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 80329 17408
rect 95063 17368 95072 17408
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95440 17368 95449 17408
rect 0 17348 80 17368
rect 6019 17116 6028 17156
rect 6068 17116 10156 17156
rect 10196 17116 11116 17156
rect 11156 17116 11308 17156
rect 11348 17116 11357 17156
rect 22723 17116 22732 17156
rect 22772 17116 23788 17156
rect 23828 17116 23837 17156
rect 27331 17116 27340 17156
rect 27380 17116 30988 17156
rect 31028 17116 31037 17156
rect 34051 17116 34060 17156
rect 34100 17116 36172 17156
rect 36212 17116 36221 17156
rect 40396 17116 41356 17156
rect 41396 17116 41405 17156
rect 40396 17072 40436 17116
rect 17251 17032 17260 17072
rect 17300 17032 17644 17072
rect 17684 17032 17693 17072
rect 18115 17032 18124 17072
rect 18164 17032 18508 17072
rect 18548 17032 18557 17072
rect 21379 17032 21388 17072
rect 21428 17032 23116 17072
rect 23156 17032 23165 17072
rect 37603 17032 37612 17072
rect 37652 17032 40396 17072
rect 40436 17032 40445 17072
rect 41251 17032 41260 17072
rect 41300 17032 42316 17072
rect 42356 17032 42700 17072
rect 42740 17032 42749 17072
rect 5443 16948 5452 16988
rect 5492 16948 7372 16988
rect 7412 16948 8236 16988
rect 8276 16948 8285 16988
rect 8419 16948 8428 16988
rect 8468 16948 10348 16988
rect 10388 16948 11884 16988
rect 11924 16948 11933 16988
rect 41347 16948 41356 16988
rect 41396 16948 41740 16988
rect 41780 16948 41789 16988
rect 12355 16780 12364 16820
rect 12404 16780 13132 16820
rect 13172 16780 13181 16820
rect 33379 16780 33388 16820
rect 33428 16780 34924 16820
rect 34964 16780 34973 16820
rect 41539 16780 41548 16820
rect 41588 16780 42412 16820
rect 42452 16780 42461 16820
rect 3103 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 3489 16652
rect 18223 16612 18232 16652
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18600 16612 18609 16652
rect 33343 16612 33352 16652
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33720 16612 33729 16652
rect 48463 16612 48472 16652
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48840 16612 48849 16652
rect 63583 16612 63592 16652
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63960 16612 63969 16652
rect 78703 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 79089 16652
rect 93823 16612 93832 16652
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 94200 16612 94209 16652
rect 0 16568 80 16588
rect 0 16528 652 16568
rect 692 16528 701 16568
rect 0 16508 80 16528
rect 9475 16192 9484 16232
rect 9524 16192 12652 16232
rect 12692 16192 12701 16232
rect 4343 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 4729 15896
rect 19463 15856 19472 15896
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19840 15856 19849 15896
rect 34583 15856 34592 15896
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34960 15856 34969 15896
rect 49703 15856 49712 15896
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 50080 15856 50089 15896
rect 64823 15856 64832 15896
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 65200 15856 65209 15896
rect 79943 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 80329 15896
rect 95063 15856 95072 15896
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95440 15856 95449 15896
rect 55939 15772 55948 15812
rect 55988 15772 57676 15812
rect 57716 15772 57725 15812
rect 0 15728 80 15748
rect 0 15688 556 15728
rect 596 15688 605 15728
rect 42595 15688 42604 15728
rect 42644 15688 44332 15728
rect 44372 15688 45100 15728
rect 45140 15688 45149 15728
rect 0 15668 80 15688
rect 48355 15604 48364 15644
rect 48404 15604 49228 15644
rect 49268 15604 49277 15644
rect 35683 15520 35692 15560
rect 35732 15520 36268 15560
rect 36308 15520 36317 15560
rect 27619 15436 27628 15476
rect 27668 15436 34060 15476
rect 34100 15436 42604 15476
rect 42644 15436 42653 15476
rect 51619 15436 51628 15476
rect 51668 15436 52780 15476
rect 52820 15436 53452 15476
rect 53492 15436 53501 15476
rect 35971 15268 35980 15308
rect 36020 15268 36748 15308
rect 36788 15268 36797 15308
rect 51427 15268 51436 15308
rect 51476 15268 52108 15308
rect 52148 15268 52157 15308
rect 3103 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 3489 15140
rect 18223 15100 18232 15140
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18600 15100 18609 15140
rect 33343 15100 33352 15140
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33720 15100 33729 15140
rect 48463 15100 48472 15140
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48840 15100 48849 15140
rect 63583 15100 63592 15140
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63960 15100 63969 15140
rect 78703 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 79089 15140
rect 93823 15100 93832 15140
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 94200 15100 94209 15140
rect 0 14888 80 14908
rect 0 14848 652 14888
rect 692 14848 701 14888
rect 21667 14848 21676 14888
rect 21716 14848 23116 14888
rect 23156 14848 23165 14888
rect 0 14828 80 14848
rect 9763 14680 9772 14720
rect 9812 14680 18892 14720
rect 18932 14680 23308 14720
rect 23348 14680 23357 14720
rect 40867 14680 40876 14720
rect 40916 14680 41548 14720
rect 41588 14680 41597 14720
rect 46051 14680 46060 14720
rect 46100 14680 46636 14720
rect 46676 14680 49612 14720
rect 49652 14680 52204 14720
rect 52244 14680 52253 14720
rect 52771 14680 52780 14720
rect 52820 14680 54796 14720
rect 54836 14680 54845 14720
rect 40195 14596 40204 14636
rect 40244 14596 40780 14636
rect 40820 14596 40829 14636
rect 51331 14596 51340 14636
rect 51380 14596 52876 14636
rect 52916 14596 52925 14636
rect 50371 14512 50380 14552
rect 50420 14512 51628 14552
rect 51668 14512 51677 14552
rect 56995 14512 57004 14552
rect 57044 14512 57964 14552
rect 58004 14512 58013 14552
rect 4343 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 4729 14384
rect 19463 14344 19472 14384
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19840 14344 19849 14384
rect 34583 14344 34592 14384
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34960 14344 34969 14384
rect 49703 14344 49712 14384
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 50080 14344 50089 14384
rect 64823 14344 64832 14384
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 65200 14344 65209 14384
rect 79943 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 80329 14384
rect 95063 14344 95072 14384
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95440 14344 95449 14384
rect 51235 14260 51244 14300
rect 51284 14260 52684 14300
rect 52724 14260 53068 14300
rect 53108 14260 53117 14300
rect 51235 14092 51244 14132
rect 51284 14092 52876 14132
rect 52916 14092 52925 14132
rect 56323 14092 56332 14132
rect 56372 14092 56812 14132
rect 56852 14092 56861 14132
rect 0 14048 80 14068
rect 0 14008 652 14048
rect 692 14008 701 14048
rect 14659 14008 14668 14048
rect 14708 14008 15148 14048
rect 15188 14008 15197 14048
rect 16387 14008 16396 14048
rect 16436 14008 18124 14048
rect 18164 14008 18173 14048
rect 18595 14008 18604 14048
rect 18644 14008 19084 14048
rect 19124 14008 19660 14048
rect 19700 14008 19709 14048
rect 32515 14008 32524 14048
rect 32564 14008 33676 14048
rect 33716 14008 33725 14048
rect 39619 14008 39628 14048
rect 39668 14008 40300 14048
rect 40340 14008 40349 14048
rect 41251 14008 41260 14048
rect 41300 14008 42124 14048
rect 42164 14008 42173 14048
rect 47875 14008 47884 14048
rect 47924 14008 49996 14048
rect 50036 14008 50420 14048
rect 0 13988 80 14008
rect 50380 13964 50420 14008
rect 18403 13924 18412 13964
rect 18452 13924 18988 13964
rect 19028 13924 19037 13964
rect 50380 13924 56716 13964
rect 56756 13924 57292 13964
rect 57332 13924 57341 13964
rect 12259 13840 12268 13880
rect 12308 13840 12844 13880
rect 12884 13840 12893 13880
rect 17347 13840 17356 13880
rect 17396 13840 18700 13880
rect 18740 13840 18749 13880
rect 23875 13840 23884 13880
rect 23924 13840 25132 13880
rect 25172 13840 25181 13880
rect 25315 13840 25324 13880
rect 25364 13840 25900 13880
rect 25940 13840 28876 13880
rect 28916 13840 28925 13880
rect 39907 13840 39916 13880
rect 39956 13840 42700 13880
rect 42740 13840 42749 13880
rect 47971 13840 47980 13880
rect 48020 13840 49612 13880
rect 49652 13840 49661 13880
rect 48355 13756 48364 13796
rect 48404 13756 50572 13796
rect 50612 13756 50621 13796
rect 3103 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 3489 13628
rect 18223 13588 18232 13628
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18600 13588 18609 13628
rect 33343 13588 33352 13628
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33720 13588 33729 13628
rect 48463 13588 48472 13628
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48840 13588 48849 13628
rect 63583 13588 63592 13628
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63960 13588 63969 13628
rect 78703 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 79089 13628
rect 93823 13588 93832 13628
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 94200 13588 94209 13628
rect 49987 13420 49996 13460
rect 50036 13420 50476 13460
rect 50516 13420 52972 13460
rect 53012 13420 53021 13460
rect 18691 13336 18700 13376
rect 18740 13336 20428 13376
rect 20468 13336 20477 13376
rect 19075 13252 19084 13292
rect 19124 13252 20236 13292
rect 20276 13252 20285 13292
rect 52195 13252 52204 13292
rect 52244 13252 52876 13292
rect 52916 13252 53836 13292
rect 53876 13252 53885 13292
rect 0 13208 80 13228
rect 0 13168 652 13208
rect 692 13168 701 13208
rect 2467 13168 2476 13208
rect 2516 13168 2956 13208
rect 2996 13168 3005 13208
rect 8035 13168 8044 13208
rect 8084 13168 9772 13208
rect 9812 13168 9821 13208
rect 11683 13168 11692 13208
rect 11732 13168 12652 13208
rect 12692 13168 13132 13208
rect 13172 13168 13181 13208
rect 19363 13168 19372 13208
rect 19412 13168 20332 13208
rect 20372 13168 20381 13208
rect 23491 13168 23500 13208
rect 23540 13168 24268 13208
rect 24308 13168 24317 13208
rect 28963 13168 28972 13208
rect 29012 13168 30508 13208
rect 30548 13168 30557 13208
rect 38467 13168 38476 13208
rect 38516 13168 39244 13208
rect 39284 13168 39532 13208
rect 39572 13168 39581 13208
rect 45283 13168 45292 13208
rect 45332 13168 47116 13208
rect 47156 13168 49132 13208
rect 49172 13168 49324 13208
rect 49364 13168 49373 13208
rect 50275 13168 50284 13208
rect 50324 13168 52300 13208
rect 52340 13168 54604 13208
rect 54644 13168 54653 13208
rect 0 13148 80 13168
rect 23299 13084 23308 13124
rect 23348 13084 28012 13124
rect 28052 13084 28061 13124
rect 27619 13000 27628 13040
rect 27668 13000 28396 13040
rect 28436 13000 28445 13040
rect 28579 13000 28588 13040
rect 28628 13000 29068 13040
rect 29108 13000 29452 13040
rect 29492 13000 32332 13040
rect 32372 13000 32381 13040
rect 45955 13000 45964 13040
rect 46004 13000 46828 13040
rect 46868 13000 46877 13040
rect 55075 13000 55084 13040
rect 55124 13000 56140 13040
rect 56180 13000 56428 13040
rect 56468 13000 57484 13040
rect 57524 13000 57533 13040
rect 4343 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 4729 12872
rect 19463 12832 19472 12872
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19840 12832 19849 12872
rect 34583 12832 34592 12872
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34960 12832 34969 12872
rect 49703 12832 49712 12872
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 50080 12832 50089 12872
rect 64823 12832 64832 12872
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 65200 12832 65209 12872
rect 79943 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 80329 12872
rect 95063 12832 95072 12872
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95440 12832 95449 12872
rect 55171 12664 55180 12704
rect 55220 12664 56428 12704
rect 56468 12664 57676 12704
rect 57716 12664 57725 12704
rect 8611 12580 8620 12620
rect 8660 12580 9196 12620
rect 9236 12580 9245 12620
rect 9859 12580 9868 12620
rect 9908 12580 11692 12620
rect 11732 12580 11741 12620
rect 18787 12580 18796 12620
rect 18836 12580 19948 12620
rect 19988 12580 19997 12620
rect 25123 12580 25132 12620
rect 25172 12580 28876 12620
rect 28916 12580 32620 12620
rect 32660 12580 35020 12620
rect 35060 12580 35069 12620
rect 55459 12580 55468 12620
rect 55508 12580 56716 12620
rect 56756 12580 56765 12620
rect 3331 12496 3340 12536
rect 3380 12496 3628 12536
rect 3668 12496 3820 12536
rect 3860 12496 3869 12536
rect 10723 12496 10732 12536
rect 10772 12496 13516 12536
rect 13556 12496 13565 12536
rect 17251 12496 17260 12536
rect 17300 12496 18508 12536
rect 18548 12496 19852 12536
rect 19892 12496 19901 12536
rect 20131 12496 20140 12536
rect 20180 12496 21292 12536
rect 21332 12496 21341 12536
rect 33475 12496 33484 12536
rect 33524 12496 36172 12536
rect 36212 12496 36221 12536
rect 2371 12412 2380 12452
rect 2420 12412 3532 12452
rect 3572 12412 3581 12452
rect 6280 12412 6604 12452
rect 6644 12412 11212 12452
rect 11252 12412 11261 12452
rect 18787 12412 18796 12452
rect 18836 12412 19660 12452
rect 19700 12412 19709 12452
rect 31171 12412 31180 12452
rect 31220 12412 32236 12452
rect 32276 12412 33772 12452
rect 33812 12412 33821 12452
rect 0 12368 80 12388
rect 6280 12368 6320 12412
rect 0 12328 652 12368
rect 692 12328 701 12368
rect 2947 12328 2956 12368
rect 2996 12328 3724 12368
rect 3764 12328 6320 12368
rect 0 12308 80 12328
rect 21955 12244 21964 12284
rect 22004 12244 23020 12284
rect 23060 12244 23069 12284
rect 3103 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 3489 12116
rect 18223 12076 18232 12116
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18600 12076 18609 12116
rect 33343 12076 33352 12116
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33720 12076 33729 12116
rect 48463 12076 48472 12116
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48840 12076 48849 12116
rect 63583 12076 63592 12116
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63960 12076 63969 12116
rect 78703 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 79089 12116
rect 93823 12076 93832 12116
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 94200 12076 94209 12116
rect 33955 11908 33964 11948
rect 34004 11908 34444 11948
rect 34484 11908 34493 11948
rect 3523 11740 3532 11780
rect 3572 11740 3916 11780
rect 3956 11740 3965 11780
rect 4003 11656 4012 11696
rect 4052 11656 5164 11696
rect 5204 11656 5213 11696
rect 16291 11656 16300 11696
rect 16340 11656 17164 11696
rect 17204 11656 17213 11696
rect 28003 11656 28012 11696
rect 28052 11656 28300 11696
rect 28340 11656 31468 11696
rect 31508 11656 31948 11696
rect 31988 11656 31997 11696
rect 32323 11656 32332 11696
rect 32372 11656 32812 11696
rect 32852 11656 32861 11696
rect 0 11528 80 11548
rect 0 11488 652 11528
rect 692 11488 701 11528
rect 3427 11488 3436 11528
rect 3476 11488 4108 11528
rect 4148 11488 4300 11528
rect 4340 11488 5356 11528
rect 5396 11488 5405 11528
rect 0 11468 80 11488
rect 4343 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 4729 11360
rect 6280 11320 7180 11360
rect 7220 11320 8716 11360
rect 8756 11320 8765 11360
rect 19463 11320 19472 11360
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19840 11320 19849 11360
rect 31363 11320 31372 11360
rect 31412 11320 31852 11360
rect 31892 11320 32812 11360
rect 32852 11320 32861 11360
rect 34583 11320 34592 11360
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34960 11320 34969 11360
rect 36163 11320 36172 11360
rect 36212 11320 38956 11360
rect 38996 11320 39005 11360
rect 49703 11320 49712 11360
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 50080 11320 50089 11360
rect 64823 11320 64832 11360
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 65200 11320 65209 11360
rect 79943 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 80329 11360
rect 95063 11320 95072 11360
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95440 11320 95449 11360
rect 6280 11276 6320 11320
rect 4195 11236 4204 11276
rect 4244 11236 6320 11276
rect 54019 11152 54028 11192
rect 54068 11152 54700 11192
rect 54740 11152 55084 11192
rect 55124 11152 55756 11192
rect 55796 11152 55805 11192
rect 40867 11068 40876 11108
rect 40916 11068 43660 11108
rect 43700 11068 43709 11108
rect 19363 10984 19372 11024
rect 19412 10984 23404 11024
rect 23444 10984 23453 11024
rect 38371 10984 38380 11024
rect 38420 10984 39916 11024
rect 39956 10984 40300 11024
rect 40340 10984 40349 11024
rect 41155 10732 41164 10772
rect 41204 10732 44332 10772
rect 44372 10732 44381 10772
rect 52771 10732 52780 10772
rect 52820 10732 53836 10772
rect 53876 10732 53885 10772
rect 0 10688 80 10708
rect 0 10648 652 10688
rect 692 10648 701 10688
rect 0 10628 80 10648
rect 3103 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 3489 10604
rect 18223 10564 18232 10604
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18600 10564 18609 10604
rect 33343 10564 33352 10604
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33720 10564 33729 10604
rect 48463 10564 48472 10604
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48840 10564 48849 10604
rect 63583 10564 63592 10604
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63960 10564 63969 10604
rect 78703 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 79089 10604
rect 93823 10564 93832 10604
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 94200 10564 94209 10604
rect 54883 10312 54892 10352
rect 54932 10312 55564 10352
rect 55604 10312 55613 10352
rect 47011 10228 47020 10268
rect 47060 10228 48460 10268
rect 48500 10228 48509 10268
rect 55747 10228 55756 10268
rect 55796 10228 55948 10268
rect 55988 10228 56620 10268
rect 56660 10228 56669 10268
rect 14275 10144 14284 10184
rect 14324 10144 16012 10184
rect 16052 10144 16061 10184
rect 20227 10144 20236 10184
rect 20276 10144 24268 10184
rect 24308 10144 24317 10184
rect 31075 10144 31084 10184
rect 31124 10144 31660 10184
rect 31700 10144 31709 10184
rect 47107 10144 47116 10184
rect 47156 10144 47884 10184
rect 47924 10144 47933 10184
rect 48547 10144 48556 10184
rect 48596 10144 49804 10184
rect 49844 10144 49853 10184
rect 50275 10144 50284 10184
rect 50324 10144 50764 10184
rect 50804 10144 50813 10184
rect 931 10060 940 10100
rect 980 10060 25420 10100
rect 25460 10060 25469 10100
rect 46531 10060 46540 10100
rect 46580 10060 47308 10100
rect 47348 10060 47357 10100
rect 0 9848 80 9868
rect 0 9808 652 9848
rect 692 9808 701 9848
rect 4343 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 4729 9848
rect 19463 9808 19472 9848
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19840 9808 19849 9848
rect 34583 9808 34592 9848
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34960 9808 34969 9848
rect 49703 9808 49712 9848
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 50080 9808 50089 9848
rect 64823 9808 64832 9848
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 65200 9808 65209 9848
rect 79943 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 80329 9848
rect 95063 9808 95072 9848
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95440 9808 95449 9848
rect 0 9788 80 9808
rect 2947 9640 2956 9680
rect 2996 9640 3340 9680
rect 3380 9640 4396 9680
rect 4436 9640 5260 9680
rect 5300 9640 5309 9680
rect 40579 9640 40588 9680
rect 40628 9640 41356 9680
rect 41396 9640 41405 9680
rect 44995 9640 45004 9680
rect 45044 9640 47212 9680
rect 47252 9640 47261 9680
rect 51811 9640 51820 9680
rect 51860 9640 53164 9680
rect 53204 9640 53213 9680
rect 3235 9556 3244 9596
rect 3284 9556 5452 9596
rect 5492 9556 5501 9596
rect 18883 9556 18892 9596
rect 18932 9556 19660 9596
rect 19700 9556 19709 9596
rect 2467 9472 2476 9512
rect 2516 9472 3148 9512
rect 3188 9472 3532 9512
rect 3572 9472 3581 9512
rect 10051 9472 10060 9512
rect 10100 9472 11212 9512
rect 11252 9472 12268 9512
rect 12308 9472 12317 9512
rect 13123 9472 13132 9512
rect 13172 9472 17164 9512
rect 17204 9472 17213 9512
rect 25507 9472 25516 9512
rect 25556 9472 26380 9512
rect 26420 9472 26764 9512
rect 26804 9472 26813 9512
rect 40195 9472 40204 9512
rect 40244 9472 41548 9512
rect 41588 9472 41597 9512
rect 47683 9472 47692 9512
rect 47732 9472 48556 9512
rect 48596 9472 48605 9512
rect 53059 9472 53068 9512
rect 53108 9472 55276 9512
rect 55316 9472 55325 9512
rect 25987 9428 26045 9429
rect 25902 9388 25996 9428
rect 26036 9388 26045 9428
rect 25987 9387 26045 9388
rect 25795 9304 25804 9344
rect 25844 9304 26188 9344
rect 26228 9304 26237 9344
rect 25987 9260 26045 9261
rect 4771 9220 4780 9260
rect 4820 9220 5548 9260
rect 5588 9220 5597 9260
rect 20140 9220 25516 9260
rect 25556 9220 25565 9260
rect 25987 9220 25996 9260
rect 26036 9220 26668 9260
rect 26708 9220 26717 9260
rect 38755 9220 38764 9260
rect 38804 9220 39532 9260
rect 39572 9220 39581 9260
rect 20140 9176 20180 9220
rect 25987 9219 26045 9220
rect 835 9136 844 9176
rect 884 9136 20180 9176
rect 3103 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3489 9092
rect 18223 9052 18232 9092
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18600 9052 18609 9092
rect 33343 9052 33352 9092
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33720 9052 33729 9092
rect 48463 9052 48472 9092
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48840 9052 48849 9092
rect 63583 9052 63592 9092
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63960 9052 63969 9092
rect 78703 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 79089 9092
rect 93823 9052 93832 9092
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 94200 9052 94209 9092
rect 0 9008 80 9028
rect 0 8968 652 9008
rect 692 8968 701 9008
rect 0 8948 80 8968
rect 25603 8884 25612 8924
rect 25652 8884 25804 8924
rect 25844 8884 25853 8924
rect 7171 8800 7180 8840
rect 7220 8800 8044 8840
rect 8084 8800 8093 8840
rect 9763 8800 9772 8840
rect 9812 8800 10636 8840
rect 10676 8800 10685 8840
rect 12355 8800 12364 8840
rect 12404 8800 12940 8840
rect 12980 8800 12989 8840
rect 17155 8800 17164 8840
rect 17204 8800 17452 8840
rect 17492 8800 19180 8840
rect 19220 8800 20236 8840
rect 20276 8800 20285 8840
rect 24931 8800 24940 8840
rect 24980 8800 26476 8840
rect 26516 8800 26525 8840
rect 38755 8800 38764 8840
rect 38804 8800 40684 8840
rect 40724 8800 41548 8840
rect 41588 8800 41597 8840
rect 2371 8716 2380 8756
rect 2420 8716 3052 8756
rect 3092 8716 3724 8756
rect 3764 8716 5164 8756
rect 5204 8716 5213 8756
rect 7747 8716 7756 8756
rect 7796 8716 10060 8756
rect 10100 8716 10109 8756
rect 10339 8716 10348 8756
rect 10388 8716 11692 8756
rect 11732 8716 11741 8756
rect 20908 8716 22252 8756
rect 22292 8716 22301 8756
rect 39043 8716 39052 8756
rect 39092 8716 40588 8756
rect 40628 8716 40637 8756
rect 20908 8672 20948 8716
rect 25987 8672 26045 8673
rect 3235 8632 3244 8672
rect 3284 8632 3628 8672
rect 3668 8632 3916 8672
rect 3956 8632 6028 8672
rect 6068 8632 6077 8672
rect 7459 8632 7468 8672
rect 7508 8632 8332 8672
rect 8372 8632 8620 8672
rect 8660 8632 9100 8672
rect 9140 8632 11212 8672
rect 11252 8632 11261 8672
rect 18787 8632 18796 8672
rect 18836 8632 19756 8672
rect 19796 8632 19805 8672
rect 20323 8632 20332 8672
rect 20372 8632 20908 8672
rect 20948 8632 20957 8672
rect 21091 8632 21100 8672
rect 21140 8632 22060 8672
rect 22100 8632 22109 8672
rect 25902 8632 25996 8672
rect 26036 8632 26045 8672
rect 45859 8632 45868 8672
rect 45908 8632 47116 8672
rect 47156 8632 47165 8672
rect 25987 8631 26045 8632
rect 19843 8548 19852 8588
rect 19892 8548 21580 8588
rect 21620 8548 22924 8588
rect 22964 8548 22973 8588
rect 20995 8464 21004 8504
rect 21044 8464 23020 8504
rect 23060 8464 23069 8504
rect 35971 8464 35980 8504
rect 36020 8464 38380 8504
rect 38420 8464 38429 8504
rect 4343 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4729 8336
rect 19463 8296 19472 8336
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19840 8296 19849 8336
rect 34583 8296 34592 8336
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34960 8296 34969 8336
rect 49703 8296 49712 8336
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 50080 8296 50089 8336
rect 64823 8296 64832 8336
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 65200 8296 65209 8336
rect 79943 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 80329 8336
rect 95063 8296 95072 8336
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95440 8296 95449 8336
rect 0 8168 80 8188
rect 0 8128 556 8168
rect 596 8128 605 8168
rect 23203 8128 23212 8168
rect 23252 8128 25708 8168
rect 25748 8128 25757 8168
rect 0 8108 80 8128
rect 27331 8044 27340 8084
rect 27380 8044 28684 8084
rect 28724 8044 28733 8084
rect 38659 8044 38668 8084
rect 38708 8044 39916 8084
rect 39956 8044 39965 8084
rect 22147 7960 22156 8000
rect 22196 7960 23116 8000
rect 23156 7960 23165 8000
rect 29635 7960 29644 8000
rect 29684 7960 30316 8000
rect 30356 7960 30365 8000
rect 37027 7960 37036 8000
rect 37076 7960 37228 8000
rect 37268 7960 50956 8000
rect 50996 7960 51724 8000
rect 51764 7960 51773 8000
rect 18691 7876 18700 7916
rect 18740 7876 19180 7916
rect 19220 7876 19948 7916
rect 19988 7876 19997 7916
rect 35587 7792 35596 7832
rect 35636 7792 38092 7832
rect 38132 7792 38141 7832
rect 31075 7708 31084 7748
rect 31124 7708 32236 7748
rect 32276 7708 32285 7748
rect 3103 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3489 7580
rect 18223 7540 18232 7580
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18600 7540 18609 7580
rect 33343 7540 33352 7580
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33720 7540 33729 7580
rect 48463 7540 48472 7580
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48840 7540 48849 7580
rect 63583 7540 63592 7580
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63960 7540 63969 7580
rect 78703 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 79089 7580
rect 93823 7540 93832 7580
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 94200 7540 94209 7580
rect 0 7328 80 7348
rect 0 7288 652 7328
rect 692 7288 701 7328
rect 20140 7288 22348 7328
rect 22388 7288 23404 7328
rect 23444 7288 26956 7328
rect 26996 7288 27005 7328
rect 0 7268 80 7288
rect 20140 7244 20180 7288
rect 16099 7204 16108 7244
rect 16148 7204 16300 7244
rect 16340 7204 16588 7244
rect 16628 7204 20180 7244
rect 26668 7204 29068 7244
rect 29108 7204 29117 7244
rect 26668 7160 26708 7204
rect 16195 7120 16204 7160
rect 16244 7120 22924 7160
rect 22964 7120 22973 7160
rect 26659 7120 26668 7160
rect 26708 7120 26717 7160
rect 28867 7120 28876 7160
rect 28916 7120 29000 7160
rect 30019 7120 30028 7160
rect 30068 7120 30220 7160
rect 30260 7120 30604 7160
rect 30644 7120 30653 7160
rect 47107 7120 47116 7160
rect 47156 7120 48748 7160
rect 48788 7120 51820 7160
rect 51860 7120 51869 7160
rect 28960 7076 29000 7120
rect 22723 7036 22732 7076
rect 22772 7036 25996 7076
rect 26036 7036 26045 7076
rect 28960 7036 32332 7076
rect 32372 7036 32780 7076
rect 35875 7036 35884 7076
rect 35924 7036 37996 7076
rect 38036 7036 38045 7076
rect 32740 6992 32780 7036
rect 23587 6952 23596 6992
rect 23636 6952 28396 6992
rect 28436 6952 28445 6992
rect 29443 6952 29452 6992
rect 29492 6952 29932 6992
rect 29972 6952 29981 6992
rect 32740 6952 33484 6992
rect 33524 6952 33533 6992
rect 38755 6952 38764 6992
rect 38804 6952 39532 6992
rect 39572 6952 40012 6992
rect 40052 6952 40061 6992
rect 4343 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4729 6824
rect 19463 6784 19472 6824
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19840 6784 19849 6824
rect 34583 6784 34592 6824
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34960 6784 34969 6824
rect 49703 6784 49712 6824
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 50080 6784 50089 6824
rect 64823 6784 64832 6824
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 65200 6784 65209 6824
rect 79943 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 80329 6824
rect 95063 6784 95072 6824
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95440 6784 95449 6824
rect 28579 6616 28588 6656
rect 28628 6616 29452 6656
rect 29492 6616 29644 6656
rect 29684 6616 29693 6656
rect 53731 6616 53740 6656
rect 53780 6616 54988 6656
rect 55028 6616 55037 6656
rect 0 6488 80 6508
rect 0 6448 652 6488
rect 692 6448 701 6488
rect 29827 6448 29836 6488
rect 29876 6448 31660 6488
rect 31700 6448 31709 6488
rect 36547 6448 36556 6488
rect 36596 6448 39340 6488
rect 39380 6448 39389 6488
rect 45187 6448 45196 6488
rect 45236 6448 46252 6488
rect 46292 6448 46444 6488
rect 46484 6448 46493 6488
rect 47395 6448 47404 6488
rect 47444 6448 47980 6488
rect 48020 6448 48029 6488
rect 51139 6448 51148 6488
rect 51188 6448 54028 6488
rect 54068 6448 54077 6488
rect 0 6428 80 6448
rect 38532 6280 38572 6320
rect 38612 6280 38621 6320
rect 38572 6236 38612 6280
rect 18115 6196 18124 6236
rect 18164 6196 18892 6236
rect 18932 6196 21580 6236
rect 21620 6196 21629 6236
rect 37699 6196 37708 6236
rect 37748 6196 38612 6236
rect 3103 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3489 6068
rect 18223 6028 18232 6068
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18600 6028 18609 6068
rect 33343 6028 33352 6068
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33720 6028 33729 6068
rect 48463 6028 48472 6068
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48840 6028 48849 6068
rect 63583 6028 63592 6068
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63960 6028 63969 6068
rect 78703 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 79089 6068
rect 93823 6028 93832 6068
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 94200 6028 94209 6068
rect 48355 5860 48364 5900
rect 48404 5860 49612 5900
rect 49652 5860 49661 5900
rect 0 5648 80 5668
rect 0 5608 652 5648
rect 692 5608 701 5648
rect 33859 5608 33868 5648
rect 33908 5608 36556 5648
rect 36596 5608 36605 5648
rect 43651 5608 43660 5648
rect 43700 5608 44812 5648
rect 44852 5608 45292 5648
rect 45332 5608 45341 5648
rect 46531 5608 46540 5648
rect 46580 5608 47212 5648
rect 47252 5608 47261 5648
rect 48643 5608 48652 5648
rect 48692 5608 51148 5648
rect 51188 5608 51197 5648
rect 56611 5608 56620 5648
rect 56660 5608 57196 5648
rect 57236 5608 57245 5648
rect 0 5588 80 5608
rect 45955 5524 45964 5564
rect 46004 5524 46636 5564
rect 46676 5524 46685 5564
rect 54403 5440 54412 5480
rect 54452 5440 55948 5480
rect 55988 5440 55997 5480
rect 4343 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4729 5312
rect 19463 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 19849 5312
rect 34583 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 34969 5312
rect 49703 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 50089 5312
rect 64823 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 65209 5312
rect 79943 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 80329 5312
rect 95063 5272 95072 5312
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95440 5272 95449 5312
rect 33379 5020 33388 5060
rect 33428 5020 34348 5060
rect 34388 5020 34397 5060
rect 47683 5020 47692 5060
rect 47732 5020 51916 5060
rect 51956 5020 51965 5060
rect 11875 4936 11884 4976
rect 11924 4936 15628 4976
rect 15668 4936 15677 4976
rect 24547 4936 24556 4976
rect 24596 4936 25612 4976
rect 25652 4936 25661 4976
rect 26851 4936 26860 4976
rect 26900 4936 28300 4976
rect 28340 4936 28349 4976
rect 41560 4936 42508 4976
rect 42548 4936 42557 4976
rect 52099 4936 52108 4976
rect 52148 4936 53068 4976
rect 53108 4936 54028 4976
rect 54068 4936 54077 4976
rect 41560 4892 41600 4936
rect 39235 4852 39244 4892
rect 39284 4852 39628 4892
rect 39668 4852 41600 4892
rect 0 4808 80 4828
rect 0 4768 652 4808
rect 692 4768 701 4808
rect 0 4748 80 4768
rect 52963 4600 52972 4640
rect 53012 4600 54796 4640
rect 54836 4600 55180 4640
rect 55220 4600 55229 4640
rect 3103 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3489 4556
rect 18223 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 18609 4556
rect 33343 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 33729 4556
rect 48463 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 48849 4556
rect 63583 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 63969 4556
rect 78703 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 79089 4556
rect 93823 4516 93832 4556
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 94200 4516 94209 4556
rect 23779 4180 23788 4220
rect 23828 4180 24364 4220
rect 24404 4180 24413 4220
rect 34435 4180 34444 4220
rect 34484 4180 38956 4220
rect 38996 4180 40204 4220
rect 40244 4180 40492 4220
rect 40532 4180 40541 4220
rect 11587 4096 11596 4136
rect 11636 4096 11884 4136
rect 11924 4096 11933 4136
rect 20035 4096 20044 4136
rect 20084 4096 20524 4136
rect 20564 4096 20573 4136
rect 27715 4096 27724 4136
rect 27764 4096 29164 4136
rect 29204 4096 34348 4136
rect 34388 4096 34397 4136
rect 40099 4096 40108 4136
rect 40148 4096 41356 4136
rect 41396 4096 41405 4136
rect 0 3968 80 3988
rect 0 3928 652 3968
rect 692 3928 701 3968
rect 33379 3928 33388 3968
rect 33428 3928 34252 3968
rect 34292 3928 34301 3968
rect 41635 3928 41644 3968
rect 41684 3928 44044 3968
rect 44084 3928 44093 3968
rect 0 3908 80 3928
rect 4343 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4729 3800
rect 19463 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 19849 3800
rect 34583 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 34969 3800
rect 37987 3760 37996 3800
rect 38036 3760 39244 3800
rect 39284 3760 40588 3800
rect 40628 3760 40637 3800
rect 45283 3760 45292 3800
rect 45332 3760 46444 3800
rect 46484 3760 48268 3800
rect 48308 3760 48317 3800
rect 49703 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 50089 3800
rect 64823 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 65209 3800
rect 79943 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 80329 3800
rect 95063 3760 95072 3800
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95440 3760 95449 3800
rect 6280 3592 21100 3632
rect 21140 3592 21149 3632
rect 21763 3592 21772 3632
rect 21812 3592 21821 3632
rect 35779 3592 35788 3632
rect 35828 3592 38284 3632
rect 38324 3592 38333 3632
rect 6280 3548 6320 3592
rect 21772 3548 21812 3592
rect 835 3508 844 3548
rect 884 3508 6320 3548
rect 11491 3508 11500 3548
rect 11540 3508 11980 3548
rect 12020 3508 12652 3548
rect 12692 3508 13036 3548
rect 13076 3508 13085 3548
rect 21772 3508 22540 3548
rect 22580 3508 25132 3548
rect 25172 3508 26860 3548
rect 26900 3508 26909 3548
rect 40291 3508 40300 3548
rect 40340 3508 41068 3548
rect 41108 3508 41117 3548
rect 52003 3508 52012 3548
rect 52052 3508 53164 3548
rect 53204 3508 53213 3548
rect 10819 3424 10828 3464
rect 10868 3424 11116 3464
rect 11156 3424 12364 3464
rect 12404 3424 12413 3464
rect 12739 3424 12748 3464
rect 12788 3424 15340 3464
rect 15380 3424 17260 3464
rect 17300 3424 18700 3464
rect 18740 3424 18892 3464
rect 18932 3424 18941 3464
rect 22627 3424 22636 3464
rect 22676 3424 23404 3464
rect 23444 3424 25996 3464
rect 26036 3424 26045 3464
rect 40003 3424 40012 3464
rect 40052 3424 40396 3464
rect 40436 3424 40972 3464
rect 41012 3424 41021 3464
rect 47107 3424 47116 3464
rect 47156 3424 47692 3464
rect 47732 3424 47741 3464
rect 51715 3424 51724 3464
rect 51764 3424 53836 3464
rect 53876 3424 55660 3464
rect 55700 3424 56044 3464
rect 56084 3424 56093 3464
rect 38371 3340 38380 3380
rect 38420 3340 39532 3380
rect 39572 3340 40204 3380
rect 40244 3340 40253 3380
rect 51427 3340 51436 3380
rect 51476 3340 51916 3380
rect 51956 3340 51965 3380
rect 643 3172 652 3212
rect 692 3172 701 3212
rect 0 3128 80 3148
rect 652 3128 692 3172
rect 0 3088 692 3128
rect 0 3068 80 3088
rect 3103 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3489 3044
rect 18223 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 18609 3044
rect 33343 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 33729 3044
rect 48463 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 48849 3044
rect 63583 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 63969 3044
rect 78703 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 79089 3044
rect 93823 3004 93832 3044
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 94200 3004 94209 3044
rect 15148 2836 17836 2876
rect 17876 2836 18028 2876
rect 18068 2836 18077 2876
rect 19843 2836 19852 2876
rect 19892 2836 21100 2876
rect 21140 2836 21149 2876
rect 46435 2836 46444 2876
rect 46484 2836 48076 2876
rect 48116 2836 48125 2876
rect 15148 2792 15188 2836
rect 7459 2752 7468 2792
rect 7508 2752 7660 2792
rect 7700 2752 10732 2792
rect 10772 2752 14476 2792
rect 14516 2752 15148 2792
rect 15188 2752 15197 2792
rect 16492 2752 17932 2792
rect 17972 2752 17981 2792
rect 52099 2752 52108 2792
rect 52148 2752 54740 2792
rect 16492 2708 16532 2752
rect 54700 2708 54740 2752
rect 835 2668 844 2708
rect 884 2668 16532 2708
rect 17635 2668 17644 2708
rect 17684 2668 17693 2708
rect 33763 2668 33772 2708
rect 33812 2668 35500 2708
rect 35540 2668 37132 2708
rect 37172 2668 39764 2708
rect 49507 2668 49516 2708
rect 49556 2668 53452 2708
rect 53492 2668 53501 2708
rect 54691 2668 54700 2708
rect 54740 2668 55852 2708
rect 55892 2668 55901 2708
rect 11011 2584 11020 2624
rect 11060 2584 11692 2624
rect 11732 2584 11741 2624
rect 12835 2584 12844 2624
rect 12884 2584 14092 2624
rect 14132 2584 14141 2624
rect 17644 2540 17684 2668
rect 39724 2624 39764 2668
rect 36739 2584 36748 2624
rect 36788 2584 38188 2624
rect 38228 2584 38237 2624
rect 39715 2584 39724 2624
rect 39764 2584 39773 2624
rect 44419 2584 44428 2624
rect 44468 2584 47308 2624
rect 47348 2584 49132 2624
rect 49172 2584 50860 2624
rect 50900 2584 50909 2624
rect 8419 2500 8428 2540
rect 8468 2500 10540 2540
rect 10580 2500 10924 2540
rect 10964 2500 10973 2540
rect 12163 2500 12172 2540
rect 12212 2500 17684 2540
rect 7075 2416 7084 2456
rect 7124 2416 7852 2456
rect 7892 2416 7901 2456
rect 0 2288 80 2308
rect 0 2248 652 2288
rect 692 2248 701 2288
rect 4343 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4729 2288
rect 19463 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 19849 2288
rect 34583 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 34969 2288
rect 49703 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 50089 2288
rect 64823 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 65209 2288
rect 79943 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 80329 2288
rect 95063 2248 95072 2288
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95440 2248 95449 2288
rect 0 2228 80 2248
rect 7267 2080 7276 2120
rect 7316 2080 8236 2120
rect 8276 2080 8285 2120
rect 8899 2080 8908 2120
rect 8948 2080 11308 2120
rect 11348 2080 11357 2120
rect 8908 2036 8948 2080
rect 8035 1996 8044 2036
rect 8084 1996 8948 2036
rect 3103 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3489 1532
rect 18223 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 18609 1532
rect 33343 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 33729 1532
rect 48463 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 48849 1532
rect 63583 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 63969 1532
rect 78703 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 79089 1532
rect 93823 1492 93832 1532
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 94200 1492 94209 1532
rect 4343 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4729 776
rect 19463 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 19849 776
rect 34583 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 34969 776
rect 49703 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 50089 776
rect 64823 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 65209 776
rect 79943 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 80329 776
rect 95063 736 95072 776
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95440 736 95449 776
<< via3 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 25996 9388 26036 9428
rect 25996 9220 26036 9260
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 25996 8632 26036 8672
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal4 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 95072 38576 95440 38585
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95072 38527 95440 38536
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 93832 37820 94200 37829
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 93832 37771 94200 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 95072 37064 95440 37073
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95072 37015 95440 37024
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 93832 36308 94200 36317
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 93832 36259 94200 36268
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 95072 35552 95440 35561
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95072 35503 95440 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 93832 34796 94200 34805
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 93832 34747 94200 34756
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 95072 34040 95440 34049
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95072 33991 95440 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 18232 33284 18600 33293
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18232 33235 18600 33244
rect 33352 33284 33720 33293
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33352 33235 33720 33244
rect 48472 33284 48840 33293
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48472 33235 48840 33244
rect 63592 33284 63960 33293
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63592 33235 63960 33244
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 93832 33284 94200 33293
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 93832 33235 94200 33244
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 19472 32528 19840 32537
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19472 32479 19840 32488
rect 34592 32528 34960 32537
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34592 32479 34960 32488
rect 49712 32528 50080 32537
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 49712 32479 50080 32488
rect 64832 32528 65200 32537
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 64832 32479 65200 32488
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 95072 32528 95440 32537
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95072 32479 95440 32488
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 18232 31772 18600 31781
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18232 31723 18600 31732
rect 33352 31772 33720 31781
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33352 31723 33720 31732
rect 48472 31772 48840 31781
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48472 31723 48840 31732
rect 63592 31772 63960 31781
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63592 31723 63960 31732
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 93832 31772 94200 31781
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 93832 31723 94200 31732
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 19472 31016 19840 31025
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19472 30967 19840 30976
rect 34592 31016 34960 31025
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34592 30967 34960 30976
rect 49712 31016 50080 31025
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 49712 30967 50080 30976
rect 64832 31016 65200 31025
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 64832 30967 65200 30976
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 95072 31016 95440 31025
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95072 30967 95440 30976
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 18232 30260 18600 30269
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18232 30211 18600 30220
rect 33352 30260 33720 30269
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33352 30211 33720 30220
rect 48472 30260 48840 30269
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48472 30211 48840 30220
rect 63592 30260 63960 30269
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63592 30211 63960 30220
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 93832 30260 94200 30269
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 93832 30211 94200 30220
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 19472 29504 19840 29513
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19472 29455 19840 29464
rect 34592 29504 34960 29513
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34592 29455 34960 29464
rect 49712 29504 50080 29513
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 49712 29455 50080 29464
rect 64832 29504 65200 29513
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 64832 29455 65200 29464
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 95072 29504 95440 29513
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95072 29455 95440 29464
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 18232 28748 18600 28757
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18232 28699 18600 28708
rect 33352 28748 33720 28757
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33352 28699 33720 28708
rect 48472 28748 48840 28757
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48472 28699 48840 28708
rect 63592 28748 63960 28757
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63592 28699 63960 28708
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 93832 28748 94200 28757
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 93832 28699 94200 28708
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 19472 27992 19840 28001
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19472 27943 19840 27952
rect 34592 27992 34960 28001
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34592 27943 34960 27952
rect 49712 27992 50080 28001
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 49712 27943 50080 27952
rect 64832 27992 65200 28001
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 64832 27943 65200 27952
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 95072 27992 95440 28001
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95072 27943 95440 27952
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 18232 27236 18600 27245
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18232 27187 18600 27196
rect 33352 27236 33720 27245
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33352 27187 33720 27196
rect 48472 27236 48840 27245
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48472 27187 48840 27196
rect 63592 27236 63960 27245
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63592 27187 63960 27196
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 93832 27236 94200 27245
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 93832 27187 94200 27196
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 19472 26480 19840 26489
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19472 26431 19840 26440
rect 34592 26480 34960 26489
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34592 26431 34960 26440
rect 49712 26480 50080 26489
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 49712 26431 50080 26440
rect 64832 26480 65200 26489
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 64832 26431 65200 26440
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 95072 26480 95440 26489
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95072 26431 95440 26440
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 18232 25724 18600 25733
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18232 25675 18600 25684
rect 33352 25724 33720 25733
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33352 25675 33720 25684
rect 48472 25724 48840 25733
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48472 25675 48840 25684
rect 63592 25724 63960 25733
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63592 25675 63960 25684
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 93832 25724 94200 25733
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 93832 25675 94200 25684
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 19472 24968 19840 24977
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19472 24919 19840 24928
rect 34592 24968 34960 24977
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34592 24919 34960 24928
rect 49712 24968 50080 24977
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 49712 24919 50080 24928
rect 64832 24968 65200 24977
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 64832 24919 65200 24928
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 95072 24968 95440 24977
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95072 24919 95440 24928
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 18232 24212 18600 24221
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18232 24163 18600 24172
rect 33352 24212 33720 24221
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33352 24163 33720 24172
rect 48472 24212 48840 24221
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48472 24163 48840 24172
rect 63592 24212 63960 24221
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63592 24163 63960 24172
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 93832 24212 94200 24221
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 93832 24163 94200 24172
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 19472 23456 19840 23465
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19472 23407 19840 23416
rect 34592 23456 34960 23465
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34592 23407 34960 23416
rect 49712 23456 50080 23465
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 49712 23407 50080 23416
rect 64832 23456 65200 23465
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 64832 23407 65200 23416
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 95072 23456 95440 23465
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95072 23407 95440 23416
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 18232 22700 18600 22709
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18232 22651 18600 22660
rect 33352 22700 33720 22709
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33352 22651 33720 22660
rect 48472 22700 48840 22709
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48472 22651 48840 22660
rect 63592 22700 63960 22709
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63592 22651 63960 22660
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 93832 22700 94200 22709
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 93832 22651 94200 22660
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 19472 21944 19840 21953
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19472 21895 19840 21904
rect 34592 21944 34960 21953
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34592 21895 34960 21904
rect 49712 21944 50080 21953
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 49712 21895 50080 21904
rect 64832 21944 65200 21953
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 64832 21895 65200 21904
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 95072 21944 95440 21953
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95072 21895 95440 21904
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 18232 21188 18600 21197
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18232 21139 18600 21148
rect 33352 21188 33720 21197
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33352 21139 33720 21148
rect 48472 21188 48840 21197
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48472 21139 48840 21148
rect 63592 21188 63960 21197
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63592 21139 63960 21148
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 93832 21188 94200 21197
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 93832 21139 94200 21148
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 19472 20432 19840 20441
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19472 20383 19840 20392
rect 34592 20432 34960 20441
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34592 20383 34960 20392
rect 49712 20432 50080 20441
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 49712 20383 50080 20392
rect 64832 20432 65200 20441
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 64832 20383 65200 20392
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 95072 20432 95440 20441
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95072 20383 95440 20392
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 18232 19676 18600 19685
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18232 19627 18600 19636
rect 33352 19676 33720 19685
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33352 19627 33720 19636
rect 48472 19676 48840 19685
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48472 19627 48840 19636
rect 63592 19676 63960 19685
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63592 19627 63960 19636
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 93832 19676 94200 19685
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 93832 19627 94200 19636
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 19472 18920 19840 18929
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19472 18871 19840 18880
rect 34592 18920 34960 18929
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34592 18871 34960 18880
rect 49712 18920 50080 18929
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 49712 18871 50080 18880
rect 64832 18920 65200 18929
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 64832 18871 65200 18880
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 95072 18920 95440 18929
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95072 18871 95440 18880
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 18232 18164 18600 18173
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18232 18115 18600 18124
rect 33352 18164 33720 18173
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33352 18115 33720 18124
rect 48472 18164 48840 18173
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48472 18115 48840 18124
rect 63592 18164 63960 18173
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63592 18115 63960 18124
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 93832 18164 94200 18173
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 93832 18115 94200 18124
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 19472 17408 19840 17417
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19472 17359 19840 17368
rect 34592 17408 34960 17417
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34592 17359 34960 17368
rect 49712 17408 50080 17417
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 49712 17359 50080 17368
rect 64832 17408 65200 17417
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 64832 17359 65200 17368
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 95072 17408 95440 17417
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95072 17359 95440 17368
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 18232 16652 18600 16661
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18232 16603 18600 16612
rect 33352 16652 33720 16661
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33352 16603 33720 16612
rect 48472 16652 48840 16661
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48472 16603 48840 16612
rect 63592 16652 63960 16661
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63592 16603 63960 16612
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 93832 16652 94200 16661
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 93832 16603 94200 16612
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 19472 15896 19840 15905
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19472 15847 19840 15856
rect 34592 15896 34960 15905
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34592 15847 34960 15856
rect 49712 15896 50080 15905
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 49712 15847 50080 15856
rect 64832 15896 65200 15905
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 64832 15847 65200 15856
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 95072 15896 95440 15905
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95072 15847 95440 15856
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 18232 15140 18600 15149
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18232 15091 18600 15100
rect 33352 15140 33720 15149
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33352 15091 33720 15100
rect 48472 15140 48840 15149
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48472 15091 48840 15100
rect 63592 15140 63960 15149
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63592 15091 63960 15100
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 93832 15140 94200 15149
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 93832 15091 94200 15100
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 19472 14384 19840 14393
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19472 14335 19840 14344
rect 34592 14384 34960 14393
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34592 14335 34960 14344
rect 49712 14384 50080 14393
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 49712 14335 50080 14344
rect 64832 14384 65200 14393
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 64832 14335 65200 14344
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 95072 14384 95440 14393
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95072 14335 95440 14344
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 18232 13628 18600 13637
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18232 13579 18600 13588
rect 33352 13628 33720 13637
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33352 13579 33720 13588
rect 48472 13628 48840 13637
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48472 13579 48840 13588
rect 63592 13628 63960 13637
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63592 13579 63960 13588
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 93832 13628 94200 13637
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 93832 13579 94200 13588
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 19472 12872 19840 12881
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19472 12823 19840 12832
rect 34592 12872 34960 12881
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34592 12823 34960 12832
rect 49712 12872 50080 12881
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 49712 12823 50080 12832
rect 64832 12872 65200 12881
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 64832 12823 65200 12832
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 95072 12872 95440 12881
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95072 12823 95440 12832
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 18232 12116 18600 12125
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18232 12067 18600 12076
rect 33352 12116 33720 12125
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33352 12067 33720 12076
rect 48472 12116 48840 12125
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48472 12067 48840 12076
rect 63592 12116 63960 12125
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63592 12067 63960 12076
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 93832 12116 94200 12125
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 93832 12067 94200 12076
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 19472 11360 19840 11369
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19472 11311 19840 11320
rect 34592 11360 34960 11369
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34592 11311 34960 11320
rect 49712 11360 50080 11369
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 49712 11311 50080 11320
rect 64832 11360 65200 11369
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 64832 11311 65200 11320
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 95072 11360 95440 11369
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95072 11311 95440 11320
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 18232 10604 18600 10613
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18232 10555 18600 10564
rect 33352 10604 33720 10613
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33352 10555 33720 10564
rect 48472 10604 48840 10613
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48472 10555 48840 10564
rect 63592 10604 63960 10613
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63592 10555 63960 10564
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 93832 10604 94200 10613
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 93832 10555 94200 10564
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 19472 9848 19840 9857
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19472 9799 19840 9808
rect 34592 9848 34960 9857
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34592 9799 34960 9808
rect 49712 9848 50080 9857
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 49712 9799 50080 9808
rect 64832 9848 65200 9857
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 64832 9799 65200 9808
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 95072 9848 95440 9857
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95072 9799 95440 9808
rect 25996 9428 26036 9437
rect 25996 9260 26036 9388
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 18232 9092 18600 9101
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18232 9043 18600 9052
rect 25996 8672 26036 9220
rect 33352 9092 33720 9101
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33352 9043 33720 9052
rect 48472 9092 48840 9101
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48472 9043 48840 9052
rect 63592 9092 63960 9101
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63592 9043 63960 9052
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 93832 9092 94200 9101
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 93832 9043 94200 9052
rect 25996 8623 26036 8632
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 19472 8336 19840 8345
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19472 8287 19840 8296
rect 34592 8336 34960 8345
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34592 8287 34960 8296
rect 49712 8336 50080 8345
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 49712 8287 50080 8296
rect 64832 8336 65200 8345
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 64832 8287 65200 8296
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 95072 8336 95440 8345
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95072 8287 95440 8296
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 18232 7580 18600 7589
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18232 7531 18600 7540
rect 33352 7580 33720 7589
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33352 7531 33720 7540
rect 48472 7580 48840 7589
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48472 7531 48840 7540
rect 63592 7580 63960 7589
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63592 7531 63960 7540
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 93832 7580 94200 7589
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 93832 7531 94200 7540
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 19472 6824 19840 6833
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19472 6775 19840 6784
rect 34592 6824 34960 6833
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34592 6775 34960 6784
rect 49712 6824 50080 6833
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 49712 6775 50080 6784
rect 64832 6824 65200 6833
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 64832 6775 65200 6784
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 95072 6824 95440 6833
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95072 6775 95440 6784
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 18232 6068 18600 6077
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18232 6019 18600 6028
rect 33352 6068 33720 6077
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33352 6019 33720 6028
rect 48472 6068 48840 6077
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48472 6019 48840 6028
rect 63592 6068 63960 6077
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63592 6019 63960 6028
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 93832 6068 94200 6077
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 93832 6019 94200 6028
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 95072 5312 95440 5321
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95072 5263 95440 5272
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 93832 4556 94200 4565
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 93832 4507 94200 4516
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 95072 3800 95440 3809
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95072 3751 95440 3760
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 93832 3044 94200 3053
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 93832 2995 94200 3004
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 95072 2288 95440 2297
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95072 2239 95440 2248
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 93832 1532 94200 1541
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 93832 1483 94200 1492
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
rect 95072 776 95440 785
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95072 727 95440 736
<< via4 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal5 >>
rect 4343 38599 4729 38618
rect 4343 38576 4409 38599
rect 4495 38576 4577 38599
rect 4663 38576 4729 38599
rect 4343 38536 4352 38576
rect 4392 38536 4409 38576
rect 4495 38536 4516 38576
rect 4556 38536 4577 38576
rect 4663 38536 4680 38576
rect 4720 38536 4729 38576
rect 4343 38513 4409 38536
rect 4495 38513 4577 38536
rect 4663 38513 4729 38536
rect 4343 38494 4729 38513
rect 19463 38599 19849 38618
rect 19463 38576 19529 38599
rect 19615 38576 19697 38599
rect 19783 38576 19849 38599
rect 19463 38536 19472 38576
rect 19512 38536 19529 38576
rect 19615 38536 19636 38576
rect 19676 38536 19697 38576
rect 19783 38536 19800 38576
rect 19840 38536 19849 38576
rect 19463 38513 19529 38536
rect 19615 38513 19697 38536
rect 19783 38513 19849 38536
rect 19463 38494 19849 38513
rect 34583 38599 34969 38618
rect 34583 38576 34649 38599
rect 34735 38576 34817 38599
rect 34903 38576 34969 38599
rect 34583 38536 34592 38576
rect 34632 38536 34649 38576
rect 34735 38536 34756 38576
rect 34796 38536 34817 38576
rect 34903 38536 34920 38576
rect 34960 38536 34969 38576
rect 34583 38513 34649 38536
rect 34735 38513 34817 38536
rect 34903 38513 34969 38536
rect 34583 38494 34969 38513
rect 49703 38599 50089 38618
rect 49703 38576 49769 38599
rect 49855 38576 49937 38599
rect 50023 38576 50089 38599
rect 49703 38536 49712 38576
rect 49752 38536 49769 38576
rect 49855 38536 49876 38576
rect 49916 38536 49937 38576
rect 50023 38536 50040 38576
rect 50080 38536 50089 38576
rect 49703 38513 49769 38536
rect 49855 38513 49937 38536
rect 50023 38513 50089 38536
rect 49703 38494 50089 38513
rect 64823 38599 65209 38618
rect 64823 38576 64889 38599
rect 64975 38576 65057 38599
rect 65143 38576 65209 38599
rect 64823 38536 64832 38576
rect 64872 38536 64889 38576
rect 64975 38536 64996 38576
rect 65036 38536 65057 38576
rect 65143 38536 65160 38576
rect 65200 38536 65209 38576
rect 64823 38513 64889 38536
rect 64975 38513 65057 38536
rect 65143 38513 65209 38536
rect 64823 38494 65209 38513
rect 79943 38599 80329 38618
rect 79943 38576 80009 38599
rect 80095 38576 80177 38599
rect 80263 38576 80329 38599
rect 79943 38536 79952 38576
rect 79992 38536 80009 38576
rect 80095 38536 80116 38576
rect 80156 38536 80177 38576
rect 80263 38536 80280 38576
rect 80320 38536 80329 38576
rect 79943 38513 80009 38536
rect 80095 38513 80177 38536
rect 80263 38513 80329 38536
rect 79943 38494 80329 38513
rect 95063 38599 95449 38618
rect 95063 38576 95129 38599
rect 95215 38576 95297 38599
rect 95383 38576 95449 38599
rect 95063 38536 95072 38576
rect 95112 38536 95129 38576
rect 95215 38536 95236 38576
rect 95276 38536 95297 38576
rect 95383 38536 95400 38576
rect 95440 38536 95449 38576
rect 95063 38513 95129 38536
rect 95215 38513 95297 38536
rect 95383 38513 95449 38536
rect 95063 38494 95449 38513
rect 3103 37843 3489 37862
rect 3103 37820 3169 37843
rect 3255 37820 3337 37843
rect 3423 37820 3489 37843
rect 3103 37780 3112 37820
rect 3152 37780 3169 37820
rect 3255 37780 3276 37820
rect 3316 37780 3337 37820
rect 3423 37780 3440 37820
rect 3480 37780 3489 37820
rect 3103 37757 3169 37780
rect 3255 37757 3337 37780
rect 3423 37757 3489 37780
rect 3103 37738 3489 37757
rect 18223 37843 18609 37862
rect 18223 37820 18289 37843
rect 18375 37820 18457 37843
rect 18543 37820 18609 37843
rect 18223 37780 18232 37820
rect 18272 37780 18289 37820
rect 18375 37780 18396 37820
rect 18436 37780 18457 37820
rect 18543 37780 18560 37820
rect 18600 37780 18609 37820
rect 18223 37757 18289 37780
rect 18375 37757 18457 37780
rect 18543 37757 18609 37780
rect 18223 37738 18609 37757
rect 33343 37843 33729 37862
rect 33343 37820 33409 37843
rect 33495 37820 33577 37843
rect 33663 37820 33729 37843
rect 33343 37780 33352 37820
rect 33392 37780 33409 37820
rect 33495 37780 33516 37820
rect 33556 37780 33577 37820
rect 33663 37780 33680 37820
rect 33720 37780 33729 37820
rect 33343 37757 33409 37780
rect 33495 37757 33577 37780
rect 33663 37757 33729 37780
rect 33343 37738 33729 37757
rect 48463 37843 48849 37862
rect 48463 37820 48529 37843
rect 48615 37820 48697 37843
rect 48783 37820 48849 37843
rect 48463 37780 48472 37820
rect 48512 37780 48529 37820
rect 48615 37780 48636 37820
rect 48676 37780 48697 37820
rect 48783 37780 48800 37820
rect 48840 37780 48849 37820
rect 48463 37757 48529 37780
rect 48615 37757 48697 37780
rect 48783 37757 48849 37780
rect 48463 37738 48849 37757
rect 63583 37843 63969 37862
rect 63583 37820 63649 37843
rect 63735 37820 63817 37843
rect 63903 37820 63969 37843
rect 63583 37780 63592 37820
rect 63632 37780 63649 37820
rect 63735 37780 63756 37820
rect 63796 37780 63817 37820
rect 63903 37780 63920 37820
rect 63960 37780 63969 37820
rect 63583 37757 63649 37780
rect 63735 37757 63817 37780
rect 63903 37757 63969 37780
rect 63583 37738 63969 37757
rect 78703 37843 79089 37862
rect 78703 37820 78769 37843
rect 78855 37820 78937 37843
rect 79023 37820 79089 37843
rect 78703 37780 78712 37820
rect 78752 37780 78769 37820
rect 78855 37780 78876 37820
rect 78916 37780 78937 37820
rect 79023 37780 79040 37820
rect 79080 37780 79089 37820
rect 78703 37757 78769 37780
rect 78855 37757 78937 37780
rect 79023 37757 79089 37780
rect 78703 37738 79089 37757
rect 93823 37843 94209 37862
rect 93823 37820 93889 37843
rect 93975 37820 94057 37843
rect 94143 37820 94209 37843
rect 93823 37780 93832 37820
rect 93872 37780 93889 37820
rect 93975 37780 93996 37820
rect 94036 37780 94057 37820
rect 94143 37780 94160 37820
rect 94200 37780 94209 37820
rect 93823 37757 93889 37780
rect 93975 37757 94057 37780
rect 94143 37757 94209 37780
rect 93823 37738 94209 37757
rect 4343 37087 4729 37106
rect 4343 37064 4409 37087
rect 4495 37064 4577 37087
rect 4663 37064 4729 37087
rect 4343 37024 4352 37064
rect 4392 37024 4409 37064
rect 4495 37024 4516 37064
rect 4556 37024 4577 37064
rect 4663 37024 4680 37064
rect 4720 37024 4729 37064
rect 4343 37001 4409 37024
rect 4495 37001 4577 37024
rect 4663 37001 4729 37024
rect 4343 36982 4729 37001
rect 19463 37087 19849 37106
rect 19463 37064 19529 37087
rect 19615 37064 19697 37087
rect 19783 37064 19849 37087
rect 19463 37024 19472 37064
rect 19512 37024 19529 37064
rect 19615 37024 19636 37064
rect 19676 37024 19697 37064
rect 19783 37024 19800 37064
rect 19840 37024 19849 37064
rect 19463 37001 19529 37024
rect 19615 37001 19697 37024
rect 19783 37001 19849 37024
rect 19463 36982 19849 37001
rect 34583 37087 34969 37106
rect 34583 37064 34649 37087
rect 34735 37064 34817 37087
rect 34903 37064 34969 37087
rect 34583 37024 34592 37064
rect 34632 37024 34649 37064
rect 34735 37024 34756 37064
rect 34796 37024 34817 37064
rect 34903 37024 34920 37064
rect 34960 37024 34969 37064
rect 34583 37001 34649 37024
rect 34735 37001 34817 37024
rect 34903 37001 34969 37024
rect 34583 36982 34969 37001
rect 49703 37087 50089 37106
rect 49703 37064 49769 37087
rect 49855 37064 49937 37087
rect 50023 37064 50089 37087
rect 49703 37024 49712 37064
rect 49752 37024 49769 37064
rect 49855 37024 49876 37064
rect 49916 37024 49937 37064
rect 50023 37024 50040 37064
rect 50080 37024 50089 37064
rect 49703 37001 49769 37024
rect 49855 37001 49937 37024
rect 50023 37001 50089 37024
rect 49703 36982 50089 37001
rect 64823 37087 65209 37106
rect 64823 37064 64889 37087
rect 64975 37064 65057 37087
rect 65143 37064 65209 37087
rect 64823 37024 64832 37064
rect 64872 37024 64889 37064
rect 64975 37024 64996 37064
rect 65036 37024 65057 37064
rect 65143 37024 65160 37064
rect 65200 37024 65209 37064
rect 64823 37001 64889 37024
rect 64975 37001 65057 37024
rect 65143 37001 65209 37024
rect 64823 36982 65209 37001
rect 79943 37087 80329 37106
rect 79943 37064 80009 37087
rect 80095 37064 80177 37087
rect 80263 37064 80329 37087
rect 79943 37024 79952 37064
rect 79992 37024 80009 37064
rect 80095 37024 80116 37064
rect 80156 37024 80177 37064
rect 80263 37024 80280 37064
rect 80320 37024 80329 37064
rect 79943 37001 80009 37024
rect 80095 37001 80177 37024
rect 80263 37001 80329 37024
rect 79943 36982 80329 37001
rect 95063 37087 95449 37106
rect 95063 37064 95129 37087
rect 95215 37064 95297 37087
rect 95383 37064 95449 37087
rect 95063 37024 95072 37064
rect 95112 37024 95129 37064
rect 95215 37024 95236 37064
rect 95276 37024 95297 37064
rect 95383 37024 95400 37064
rect 95440 37024 95449 37064
rect 95063 37001 95129 37024
rect 95215 37001 95297 37024
rect 95383 37001 95449 37024
rect 95063 36982 95449 37001
rect 3103 36331 3489 36350
rect 3103 36308 3169 36331
rect 3255 36308 3337 36331
rect 3423 36308 3489 36331
rect 3103 36268 3112 36308
rect 3152 36268 3169 36308
rect 3255 36268 3276 36308
rect 3316 36268 3337 36308
rect 3423 36268 3440 36308
rect 3480 36268 3489 36308
rect 3103 36245 3169 36268
rect 3255 36245 3337 36268
rect 3423 36245 3489 36268
rect 3103 36226 3489 36245
rect 18223 36331 18609 36350
rect 18223 36308 18289 36331
rect 18375 36308 18457 36331
rect 18543 36308 18609 36331
rect 18223 36268 18232 36308
rect 18272 36268 18289 36308
rect 18375 36268 18396 36308
rect 18436 36268 18457 36308
rect 18543 36268 18560 36308
rect 18600 36268 18609 36308
rect 18223 36245 18289 36268
rect 18375 36245 18457 36268
rect 18543 36245 18609 36268
rect 18223 36226 18609 36245
rect 33343 36331 33729 36350
rect 33343 36308 33409 36331
rect 33495 36308 33577 36331
rect 33663 36308 33729 36331
rect 33343 36268 33352 36308
rect 33392 36268 33409 36308
rect 33495 36268 33516 36308
rect 33556 36268 33577 36308
rect 33663 36268 33680 36308
rect 33720 36268 33729 36308
rect 33343 36245 33409 36268
rect 33495 36245 33577 36268
rect 33663 36245 33729 36268
rect 33343 36226 33729 36245
rect 48463 36331 48849 36350
rect 48463 36308 48529 36331
rect 48615 36308 48697 36331
rect 48783 36308 48849 36331
rect 48463 36268 48472 36308
rect 48512 36268 48529 36308
rect 48615 36268 48636 36308
rect 48676 36268 48697 36308
rect 48783 36268 48800 36308
rect 48840 36268 48849 36308
rect 48463 36245 48529 36268
rect 48615 36245 48697 36268
rect 48783 36245 48849 36268
rect 48463 36226 48849 36245
rect 63583 36331 63969 36350
rect 63583 36308 63649 36331
rect 63735 36308 63817 36331
rect 63903 36308 63969 36331
rect 63583 36268 63592 36308
rect 63632 36268 63649 36308
rect 63735 36268 63756 36308
rect 63796 36268 63817 36308
rect 63903 36268 63920 36308
rect 63960 36268 63969 36308
rect 63583 36245 63649 36268
rect 63735 36245 63817 36268
rect 63903 36245 63969 36268
rect 63583 36226 63969 36245
rect 78703 36331 79089 36350
rect 78703 36308 78769 36331
rect 78855 36308 78937 36331
rect 79023 36308 79089 36331
rect 78703 36268 78712 36308
rect 78752 36268 78769 36308
rect 78855 36268 78876 36308
rect 78916 36268 78937 36308
rect 79023 36268 79040 36308
rect 79080 36268 79089 36308
rect 78703 36245 78769 36268
rect 78855 36245 78937 36268
rect 79023 36245 79089 36268
rect 78703 36226 79089 36245
rect 93823 36331 94209 36350
rect 93823 36308 93889 36331
rect 93975 36308 94057 36331
rect 94143 36308 94209 36331
rect 93823 36268 93832 36308
rect 93872 36268 93889 36308
rect 93975 36268 93996 36308
rect 94036 36268 94057 36308
rect 94143 36268 94160 36308
rect 94200 36268 94209 36308
rect 93823 36245 93889 36268
rect 93975 36245 94057 36268
rect 94143 36245 94209 36268
rect 93823 36226 94209 36245
rect 4343 35575 4729 35594
rect 4343 35552 4409 35575
rect 4495 35552 4577 35575
rect 4663 35552 4729 35575
rect 4343 35512 4352 35552
rect 4392 35512 4409 35552
rect 4495 35512 4516 35552
rect 4556 35512 4577 35552
rect 4663 35512 4680 35552
rect 4720 35512 4729 35552
rect 4343 35489 4409 35512
rect 4495 35489 4577 35512
rect 4663 35489 4729 35512
rect 4343 35470 4729 35489
rect 19463 35575 19849 35594
rect 19463 35552 19529 35575
rect 19615 35552 19697 35575
rect 19783 35552 19849 35575
rect 19463 35512 19472 35552
rect 19512 35512 19529 35552
rect 19615 35512 19636 35552
rect 19676 35512 19697 35552
rect 19783 35512 19800 35552
rect 19840 35512 19849 35552
rect 19463 35489 19529 35512
rect 19615 35489 19697 35512
rect 19783 35489 19849 35512
rect 19463 35470 19849 35489
rect 34583 35575 34969 35594
rect 34583 35552 34649 35575
rect 34735 35552 34817 35575
rect 34903 35552 34969 35575
rect 34583 35512 34592 35552
rect 34632 35512 34649 35552
rect 34735 35512 34756 35552
rect 34796 35512 34817 35552
rect 34903 35512 34920 35552
rect 34960 35512 34969 35552
rect 34583 35489 34649 35512
rect 34735 35489 34817 35512
rect 34903 35489 34969 35512
rect 34583 35470 34969 35489
rect 49703 35575 50089 35594
rect 49703 35552 49769 35575
rect 49855 35552 49937 35575
rect 50023 35552 50089 35575
rect 49703 35512 49712 35552
rect 49752 35512 49769 35552
rect 49855 35512 49876 35552
rect 49916 35512 49937 35552
rect 50023 35512 50040 35552
rect 50080 35512 50089 35552
rect 49703 35489 49769 35512
rect 49855 35489 49937 35512
rect 50023 35489 50089 35512
rect 49703 35470 50089 35489
rect 64823 35575 65209 35594
rect 64823 35552 64889 35575
rect 64975 35552 65057 35575
rect 65143 35552 65209 35575
rect 64823 35512 64832 35552
rect 64872 35512 64889 35552
rect 64975 35512 64996 35552
rect 65036 35512 65057 35552
rect 65143 35512 65160 35552
rect 65200 35512 65209 35552
rect 64823 35489 64889 35512
rect 64975 35489 65057 35512
rect 65143 35489 65209 35512
rect 64823 35470 65209 35489
rect 79943 35575 80329 35594
rect 79943 35552 80009 35575
rect 80095 35552 80177 35575
rect 80263 35552 80329 35575
rect 79943 35512 79952 35552
rect 79992 35512 80009 35552
rect 80095 35512 80116 35552
rect 80156 35512 80177 35552
rect 80263 35512 80280 35552
rect 80320 35512 80329 35552
rect 79943 35489 80009 35512
rect 80095 35489 80177 35512
rect 80263 35489 80329 35512
rect 79943 35470 80329 35489
rect 95063 35575 95449 35594
rect 95063 35552 95129 35575
rect 95215 35552 95297 35575
rect 95383 35552 95449 35575
rect 95063 35512 95072 35552
rect 95112 35512 95129 35552
rect 95215 35512 95236 35552
rect 95276 35512 95297 35552
rect 95383 35512 95400 35552
rect 95440 35512 95449 35552
rect 95063 35489 95129 35512
rect 95215 35489 95297 35512
rect 95383 35489 95449 35512
rect 95063 35470 95449 35489
rect 3103 34819 3489 34838
rect 3103 34796 3169 34819
rect 3255 34796 3337 34819
rect 3423 34796 3489 34819
rect 3103 34756 3112 34796
rect 3152 34756 3169 34796
rect 3255 34756 3276 34796
rect 3316 34756 3337 34796
rect 3423 34756 3440 34796
rect 3480 34756 3489 34796
rect 3103 34733 3169 34756
rect 3255 34733 3337 34756
rect 3423 34733 3489 34756
rect 3103 34714 3489 34733
rect 18223 34819 18609 34838
rect 18223 34796 18289 34819
rect 18375 34796 18457 34819
rect 18543 34796 18609 34819
rect 18223 34756 18232 34796
rect 18272 34756 18289 34796
rect 18375 34756 18396 34796
rect 18436 34756 18457 34796
rect 18543 34756 18560 34796
rect 18600 34756 18609 34796
rect 18223 34733 18289 34756
rect 18375 34733 18457 34756
rect 18543 34733 18609 34756
rect 18223 34714 18609 34733
rect 33343 34819 33729 34838
rect 33343 34796 33409 34819
rect 33495 34796 33577 34819
rect 33663 34796 33729 34819
rect 33343 34756 33352 34796
rect 33392 34756 33409 34796
rect 33495 34756 33516 34796
rect 33556 34756 33577 34796
rect 33663 34756 33680 34796
rect 33720 34756 33729 34796
rect 33343 34733 33409 34756
rect 33495 34733 33577 34756
rect 33663 34733 33729 34756
rect 33343 34714 33729 34733
rect 48463 34819 48849 34838
rect 48463 34796 48529 34819
rect 48615 34796 48697 34819
rect 48783 34796 48849 34819
rect 48463 34756 48472 34796
rect 48512 34756 48529 34796
rect 48615 34756 48636 34796
rect 48676 34756 48697 34796
rect 48783 34756 48800 34796
rect 48840 34756 48849 34796
rect 48463 34733 48529 34756
rect 48615 34733 48697 34756
rect 48783 34733 48849 34756
rect 48463 34714 48849 34733
rect 63583 34819 63969 34838
rect 63583 34796 63649 34819
rect 63735 34796 63817 34819
rect 63903 34796 63969 34819
rect 63583 34756 63592 34796
rect 63632 34756 63649 34796
rect 63735 34756 63756 34796
rect 63796 34756 63817 34796
rect 63903 34756 63920 34796
rect 63960 34756 63969 34796
rect 63583 34733 63649 34756
rect 63735 34733 63817 34756
rect 63903 34733 63969 34756
rect 63583 34714 63969 34733
rect 78703 34819 79089 34838
rect 78703 34796 78769 34819
rect 78855 34796 78937 34819
rect 79023 34796 79089 34819
rect 78703 34756 78712 34796
rect 78752 34756 78769 34796
rect 78855 34756 78876 34796
rect 78916 34756 78937 34796
rect 79023 34756 79040 34796
rect 79080 34756 79089 34796
rect 78703 34733 78769 34756
rect 78855 34733 78937 34756
rect 79023 34733 79089 34756
rect 78703 34714 79089 34733
rect 93823 34819 94209 34838
rect 93823 34796 93889 34819
rect 93975 34796 94057 34819
rect 94143 34796 94209 34819
rect 93823 34756 93832 34796
rect 93872 34756 93889 34796
rect 93975 34756 93996 34796
rect 94036 34756 94057 34796
rect 94143 34756 94160 34796
rect 94200 34756 94209 34796
rect 93823 34733 93889 34756
rect 93975 34733 94057 34756
rect 94143 34733 94209 34756
rect 93823 34714 94209 34733
rect 4343 34063 4729 34082
rect 4343 34040 4409 34063
rect 4495 34040 4577 34063
rect 4663 34040 4729 34063
rect 4343 34000 4352 34040
rect 4392 34000 4409 34040
rect 4495 34000 4516 34040
rect 4556 34000 4577 34040
rect 4663 34000 4680 34040
rect 4720 34000 4729 34040
rect 4343 33977 4409 34000
rect 4495 33977 4577 34000
rect 4663 33977 4729 34000
rect 4343 33958 4729 33977
rect 19463 34063 19849 34082
rect 19463 34040 19529 34063
rect 19615 34040 19697 34063
rect 19783 34040 19849 34063
rect 19463 34000 19472 34040
rect 19512 34000 19529 34040
rect 19615 34000 19636 34040
rect 19676 34000 19697 34040
rect 19783 34000 19800 34040
rect 19840 34000 19849 34040
rect 19463 33977 19529 34000
rect 19615 33977 19697 34000
rect 19783 33977 19849 34000
rect 19463 33958 19849 33977
rect 34583 34063 34969 34082
rect 34583 34040 34649 34063
rect 34735 34040 34817 34063
rect 34903 34040 34969 34063
rect 34583 34000 34592 34040
rect 34632 34000 34649 34040
rect 34735 34000 34756 34040
rect 34796 34000 34817 34040
rect 34903 34000 34920 34040
rect 34960 34000 34969 34040
rect 34583 33977 34649 34000
rect 34735 33977 34817 34000
rect 34903 33977 34969 34000
rect 34583 33958 34969 33977
rect 49703 34063 50089 34082
rect 49703 34040 49769 34063
rect 49855 34040 49937 34063
rect 50023 34040 50089 34063
rect 49703 34000 49712 34040
rect 49752 34000 49769 34040
rect 49855 34000 49876 34040
rect 49916 34000 49937 34040
rect 50023 34000 50040 34040
rect 50080 34000 50089 34040
rect 49703 33977 49769 34000
rect 49855 33977 49937 34000
rect 50023 33977 50089 34000
rect 49703 33958 50089 33977
rect 64823 34063 65209 34082
rect 64823 34040 64889 34063
rect 64975 34040 65057 34063
rect 65143 34040 65209 34063
rect 64823 34000 64832 34040
rect 64872 34000 64889 34040
rect 64975 34000 64996 34040
rect 65036 34000 65057 34040
rect 65143 34000 65160 34040
rect 65200 34000 65209 34040
rect 64823 33977 64889 34000
rect 64975 33977 65057 34000
rect 65143 33977 65209 34000
rect 64823 33958 65209 33977
rect 79943 34063 80329 34082
rect 79943 34040 80009 34063
rect 80095 34040 80177 34063
rect 80263 34040 80329 34063
rect 79943 34000 79952 34040
rect 79992 34000 80009 34040
rect 80095 34000 80116 34040
rect 80156 34000 80177 34040
rect 80263 34000 80280 34040
rect 80320 34000 80329 34040
rect 79943 33977 80009 34000
rect 80095 33977 80177 34000
rect 80263 33977 80329 34000
rect 79943 33958 80329 33977
rect 95063 34063 95449 34082
rect 95063 34040 95129 34063
rect 95215 34040 95297 34063
rect 95383 34040 95449 34063
rect 95063 34000 95072 34040
rect 95112 34000 95129 34040
rect 95215 34000 95236 34040
rect 95276 34000 95297 34040
rect 95383 34000 95400 34040
rect 95440 34000 95449 34040
rect 95063 33977 95129 34000
rect 95215 33977 95297 34000
rect 95383 33977 95449 34000
rect 95063 33958 95449 33977
rect 3103 33307 3489 33326
rect 3103 33284 3169 33307
rect 3255 33284 3337 33307
rect 3423 33284 3489 33307
rect 3103 33244 3112 33284
rect 3152 33244 3169 33284
rect 3255 33244 3276 33284
rect 3316 33244 3337 33284
rect 3423 33244 3440 33284
rect 3480 33244 3489 33284
rect 3103 33221 3169 33244
rect 3255 33221 3337 33244
rect 3423 33221 3489 33244
rect 3103 33202 3489 33221
rect 18223 33307 18609 33326
rect 18223 33284 18289 33307
rect 18375 33284 18457 33307
rect 18543 33284 18609 33307
rect 18223 33244 18232 33284
rect 18272 33244 18289 33284
rect 18375 33244 18396 33284
rect 18436 33244 18457 33284
rect 18543 33244 18560 33284
rect 18600 33244 18609 33284
rect 18223 33221 18289 33244
rect 18375 33221 18457 33244
rect 18543 33221 18609 33244
rect 18223 33202 18609 33221
rect 33343 33307 33729 33326
rect 33343 33284 33409 33307
rect 33495 33284 33577 33307
rect 33663 33284 33729 33307
rect 33343 33244 33352 33284
rect 33392 33244 33409 33284
rect 33495 33244 33516 33284
rect 33556 33244 33577 33284
rect 33663 33244 33680 33284
rect 33720 33244 33729 33284
rect 33343 33221 33409 33244
rect 33495 33221 33577 33244
rect 33663 33221 33729 33244
rect 33343 33202 33729 33221
rect 48463 33307 48849 33326
rect 48463 33284 48529 33307
rect 48615 33284 48697 33307
rect 48783 33284 48849 33307
rect 48463 33244 48472 33284
rect 48512 33244 48529 33284
rect 48615 33244 48636 33284
rect 48676 33244 48697 33284
rect 48783 33244 48800 33284
rect 48840 33244 48849 33284
rect 48463 33221 48529 33244
rect 48615 33221 48697 33244
rect 48783 33221 48849 33244
rect 48463 33202 48849 33221
rect 63583 33307 63969 33326
rect 63583 33284 63649 33307
rect 63735 33284 63817 33307
rect 63903 33284 63969 33307
rect 63583 33244 63592 33284
rect 63632 33244 63649 33284
rect 63735 33244 63756 33284
rect 63796 33244 63817 33284
rect 63903 33244 63920 33284
rect 63960 33244 63969 33284
rect 63583 33221 63649 33244
rect 63735 33221 63817 33244
rect 63903 33221 63969 33244
rect 63583 33202 63969 33221
rect 78703 33307 79089 33326
rect 78703 33284 78769 33307
rect 78855 33284 78937 33307
rect 79023 33284 79089 33307
rect 78703 33244 78712 33284
rect 78752 33244 78769 33284
rect 78855 33244 78876 33284
rect 78916 33244 78937 33284
rect 79023 33244 79040 33284
rect 79080 33244 79089 33284
rect 78703 33221 78769 33244
rect 78855 33221 78937 33244
rect 79023 33221 79089 33244
rect 78703 33202 79089 33221
rect 93823 33307 94209 33326
rect 93823 33284 93889 33307
rect 93975 33284 94057 33307
rect 94143 33284 94209 33307
rect 93823 33244 93832 33284
rect 93872 33244 93889 33284
rect 93975 33244 93996 33284
rect 94036 33244 94057 33284
rect 94143 33244 94160 33284
rect 94200 33244 94209 33284
rect 93823 33221 93889 33244
rect 93975 33221 94057 33244
rect 94143 33221 94209 33244
rect 93823 33202 94209 33221
rect 4343 32551 4729 32570
rect 4343 32528 4409 32551
rect 4495 32528 4577 32551
rect 4663 32528 4729 32551
rect 4343 32488 4352 32528
rect 4392 32488 4409 32528
rect 4495 32488 4516 32528
rect 4556 32488 4577 32528
rect 4663 32488 4680 32528
rect 4720 32488 4729 32528
rect 4343 32465 4409 32488
rect 4495 32465 4577 32488
rect 4663 32465 4729 32488
rect 4343 32446 4729 32465
rect 19463 32551 19849 32570
rect 19463 32528 19529 32551
rect 19615 32528 19697 32551
rect 19783 32528 19849 32551
rect 19463 32488 19472 32528
rect 19512 32488 19529 32528
rect 19615 32488 19636 32528
rect 19676 32488 19697 32528
rect 19783 32488 19800 32528
rect 19840 32488 19849 32528
rect 19463 32465 19529 32488
rect 19615 32465 19697 32488
rect 19783 32465 19849 32488
rect 19463 32446 19849 32465
rect 34583 32551 34969 32570
rect 34583 32528 34649 32551
rect 34735 32528 34817 32551
rect 34903 32528 34969 32551
rect 34583 32488 34592 32528
rect 34632 32488 34649 32528
rect 34735 32488 34756 32528
rect 34796 32488 34817 32528
rect 34903 32488 34920 32528
rect 34960 32488 34969 32528
rect 34583 32465 34649 32488
rect 34735 32465 34817 32488
rect 34903 32465 34969 32488
rect 34583 32446 34969 32465
rect 49703 32551 50089 32570
rect 49703 32528 49769 32551
rect 49855 32528 49937 32551
rect 50023 32528 50089 32551
rect 49703 32488 49712 32528
rect 49752 32488 49769 32528
rect 49855 32488 49876 32528
rect 49916 32488 49937 32528
rect 50023 32488 50040 32528
rect 50080 32488 50089 32528
rect 49703 32465 49769 32488
rect 49855 32465 49937 32488
rect 50023 32465 50089 32488
rect 49703 32446 50089 32465
rect 64823 32551 65209 32570
rect 64823 32528 64889 32551
rect 64975 32528 65057 32551
rect 65143 32528 65209 32551
rect 64823 32488 64832 32528
rect 64872 32488 64889 32528
rect 64975 32488 64996 32528
rect 65036 32488 65057 32528
rect 65143 32488 65160 32528
rect 65200 32488 65209 32528
rect 64823 32465 64889 32488
rect 64975 32465 65057 32488
rect 65143 32465 65209 32488
rect 64823 32446 65209 32465
rect 79943 32551 80329 32570
rect 79943 32528 80009 32551
rect 80095 32528 80177 32551
rect 80263 32528 80329 32551
rect 79943 32488 79952 32528
rect 79992 32488 80009 32528
rect 80095 32488 80116 32528
rect 80156 32488 80177 32528
rect 80263 32488 80280 32528
rect 80320 32488 80329 32528
rect 79943 32465 80009 32488
rect 80095 32465 80177 32488
rect 80263 32465 80329 32488
rect 79943 32446 80329 32465
rect 95063 32551 95449 32570
rect 95063 32528 95129 32551
rect 95215 32528 95297 32551
rect 95383 32528 95449 32551
rect 95063 32488 95072 32528
rect 95112 32488 95129 32528
rect 95215 32488 95236 32528
rect 95276 32488 95297 32528
rect 95383 32488 95400 32528
rect 95440 32488 95449 32528
rect 95063 32465 95129 32488
rect 95215 32465 95297 32488
rect 95383 32465 95449 32488
rect 95063 32446 95449 32465
rect 3103 31795 3489 31814
rect 3103 31772 3169 31795
rect 3255 31772 3337 31795
rect 3423 31772 3489 31795
rect 3103 31732 3112 31772
rect 3152 31732 3169 31772
rect 3255 31732 3276 31772
rect 3316 31732 3337 31772
rect 3423 31732 3440 31772
rect 3480 31732 3489 31772
rect 3103 31709 3169 31732
rect 3255 31709 3337 31732
rect 3423 31709 3489 31732
rect 3103 31690 3489 31709
rect 18223 31795 18609 31814
rect 18223 31772 18289 31795
rect 18375 31772 18457 31795
rect 18543 31772 18609 31795
rect 18223 31732 18232 31772
rect 18272 31732 18289 31772
rect 18375 31732 18396 31772
rect 18436 31732 18457 31772
rect 18543 31732 18560 31772
rect 18600 31732 18609 31772
rect 18223 31709 18289 31732
rect 18375 31709 18457 31732
rect 18543 31709 18609 31732
rect 18223 31690 18609 31709
rect 33343 31795 33729 31814
rect 33343 31772 33409 31795
rect 33495 31772 33577 31795
rect 33663 31772 33729 31795
rect 33343 31732 33352 31772
rect 33392 31732 33409 31772
rect 33495 31732 33516 31772
rect 33556 31732 33577 31772
rect 33663 31732 33680 31772
rect 33720 31732 33729 31772
rect 33343 31709 33409 31732
rect 33495 31709 33577 31732
rect 33663 31709 33729 31732
rect 33343 31690 33729 31709
rect 48463 31795 48849 31814
rect 48463 31772 48529 31795
rect 48615 31772 48697 31795
rect 48783 31772 48849 31795
rect 48463 31732 48472 31772
rect 48512 31732 48529 31772
rect 48615 31732 48636 31772
rect 48676 31732 48697 31772
rect 48783 31732 48800 31772
rect 48840 31732 48849 31772
rect 48463 31709 48529 31732
rect 48615 31709 48697 31732
rect 48783 31709 48849 31732
rect 48463 31690 48849 31709
rect 63583 31795 63969 31814
rect 63583 31772 63649 31795
rect 63735 31772 63817 31795
rect 63903 31772 63969 31795
rect 63583 31732 63592 31772
rect 63632 31732 63649 31772
rect 63735 31732 63756 31772
rect 63796 31732 63817 31772
rect 63903 31732 63920 31772
rect 63960 31732 63969 31772
rect 63583 31709 63649 31732
rect 63735 31709 63817 31732
rect 63903 31709 63969 31732
rect 63583 31690 63969 31709
rect 78703 31795 79089 31814
rect 78703 31772 78769 31795
rect 78855 31772 78937 31795
rect 79023 31772 79089 31795
rect 78703 31732 78712 31772
rect 78752 31732 78769 31772
rect 78855 31732 78876 31772
rect 78916 31732 78937 31772
rect 79023 31732 79040 31772
rect 79080 31732 79089 31772
rect 78703 31709 78769 31732
rect 78855 31709 78937 31732
rect 79023 31709 79089 31732
rect 78703 31690 79089 31709
rect 93823 31795 94209 31814
rect 93823 31772 93889 31795
rect 93975 31772 94057 31795
rect 94143 31772 94209 31795
rect 93823 31732 93832 31772
rect 93872 31732 93889 31772
rect 93975 31732 93996 31772
rect 94036 31732 94057 31772
rect 94143 31732 94160 31772
rect 94200 31732 94209 31772
rect 93823 31709 93889 31732
rect 93975 31709 94057 31732
rect 94143 31709 94209 31732
rect 93823 31690 94209 31709
rect 4343 31039 4729 31058
rect 4343 31016 4409 31039
rect 4495 31016 4577 31039
rect 4663 31016 4729 31039
rect 4343 30976 4352 31016
rect 4392 30976 4409 31016
rect 4495 30976 4516 31016
rect 4556 30976 4577 31016
rect 4663 30976 4680 31016
rect 4720 30976 4729 31016
rect 4343 30953 4409 30976
rect 4495 30953 4577 30976
rect 4663 30953 4729 30976
rect 4343 30934 4729 30953
rect 19463 31039 19849 31058
rect 19463 31016 19529 31039
rect 19615 31016 19697 31039
rect 19783 31016 19849 31039
rect 19463 30976 19472 31016
rect 19512 30976 19529 31016
rect 19615 30976 19636 31016
rect 19676 30976 19697 31016
rect 19783 30976 19800 31016
rect 19840 30976 19849 31016
rect 19463 30953 19529 30976
rect 19615 30953 19697 30976
rect 19783 30953 19849 30976
rect 19463 30934 19849 30953
rect 34583 31039 34969 31058
rect 34583 31016 34649 31039
rect 34735 31016 34817 31039
rect 34903 31016 34969 31039
rect 34583 30976 34592 31016
rect 34632 30976 34649 31016
rect 34735 30976 34756 31016
rect 34796 30976 34817 31016
rect 34903 30976 34920 31016
rect 34960 30976 34969 31016
rect 34583 30953 34649 30976
rect 34735 30953 34817 30976
rect 34903 30953 34969 30976
rect 34583 30934 34969 30953
rect 49703 31039 50089 31058
rect 49703 31016 49769 31039
rect 49855 31016 49937 31039
rect 50023 31016 50089 31039
rect 49703 30976 49712 31016
rect 49752 30976 49769 31016
rect 49855 30976 49876 31016
rect 49916 30976 49937 31016
rect 50023 30976 50040 31016
rect 50080 30976 50089 31016
rect 49703 30953 49769 30976
rect 49855 30953 49937 30976
rect 50023 30953 50089 30976
rect 49703 30934 50089 30953
rect 64823 31039 65209 31058
rect 64823 31016 64889 31039
rect 64975 31016 65057 31039
rect 65143 31016 65209 31039
rect 64823 30976 64832 31016
rect 64872 30976 64889 31016
rect 64975 30976 64996 31016
rect 65036 30976 65057 31016
rect 65143 30976 65160 31016
rect 65200 30976 65209 31016
rect 64823 30953 64889 30976
rect 64975 30953 65057 30976
rect 65143 30953 65209 30976
rect 64823 30934 65209 30953
rect 79943 31039 80329 31058
rect 79943 31016 80009 31039
rect 80095 31016 80177 31039
rect 80263 31016 80329 31039
rect 79943 30976 79952 31016
rect 79992 30976 80009 31016
rect 80095 30976 80116 31016
rect 80156 30976 80177 31016
rect 80263 30976 80280 31016
rect 80320 30976 80329 31016
rect 79943 30953 80009 30976
rect 80095 30953 80177 30976
rect 80263 30953 80329 30976
rect 79943 30934 80329 30953
rect 95063 31039 95449 31058
rect 95063 31016 95129 31039
rect 95215 31016 95297 31039
rect 95383 31016 95449 31039
rect 95063 30976 95072 31016
rect 95112 30976 95129 31016
rect 95215 30976 95236 31016
rect 95276 30976 95297 31016
rect 95383 30976 95400 31016
rect 95440 30976 95449 31016
rect 95063 30953 95129 30976
rect 95215 30953 95297 30976
rect 95383 30953 95449 30976
rect 95063 30934 95449 30953
rect 3103 30283 3489 30302
rect 3103 30260 3169 30283
rect 3255 30260 3337 30283
rect 3423 30260 3489 30283
rect 3103 30220 3112 30260
rect 3152 30220 3169 30260
rect 3255 30220 3276 30260
rect 3316 30220 3337 30260
rect 3423 30220 3440 30260
rect 3480 30220 3489 30260
rect 3103 30197 3169 30220
rect 3255 30197 3337 30220
rect 3423 30197 3489 30220
rect 3103 30178 3489 30197
rect 18223 30283 18609 30302
rect 18223 30260 18289 30283
rect 18375 30260 18457 30283
rect 18543 30260 18609 30283
rect 18223 30220 18232 30260
rect 18272 30220 18289 30260
rect 18375 30220 18396 30260
rect 18436 30220 18457 30260
rect 18543 30220 18560 30260
rect 18600 30220 18609 30260
rect 18223 30197 18289 30220
rect 18375 30197 18457 30220
rect 18543 30197 18609 30220
rect 18223 30178 18609 30197
rect 33343 30283 33729 30302
rect 33343 30260 33409 30283
rect 33495 30260 33577 30283
rect 33663 30260 33729 30283
rect 33343 30220 33352 30260
rect 33392 30220 33409 30260
rect 33495 30220 33516 30260
rect 33556 30220 33577 30260
rect 33663 30220 33680 30260
rect 33720 30220 33729 30260
rect 33343 30197 33409 30220
rect 33495 30197 33577 30220
rect 33663 30197 33729 30220
rect 33343 30178 33729 30197
rect 48463 30283 48849 30302
rect 48463 30260 48529 30283
rect 48615 30260 48697 30283
rect 48783 30260 48849 30283
rect 48463 30220 48472 30260
rect 48512 30220 48529 30260
rect 48615 30220 48636 30260
rect 48676 30220 48697 30260
rect 48783 30220 48800 30260
rect 48840 30220 48849 30260
rect 48463 30197 48529 30220
rect 48615 30197 48697 30220
rect 48783 30197 48849 30220
rect 48463 30178 48849 30197
rect 63583 30283 63969 30302
rect 63583 30260 63649 30283
rect 63735 30260 63817 30283
rect 63903 30260 63969 30283
rect 63583 30220 63592 30260
rect 63632 30220 63649 30260
rect 63735 30220 63756 30260
rect 63796 30220 63817 30260
rect 63903 30220 63920 30260
rect 63960 30220 63969 30260
rect 63583 30197 63649 30220
rect 63735 30197 63817 30220
rect 63903 30197 63969 30220
rect 63583 30178 63969 30197
rect 78703 30283 79089 30302
rect 78703 30260 78769 30283
rect 78855 30260 78937 30283
rect 79023 30260 79089 30283
rect 78703 30220 78712 30260
rect 78752 30220 78769 30260
rect 78855 30220 78876 30260
rect 78916 30220 78937 30260
rect 79023 30220 79040 30260
rect 79080 30220 79089 30260
rect 78703 30197 78769 30220
rect 78855 30197 78937 30220
rect 79023 30197 79089 30220
rect 78703 30178 79089 30197
rect 93823 30283 94209 30302
rect 93823 30260 93889 30283
rect 93975 30260 94057 30283
rect 94143 30260 94209 30283
rect 93823 30220 93832 30260
rect 93872 30220 93889 30260
rect 93975 30220 93996 30260
rect 94036 30220 94057 30260
rect 94143 30220 94160 30260
rect 94200 30220 94209 30260
rect 93823 30197 93889 30220
rect 93975 30197 94057 30220
rect 94143 30197 94209 30220
rect 93823 30178 94209 30197
rect 4343 29527 4729 29546
rect 4343 29504 4409 29527
rect 4495 29504 4577 29527
rect 4663 29504 4729 29527
rect 4343 29464 4352 29504
rect 4392 29464 4409 29504
rect 4495 29464 4516 29504
rect 4556 29464 4577 29504
rect 4663 29464 4680 29504
rect 4720 29464 4729 29504
rect 4343 29441 4409 29464
rect 4495 29441 4577 29464
rect 4663 29441 4729 29464
rect 4343 29422 4729 29441
rect 19463 29527 19849 29546
rect 19463 29504 19529 29527
rect 19615 29504 19697 29527
rect 19783 29504 19849 29527
rect 19463 29464 19472 29504
rect 19512 29464 19529 29504
rect 19615 29464 19636 29504
rect 19676 29464 19697 29504
rect 19783 29464 19800 29504
rect 19840 29464 19849 29504
rect 19463 29441 19529 29464
rect 19615 29441 19697 29464
rect 19783 29441 19849 29464
rect 19463 29422 19849 29441
rect 34583 29527 34969 29546
rect 34583 29504 34649 29527
rect 34735 29504 34817 29527
rect 34903 29504 34969 29527
rect 34583 29464 34592 29504
rect 34632 29464 34649 29504
rect 34735 29464 34756 29504
rect 34796 29464 34817 29504
rect 34903 29464 34920 29504
rect 34960 29464 34969 29504
rect 34583 29441 34649 29464
rect 34735 29441 34817 29464
rect 34903 29441 34969 29464
rect 34583 29422 34969 29441
rect 49703 29527 50089 29546
rect 49703 29504 49769 29527
rect 49855 29504 49937 29527
rect 50023 29504 50089 29527
rect 49703 29464 49712 29504
rect 49752 29464 49769 29504
rect 49855 29464 49876 29504
rect 49916 29464 49937 29504
rect 50023 29464 50040 29504
rect 50080 29464 50089 29504
rect 49703 29441 49769 29464
rect 49855 29441 49937 29464
rect 50023 29441 50089 29464
rect 49703 29422 50089 29441
rect 64823 29527 65209 29546
rect 64823 29504 64889 29527
rect 64975 29504 65057 29527
rect 65143 29504 65209 29527
rect 64823 29464 64832 29504
rect 64872 29464 64889 29504
rect 64975 29464 64996 29504
rect 65036 29464 65057 29504
rect 65143 29464 65160 29504
rect 65200 29464 65209 29504
rect 64823 29441 64889 29464
rect 64975 29441 65057 29464
rect 65143 29441 65209 29464
rect 64823 29422 65209 29441
rect 79943 29527 80329 29546
rect 79943 29504 80009 29527
rect 80095 29504 80177 29527
rect 80263 29504 80329 29527
rect 79943 29464 79952 29504
rect 79992 29464 80009 29504
rect 80095 29464 80116 29504
rect 80156 29464 80177 29504
rect 80263 29464 80280 29504
rect 80320 29464 80329 29504
rect 79943 29441 80009 29464
rect 80095 29441 80177 29464
rect 80263 29441 80329 29464
rect 79943 29422 80329 29441
rect 95063 29527 95449 29546
rect 95063 29504 95129 29527
rect 95215 29504 95297 29527
rect 95383 29504 95449 29527
rect 95063 29464 95072 29504
rect 95112 29464 95129 29504
rect 95215 29464 95236 29504
rect 95276 29464 95297 29504
rect 95383 29464 95400 29504
rect 95440 29464 95449 29504
rect 95063 29441 95129 29464
rect 95215 29441 95297 29464
rect 95383 29441 95449 29464
rect 95063 29422 95449 29441
rect 3103 28771 3489 28790
rect 3103 28748 3169 28771
rect 3255 28748 3337 28771
rect 3423 28748 3489 28771
rect 3103 28708 3112 28748
rect 3152 28708 3169 28748
rect 3255 28708 3276 28748
rect 3316 28708 3337 28748
rect 3423 28708 3440 28748
rect 3480 28708 3489 28748
rect 3103 28685 3169 28708
rect 3255 28685 3337 28708
rect 3423 28685 3489 28708
rect 3103 28666 3489 28685
rect 18223 28771 18609 28790
rect 18223 28748 18289 28771
rect 18375 28748 18457 28771
rect 18543 28748 18609 28771
rect 18223 28708 18232 28748
rect 18272 28708 18289 28748
rect 18375 28708 18396 28748
rect 18436 28708 18457 28748
rect 18543 28708 18560 28748
rect 18600 28708 18609 28748
rect 18223 28685 18289 28708
rect 18375 28685 18457 28708
rect 18543 28685 18609 28708
rect 18223 28666 18609 28685
rect 33343 28771 33729 28790
rect 33343 28748 33409 28771
rect 33495 28748 33577 28771
rect 33663 28748 33729 28771
rect 33343 28708 33352 28748
rect 33392 28708 33409 28748
rect 33495 28708 33516 28748
rect 33556 28708 33577 28748
rect 33663 28708 33680 28748
rect 33720 28708 33729 28748
rect 33343 28685 33409 28708
rect 33495 28685 33577 28708
rect 33663 28685 33729 28708
rect 33343 28666 33729 28685
rect 48463 28771 48849 28790
rect 48463 28748 48529 28771
rect 48615 28748 48697 28771
rect 48783 28748 48849 28771
rect 48463 28708 48472 28748
rect 48512 28708 48529 28748
rect 48615 28708 48636 28748
rect 48676 28708 48697 28748
rect 48783 28708 48800 28748
rect 48840 28708 48849 28748
rect 48463 28685 48529 28708
rect 48615 28685 48697 28708
rect 48783 28685 48849 28708
rect 48463 28666 48849 28685
rect 63583 28771 63969 28790
rect 63583 28748 63649 28771
rect 63735 28748 63817 28771
rect 63903 28748 63969 28771
rect 63583 28708 63592 28748
rect 63632 28708 63649 28748
rect 63735 28708 63756 28748
rect 63796 28708 63817 28748
rect 63903 28708 63920 28748
rect 63960 28708 63969 28748
rect 63583 28685 63649 28708
rect 63735 28685 63817 28708
rect 63903 28685 63969 28708
rect 63583 28666 63969 28685
rect 78703 28771 79089 28790
rect 78703 28748 78769 28771
rect 78855 28748 78937 28771
rect 79023 28748 79089 28771
rect 78703 28708 78712 28748
rect 78752 28708 78769 28748
rect 78855 28708 78876 28748
rect 78916 28708 78937 28748
rect 79023 28708 79040 28748
rect 79080 28708 79089 28748
rect 78703 28685 78769 28708
rect 78855 28685 78937 28708
rect 79023 28685 79089 28708
rect 78703 28666 79089 28685
rect 93823 28771 94209 28790
rect 93823 28748 93889 28771
rect 93975 28748 94057 28771
rect 94143 28748 94209 28771
rect 93823 28708 93832 28748
rect 93872 28708 93889 28748
rect 93975 28708 93996 28748
rect 94036 28708 94057 28748
rect 94143 28708 94160 28748
rect 94200 28708 94209 28748
rect 93823 28685 93889 28708
rect 93975 28685 94057 28708
rect 94143 28685 94209 28708
rect 93823 28666 94209 28685
rect 4343 28015 4729 28034
rect 4343 27992 4409 28015
rect 4495 27992 4577 28015
rect 4663 27992 4729 28015
rect 4343 27952 4352 27992
rect 4392 27952 4409 27992
rect 4495 27952 4516 27992
rect 4556 27952 4577 27992
rect 4663 27952 4680 27992
rect 4720 27952 4729 27992
rect 4343 27929 4409 27952
rect 4495 27929 4577 27952
rect 4663 27929 4729 27952
rect 4343 27910 4729 27929
rect 19463 28015 19849 28034
rect 19463 27992 19529 28015
rect 19615 27992 19697 28015
rect 19783 27992 19849 28015
rect 19463 27952 19472 27992
rect 19512 27952 19529 27992
rect 19615 27952 19636 27992
rect 19676 27952 19697 27992
rect 19783 27952 19800 27992
rect 19840 27952 19849 27992
rect 19463 27929 19529 27952
rect 19615 27929 19697 27952
rect 19783 27929 19849 27952
rect 19463 27910 19849 27929
rect 34583 28015 34969 28034
rect 34583 27992 34649 28015
rect 34735 27992 34817 28015
rect 34903 27992 34969 28015
rect 34583 27952 34592 27992
rect 34632 27952 34649 27992
rect 34735 27952 34756 27992
rect 34796 27952 34817 27992
rect 34903 27952 34920 27992
rect 34960 27952 34969 27992
rect 34583 27929 34649 27952
rect 34735 27929 34817 27952
rect 34903 27929 34969 27952
rect 34583 27910 34969 27929
rect 49703 28015 50089 28034
rect 49703 27992 49769 28015
rect 49855 27992 49937 28015
rect 50023 27992 50089 28015
rect 49703 27952 49712 27992
rect 49752 27952 49769 27992
rect 49855 27952 49876 27992
rect 49916 27952 49937 27992
rect 50023 27952 50040 27992
rect 50080 27952 50089 27992
rect 49703 27929 49769 27952
rect 49855 27929 49937 27952
rect 50023 27929 50089 27952
rect 49703 27910 50089 27929
rect 64823 28015 65209 28034
rect 64823 27992 64889 28015
rect 64975 27992 65057 28015
rect 65143 27992 65209 28015
rect 64823 27952 64832 27992
rect 64872 27952 64889 27992
rect 64975 27952 64996 27992
rect 65036 27952 65057 27992
rect 65143 27952 65160 27992
rect 65200 27952 65209 27992
rect 64823 27929 64889 27952
rect 64975 27929 65057 27952
rect 65143 27929 65209 27952
rect 64823 27910 65209 27929
rect 79943 28015 80329 28034
rect 79943 27992 80009 28015
rect 80095 27992 80177 28015
rect 80263 27992 80329 28015
rect 79943 27952 79952 27992
rect 79992 27952 80009 27992
rect 80095 27952 80116 27992
rect 80156 27952 80177 27992
rect 80263 27952 80280 27992
rect 80320 27952 80329 27992
rect 79943 27929 80009 27952
rect 80095 27929 80177 27952
rect 80263 27929 80329 27952
rect 79943 27910 80329 27929
rect 95063 28015 95449 28034
rect 95063 27992 95129 28015
rect 95215 27992 95297 28015
rect 95383 27992 95449 28015
rect 95063 27952 95072 27992
rect 95112 27952 95129 27992
rect 95215 27952 95236 27992
rect 95276 27952 95297 27992
rect 95383 27952 95400 27992
rect 95440 27952 95449 27992
rect 95063 27929 95129 27952
rect 95215 27929 95297 27952
rect 95383 27929 95449 27952
rect 95063 27910 95449 27929
rect 3103 27259 3489 27278
rect 3103 27236 3169 27259
rect 3255 27236 3337 27259
rect 3423 27236 3489 27259
rect 3103 27196 3112 27236
rect 3152 27196 3169 27236
rect 3255 27196 3276 27236
rect 3316 27196 3337 27236
rect 3423 27196 3440 27236
rect 3480 27196 3489 27236
rect 3103 27173 3169 27196
rect 3255 27173 3337 27196
rect 3423 27173 3489 27196
rect 3103 27154 3489 27173
rect 18223 27259 18609 27278
rect 18223 27236 18289 27259
rect 18375 27236 18457 27259
rect 18543 27236 18609 27259
rect 18223 27196 18232 27236
rect 18272 27196 18289 27236
rect 18375 27196 18396 27236
rect 18436 27196 18457 27236
rect 18543 27196 18560 27236
rect 18600 27196 18609 27236
rect 18223 27173 18289 27196
rect 18375 27173 18457 27196
rect 18543 27173 18609 27196
rect 18223 27154 18609 27173
rect 33343 27259 33729 27278
rect 33343 27236 33409 27259
rect 33495 27236 33577 27259
rect 33663 27236 33729 27259
rect 33343 27196 33352 27236
rect 33392 27196 33409 27236
rect 33495 27196 33516 27236
rect 33556 27196 33577 27236
rect 33663 27196 33680 27236
rect 33720 27196 33729 27236
rect 33343 27173 33409 27196
rect 33495 27173 33577 27196
rect 33663 27173 33729 27196
rect 33343 27154 33729 27173
rect 48463 27259 48849 27278
rect 48463 27236 48529 27259
rect 48615 27236 48697 27259
rect 48783 27236 48849 27259
rect 48463 27196 48472 27236
rect 48512 27196 48529 27236
rect 48615 27196 48636 27236
rect 48676 27196 48697 27236
rect 48783 27196 48800 27236
rect 48840 27196 48849 27236
rect 48463 27173 48529 27196
rect 48615 27173 48697 27196
rect 48783 27173 48849 27196
rect 48463 27154 48849 27173
rect 63583 27259 63969 27278
rect 63583 27236 63649 27259
rect 63735 27236 63817 27259
rect 63903 27236 63969 27259
rect 63583 27196 63592 27236
rect 63632 27196 63649 27236
rect 63735 27196 63756 27236
rect 63796 27196 63817 27236
rect 63903 27196 63920 27236
rect 63960 27196 63969 27236
rect 63583 27173 63649 27196
rect 63735 27173 63817 27196
rect 63903 27173 63969 27196
rect 63583 27154 63969 27173
rect 78703 27259 79089 27278
rect 78703 27236 78769 27259
rect 78855 27236 78937 27259
rect 79023 27236 79089 27259
rect 78703 27196 78712 27236
rect 78752 27196 78769 27236
rect 78855 27196 78876 27236
rect 78916 27196 78937 27236
rect 79023 27196 79040 27236
rect 79080 27196 79089 27236
rect 78703 27173 78769 27196
rect 78855 27173 78937 27196
rect 79023 27173 79089 27196
rect 78703 27154 79089 27173
rect 93823 27259 94209 27278
rect 93823 27236 93889 27259
rect 93975 27236 94057 27259
rect 94143 27236 94209 27259
rect 93823 27196 93832 27236
rect 93872 27196 93889 27236
rect 93975 27196 93996 27236
rect 94036 27196 94057 27236
rect 94143 27196 94160 27236
rect 94200 27196 94209 27236
rect 93823 27173 93889 27196
rect 93975 27173 94057 27196
rect 94143 27173 94209 27196
rect 93823 27154 94209 27173
rect 4343 26503 4729 26522
rect 4343 26480 4409 26503
rect 4495 26480 4577 26503
rect 4663 26480 4729 26503
rect 4343 26440 4352 26480
rect 4392 26440 4409 26480
rect 4495 26440 4516 26480
rect 4556 26440 4577 26480
rect 4663 26440 4680 26480
rect 4720 26440 4729 26480
rect 4343 26417 4409 26440
rect 4495 26417 4577 26440
rect 4663 26417 4729 26440
rect 4343 26398 4729 26417
rect 19463 26503 19849 26522
rect 19463 26480 19529 26503
rect 19615 26480 19697 26503
rect 19783 26480 19849 26503
rect 19463 26440 19472 26480
rect 19512 26440 19529 26480
rect 19615 26440 19636 26480
rect 19676 26440 19697 26480
rect 19783 26440 19800 26480
rect 19840 26440 19849 26480
rect 19463 26417 19529 26440
rect 19615 26417 19697 26440
rect 19783 26417 19849 26440
rect 19463 26398 19849 26417
rect 34583 26503 34969 26522
rect 34583 26480 34649 26503
rect 34735 26480 34817 26503
rect 34903 26480 34969 26503
rect 34583 26440 34592 26480
rect 34632 26440 34649 26480
rect 34735 26440 34756 26480
rect 34796 26440 34817 26480
rect 34903 26440 34920 26480
rect 34960 26440 34969 26480
rect 34583 26417 34649 26440
rect 34735 26417 34817 26440
rect 34903 26417 34969 26440
rect 34583 26398 34969 26417
rect 49703 26503 50089 26522
rect 49703 26480 49769 26503
rect 49855 26480 49937 26503
rect 50023 26480 50089 26503
rect 49703 26440 49712 26480
rect 49752 26440 49769 26480
rect 49855 26440 49876 26480
rect 49916 26440 49937 26480
rect 50023 26440 50040 26480
rect 50080 26440 50089 26480
rect 49703 26417 49769 26440
rect 49855 26417 49937 26440
rect 50023 26417 50089 26440
rect 49703 26398 50089 26417
rect 64823 26503 65209 26522
rect 64823 26480 64889 26503
rect 64975 26480 65057 26503
rect 65143 26480 65209 26503
rect 64823 26440 64832 26480
rect 64872 26440 64889 26480
rect 64975 26440 64996 26480
rect 65036 26440 65057 26480
rect 65143 26440 65160 26480
rect 65200 26440 65209 26480
rect 64823 26417 64889 26440
rect 64975 26417 65057 26440
rect 65143 26417 65209 26440
rect 64823 26398 65209 26417
rect 79943 26503 80329 26522
rect 79943 26480 80009 26503
rect 80095 26480 80177 26503
rect 80263 26480 80329 26503
rect 79943 26440 79952 26480
rect 79992 26440 80009 26480
rect 80095 26440 80116 26480
rect 80156 26440 80177 26480
rect 80263 26440 80280 26480
rect 80320 26440 80329 26480
rect 79943 26417 80009 26440
rect 80095 26417 80177 26440
rect 80263 26417 80329 26440
rect 79943 26398 80329 26417
rect 95063 26503 95449 26522
rect 95063 26480 95129 26503
rect 95215 26480 95297 26503
rect 95383 26480 95449 26503
rect 95063 26440 95072 26480
rect 95112 26440 95129 26480
rect 95215 26440 95236 26480
rect 95276 26440 95297 26480
rect 95383 26440 95400 26480
rect 95440 26440 95449 26480
rect 95063 26417 95129 26440
rect 95215 26417 95297 26440
rect 95383 26417 95449 26440
rect 95063 26398 95449 26417
rect 3103 25747 3489 25766
rect 3103 25724 3169 25747
rect 3255 25724 3337 25747
rect 3423 25724 3489 25747
rect 3103 25684 3112 25724
rect 3152 25684 3169 25724
rect 3255 25684 3276 25724
rect 3316 25684 3337 25724
rect 3423 25684 3440 25724
rect 3480 25684 3489 25724
rect 3103 25661 3169 25684
rect 3255 25661 3337 25684
rect 3423 25661 3489 25684
rect 3103 25642 3489 25661
rect 18223 25747 18609 25766
rect 18223 25724 18289 25747
rect 18375 25724 18457 25747
rect 18543 25724 18609 25747
rect 18223 25684 18232 25724
rect 18272 25684 18289 25724
rect 18375 25684 18396 25724
rect 18436 25684 18457 25724
rect 18543 25684 18560 25724
rect 18600 25684 18609 25724
rect 18223 25661 18289 25684
rect 18375 25661 18457 25684
rect 18543 25661 18609 25684
rect 18223 25642 18609 25661
rect 33343 25747 33729 25766
rect 33343 25724 33409 25747
rect 33495 25724 33577 25747
rect 33663 25724 33729 25747
rect 33343 25684 33352 25724
rect 33392 25684 33409 25724
rect 33495 25684 33516 25724
rect 33556 25684 33577 25724
rect 33663 25684 33680 25724
rect 33720 25684 33729 25724
rect 33343 25661 33409 25684
rect 33495 25661 33577 25684
rect 33663 25661 33729 25684
rect 33343 25642 33729 25661
rect 48463 25747 48849 25766
rect 48463 25724 48529 25747
rect 48615 25724 48697 25747
rect 48783 25724 48849 25747
rect 48463 25684 48472 25724
rect 48512 25684 48529 25724
rect 48615 25684 48636 25724
rect 48676 25684 48697 25724
rect 48783 25684 48800 25724
rect 48840 25684 48849 25724
rect 48463 25661 48529 25684
rect 48615 25661 48697 25684
rect 48783 25661 48849 25684
rect 48463 25642 48849 25661
rect 63583 25747 63969 25766
rect 63583 25724 63649 25747
rect 63735 25724 63817 25747
rect 63903 25724 63969 25747
rect 63583 25684 63592 25724
rect 63632 25684 63649 25724
rect 63735 25684 63756 25724
rect 63796 25684 63817 25724
rect 63903 25684 63920 25724
rect 63960 25684 63969 25724
rect 63583 25661 63649 25684
rect 63735 25661 63817 25684
rect 63903 25661 63969 25684
rect 63583 25642 63969 25661
rect 78703 25747 79089 25766
rect 78703 25724 78769 25747
rect 78855 25724 78937 25747
rect 79023 25724 79089 25747
rect 78703 25684 78712 25724
rect 78752 25684 78769 25724
rect 78855 25684 78876 25724
rect 78916 25684 78937 25724
rect 79023 25684 79040 25724
rect 79080 25684 79089 25724
rect 78703 25661 78769 25684
rect 78855 25661 78937 25684
rect 79023 25661 79089 25684
rect 78703 25642 79089 25661
rect 93823 25747 94209 25766
rect 93823 25724 93889 25747
rect 93975 25724 94057 25747
rect 94143 25724 94209 25747
rect 93823 25684 93832 25724
rect 93872 25684 93889 25724
rect 93975 25684 93996 25724
rect 94036 25684 94057 25724
rect 94143 25684 94160 25724
rect 94200 25684 94209 25724
rect 93823 25661 93889 25684
rect 93975 25661 94057 25684
rect 94143 25661 94209 25684
rect 93823 25642 94209 25661
rect 4343 24991 4729 25010
rect 4343 24968 4409 24991
rect 4495 24968 4577 24991
rect 4663 24968 4729 24991
rect 4343 24928 4352 24968
rect 4392 24928 4409 24968
rect 4495 24928 4516 24968
rect 4556 24928 4577 24968
rect 4663 24928 4680 24968
rect 4720 24928 4729 24968
rect 4343 24905 4409 24928
rect 4495 24905 4577 24928
rect 4663 24905 4729 24928
rect 4343 24886 4729 24905
rect 19463 24991 19849 25010
rect 19463 24968 19529 24991
rect 19615 24968 19697 24991
rect 19783 24968 19849 24991
rect 19463 24928 19472 24968
rect 19512 24928 19529 24968
rect 19615 24928 19636 24968
rect 19676 24928 19697 24968
rect 19783 24928 19800 24968
rect 19840 24928 19849 24968
rect 19463 24905 19529 24928
rect 19615 24905 19697 24928
rect 19783 24905 19849 24928
rect 19463 24886 19849 24905
rect 34583 24991 34969 25010
rect 34583 24968 34649 24991
rect 34735 24968 34817 24991
rect 34903 24968 34969 24991
rect 34583 24928 34592 24968
rect 34632 24928 34649 24968
rect 34735 24928 34756 24968
rect 34796 24928 34817 24968
rect 34903 24928 34920 24968
rect 34960 24928 34969 24968
rect 34583 24905 34649 24928
rect 34735 24905 34817 24928
rect 34903 24905 34969 24928
rect 34583 24886 34969 24905
rect 49703 24991 50089 25010
rect 49703 24968 49769 24991
rect 49855 24968 49937 24991
rect 50023 24968 50089 24991
rect 49703 24928 49712 24968
rect 49752 24928 49769 24968
rect 49855 24928 49876 24968
rect 49916 24928 49937 24968
rect 50023 24928 50040 24968
rect 50080 24928 50089 24968
rect 49703 24905 49769 24928
rect 49855 24905 49937 24928
rect 50023 24905 50089 24928
rect 49703 24886 50089 24905
rect 64823 24991 65209 25010
rect 64823 24968 64889 24991
rect 64975 24968 65057 24991
rect 65143 24968 65209 24991
rect 64823 24928 64832 24968
rect 64872 24928 64889 24968
rect 64975 24928 64996 24968
rect 65036 24928 65057 24968
rect 65143 24928 65160 24968
rect 65200 24928 65209 24968
rect 64823 24905 64889 24928
rect 64975 24905 65057 24928
rect 65143 24905 65209 24928
rect 64823 24886 65209 24905
rect 79943 24991 80329 25010
rect 79943 24968 80009 24991
rect 80095 24968 80177 24991
rect 80263 24968 80329 24991
rect 79943 24928 79952 24968
rect 79992 24928 80009 24968
rect 80095 24928 80116 24968
rect 80156 24928 80177 24968
rect 80263 24928 80280 24968
rect 80320 24928 80329 24968
rect 79943 24905 80009 24928
rect 80095 24905 80177 24928
rect 80263 24905 80329 24928
rect 79943 24886 80329 24905
rect 95063 24991 95449 25010
rect 95063 24968 95129 24991
rect 95215 24968 95297 24991
rect 95383 24968 95449 24991
rect 95063 24928 95072 24968
rect 95112 24928 95129 24968
rect 95215 24928 95236 24968
rect 95276 24928 95297 24968
rect 95383 24928 95400 24968
rect 95440 24928 95449 24968
rect 95063 24905 95129 24928
rect 95215 24905 95297 24928
rect 95383 24905 95449 24928
rect 95063 24886 95449 24905
rect 3103 24235 3489 24254
rect 3103 24212 3169 24235
rect 3255 24212 3337 24235
rect 3423 24212 3489 24235
rect 3103 24172 3112 24212
rect 3152 24172 3169 24212
rect 3255 24172 3276 24212
rect 3316 24172 3337 24212
rect 3423 24172 3440 24212
rect 3480 24172 3489 24212
rect 3103 24149 3169 24172
rect 3255 24149 3337 24172
rect 3423 24149 3489 24172
rect 3103 24130 3489 24149
rect 18223 24235 18609 24254
rect 18223 24212 18289 24235
rect 18375 24212 18457 24235
rect 18543 24212 18609 24235
rect 18223 24172 18232 24212
rect 18272 24172 18289 24212
rect 18375 24172 18396 24212
rect 18436 24172 18457 24212
rect 18543 24172 18560 24212
rect 18600 24172 18609 24212
rect 18223 24149 18289 24172
rect 18375 24149 18457 24172
rect 18543 24149 18609 24172
rect 18223 24130 18609 24149
rect 33343 24235 33729 24254
rect 33343 24212 33409 24235
rect 33495 24212 33577 24235
rect 33663 24212 33729 24235
rect 33343 24172 33352 24212
rect 33392 24172 33409 24212
rect 33495 24172 33516 24212
rect 33556 24172 33577 24212
rect 33663 24172 33680 24212
rect 33720 24172 33729 24212
rect 33343 24149 33409 24172
rect 33495 24149 33577 24172
rect 33663 24149 33729 24172
rect 33343 24130 33729 24149
rect 48463 24235 48849 24254
rect 48463 24212 48529 24235
rect 48615 24212 48697 24235
rect 48783 24212 48849 24235
rect 48463 24172 48472 24212
rect 48512 24172 48529 24212
rect 48615 24172 48636 24212
rect 48676 24172 48697 24212
rect 48783 24172 48800 24212
rect 48840 24172 48849 24212
rect 48463 24149 48529 24172
rect 48615 24149 48697 24172
rect 48783 24149 48849 24172
rect 48463 24130 48849 24149
rect 63583 24235 63969 24254
rect 63583 24212 63649 24235
rect 63735 24212 63817 24235
rect 63903 24212 63969 24235
rect 63583 24172 63592 24212
rect 63632 24172 63649 24212
rect 63735 24172 63756 24212
rect 63796 24172 63817 24212
rect 63903 24172 63920 24212
rect 63960 24172 63969 24212
rect 63583 24149 63649 24172
rect 63735 24149 63817 24172
rect 63903 24149 63969 24172
rect 63583 24130 63969 24149
rect 78703 24235 79089 24254
rect 78703 24212 78769 24235
rect 78855 24212 78937 24235
rect 79023 24212 79089 24235
rect 78703 24172 78712 24212
rect 78752 24172 78769 24212
rect 78855 24172 78876 24212
rect 78916 24172 78937 24212
rect 79023 24172 79040 24212
rect 79080 24172 79089 24212
rect 78703 24149 78769 24172
rect 78855 24149 78937 24172
rect 79023 24149 79089 24172
rect 78703 24130 79089 24149
rect 93823 24235 94209 24254
rect 93823 24212 93889 24235
rect 93975 24212 94057 24235
rect 94143 24212 94209 24235
rect 93823 24172 93832 24212
rect 93872 24172 93889 24212
rect 93975 24172 93996 24212
rect 94036 24172 94057 24212
rect 94143 24172 94160 24212
rect 94200 24172 94209 24212
rect 93823 24149 93889 24172
rect 93975 24149 94057 24172
rect 94143 24149 94209 24172
rect 93823 24130 94209 24149
rect 4343 23479 4729 23498
rect 4343 23456 4409 23479
rect 4495 23456 4577 23479
rect 4663 23456 4729 23479
rect 4343 23416 4352 23456
rect 4392 23416 4409 23456
rect 4495 23416 4516 23456
rect 4556 23416 4577 23456
rect 4663 23416 4680 23456
rect 4720 23416 4729 23456
rect 4343 23393 4409 23416
rect 4495 23393 4577 23416
rect 4663 23393 4729 23416
rect 4343 23374 4729 23393
rect 19463 23479 19849 23498
rect 19463 23456 19529 23479
rect 19615 23456 19697 23479
rect 19783 23456 19849 23479
rect 19463 23416 19472 23456
rect 19512 23416 19529 23456
rect 19615 23416 19636 23456
rect 19676 23416 19697 23456
rect 19783 23416 19800 23456
rect 19840 23416 19849 23456
rect 19463 23393 19529 23416
rect 19615 23393 19697 23416
rect 19783 23393 19849 23416
rect 19463 23374 19849 23393
rect 34583 23479 34969 23498
rect 34583 23456 34649 23479
rect 34735 23456 34817 23479
rect 34903 23456 34969 23479
rect 34583 23416 34592 23456
rect 34632 23416 34649 23456
rect 34735 23416 34756 23456
rect 34796 23416 34817 23456
rect 34903 23416 34920 23456
rect 34960 23416 34969 23456
rect 34583 23393 34649 23416
rect 34735 23393 34817 23416
rect 34903 23393 34969 23416
rect 34583 23374 34969 23393
rect 49703 23479 50089 23498
rect 49703 23456 49769 23479
rect 49855 23456 49937 23479
rect 50023 23456 50089 23479
rect 49703 23416 49712 23456
rect 49752 23416 49769 23456
rect 49855 23416 49876 23456
rect 49916 23416 49937 23456
rect 50023 23416 50040 23456
rect 50080 23416 50089 23456
rect 49703 23393 49769 23416
rect 49855 23393 49937 23416
rect 50023 23393 50089 23416
rect 49703 23374 50089 23393
rect 64823 23479 65209 23498
rect 64823 23456 64889 23479
rect 64975 23456 65057 23479
rect 65143 23456 65209 23479
rect 64823 23416 64832 23456
rect 64872 23416 64889 23456
rect 64975 23416 64996 23456
rect 65036 23416 65057 23456
rect 65143 23416 65160 23456
rect 65200 23416 65209 23456
rect 64823 23393 64889 23416
rect 64975 23393 65057 23416
rect 65143 23393 65209 23416
rect 64823 23374 65209 23393
rect 79943 23479 80329 23498
rect 79943 23456 80009 23479
rect 80095 23456 80177 23479
rect 80263 23456 80329 23479
rect 79943 23416 79952 23456
rect 79992 23416 80009 23456
rect 80095 23416 80116 23456
rect 80156 23416 80177 23456
rect 80263 23416 80280 23456
rect 80320 23416 80329 23456
rect 79943 23393 80009 23416
rect 80095 23393 80177 23416
rect 80263 23393 80329 23416
rect 79943 23374 80329 23393
rect 95063 23479 95449 23498
rect 95063 23456 95129 23479
rect 95215 23456 95297 23479
rect 95383 23456 95449 23479
rect 95063 23416 95072 23456
rect 95112 23416 95129 23456
rect 95215 23416 95236 23456
rect 95276 23416 95297 23456
rect 95383 23416 95400 23456
rect 95440 23416 95449 23456
rect 95063 23393 95129 23416
rect 95215 23393 95297 23416
rect 95383 23393 95449 23416
rect 95063 23374 95449 23393
rect 3103 22723 3489 22742
rect 3103 22700 3169 22723
rect 3255 22700 3337 22723
rect 3423 22700 3489 22723
rect 3103 22660 3112 22700
rect 3152 22660 3169 22700
rect 3255 22660 3276 22700
rect 3316 22660 3337 22700
rect 3423 22660 3440 22700
rect 3480 22660 3489 22700
rect 3103 22637 3169 22660
rect 3255 22637 3337 22660
rect 3423 22637 3489 22660
rect 3103 22618 3489 22637
rect 18223 22723 18609 22742
rect 18223 22700 18289 22723
rect 18375 22700 18457 22723
rect 18543 22700 18609 22723
rect 18223 22660 18232 22700
rect 18272 22660 18289 22700
rect 18375 22660 18396 22700
rect 18436 22660 18457 22700
rect 18543 22660 18560 22700
rect 18600 22660 18609 22700
rect 18223 22637 18289 22660
rect 18375 22637 18457 22660
rect 18543 22637 18609 22660
rect 18223 22618 18609 22637
rect 33343 22723 33729 22742
rect 33343 22700 33409 22723
rect 33495 22700 33577 22723
rect 33663 22700 33729 22723
rect 33343 22660 33352 22700
rect 33392 22660 33409 22700
rect 33495 22660 33516 22700
rect 33556 22660 33577 22700
rect 33663 22660 33680 22700
rect 33720 22660 33729 22700
rect 33343 22637 33409 22660
rect 33495 22637 33577 22660
rect 33663 22637 33729 22660
rect 33343 22618 33729 22637
rect 48463 22723 48849 22742
rect 48463 22700 48529 22723
rect 48615 22700 48697 22723
rect 48783 22700 48849 22723
rect 48463 22660 48472 22700
rect 48512 22660 48529 22700
rect 48615 22660 48636 22700
rect 48676 22660 48697 22700
rect 48783 22660 48800 22700
rect 48840 22660 48849 22700
rect 48463 22637 48529 22660
rect 48615 22637 48697 22660
rect 48783 22637 48849 22660
rect 48463 22618 48849 22637
rect 63583 22723 63969 22742
rect 63583 22700 63649 22723
rect 63735 22700 63817 22723
rect 63903 22700 63969 22723
rect 63583 22660 63592 22700
rect 63632 22660 63649 22700
rect 63735 22660 63756 22700
rect 63796 22660 63817 22700
rect 63903 22660 63920 22700
rect 63960 22660 63969 22700
rect 63583 22637 63649 22660
rect 63735 22637 63817 22660
rect 63903 22637 63969 22660
rect 63583 22618 63969 22637
rect 78703 22723 79089 22742
rect 78703 22700 78769 22723
rect 78855 22700 78937 22723
rect 79023 22700 79089 22723
rect 78703 22660 78712 22700
rect 78752 22660 78769 22700
rect 78855 22660 78876 22700
rect 78916 22660 78937 22700
rect 79023 22660 79040 22700
rect 79080 22660 79089 22700
rect 78703 22637 78769 22660
rect 78855 22637 78937 22660
rect 79023 22637 79089 22660
rect 78703 22618 79089 22637
rect 93823 22723 94209 22742
rect 93823 22700 93889 22723
rect 93975 22700 94057 22723
rect 94143 22700 94209 22723
rect 93823 22660 93832 22700
rect 93872 22660 93889 22700
rect 93975 22660 93996 22700
rect 94036 22660 94057 22700
rect 94143 22660 94160 22700
rect 94200 22660 94209 22700
rect 93823 22637 93889 22660
rect 93975 22637 94057 22660
rect 94143 22637 94209 22660
rect 93823 22618 94209 22637
rect 4343 21967 4729 21986
rect 4343 21944 4409 21967
rect 4495 21944 4577 21967
rect 4663 21944 4729 21967
rect 4343 21904 4352 21944
rect 4392 21904 4409 21944
rect 4495 21904 4516 21944
rect 4556 21904 4577 21944
rect 4663 21904 4680 21944
rect 4720 21904 4729 21944
rect 4343 21881 4409 21904
rect 4495 21881 4577 21904
rect 4663 21881 4729 21904
rect 4343 21862 4729 21881
rect 19463 21967 19849 21986
rect 19463 21944 19529 21967
rect 19615 21944 19697 21967
rect 19783 21944 19849 21967
rect 19463 21904 19472 21944
rect 19512 21904 19529 21944
rect 19615 21904 19636 21944
rect 19676 21904 19697 21944
rect 19783 21904 19800 21944
rect 19840 21904 19849 21944
rect 19463 21881 19529 21904
rect 19615 21881 19697 21904
rect 19783 21881 19849 21904
rect 19463 21862 19849 21881
rect 34583 21967 34969 21986
rect 34583 21944 34649 21967
rect 34735 21944 34817 21967
rect 34903 21944 34969 21967
rect 34583 21904 34592 21944
rect 34632 21904 34649 21944
rect 34735 21904 34756 21944
rect 34796 21904 34817 21944
rect 34903 21904 34920 21944
rect 34960 21904 34969 21944
rect 34583 21881 34649 21904
rect 34735 21881 34817 21904
rect 34903 21881 34969 21904
rect 34583 21862 34969 21881
rect 49703 21967 50089 21986
rect 49703 21944 49769 21967
rect 49855 21944 49937 21967
rect 50023 21944 50089 21967
rect 49703 21904 49712 21944
rect 49752 21904 49769 21944
rect 49855 21904 49876 21944
rect 49916 21904 49937 21944
rect 50023 21904 50040 21944
rect 50080 21904 50089 21944
rect 49703 21881 49769 21904
rect 49855 21881 49937 21904
rect 50023 21881 50089 21904
rect 49703 21862 50089 21881
rect 64823 21967 65209 21986
rect 64823 21944 64889 21967
rect 64975 21944 65057 21967
rect 65143 21944 65209 21967
rect 64823 21904 64832 21944
rect 64872 21904 64889 21944
rect 64975 21904 64996 21944
rect 65036 21904 65057 21944
rect 65143 21904 65160 21944
rect 65200 21904 65209 21944
rect 64823 21881 64889 21904
rect 64975 21881 65057 21904
rect 65143 21881 65209 21904
rect 64823 21862 65209 21881
rect 79943 21967 80329 21986
rect 79943 21944 80009 21967
rect 80095 21944 80177 21967
rect 80263 21944 80329 21967
rect 79943 21904 79952 21944
rect 79992 21904 80009 21944
rect 80095 21904 80116 21944
rect 80156 21904 80177 21944
rect 80263 21904 80280 21944
rect 80320 21904 80329 21944
rect 79943 21881 80009 21904
rect 80095 21881 80177 21904
rect 80263 21881 80329 21904
rect 79943 21862 80329 21881
rect 95063 21967 95449 21986
rect 95063 21944 95129 21967
rect 95215 21944 95297 21967
rect 95383 21944 95449 21967
rect 95063 21904 95072 21944
rect 95112 21904 95129 21944
rect 95215 21904 95236 21944
rect 95276 21904 95297 21944
rect 95383 21904 95400 21944
rect 95440 21904 95449 21944
rect 95063 21881 95129 21904
rect 95215 21881 95297 21904
rect 95383 21881 95449 21904
rect 95063 21862 95449 21881
rect 3103 21211 3489 21230
rect 3103 21188 3169 21211
rect 3255 21188 3337 21211
rect 3423 21188 3489 21211
rect 3103 21148 3112 21188
rect 3152 21148 3169 21188
rect 3255 21148 3276 21188
rect 3316 21148 3337 21188
rect 3423 21148 3440 21188
rect 3480 21148 3489 21188
rect 3103 21125 3169 21148
rect 3255 21125 3337 21148
rect 3423 21125 3489 21148
rect 3103 21106 3489 21125
rect 18223 21211 18609 21230
rect 18223 21188 18289 21211
rect 18375 21188 18457 21211
rect 18543 21188 18609 21211
rect 18223 21148 18232 21188
rect 18272 21148 18289 21188
rect 18375 21148 18396 21188
rect 18436 21148 18457 21188
rect 18543 21148 18560 21188
rect 18600 21148 18609 21188
rect 18223 21125 18289 21148
rect 18375 21125 18457 21148
rect 18543 21125 18609 21148
rect 18223 21106 18609 21125
rect 33343 21211 33729 21230
rect 33343 21188 33409 21211
rect 33495 21188 33577 21211
rect 33663 21188 33729 21211
rect 33343 21148 33352 21188
rect 33392 21148 33409 21188
rect 33495 21148 33516 21188
rect 33556 21148 33577 21188
rect 33663 21148 33680 21188
rect 33720 21148 33729 21188
rect 33343 21125 33409 21148
rect 33495 21125 33577 21148
rect 33663 21125 33729 21148
rect 33343 21106 33729 21125
rect 48463 21211 48849 21230
rect 48463 21188 48529 21211
rect 48615 21188 48697 21211
rect 48783 21188 48849 21211
rect 48463 21148 48472 21188
rect 48512 21148 48529 21188
rect 48615 21148 48636 21188
rect 48676 21148 48697 21188
rect 48783 21148 48800 21188
rect 48840 21148 48849 21188
rect 48463 21125 48529 21148
rect 48615 21125 48697 21148
rect 48783 21125 48849 21148
rect 48463 21106 48849 21125
rect 63583 21211 63969 21230
rect 63583 21188 63649 21211
rect 63735 21188 63817 21211
rect 63903 21188 63969 21211
rect 63583 21148 63592 21188
rect 63632 21148 63649 21188
rect 63735 21148 63756 21188
rect 63796 21148 63817 21188
rect 63903 21148 63920 21188
rect 63960 21148 63969 21188
rect 63583 21125 63649 21148
rect 63735 21125 63817 21148
rect 63903 21125 63969 21148
rect 63583 21106 63969 21125
rect 78703 21211 79089 21230
rect 78703 21188 78769 21211
rect 78855 21188 78937 21211
rect 79023 21188 79089 21211
rect 78703 21148 78712 21188
rect 78752 21148 78769 21188
rect 78855 21148 78876 21188
rect 78916 21148 78937 21188
rect 79023 21148 79040 21188
rect 79080 21148 79089 21188
rect 78703 21125 78769 21148
rect 78855 21125 78937 21148
rect 79023 21125 79089 21148
rect 78703 21106 79089 21125
rect 93823 21211 94209 21230
rect 93823 21188 93889 21211
rect 93975 21188 94057 21211
rect 94143 21188 94209 21211
rect 93823 21148 93832 21188
rect 93872 21148 93889 21188
rect 93975 21148 93996 21188
rect 94036 21148 94057 21188
rect 94143 21148 94160 21188
rect 94200 21148 94209 21188
rect 93823 21125 93889 21148
rect 93975 21125 94057 21148
rect 94143 21125 94209 21148
rect 93823 21106 94209 21125
rect 4343 20455 4729 20474
rect 4343 20432 4409 20455
rect 4495 20432 4577 20455
rect 4663 20432 4729 20455
rect 4343 20392 4352 20432
rect 4392 20392 4409 20432
rect 4495 20392 4516 20432
rect 4556 20392 4577 20432
rect 4663 20392 4680 20432
rect 4720 20392 4729 20432
rect 4343 20369 4409 20392
rect 4495 20369 4577 20392
rect 4663 20369 4729 20392
rect 4343 20350 4729 20369
rect 19463 20455 19849 20474
rect 19463 20432 19529 20455
rect 19615 20432 19697 20455
rect 19783 20432 19849 20455
rect 19463 20392 19472 20432
rect 19512 20392 19529 20432
rect 19615 20392 19636 20432
rect 19676 20392 19697 20432
rect 19783 20392 19800 20432
rect 19840 20392 19849 20432
rect 19463 20369 19529 20392
rect 19615 20369 19697 20392
rect 19783 20369 19849 20392
rect 19463 20350 19849 20369
rect 34583 20455 34969 20474
rect 34583 20432 34649 20455
rect 34735 20432 34817 20455
rect 34903 20432 34969 20455
rect 34583 20392 34592 20432
rect 34632 20392 34649 20432
rect 34735 20392 34756 20432
rect 34796 20392 34817 20432
rect 34903 20392 34920 20432
rect 34960 20392 34969 20432
rect 34583 20369 34649 20392
rect 34735 20369 34817 20392
rect 34903 20369 34969 20392
rect 34583 20350 34969 20369
rect 49703 20455 50089 20474
rect 49703 20432 49769 20455
rect 49855 20432 49937 20455
rect 50023 20432 50089 20455
rect 49703 20392 49712 20432
rect 49752 20392 49769 20432
rect 49855 20392 49876 20432
rect 49916 20392 49937 20432
rect 50023 20392 50040 20432
rect 50080 20392 50089 20432
rect 49703 20369 49769 20392
rect 49855 20369 49937 20392
rect 50023 20369 50089 20392
rect 49703 20350 50089 20369
rect 64823 20455 65209 20474
rect 64823 20432 64889 20455
rect 64975 20432 65057 20455
rect 65143 20432 65209 20455
rect 64823 20392 64832 20432
rect 64872 20392 64889 20432
rect 64975 20392 64996 20432
rect 65036 20392 65057 20432
rect 65143 20392 65160 20432
rect 65200 20392 65209 20432
rect 64823 20369 64889 20392
rect 64975 20369 65057 20392
rect 65143 20369 65209 20392
rect 64823 20350 65209 20369
rect 79943 20455 80329 20474
rect 79943 20432 80009 20455
rect 80095 20432 80177 20455
rect 80263 20432 80329 20455
rect 79943 20392 79952 20432
rect 79992 20392 80009 20432
rect 80095 20392 80116 20432
rect 80156 20392 80177 20432
rect 80263 20392 80280 20432
rect 80320 20392 80329 20432
rect 79943 20369 80009 20392
rect 80095 20369 80177 20392
rect 80263 20369 80329 20392
rect 79943 20350 80329 20369
rect 95063 20455 95449 20474
rect 95063 20432 95129 20455
rect 95215 20432 95297 20455
rect 95383 20432 95449 20455
rect 95063 20392 95072 20432
rect 95112 20392 95129 20432
rect 95215 20392 95236 20432
rect 95276 20392 95297 20432
rect 95383 20392 95400 20432
rect 95440 20392 95449 20432
rect 95063 20369 95129 20392
rect 95215 20369 95297 20392
rect 95383 20369 95449 20392
rect 95063 20350 95449 20369
rect 3103 19699 3489 19718
rect 3103 19676 3169 19699
rect 3255 19676 3337 19699
rect 3423 19676 3489 19699
rect 3103 19636 3112 19676
rect 3152 19636 3169 19676
rect 3255 19636 3276 19676
rect 3316 19636 3337 19676
rect 3423 19636 3440 19676
rect 3480 19636 3489 19676
rect 3103 19613 3169 19636
rect 3255 19613 3337 19636
rect 3423 19613 3489 19636
rect 3103 19594 3489 19613
rect 18223 19699 18609 19718
rect 18223 19676 18289 19699
rect 18375 19676 18457 19699
rect 18543 19676 18609 19699
rect 18223 19636 18232 19676
rect 18272 19636 18289 19676
rect 18375 19636 18396 19676
rect 18436 19636 18457 19676
rect 18543 19636 18560 19676
rect 18600 19636 18609 19676
rect 18223 19613 18289 19636
rect 18375 19613 18457 19636
rect 18543 19613 18609 19636
rect 18223 19594 18609 19613
rect 33343 19699 33729 19718
rect 33343 19676 33409 19699
rect 33495 19676 33577 19699
rect 33663 19676 33729 19699
rect 33343 19636 33352 19676
rect 33392 19636 33409 19676
rect 33495 19636 33516 19676
rect 33556 19636 33577 19676
rect 33663 19636 33680 19676
rect 33720 19636 33729 19676
rect 33343 19613 33409 19636
rect 33495 19613 33577 19636
rect 33663 19613 33729 19636
rect 33343 19594 33729 19613
rect 48463 19699 48849 19718
rect 48463 19676 48529 19699
rect 48615 19676 48697 19699
rect 48783 19676 48849 19699
rect 48463 19636 48472 19676
rect 48512 19636 48529 19676
rect 48615 19636 48636 19676
rect 48676 19636 48697 19676
rect 48783 19636 48800 19676
rect 48840 19636 48849 19676
rect 48463 19613 48529 19636
rect 48615 19613 48697 19636
rect 48783 19613 48849 19636
rect 48463 19594 48849 19613
rect 63583 19699 63969 19718
rect 63583 19676 63649 19699
rect 63735 19676 63817 19699
rect 63903 19676 63969 19699
rect 63583 19636 63592 19676
rect 63632 19636 63649 19676
rect 63735 19636 63756 19676
rect 63796 19636 63817 19676
rect 63903 19636 63920 19676
rect 63960 19636 63969 19676
rect 63583 19613 63649 19636
rect 63735 19613 63817 19636
rect 63903 19613 63969 19636
rect 63583 19594 63969 19613
rect 78703 19699 79089 19718
rect 78703 19676 78769 19699
rect 78855 19676 78937 19699
rect 79023 19676 79089 19699
rect 78703 19636 78712 19676
rect 78752 19636 78769 19676
rect 78855 19636 78876 19676
rect 78916 19636 78937 19676
rect 79023 19636 79040 19676
rect 79080 19636 79089 19676
rect 78703 19613 78769 19636
rect 78855 19613 78937 19636
rect 79023 19613 79089 19636
rect 78703 19594 79089 19613
rect 93823 19699 94209 19718
rect 93823 19676 93889 19699
rect 93975 19676 94057 19699
rect 94143 19676 94209 19699
rect 93823 19636 93832 19676
rect 93872 19636 93889 19676
rect 93975 19636 93996 19676
rect 94036 19636 94057 19676
rect 94143 19636 94160 19676
rect 94200 19636 94209 19676
rect 93823 19613 93889 19636
rect 93975 19613 94057 19636
rect 94143 19613 94209 19636
rect 93823 19594 94209 19613
rect 4343 18943 4729 18962
rect 4343 18920 4409 18943
rect 4495 18920 4577 18943
rect 4663 18920 4729 18943
rect 4343 18880 4352 18920
rect 4392 18880 4409 18920
rect 4495 18880 4516 18920
rect 4556 18880 4577 18920
rect 4663 18880 4680 18920
rect 4720 18880 4729 18920
rect 4343 18857 4409 18880
rect 4495 18857 4577 18880
rect 4663 18857 4729 18880
rect 4343 18838 4729 18857
rect 19463 18943 19849 18962
rect 19463 18920 19529 18943
rect 19615 18920 19697 18943
rect 19783 18920 19849 18943
rect 19463 18880 19472 18920
rect 19512 18880 19529 18920
rect 19615 18880 19636 18920
rect 19676 18880 19697 18920
rect 19783 18880 19800 18920
rect 19840 18880 19849 18920
rect 19463 18857 19529 18880
rect 19615 18857 19697 18880
rect 19783 18857 19849 18880
rect 19463 18838 19849 18857
rect 34583 18943 34969 18962
rect 34583 18920 34649 18943
rect 34735 18920 34817 18943
rect 34903 18920 34969 18943
rect 34583 18880 34592 18920
rect 34632 18880 34649 18920
rect 34735 18880 34756 18920
rect 34796 18880 34817 18920
rect 34903 18880 34920 18920
rect 34960 18880 34969 18920
rect 34583 18857 34649 18880
rect 34735 18857 34817 18880
rect 34903 18857 34969 18880
rect 34583 18838 34969 18857
rect 49703 18943 50089 18962
rect 49703 18920 49769 18943
rect 49855 18920 49937 18943
rect 50023 18920 50089 18943
rect 49703 18880 49712 18920
rect 49752 18880 49769 18920
rect 49855 18880 49876 18920
rect 49916 18880 49937 18920
rect 50023 18880 50040 18920
rect 50080 18880 50089 18920
rect 49703 18857 49769 18880
rect 49855 18857 49937 18880
rect 50023 18857 50089 18880
rect 49703 18838 50089 18857
rect 64823 18943 65209 18962
rect 64823 18920 64889 18943
rect 64975 18920 65057 18943
rect 65143 18920 65209 18943
rect 64823 18880 64832 18920
rect 64872 18880 64889 18920
rect 64975 18880 64996 18920
rect 65036 18880 65057 18920
rect 65143 18880 65160 18920
rect 65200 18880 65209 18920
rect 64823 18857 64889 18880
rect 64975 18857 65057 18880
rect 65143 18857 65209 18880
rect 64823 18838 65209 18857
rect 79943 18943 80329 18962
rect 79943 18920 80009 18943
rect 80095 18920 80177 18943
rect 80263 18920 80329 18943
rect 79943 18880 79952 18920
rect 79992 18880 80009 18920
rect 80095 18880 80116 18920
rect 80156 18880 80177 18920
rect 80263 18880 80280 18920
rect 80320 18880 80329 18920
rect 79943 18857 80009 18880
rect 80095 18857 80177 18880
rect 80263 18857 80329 18880
rect 79943 18838 80329 18857
rect 95063 18943 95449 18962
rect 95063 18920 95129 18943
rect 95215 18920 95297 18943
rect 95383 18920 95449 18943
rect 95063 18880 95072 18920
rect 95112 18880 95129 18920
rect 95215 18880 95236 18920
rect 95276 18880 95297 18920
rect 95383 18880 95400 18920
rect 95440 18880 95449 18920
rect 95063 18857 95129 18880
rect 95215 18857 95297 18880
rect 95383 18857 95449 18880
rect 95063 18838 95449 18857
rect 3103 18187 3489 18206
rect 3103 18164 3169 18187
rect 3255 18164 3337 18187
rect 3423 18164 3489 18187
rect 3103 18124 3112 18164
rect 3152 18124 3169 18164
rect 3255 18124 3276 18164
rect 3316 18124 3337 18164
rect 3423 18124 3440 18164
rect 3480 18124 3489 18164
rect 3103 18101 3169 18124
rect 3255 18101 3337 18124
rect 3423 18101 3489 18124
rect 3103 18082 3489 18101
rect 18223 18187 18609 18206
rect 18223 18164 18289 18187
rect 18375 18164 18457 18187
rect 18543 18164 18609 18187
rect 18223 18124 18232 18164
rect 18272 18124 18289 18164
rect 18375 18124 18396 18164
rect 18436 18124 18457 18164
rect 18543 18124 18560 18164
rect 18600 18124 18609 18164
rect 18223 18101 18289 18124
rect 18375 18101 18457 18124
rect 18543 18101 18609 18124
rect 18223 18082 18609 18101
rect 33343 18187 33729 18206
rect 33343 18164 33409 18187
rect 33495 18164 33577 18187
rect 33663 18164 33729 18187
rect 33343 18124 33352 18164
rect 33392 18124 33409 18164
rect 33495 18124 33516 18164
rect 33556 18124 33577 18164
rect 33663 18124 33680 18164
rect 33720 18124 33729 18164
rect 33343 18101 33409 18124
rect 33495 18101 33577 18124
rect 33663 18101 33729 18124
rect 33343 18082 33729 18101
rect 48463 18187 48849 18206
rect 48463 18164 48529 18187
rect 48615 18164 48697 18187
rect 48783 18164 48849 18187
rect 48463 18124 48472 18164
rect 48512 18124 48529 18164
rect 48615 18124 48636 18164
rect 48676 18124 48697 18164
rect 48783 18124 48800 18164
rect 48840 18124 48849 18164
rect 48463 18101 48529 18124
rect 48615 18101 48697 18124
rect 48783 18101 48849 18124
rect 48463 18082 48849 18101
rect 63583 18187 63969 18206
rect 63583 18164 63649 18187
rect 63735 18164 63817 18187
rect 63903 18164 63969 18187
rect 63583 18124 63592 18164
rect 63632 18124 63649 18164
rect 63735 18124 63756 18164
rect 63796 18124 63817 18164
rect 63903 18124 63920 18164
rect 63960 18124 63969 18164
rect 63583 18101 63649 18124
rect 63735 18101 63817 18124
rect 63903 18101 63969 18124
rect 63583 18082 63969 18101
rect 78703 18187 79089 18206
rect 78703 18164 78769 18187
rect 78855 18164 78937 18187
rect 79023 18164 79089 18187
rect 78703 18124 78712 18164
rect 78752 18124 78769 18164
rect 78855 18124 78876 18164
rect 78916 18124 78937 18164
rect 79023 18124 79040 18164
rect 79080 18124 79089 18164
rect 78703 18101 78769 18124
rect 78855 18101 78937 18124
rect 79023 18101 79089 18124
rect 78703 18082 79089 18101
rect 93823 18187 94209 18206
rect 93823 18164 93889 18187
rect 93975 18164 94057 18187
rect 94143 18164 94209 18187
rect 93823 18124 93832 18164
rect 93872 18124 93889 18164
rect 93975 18124 93996 18164
rect 94036 18124 94057 18164
rect 94143 18124 94160 18164
rect 94200 18124 94209 18164
rect 93823 18101 93889 18124
rect 93975 18101 94057 18124
rect 94143 18101 94209 18124
rect 93823 18082 94209 18101
rect 4343 17431 4729 17450
rect 4343 17408 4409 17431
rect 4495 17408 4577 17431
rect 4663 17408 4729 17431
rect 4343 17368 4352 17408
rect 4392 17368 4409 17408
rect 4495 17368 4516 17408
rect 4556 17368 4577 17408
rect 4663 17368 4680 17408
rect 4720 17368 4729 17408
rect 4343 17345 4409 17368
rect 4495 17345 4577 17368
rect 4663 17345 4729 17368
rect 4343 17326 4729 17345
rect 19463 17431 19849 17450
rect 19463 17408 19529 17431
rect 19615 17408 19697 17431
rect 19783 17408 19849 17431
rect 19463 17368 19472 17408
rect 19512 17368 19529 17408
rect 19615 17368 19636 17408
rect 19676 17368 19697 17408
rect 19783 17368 19800 17408
rect 19840 17368 19849 17408
rect 19463 17345 19529 17368
rect 19615 17345 19697 17368
rect 19783 17345 19849 17368
rect 19463 17326 19849 17345
rect 34583 17431 34969 17450
rect 34583 17408 34649 17431
rect 34735 17408 34817 17431
rect 34903 17408 34969 17431
rect 34583 17368 34592 17408
rect 34632 17368 34649 17408
rect 34735 17368 34756 17408
rect 34796 17368 34817 17408
rect 34903 17368 34920 17408
rect 34960 17368 34969 17408
rect 34583 17345 34649 17368
rect 34735 17345 34817 17368
rect 34903 17345 34969 17368
rect 34583 17326 34969 17345
rect 49703 17431 50089 17450
rect 49703 17408 49769 17431
rect 49855 17408 49937 17431
rect 50023 17408 50089 17431
rect 49703 17368 49712 17408
rect 49752 17368 49769 17408
rect 49855 17368 49876 17408
rect 49916 17368 49937 17408
rect 50023 17368 50040 17408
rect 50080 17368 50089 17408
rect 49703 17345 49769 17368
rect 49855 17345 49937 17368
rect 50023 17345 50089 17368
rect 49703 17326 50089 17345
rect 64823 17431 65209 17450
rect 64823 17408 64889 17431
rect 64975 17408 65057 17431
rect 65143 17408 65209 17431
rect 64823 17368 64832 17408
rect 64872 17368 64889 17408
rect 64975 17368 64996 17408
rect 65036 17368 65057 17408
rect 65143 17368 65160 17408
rect 65200 17368 65209 17408
rect 64823 17345 64889 17368
rect 64975 17345 65057 17368
rect 65143 17345 65209 17368
rect 64823 17326 65209 17345
rect 79943 17431 80329 17450
rect 79943 17408 80009 17431
rect 80095 17408 80177 17431
rect 80263 17408 80329 17431
rect 79943 17368 79952 17408
rect 79992 17368 80009 17408
rect 80095 17368 80116 17408
rect 80156 17368 80177 17408
rect 80263 17368 80280 17408
rect 80320 17368 80329 17408
rect 79943 17345 80009 17368
rect 80095 17345 80177 17368
rect 80263 17345 80329 17368
rect 79943 17326 80329 17345
rect 95063 17431 95449 17450
rect 95063 17408 95129 17431
rect 95215 17408 95297 17431
rect 95383 17408 95449 17431
rect 95063 17368 95072 17408
rect 95112 17368 95129 17408
rect 95215 17368 95236 17408
rect 95276 17368 95297 17408
rect 95383 17368 95400 17408
rect 95440 17368 95449 17408
rect 95063 17345 95129 17368
rect 95215 17345 95297 17368
rect 95383 17345 95449 17368
rect 95063 17326 95449 17345
rect 3103 16675 3489 16694
rect 3103 16652 3169 16675
rect 3255 16652 3337 16675
rect 3423 16652 3489 16675
rect 3103 16612 3112 16652
rect 3152 16612 3169 16652
rect 3255 16612 3276 16652
rect 3316 16612 3337 16652
rect 3423 16612 3440 16652
rect 3480 16612 3489 16652
rect 3103 16589 3169 16612
rect 3255 16589 3337 16612
rect 3423 16589 3489 16612
rect 3103 16570 3489 16589
rect 18223 16675 18609 16694
rect 18223 16652 18289 16675
rect 18375 16652 18457 16675
rect 18543 16652 18609 16675
rect 18223 16612 18232 16652
rect 18272 16612 18289 16652
rect 18375 16612 18396 16652
rect 18436 16612 18457 16652
rect 18543 16612 18560 16652
rect 18600 16612 18609 16652
rect 18223 16589 18289 16612
rect 18375 16589 18457 16612
rect 18543 16589 18609 16612
rect 18223 16570 18609 16589
rect 33343 16675 33729 16694
rect 33343 16652 33409 16675
rect 33495 16652 33577 16675
rect 33663 16652 33729 16675
rect 33343 16612 33352 16652
rect 33392 16612 33409 16652
rect 33495 16612 33516 16652
rect 33556 16612 33577 16652
rect 33663 16612 33680 16652
rect 33720 16612 33729 16652
rect 33343 16589 33409 16612
rect 33495 16589 33577 16612
rect 33663 16589 33729 16612
rect 33343 16570 33729 16589
rect 48463 16675 48849 16694
rect 48463 16652 48529 16675
rect 48615 16652 48697 16675
rect 48783 16652 48849 16675
rect 48463 16612 48472 16652
rect 48512 16612 48529 16652
rect 48615 16612 48636 16652
rect 48676 16612 48697 16652
rect 48783 16612 48800 16652
rect 48840 16612 48849 16652
rect 48463 16589 48529 16612
rect 48615 16589 48697 16612
rect 48783 16589 48849 16612
rect 48463 16570 48849 16589
rect 63583 16675 63969 16694
rect 63583 16652 63649 16675
rect 63735 16652 63817 16675
rect 63903 16652 63969 16675
rect 63583 16612 63592 16652
rect 63632 16612 63649 16652
rect 63735 16612 63756 16652
rect 63796 16612 63817 16652
rect 63903 16612 63920 16652
rect 63960 16612 63969 16652
rect 63583 16589 63649 16612
rect 63735 16589 63817 16612
rect 63903 16589 63969 16612
rect 63583 16570 63969 16589
rect 78703 16675 79089 16694
rect 78703 16652 78769 16675
rect 78855 16652 78937 16675
rect 79023 16652 79089 16675
rect 78703 16612 78712 16652
rect 78752 16612 78769 16652
rect 78855 16612 78876 16652
rect 78916 16612 78937 16652
rect 79023 16612 79040 16652
rect 79080 16612 79089 16652
rect 78703 16589 78769 16612
rect 78855 16589 78937 16612
rect 79023 16589 79089 16612
rect 78703 16570 79089 16589
rect 93823 16675 94209 16694
rect 93823 16652 93889 16675
rect 93975 16652 94057 16675
rect 94143 16652 94209 16675
rect 93823 16612 93832 16652
rect 93872 16612 93889 16652
rect 93975 16612 93996 16652
rect 94036 16612 94057 16652
rect 94143 16612 94160 16652
rect 94200 16612 94209 16652
rect 93823 16589 93889 16612
rect 93975 16589 94057 16612
rect 94143 16589 94209 16612
rect 93823 16570 94209 16589
rect 4343 15919 4729 15938
rect 4343 15896 4409 15919
rect 4495 15896 4577 15919
rect 4663 15896 4729 15919
rect 4343 15856 4352 15896
rect 4392 15856 4409 15896
rect 4495 15856 4516 15896
rect 4556 15856 4577 15896
rect 4663 15856 4680 15896
rect 4720 15856 4729 15896
rect 4343 15833 4409 15856
rect 4495 15833 4577 15856
rect 4663 15833 4729 15856
rect 4343 15814 4729 15833
rect 19463 15919 19849 15938
rect 19463 15896 19529 15919
rect 19615 15896 19697 15919
rect 19783 15896 19849 15919
rect 19463 15856 19472 15896
rect 19512 15856 19529 15896
rect 19615 15856 19636 15896
rect 19676 15856 19697 15896
rect 19783 15856 19800 15896
rect 19840 15856 19849 15896
rect 19463 15833 19529 15856
rect 19615 15833 19697 15856
rect 19783 15833 19849 15856
rect 19463 15814 19849 15833
rect 34583 15919 34969 15938
rect 34583 15896 34649 15919
rect 34735 15896 34817 15919
rect 34903 15896 34969 15919
rect 34583 15856 34592 15896
rect 34632 15856 34649 15896
rect 34735 15856 34756 15896
rect 34796 15856 34817 15896
rect 34903 15856 34920 15896
rect 34960 15856 34969 15896
rect 34583 15833 34649 15856
rect 34735 15833 34817 15856
rect 34903 15833 34969 15856
rect 34583 15814 34969 15833
rect 49703 15919 50089 15938
rect 49703 15896 49769 15919
rect 49855 15896 49937 15919
rect 50023 15896 50089 15919
rect 49703 15856 49712 15896
rect 49752 15856 49769 15896
rect 49855 15856 49876 15896
rect 49916 15856 49937 15896
rect 50023 15856 50040 15896
rect 50080 15856 50089 15896
rect 49703 15833 49769 15856
rect 49855 15833 49937 15856
rect 50023 15833 50089 15856
rect 49703 15814 50089 15833
rect 64823 15919 65209 15938
rect 64823 15896 64889 15919
rect 64975 15896 65057 15919
rect 65143 15896 65209 15919
rect 64823 15856 64832 15896
rect 64872 15856 64889 15896
rect 64975 15856 64996 15896
rect 65036 15856 65057 15896
rect 65143 15856 65160 15896
rect 65200 15856 65209 15896
rect 64823 15833 64889 15856
rect 64975 15833 65057 15856
rect 65143 15833 65209 15856
rect 64823 15814 65209 15833
rect 79943 15919 80329 15938
rect 79943 15896 80009 15919
rect 80095 15896 80177 15919
rect 80263 15896 80329 15919
rect 79943 15856 79952 15896
rect 79992 15856 80009 15896
rect 80095 15856 80116 15896
rect 80156 15856 80177 15896
rect 80263 15856 80280 15896
rect 80320 15856 80329 15896
rect 79943 15833 80009 15856
rect 80095 15833 80177 15856
rect 80263 15833 80329 15856
rect 79943 15814 80329 15833
rect 95063 15919 95449 15938
rect 95063 15896 95129 15919
rect 95215 15896 95297 15919
rect 95383 15896 95449 15919
rect 95063 15856 95072 15896
rect 95112 15856 95129 15896
rect 95215 15856 95236 15896
rect 95276 15856 95297 15896
rect 95383 15856 95400 15896
rect 95440 15856 95449 15896
rect 95063 15833 95129 15856
rect 95215 15833 95297 15856
rect 95383 15833 95449 15856
rect 95063 15814 95449 15833
rect 3103 15163 3489 15182
rect 3103 15140 3169 15163
rect 3255 15140 3337 15163
rect 3423 15140 3489 15163
rect 3103 15100 3112 15140
rect 3152 15100 3169 15140
rect 3255 15100 3276 15140
rect 3316 15100 3337 15140
rect 3423 15100 3440 15140
rect 3480 15100 3489 15140
rect 3103 15077 3169 15100
rect 3255 15077 3337 15100
rect 3423 15077 3489 15100
rect 3103 15058 3489 15077
rect 18223 15163 18609 15182
rect 18223 15140 18289 15163
rect 18375 15140 18457 15163
rect 18543 15140 18609 15163
rect 18223 15100 18232 15140
rect 18272 15100 18289 15140
rect 18375 15100 18396 15140
rect 18436 15100 18457 15140
rect 18543 15100 18560 15140
rect 18600 15100 18609 15140
rect 18223 15077 18289 15100
rect 18375 15077 18457 15100
rect 18543 15077 18609 15100
rect 18223 15058 18609 15077
rect 33343 15163 33729 15182
rect 33343 15140 33409 15163
rect 33495 15140 33577 15163
rect 33663 15140 33729 15163
rect 33343 15100 33352 15140
rect 33392 15100 33409 15140
rect 33495 15100 33516 15140
rect 33556 15100 33577 15140
rect 33663 15100 33680 15140
rect 33720 15100 33729 15140
rect 33343 15077 33409 15100
rect 33495 15077 33577 15100
rect 33663 15077 33729 15100
rect 33343 15058 33729 15077
rect 48463 15163 48849 15182
rect 48463 15140 48529 15163
rect 48615 15140 48697 15163
rect 48783 15140 48849 15163
rect 48463 15100 48472 15140
rect 48512 15100 48529 15140
rect 48615 15100 48636 15140
rect 48676 15100 48697 15140
rect 48783 15100 48800 15140
rect 48840 15100 48849 15140
rect 48463 15077 48529 15100
rect 48615 15077 48697 15100
rect 48783 15077 48849 15100
rect 48463 15058 48849 15077
rect 63583 15163 63969 15182
rect 63583 15140 63649 15163
rect 63735 15140 63817 15163
rect 63903 15140 63969 15163
rect 63583 15100 63592 15140
rect 63632 15100 63649 15140
rect 63735 15100 63756 15140
rect 63796 15100 63817 15140
rect 63903 15100 63920 15140
rect 63960 15100 63969 15140
rect 63583 15077 63649 15100
rect 63735 15077 63817 15100
rect 63903 15077 63969 15100
rect 63583 15058 63969 15077
rect 78703 15163 79089 15182
rect 78703 15140 78769 15163
rect 78855 15140 78937 15163
rect 79023 15140 79089 15163
rect 78703 15100 78712 15140
rect 78752 15100 78769 15140
rect 78855 15100 78876 15140
rect 78916 15100 78937 15140
rect 79023 15100 79040 15140
rect 79080 15100 79089 15140
rect 78703 15077 78769 15100
rect 78855 15077 78937 15100
rect 79023 15077 79089 15100
rect 78703 15058 79089 15077
rect 93823 15163 94209 15182
rect 93823 15140 93889 15163
rect 93975 15140 94057 15163
rect 94143 15140 94209 15163
rect 93823 15100 93832 15140
rect 93872 15100 93889 15140
rect 93975 15100 93996 15140
rect 94036 15100 94057 15140
rect 94143 15100 94160 15140
rect 94200 15100 94209 15140
rect 93823 15077 93889 15100
rect 93975 15077 94057 15100
rect 94143 15077 94209 15100
rect 93823 15058 94209 15077
rect 4343 14407 4729 14426
rect 4343 14384 4409 14407
rect 4495 14384 4577 14407
rect 4663 14384 4729 14407
rect 4343 14344 4352 14384
rect 4392 14344 4409 14384
rect 4495 14344 4516 14384
rect 4556 14344 4577 14384
rect 4663 14344 4680 14384
rect 4720 14344 4729 14384
rect 4343 14321 4409 14344
rect 4495 14321 4577 14344
rect 4663 14321 4729 14344
rect 4343 14302 4729 14321
rect 19463 14407 19849 14426
rect 19463 14384 19529 14407
rect 19615 14384 19697 14407
rect 19783 14384 19849 14407
rect 19463 14344 19472 14384
rect 19512 14344 19529 14384
rect 19615 14344 19636 14384
rect 19676 14344 19697 14384
rect 19783 14344 19800 14384
rect 19840 14344 19849 14384
rect 19463 14321 19529 14344
rect 19615 14321 19697 14344
rect 19783 14321 19849 14344
rect 19463 14302 19849 14321
rect 34583 14407 34969 14426
rect 34583 14384 34649 14407
rect 34735 14384 34817 14407
rect 34903 14384 34969 14407
rect 34583 14344 34592 14384
rect 34632 14344 34649 14384
rect 34735 14344 34756 14384
rect 34796 14344 34817 14384
rect 34903 14344 34920 14384
rect 34960 14344 34969 14384
rect 34583 14321 34649 14344
rect 34735 14321 34817 14344
rect 34903 14321 34969 14344
rect 34583 14302 34969 14321
rect 49703 14407 50089 14426
rect 49703 14384 49769 14407
rect 49855 14384 49937 14407
rect 50023 14384 50089 14407
rect 49703 14344 49712 14384
rect 49752 14344 49769 14384
rect 49855 14344 49876 14384
rect 49916 14344 49937 14384
rect 50023 14344 50040 14384
rect 50080 14344 50089 14384
rect 49703 14321 49769 14344
rect 49855 14321 49937 14344
rect 50023 14321 50089 14344
rect 49703 14302 50089 14321
rect 64823 14407 65209 14426
rect 64823 14384 64889 14407
rect 64975 14384 65057 14407
rect 65143 14384 65209 14407
rect 64823 14344 64832 14384
rect 64872 14344 64889 14384
rect 64975 14344 64996 14384
rect 65036 14344 65057 14384
rect 65143 14344 65160 14384
rect 65200 14344 65209 14384
rect 64823 14321 64889 14344
rect 64975 14321 65057 14344
rect 65143 14321 65209 14344
rect 64823 14302 65209 14321
rect 79943 14407 80329 14426
rect 79943 14384 80009 14407
rect 80095 14384 80177 14407
rect 80263 14384 80329 14407
rect 79943 14344 79952 14384
rect 79992 14344 80009 14384
rect 80095 14344 80116 14384
rect 80156 14344 80177 14384
rect 80263 14344 80280 14384
rect 80320 14344 80329 14384
rect 79943 14321 80009 14344
rect 80095 14321 80177 14344
rect 80263 14321 80329 14344
rect 79943 14302 80329 14321
rect 95063 14407 95449 14426
rect 95063 14384 95129 14407
rect 95215 14384 95297 14407
rect 95383 14384 95449 14407
rect 95063 14344 95072 14384
rect 95112 14344 95129 14384
rect 95215 14344 95236 14384
rect 95276 14344 95297 14384
rect 95383 14344 95400 14384
rect 95440 14344 95449 14384
rect 95063 14321 95129 14344
rect 95215 14321 95297 14344
rect 95383 14321 95449 14344
rect 95063 14302 95449 14321
rect 3103 13651 3489 13670
rect 3103 13628 3169 13651
rect 3255 13628 3337 13651
rect 3423 13628 3489 13651
rect 3103 13588 3112 13628
rect 3152 13588 3169 13628
rect 3255 13588 3276 13628
rect 3316 13588 3337 13628
rect 3423 13588 3440 13628
rect 3480 13588 3489 13628
rect 3103 13565 3169 13588
rect 3255 13565 3337 13588
rect 3423 13565 3489 13588
rect 3103 13546 3489 13565
rect 18223 13651 18609 13670
rect 18223 13628 18289 13651
rect 18375 13628 18457 13651
rect 18543 13628 18609 13651
rect 18223 13588 18232 13628
rect 18272 13588 18289 13628
rect 18375 13588 18396 13628
rect 18436 13588 18457 13628
rect 18543 13588 18560 13628
rect 18600 13588 18609 13628
rect 18223 13565 18289 13588
rect 18375 13565 18457 13588
rect 18543 13565 18609 13588
rect 18223 13546 18609 13565
rect 33343 13651 33729 13670
rect 33343 13628 33409 13651
rect 33495 13628 33577 13651
rect 33663 13628 33729 13651
rect 33343 13588 33352 13628
rect 33392 13588 33409 13628
rect 33495 13588 33516 13628
rect 33556 13588 33577 13628
rect 33663 13588 33680 13628
rect 33720 13588 33729 13628
rect 33343 13565 33409 13588
rect 33495 13565 33577 13588
rect 33663 13565 33729 13588
rect 33343 13546 33729 13565
rect 48463 13651 48849 13670
rect 48463 13628 48529 13651
rect 48615 13628 48697 13651
rect 48783 13628 48849 13651
rect 48463 13588 48472 13628
rect 48512 13588 48529 13628
rect 48615 13588 48636 13628
rect 48676 13588 48697 13628
rect 48783 13588 48800 13628
rect 48840 13588 48849 13628
rect 48463 13565 48529 13588
rect 48615 13565 48697 13588
rect 48783 13565 48849 13588
rect 48463 13546 48849 13565
rect 63583 13651 63969 13670
rect 63583 13628 63649 13651
rect 63735 13628 63817 13651
rect 63903 13628 63969 13651
rect 63583 13588 63592 13628
rect 63632 13588 63649 13628
rect 63735 13588 63756 13628
rect 63796 13588 63817 13628
rect 63903 13588 63920 13628
rect 63960 13588 63969 13628
rect 63583 13565 63649 13588
rect 63735 13565 63817 13588
rect 63903 13565 63969 13588
rect 63583 13546 63969 13565
rect 78703 13651 79089 13670
rect 78703 13628 78769 13651
rect 78855 13628 78937 13651
rect 79023 13628 79089 13651
rect 78703 13588 78712 13628
rect 78752 13588 78769 13628
rect 78855 13588 78876 13628
rect 78916 13588 78937 13628
rect 79023 13588 79040 13628
rect 79080 13588 79089 13628
rect 78703 13565 78769 13588
rect 78855 13565 78937 13588
rect 79023 13565 79089 13588
rect 78703 13546 79089 13565
rect 93823 13651 94209 13670
rect 93823 13628 93889 13651
rect 93975 13628 94057 13651
rect 94143 13628 94209 13651
rect 93823 13588 93832 13628
rect 93872 13588 93889 13628
rect 93975 13588 93996 13628
rect 94036 13588 94057 13628
rect 94143 13588 94160 13628
rect 94200 13588 94209 13628
rect 93823 13565 93889 13588
rect 93975 13565 94057 13588
rect 94143 13565 94209 13588
rect 93823 13546 94209 13565
rect 4343 12895 4729 12914
rect 4343 12872 4409 12895
rect 4495 12872 4577 12895
rect 4663 12872 4729 12895
rect 4343 12832 4352 12872
rect 4392 12832 4409 12872
rect 4495 12832 4516 12872
rect 4556 12832 4577 12872
rect 4663 12832 4680 12872
rect 4720 12832 4729 12872
rect 4343 12809 4409 12832
rect 4495 12809 4577 12832
rect 4663 12809 4729 12832
rect 4343 12790 4729 12809
rect 19463 12895 19849 12914
rect 19463 12872 19529 12895
rect 19615 12872 19697 12895
rect 19783 12872 19849 12895
rect 19463 12832 19472 12872
rect 19512 12832 19529 12872
rect 19615 12832 19636 12872
rect 19676 12832 19697 12872
rect 19783 12832 19800 12872
rect 19840 12832 19849 12872
rect 19463 12809 19529 12832
rect 19615 12809 19697 12832
rect 19783 12809 19849 12832
rect 19463 12790 19849 12809
rect 34583 12895 34969 12914
rect 34583 12872 34649 12895
rect 34735 12872 34817 12895
rect 34903 12872 34969 12895
rect 34583 12832 34592 12872
rect 34632 12832 34649 12872
rect 34735 12832 34756 12872
rect 34796 12832 34817 12872
rect 34903 12832 34920 12872
rect 34960 12832 34969 12872
rect 34583 12809 34649 12832
rect 34735 12809 34817 12832
rect 34903 12809 34969 12832
rect 34583 12790 34969 12809
rect 49703 12895 50089 12914
rect 49703 12872 49769 12895
rect 49855 12872 49937 12895
rect 50023 12872 50089 12895
rect 49703 12832 49712 12872
rect 49752 12832 49769 12872
rect 49855 12832 49876 12872
rect 49916 12832 49937 12872
rect 50023 12832 50040 12872
rect 50080 12832 50089 12872
rect 49703 12809 49769 12832
rect 49855 12809 49937 12832
rect 50023 12809 50089 12832
rect 49703 12790 50089 12809
rect 64823 12895 65209 12914
rect 64823 12872 64889 12895
rect 64975 12872 65057 12895
rect 65143 12872 65209 12895
rect 64823 12832 64832 12872
rect 64872 12832 64889 12872
rect 64975 12832 64996 12872
rect 65036 12832 65057 12872
rect 65143 12832 65160 12872
rect 65200 12832 65209 12872
rect 64823 12809 64889 12832
rect 64975 12809 65057 12832
rect 65143 12809 65209 12832
rect 64823 12790 65209 12809
rect 79943 12895 80329 12914
rect 79943 12872 80009 12895
rect 80095 12872 80177 12895
rect 80263 12872 80329 12895
rect 79943 12832 79952 12872
rect 79992 12832 80009 12872
rect 80095 12832 80116 12872
rect 80156 12832 80177 12872
rect 80263 12832 80280 12872
rect 80320 12832 80329 12872
rect 79943 12809 80009 12832
rect 80095 12809 80177 12832
rect 80263 12809 80329 12832
rect 79943 12790 80329 12809
rect 95063 12895 95449 12914
rect 95063 12872 95129 12895
rect 95215 12872 95297 12895
rect 95383 12872 95449 12895
rect 95063 12832 95072 12872
rect 95112 12832 95129 12872
rect 95215 12832 95236 12872
rect 95276 12832 95297 12872
rect 95383 12832 95400 12872
rect 95440 12832 95449 12872
rect 95063 12809 95129 12832
rect 95215 12809 95297 12832
rect 95383 12809 95449 12832
rect 95063 12790 95449 12809
rect 3103 12139 3489 12158
rect 3103 12116 3169 12139
rect 3255 12116 3337 12139
rect 3423 12116 3489 12139
rect 3103 12076 3112 12116
rect 3152 12076 3169 12116
rect 3255 12076 3276 12116
rect 3316 12076 3337 12116
rect 3423 12076 3440 12116
rect 3480 12076 3489 12116
rect 3103 12053 3169 12076
rect 3255 12053 3337 12076
rect 3423 12053 3489 12076
rect 3103 12034 3489 12053
rect 18223 12139 18609 12158
rect 18223 12116 18289 12139
rect 18375 12116 18457 12139
rect 18543 12116 18609 12139
rect 18223 12076 18232 12116
rect 18272 12076 18289 12116
rect 18375 12076 18396 12116
rect 18436 12076 18457 12116
rect 18543 12076 18560 12116
rect 18600 12076 18609 12116
rect 18223 12053 18289 12076
rect 18375 12053 18457 12076
rect 18543 12053 18609 12076
rect 18223 12034 18609 12053
rect 33343 12139 33729 12158
rect 33343 12116 33409 12139
rect 33495 12116 33577 12139
rect 33663 12116 33729 12139
rect 33343 12076 33352 12116
rect 33392 12076 33409 12116
rect 33495 12076 33516 12116
rect 33556 12076 33577 12116
rect 33663 12076 33680 12116
rect 33720 12076 33729 12116
rect 33343 12053 33409 12076
rect 33495 12053 33577 12076
rect 33663 12053 33729 12076
rect 33343 12034 33729 12053
rect 48463 12139 48849 12158
rect 48463 12116 48529 12139
rect 48615 12116 48697 12139
rect 48783 12116 48849 12139
rect 48463 12076 48472 12116
rect 48512 12076 48529 12116
rect 48615 12076 48636 12116
rect 48676 12076 48697 12116
rect 48783 12076 48800 12116
rect 48840 12076 48849 12116
rect 48463 12053 48529 12076
rect 48615 12053 48697 12076
rect 48783 12053 48849 12076
rect 48463 12034 48849 12053
rect 63583 12139 63969 12158
rect 63583 12116 63649 12139
rect 63735 12116 63817 12139
rect 63903 12116 63969 12139
rect 63583 12076 63592 12116
rect 63632 12076 63649 12116
rect 63735 12076 63756 12116
rect 63796 12076 63817 12116
rect 63903 12076 63920 12116
rect 63960 12076 63969 12116
rect 63583 12053 63649 12076
rect 63735 12053 63817 12076
rect 63903 12053 63969 12076
rect 63583 12034 63969 12053
rect 78703 12139 79089 12158
rect 78703 12116 78769 12139
rect 78855 12116 78937 12139
rect 79023 12116 79089 12139
rect 78703 12076 78712 12116
rect 78752 12076 78769 12116
rect 78855 12076 78876 12116
rect 78916 12076 78937 12116
rect 79023 12076 79040 12116
rect 79080 12076 79089 12116
rect 78703 12053 78769 12076
rect 78855 12053 78937 12076
rect 79023 12053 79089 12076
rect 78703 12034 79089 12053
rect 93823 12139 94209 12158
rect 93823 12116 93889 12139
rect 93975 12116 94057 12139
rect 94143 12116 94209 12139
rect 93823 12076 93832 12116
rect 93872 12076 93889 12116
rect 93975 12076 93996 12116
rect 94036 12076 94057 12116
rect 94143 12076 94160 12116
rect 94200 12076 94209 12116
rect 93823 12053 93889 12076
rect 93975 12053 94057 12076
rect 94143 12053 94209 12076
rect 93823 12034 94209 12053
rect 4343 11383 4729 11402
rect 4343 11360 4409 11383
rect 4495 11360 4577 11383
rect 4663 11360 4729 11383
rect 4343 11320 4352 11360
rect 4392 11320 4409 11360
rect 4495 11320 4516 11360
rect 4556 11320 4577 11360
rect 4663 11320 4680 11360
rect 4720 11320 4729 11360
rect 4343 11297 4409 11320
rect 4495 11297 4577 11320
rect 4663 11297 4729 11320
rect 4343 11278 4729 11297
rect 19463 11383 19849 11402
rect 19463 11360 19529 11383
rect 19615 11360 19697 11383
rect 19783 11360 19849 11383
rect 19463 11320 19472 11360
rect 19512 11320 19529 11360
rect 19615 11320 19636 11360
rect 19676 11320 19697 11360
rect 19783 11320 19800 11360
rect 19840 11320 19849 11360
rect 19463 11297 19529 11320
rect 19615 11297 19697 11320
rect 19783 11297 19849 11320
rect 19463 11278 19849 11297
rect 34583 11383 34969 11402
rect 34583 11360 34649 11383
rect 34735 11360 34817 11383
rect 34903 11360 34969 11383
rect 34583 11320 34592 11360
rect 34632 11320 34649 11360
rect 34735 11320 34756 11360
rect 34796 11320 34817 11360
rect 34903 11320 34920 11360
rect 34960 11320 34969 11360
rect 34583 11297 34649 11320
rect 34735 11297 34817 11320
rect 34903 11297 34969 11320
rect 34583 11278 34969 11297
rect 49703 11383 50089 11402
rect 49703 11360 49769 11383
rect 49855 11360 49937 11383
rect 50023 11360 50089 11383
rect 49703 11320 49712 11360
rect 49752 11320 49769 11360
rect 49855 11320 49876 11360
rect 49916 11320 49937 11360
rect 50023 11320 50040 11360
rect 50080 11320 50089 11360
rect 49703 11297 49769 11320
rect 49855 11297 49937 11320
rect 50023 11297 50089 11320
rect 49703 11278 50089 11297
rect 64823 11383 65209 11402
rect 64823 11360 64889 11383
rect 64975 11360 65057 11383
rect 65143 11360 65209 11383
rect 64823 11320 64832 11360
rect 64872 11320 64889 11360
rect 64975 11320 64996 11360
rect 65036 11320 65057 11360
rect 65143 11320 65160 11360
rect 65200 11320 65209 11360
rect 64823 11297 64889 11320
rect 64975 11297 65057 11320
rect 65143 11297 65209 11320
rect 64823 11278 65209 11297
rect 79943 11383 80329 11402
rect 79943 11360 80009 11383
rect 80095 11360 80177 11383
rect 80263 11360 80329 11383
rect 79943 11320 79952 11360
rect 79992 11320 80009 11360
rect 80095 11320 80116 11360
rect 80156 11320 80177 11360
rect 80263 11320 80280 11360
rect 80320 11320 80329 11360
rect 79943 11297 80009 11320
rect 80095 11297 80177 11320
rect 80263 11297 80329 11320
rect 79943 11278 80329 11297
rect 95063 11383 95449 11402
rect 95063 11360 95129 11383
rect 95215 11360 95297 11383
rect 95383 11360 95449 11383
rect 95063 11320 95072 11360
rect 95112 11320 95129 11360
rect 95215 11320 95236 11360
rect 95276 11320 95297 11360
rect 95383 11320 95400 11360
rect 95440 11320 95449 11360
rect 95063 11297 95129 11320
rect 95215 11297 95297 11320
rect 95383 11297 95449 11320
rect 95063 11278 95449 11297
rect 3103 10627 3489 10646
rect 3103 10604 3169 10627
rect 3255 10604 3337 10627
rect 3423 10604 3489 10627
rect 3103 10564 3112 10604
rect 3152 10564 3169 10604
rect 3255 10564 3276 10604
rect 3316 10564 3337 10604
rect 3423 10564 3440 10604
rect 3480 10564 3489 10604
rect 3103 10541 3169 10564
rect 3255 10541 3337 10564
rect 3423 10541 3489 10564
rect 3103 10522 3489 10541
rect 18223 10627 18609 10646
rect 18223 10604 18289 10627
rect 18375 10604 18457 10627
rect 18543 10604 18609 10627
rect 18223 10564 18232 10604
rect 18272 10564 18289 10604
rect 18375 10564 18396 10604
rect 18436 10564 18457 10604
rect 18543 10564 18560 10604
rect 18600 10564 18609 10604
rect 18223 10541 18289 10564
rect 18375 10541 18457 10564
rect 18543 10541 18609 10564
rect 18223 10522 18609 10541
rect 33343 10627 33729 10646
rect 33343 10604 33409 10627
rect 33495 10604 33577 10627
rect 33663 10604 33729 10627
rect 33343 10564 33352 10604
rect 33392 10564 33409 10604
rect 33495 10564 33516 10604
rect 33556 10564 33577 10604
rect 33663 10564 33680 10604
rect 33720 10564 33729 10604
rect 33343 10541 33409 10564
rect 33495 10541 33577 10564
rect 33663 10541 33729 10564
rect 33343 10522 33729 10541
rect 48463 10627 48849 10646
rect 48463 10604 48529 10627
rect 48615 10604 48697 10627
rect 48783 10604 48849 10627
rect 48463 10564 48472 10604
rect 48512 10564 48529 10604
rect 48615 10564 48636 10604
rect 48676 10564 48697 10604
rect 48783 10564 48800 10604
rect 48840 10564 48849 10604
rect 48463 10541 48529 10564
rect 48615 10541 48697 10564
rect 48783 10541 48849 10564
rect 48463 10522 48849 10541
rect 63583 10627 63969 10646
rect 63583 10604 63649 10627
rect 63735 10604 63817 10627
rect 63903 10604 63969 10627
rect 63583 10564 63592 10604
rect 63632 10564 63649 10604
rect 63735 10564 63756 10604
rect 63796 10564 63817 10604
rect 63903 10564 63920 10604
rect 63960 10564 63969 10604
rect 63583 10541 63649 10564
rect 63735 10541 63817 10564
rect 63903 10541 63969 10564
rect 63583 10522 63969 10541
rect 78703 10627 79089 10646
rect 78703 10604 78769 10627
rect 78855 10604 78937 10627
rect 79023 10604 79089 10627
rect 78703 10564 78712 10604
rect 78752 10564 78769 10604
rect 78855 10564 78876 10604
rect 78916 10564 78937 10604
rect 79023 10564 79040 10604
rect 79080 10564 79089 10604
rect 78703 10541 78769 10564
rect 78855 10541 78937 10564
rect 79023 10541 79089 10564
rect 78703 10522 79089 10541
rect 93823 10627 94209 10646
rect 93823 10604 93889 10627
rect 93975 10604 94057 10627
rect 94143 10604 94209 10627
rect 93823 10564 93832 10604
rect 93872 10564 93889 10604
rect 93975 10564 93996 10604
rect 94036 10564 94057 10604
rect 94143 10564 94160 10604
rect 94200 10564 94209 10604
rect 93823 10541 93889 10564
rect 93975 10541 94057 10564
rect 94143 10541 94209 10564
rect 93823 10522 94209 10541
rect 4343 9871 4729 9890
rect 4343 9848 4409 9871
rect 4495 9848 4577 9871
rect 4663 9848 4729 9871
rect 4343 9808 4352 9848
rect 4392 9808 4409 9848
rect 4495 9808 4516 9848
rect 4556 9808 4577 9848
rect 4663 9808 4680 9848
rect 4720 9808 4729 9848
rect 4343 9785 4409 9808
rect 4495 9785 4577 9808
rect 4663 9785 4729 9808
rect 4343 9766 4729 9785
rect 19463 9871 19849 9890
rect 19463 9848 19529 9871
rect 19615 9848 19697 9871
rect 19783 9848 19849 9871
rect 19463 9808 19472 9848
rect 19512 9808 19529 9848
rect 19615 9808 19636 9848
rect 19676 9808 19697 9848
rect 19783 9808 19800 9848
rect 19840 9808 19849 9848
rect 19463 9785 19529 9808
rect 19615 9785 19697 9808
rect 19783 9785 19849 9808
rect 19463 9766 19849 9785
rect 34583 9871 34969 9890
rect 34583 9848 34649 9871
rect 34735 9848 34817 9871
rect 34903 9848 34969 9871
rect 34583 9808 34592 9848
rect 34632 9808 34649 9848
rect 34735 9808 34756 9848
rect 34796 9808 34817 9848
rect 34903 9808 34920 9848
rect 34960 9808 34969 9848
rect 34583 9785 34649 9808
rect 34735 9785 34817 9808
rect 34903 9785 34969 9808
rect 34583 9766 34969 9785
rect 49703 9871 50089 9890
rect 49703 9848 49769 9871
rect 49855 9848 49937 9871
rect 50023 9848 50089 9871
rect 49703 9808 49712 9848
rect 49752 9808 49769 9848
rect 49855 9808 49876 9848
rect 49916 9808 49937 9848
rect 50023 9808 50040 9848
rect 50080 9808 50089 9848
rect 49703 9785 49769 9808
rect 49855 9785 49937 9808
rect 50023 9785 50089 9808
rect 49703 9766 50089 9785
rect 64823 9871 65209 9890
rect 64823 9848 64889 9871
rect 64975 9848 65057 9871
rect 65143 9848 65209 9871
rect 64823 9808 64832 9848
rect 64872 9808 64889 9848
rect 64975 9808 64996 9848
rect 65036 9808 65057 9848
rect 65143 9808 65160 9848
rect 65200 9808 65209 9848
rect 64823 9785 64889 9808
rect 64975 9785 65057 9808
rect 65143 9785 65209 9808
rect 64823 9766 65209 9785
rect 79943 9871 80329 9890
rect 79943 9848 80009 9871
rect 80095 9848 80177 9871
rect 80263 9848 80329 9871
rect 79943 9808 79952 9848
rect 79992 9808 80009 9848
rect 80095 9808 80116 9848
rect 80156 9808 80177 9848
rect 80263 9808 80280 9848
rect 80320 9808 80329 9848
rect 79943 9785 80009 9808
rect 80095 9785 80177 9808
rect 80263 9785 80329 9808
rect 79943 9766 80329 9785
rect 95063 9871 95449 9890
rect 95063 9848 95129 9871
rect 95215 9848 95297 9871
rect 95383 9848 95449 9871
rect 95063 9808 95072 9848
rect 95112 9808 95129 9848
rect 95215 9808 95236 9848
rect 95276 9808 95297 9848
rect 95383 9808 95400 9848
rect 95440 9808 95449 9848
rect 95063 9785 95129 9808
rect 95215 9785 95297 9808
rect 95383 9785 95449 9808
rect 95063 9766 95449 9785
rect 3103 9115 3489 9134
rect 3103 9092 3169 9115
rect 3255 9092 3337 9115
rect 3423 9092 3489 9115
rect 3103 9052 3112 9092
rect 3152 9052 3169 9092
rect 3255 9052 3276 9092
rect 3316 9052 3337 9092
rect 3423 9052 3440 9092
rect 3480 9052 3489 9092
rect 3103 9029 3169 9052
rect 3255 9029 3337 9052
rect 3423 9029 3489 9052
rect 3103 9010 3489 9029
rect 18223 9115 18609 9134
rect 18223 9092 18289 9115
rect 18375 9092 18457 9115
rect 18543 9092 18609 9115
rect 18223 9052 18232 9092
rect 18272 9052 18289 9092
rect 18375 9052 18396 9092
rect 18436 9052 18457 9092
rect 18543 9052 18560 9092
rect 18600 9052 18609 9092
rect 18223 9029 18289 9052
rect 18375 9029 18457 9052
rect 18543 9029 18609 9052
rect 18223 9010 18609 9029
rect 33343 9115 33729 9134
rect 33343 9092 33409 9115
rect 33495 9092 33577 9115
rect 33663 9092 33729 9115
rect 33343 9052 33352 9092
rect 33392 9052 33409 9092
rect 33495 9052 33516 9092
rect 33556 9052 33577 9092
rect 33663 9052 33680 9092
rect 33720 9052 33729 9092
rect 33343 9029 33409 9052
rect 33495 9029 33577 9052
rect 33663 9029 33729 9052
rect 33343 9010 33729 9029
rect 48463 9115 48849 9134
rect 48463 9092 48529 9115
rect 48615 9092 48697 9115
rect 48783 9092 48849 9115
rect 48463 9052 48472 9092
rect 48512 9052 48529 9092
rect 48615 9052 48636 9092
rect 48676 9052 48697 9092
rect 48783 9052 48800 9092
rect 48840 9052 48849 9092
rect 48463 9029 48529 9052
rect 48615 9029 48697 9052
rect 48783 9029 48849 9052
rect 48463 9010 48849 9029
rect 63583 9115 63969 9134
rect 63583 9092 63649 9115
rect 63735 9092 63817 9115
rect 63903 9092 63969 9115
rect 63583 9052 63592 9092
rect 63632 9052 63649 9092
rect 63735 9052 63756 9092
rect 63796 9052 63817 9092
rect 63903 9052 63920 9092
rect 63960 9052 63969 9092
rect 63583 9029 63649 9052
rect 63735 9029 63817 9052
rect 63903 9029 63969 9052
rect 63583 9010 63969 9029
rect 78703 9115 79089 9134
rect 78703 9092 78769 9115
rect 78855 9092 78937 9115
rect 79023 9092 79089 9115
rect 78703 9052 78712 9092
rect 78752 9052 78769 9092
rect 78855 9052 78876 9092
rect 78916 9052 78937 9092
rect 79023 9052 79040 9092
rect 79080 9052 79089 9092
rect 78703 9029 78769 9052
rect 78855 9029 78937 9052
rect 79023 9029 79089 9052
rect 78703 9010 79089 9029
rect 93823 9115 94209 9134
rect 93823 9092 93889 9115
rect 93975 9092 94057 9115
rect 94143 9092 94209 9115
rect 93823 9052 93832 9092
rect 93872 9052 93889 9092
rect 93975 9052 93996 9092
rect 94036 9052 94057 9092
rect 94143 9052 94160 9092
rect 94200 9052 94209 9092
rect 93823 9029 93889 9052
rect 93975 9029 94057 9052
rect 94143 9029 94209 9052
rect 93823 9010 94209 9029
rect 4343 8359 4729 8378
rect 4343 8336 4409 8359
rect 4495 8336 4577 8359
rect 4663 8336 4729 8359
rect 4343 8296 4352 8336
rect 4392 8296 4409 8336
rect 4495 8296 4516 8336
rect 4556 8296 4577 8336
rect 4663 8296 4680 8336
rect 4720 8296 4729 8336
rect 4343 8273 4409 8296
rect 4495 8273 4577 8296
rect 4663 8273 4729 8296
rect 4343 8254 4729 8273
rect 19463 8359 19849 8378
rect 19463 8336 19529 8359
rect 19615 8336 19697 8359
rect 19783 8336 19849 8359
rect 19463 8296 19472 8336
rect 19512 8296 19529 8336
rect 19615 8296 19636 8336
rect 19676 8296 19697 8336
rect 19783 8296 19800 8336
rect 19840 8296 19849 8336
rect 19463 8273 19529 8296
rect 19615 8273 19697 8296
rect 19783 8273 19849 8296
rect 19463 8254 19849 8273
rect 34583 8359 34969 8378
rect 34583 8336 34649 8359
rect 34735 8336 34817 8359
rect 34903 8336 34969 8359
rect 34583 8296 34592 8336
rect 34632 8296 34649 8336
rect 34735 8296 34756 8336
rect 34796 8296 34817 8336
rect 34903 8296 34920 8336
rect 34960 8296 34969 8336
rect 34583 8273 34649 8296
rect 34735 8273 34817 8296
rect 34903 8273 34969 8296
rect 34583 8254 34969 8273
rect 49703 8359 50089 8378
rect 49703 8336 49769 8359
rect 49855 8336 49937 8359
rect 50023 8336 50089 8359
rect 49703 8296 49712 8336
rect 49752 8296 49769 8336
rect 49855 8296 49876 8336
rect 49916 8296 49937 8336
rect 50023 8296 50040 8336
rect 50080 8296 50089 8336
rect 49703 8273 49769 8296
rect 49855 8273 49937 8296
rect 50023 8273 50089 8296
rect 49703 8254 50089 8273
rect 64823 8359 65209 8378
rect 64823 8336 64889 8359
rect 64975 8336 65057 8359
rect 65143 8336 65209 8359
rect 64823 8296 64832 8336
rect 64872 8296 64889 8336
rect 64975 8296 64996 8336
rect 65036 8296 65057 8336
rect 65143 8296 65160 8336
rect 65200 8296 65209 8336
rect 64823 8273 64889 8296
rect 64975 8273 65057 8296
rect 65143 8273 65209 8296
rect 64823 8254 65209 8273
rect 79943 8359 80329 8378
rect 79943 8336 80009 8359
rect 80095 8336 80177 8359
rect 80263 8336 80329 8359
rect 79943 8296 79952 8336
rect 79992 8296 80009 8336
rect 80095 8296 80116 8336
rect 80156 8296 80177 8336
rect 80263 8296 80280 8336
rect 80320 8296 80329 8336
rect 79943 8273 80009 8296
rect 80095 8273 80177 8296
rect 80263 8273 80329 8296
rect 79943 8254 80329 8273
rect 95063 8359 95449 8378
rect 95063 8336 95129 8359
rect 95215 8336 95297 8359
rect 95383 8336 95449 8359
rect 95063 8296 95072 8336
rect 95112 8296 95129 8336
rect 95215 8296 95236 8336
rect 95276 8296 95297 8336
rect 95383 8296 95400 8336
rect 95440 8296 95449 8336
rect 95063 8273 95129 8296
rect 95215 8273 95297 8296
rect 95383 8273 95449 8296
rect 95063 8254 95449 8273
rect 3103 7603 3489 7622
rect 3103 7580 3169 7603
rect 3255 7580 3337 7603
rect 3423 7580 3489 7603
rect 3103 7540 3112 7580
rect 3152 7540 3169 7580
rect 3255 7540 3276 7580
rect 3316 7540 3337 7580
rect 3423 7540 3440 7580
rect 3480 7540 3489 7580
rect 3103 7517 3169 7540
rect 3255 7517 3337 7540
rect 3423 7517 3489 7540
rect 3103 7498 3489 7517
rect 18223 7603 18609 7622
rect 18223 7580 18289 7603
rect 18375 7580 18457 7603
rect 18543 7580 18609 7603
rect 18223 7540 18232 7580
rect 18272 7540 18289 7580
rect 18375 7540 18396 7580
rect 18436 7540 18457 7580
rect 18543 7540 18560 7580
rect 18600 7540 18609 7580
rect 18223 7517 18289 7540
rect 18375 7517 18457 7540
rect 18543 7517 18609 7540
rect 18223 7498 18609 7517
rect 33343 7603 33729 7622
rect 33343 7580 33409 7603
rect 33495 7580 33577 7603
rect 33663 7580 33729 7603
rect 33343 7540 33352 7580
rect 33392 7540 33409 7580
rect 33495 7540 33516 7580
rect 33556 7540 33577 7580
rect 33663 7540 33680 7580
rect 33720 7540 33729 7580
rect 33343 7517 33409 7540
rect 33495 7517 33577 7540
rect 33663 7517 33729 7540
rect 33343 7498 33729 7517
rect 48463 7603 48849 7622
rect 48463 7580 48529 7603
rect 48615 7580 48697 7603
rect 48783 7580 48849 7603
rect 48463 7540 48472 7580
rect 48512 7540 48529 7580
rect 48615 7540 48636 7580
rect 48676 7540 48697 7580
rect 48783 7540 48800 7580
rect 48840 7540 48849 7580
rect 48463 7517 48529 7540
rect 48615 7517 48697 7540
rect 48783 7517 48849 7540
rect 48463 7498 48849 7517
rect 63583 7603 63969 7622
rect 63583 7580 63649 7603
rect 63735 7580 63817 7603
rect 63903 7580 63969 7603
rect 63583 7540 63592 7580
rect 63632 7540 63649 7580
rect 63735 7540 63756 7580
rect 63796 7540 63817 7580
rect 63903 7540 63920 7580
rect 63960 7540 63969 7580
rect 63583 7517 63649 7540
rect 63735 7517 63817 7540
rect 63903 7517 63969 7540
rect 63583 7498 63969 7517
rect 78703 7603 79089 7622
rect 78703 7580 78769 7603
rect 78855 7580 78937 7603
rect 79023 7580 79089 7603
rect 78703 7540 78712 7580
rect 78752 7540 78769 7580
rect 78855 7540 78876 7580
rect 78916 7540 78937 7580
rect 79023 7540 79040 7580
rect 79080 7540 79089 7580
rect 78703 7517 78769 7540
rect 78855 7517 78937 7540
rect 79023 7517 79089 7540
rect 78703 7498 79089 7517
rect 93823 7603 94209 7622
rect 93823 7580 93889 7603
rect 93975 7580 94057 7603
rect 94143 7580 94209 7603
rect 93823 7540 93832 7580
rect 93872 7540 93889 7580
rect 93975 7540 93996 7580
rect 94036 7540 94057 7580
rect 94143 7540 94160 7580
rect 94200 7540 94209 7580
rect 93823 7517 93889 7540
rect 93975 7517 94057 7540
rect 94143 7517 94209 7540
rect 93823 7498 94209 7517
rect 4343 6847 4729 6866
rect 4343 6824 4409 6847
rect 4495 6824 4577 6847
rect 4663 6824 4729 6847
rect 4343 6784 4352 6824
rect 4392 6784 4409 6824
rect 4495 6784 4516 6824
rect 4556 6784 4577 6824
rect 4663 6784 4680 6824
rect 4720 6784 4729 6824
rect 4343 6761 4409 6784
rect 4495 6761 4577 6784
rect 4663 6761 4729 6784
rect 4343 6742 4729 6761
rect 19463 6847 19849 6866
rect 19463 6824 19529 6847
rect 19615 6824 19697 6847
rect 19783 6824 19849 6847
rect 19463 6784 19472 6824
rect 19512 6784 19529 6824
rect 19615 6784 19636 6824
rect 19676 6784 19697 6824
rect 19783 6784 19800 6824
rect 19840 6784 19849 6824
rect 19463 6761 19529 6784
rect 19615 6761 19697 6784
rect 19783 6761 19849 6784
rect 19463 6742 19849 6761
rect 34583 6847 34969 6866
rect 34583 6824 34649 6847
rect 34735 6824 34817 6847
rect 34903 6824 34969 6847
rect 34583 6784 34592 6824
rect 34632 6784 34649 6824
rect 34735 6784 34756 6824
rect 34796 6784 34817 6824
rect 34903 6784 34920 6824
rect 34960 6784 34969 6824
rect 34583 6761 34649 6784
rect 34735 6761 34817 6784
rect 34903 6761 34969 6784
rect 34583 6742 34969 6761
rect 49703 6847 50089 6866
rect 49703 6824 49769 6847
rect 49855 6824 49937 6847
rect 50023 6824 50089 6847
rect 49703 6784 49712 6824
rect 49752 6784 49769 6824
rect 49855 6784 49876 6824
rect 49916 6784 49937 6824
rect 50023 6784 50040 6824
rect 50080 6784 50089 6824
rect 49703 6761 49769 6784
rect 49855 6761 49937 6784
rect 50023 6761 50089 6784
rect 49703 6742 50089 6761
rect 64823 6847 65209 6866
rect 64823 6824 64889 6847
rect 64975 6824 65057 6847
rect 65143 6824 65209 6847
rect 64823 6784 64832 6824
rect 64872 6784 64889 6824
rect 64975 6784 64996 6824
rect 65036 6784 65057 6824
rect 65143 6784 65160 6824
rect 65200 6784 65209 6824
rect 64823 6761 64889 6784
rect 64975 6761 65057 6784
rect 65143 6761 65209 6784
rect 64823 6742 65209 6761
rect 79943 6847 80329 6866
rect 79943 6824 80009 6847
rect 80095 6824 80177 6847
rect 80263 6824 80329 6847
rect 79943 6784 79952 6824
rect 79992 6784 80009 6824
rect 80095 6784 80116 6824
rect 80156 6784 80177 6824
rect 80263 6784 80280 6824
rect 80320 6784 80329 6824
rect 79943 6761 80009 6784
rect 80095 6761 80177 6784
rect 80263 6761 80329 6784
rect 79943 6742 80329 6761
rect 95063 6847 95449 6866
rect 95063 6824 95129 6847
rect 95215 6824 95297 6847
rect 95383 6824 95449 6847
rect 95063 6784 95072 6824
rect 95112 6784 95129 6824
rect 95215 6784 95236 6824
rect 95276 6784 95297 6824
rect 95383 6784 95400 6824
rect 95440 6784 95449 6824
rect 95063 6761 95129 6784
rect 95215 6761 95297 6784
rect 95383 6761 95449 6784
rect 95063 6742 95449 6761
rect 3103 6091 3489 6110
rect 3103 6068 3169 6091
rect 3255 6068 3337 6091
rect 3423 6068 3489 6091
rect 3103 6028 3112 6068
rect 3152 6028 3169 6068
rect 3255 6028 3276 6068
rect 3316 6028 3337 6068
rect 3423 6028 3440 6068
rect 3480 6028 3489 6068
rect 3103 6005 3169 6028
rect 3255 6005 3337 6028
rect 3423 6005 3489 6028
rect 3103 5986 3489 6005
rect 18223 6091 18609 6110
rect 18223 6068 18289 6091
rect 18375 6068 18457 6091
rect 18543 6068 18609 6091
rect 18223 6028 18232 6068
rect 18272 6028 18289 6068
rect 18375 6028 18396 6068
rect 18436 6028 18457 6068
rect 18543 6028 18560 6068
rect 18600 6028 18609 6068
rect 18223 6005 18289 6028
rect 18375 6005 18457 6028
rect 18543 6005 18609 6028
rect 18223 5986 18609 6005
rect 33343 6091 33729 6110
rect 33343 6068 33409 6091
rect 33495 6068 33577 6091
rect 33663 6068 33729 6091
rect 33343 6028 33352 6068
rect 33392 6028 33409 6068
rect 33495 6028 33516 6068
rect 33556 6028 33577 6068
rect 33663 6028 33680 6068
rect 33720 6028 33729 6068
rect 33343 6005 33409 6028
rect 33495 6005 33577 6028
rect 33663 6005 33729 6028
rect 33343 5986 33729 6005
rect 48463 6091 48849 6110
rect 48463 6068 48529 6091
rect 48615 6068 48697 6091
rect 48783 6068 48849 6091
rect 48463 6028 48472 6068
rect 48512 6028 48529 6068
rect 48615 6028 48636 6068
rect 48676 6028 48697 6068
rect 48783 6028 48800 6068
rect 48840 6028 48849 6068
rect 48463 6005 48529 6028
rect 48615 6005 48697 6028
rect 48783 6005 48849 6028
rect 48463 5986 48849 6005
rect 63583 6091 63969 6110
rect 63583 6068 63649 6091
rect 63735 6068 63817 6091
rect 63903 6068 63969 6091
rect 63583 6028 63592 6068
rect 63632 6028 63649 6068
rect 63735 6028 63756 6068
rect 63796 6028 63817 6068
rect 63903 6028 63920 6068
rect 63960 6028 63969 6068
rect 63583 6005 63649 6028
rect 63735 6005 63817 6028
rect 63903 6005 63969 6028
rect 63583 5986 63969 6005
rect 78703 6091 79089 6110
rect 78703 6068 78769 6091
rect 78855 6068 78937 6091
rect 79023 6068 79089 6091
rect 78703 6028 78712 6068
rect 78752 6028 78769 6068
rect 78855 6028 78876 6068
rect 78916 6028 78937 6068
rect 79023 6028 79040 6068
rect 79080 6028 79089 6068
rect 78703 6005 78769 6028
rect 78855 6005 78937 6028
rect 79023 6005 79089 6028
rect 78703 5986 79089 6005
rect 93823 6091 94209 6110
rect 93823 6068 93889 6091
rect 93975 6068 94057 6091
rect 94143 6068 94209 6091
rect 93823 6028 93832 6068
rect 93872 6028 93889 6068
rect 93975 6028 93996 6068
rect 94036 6028 94057 6068
rect 94143 6028 94160 6068
rect 94200 6028 94209 6068
rect 93823 6005 93889 6028
rect 93975 6005 94057 6028
rect 94143 6005 94209 6028
rect 93823 5986 94209 6005
rect 4343 5335 4729 5354
rect 4343 5312 4409 5335
rect 4495 5312 4577 5335
rect 4663 5312 4729 5335
rect 4343 5272 4352 5312
rect 4392 5272 4409 5312
rect 4495 5272 4516 5312
rect 4556 5272 4577 5312
rect 4663 5272 4680 5312
rect 4720 5272 4729 5312
rect 4343 5249 4409 5272
rect 4495 5249 4577 5272
rect 4663 5249 4729 5272
rect 4343 5230 4729 5249
rect 19463 5335 19849 5354
rect 19463 5312 19529 5335
rect 19615 5312 19697 5335
rect 19783 5312 19849 5335
rect 19463 5272 19472 5312
rect 19512 5272 19529 5312
rect 19615 5272 19636 5312
rect 19676 5272 19697 5312
rect 19783 5272 19800 5312
rect 19840 5272 19849 5312
rect 19463 5249 19529 5272
rect 19615 5249 19697 5272
rect 19783 5249 19849 5272
rect 19463 5230 19849 5249
rect 34583 5335 34969 5354
rect 34583 5312 34649 5335
rect 34735 5312 34817 5335
rect 34903 5312 34969 5335
rect 34583 5272 34592 5312
rect 34632 5272 34649 5312
rect 34735 5272 34756 5312
rect 34796 5272 34817 5312
rect 34903 5272 34920 5312
rect 34960 5272 34969 5312
rect 34583 5249 34649 5272
rect 34735 5249 34817 5272
rect 34903 5249 34969 5272
rect 34583 5230 34969 5249
rect 49703 5335 50089 5354
rect 49703 5312 49769 5335
rect 49855 5312 49937 5335
rect 50023 5312 50089 5335
rect 49703 5272 49712 5312
rect 49752 5272 49769 5312
rect 49855 5272 49876 5312
rect 49916 5272 49937 5312
rect 50023 5272 50040 5312
rect 50080 5272 50089 5312
rect 49703 5249 49769 5272
rect 49855 5249 49937 5272
rect 50023 5249 50089 5272
rect 49703 5230 50089 5249
rect 64823 5335 65209 5354
rect 64823 5312 64889 5335
rect 64975 5312 65057 5335
rect 65143 5312 65209 5335
rect 64823 5272 64832 5312
rect 64872 5272 64889 5312
rect 64975 5272 64996 5312
rect 65036 5272 65057 5312
rect 65143 5272 65160 5312
rect 65200 5272 65209 5312
rect 64823 5249 64889 5272
rect 64975 5249 65057 5272
rect 65143 5249 65209 5272
rect 64823 5230 65209 5249
rect 79943 5335 80329 5354
rect 79943 5312 80009 5335
rect 80095 5312 80177 5335
rect 80263 5312 80329 5335
rect 79943 5272 79952 5312
rect 79992 5272 80009 5312
rect 80095 5272 80116 5312
rect 80156 5272 80177 5312
rect 80263 5272 80280 5312
rect 80320 5272 80329 5312
rect 79943 5249 80009 5272
rect 80095 5249 80177 5272
rect 80263 5249 80329 5272
rect 79943 5230 80329 5249
rect 95063 5335 95449 5354
rect 95063 5312 95129 5335
rect 95215 5312 95297 5335
rect 95383 5312 95449 5335
rect 95063 5272 95072 5312
rect 95112 5272 95129 5312
rect 95215 5272 95236 5312
rect 95276 5272 95297 5312
rect 95383 5272 95400 5312
rect 95440 5272 95449 5312
rect 95063 5249 95129 5272
rect 95215 5249 95297 5272
rect 95383 5249 95449 5272
rect 95063 5230 95449 5249
rect 3103 4579 3489 4598
rect 3103 4556 3169 4579
rect 3255 4556 3337 4579
rect 3423 4556 3489 4579
rect 3103 4516 3112 4556
rect 3152 4516 3169 4556
rect 3255 4516 3276 4556
rect 3316 4516 3337 4556
rect 3423 4516 3440 4556
rect 3480 4516 3489 4556
rect 3103 4493 3169 4516
rect 3255 4493 3337 4516
rect 3423 4493 3489 4516
rect 3103 4474 3489 4493
rect 18223 4579 18609 4598
rect 18223 4556 18289 4579
rect 18375 4556 18457 4579
rect 18543 4556 18609 4579
rect 18223 4516 18232 4556
rect 18272 4516 18289 4556
rect 18375 4516 18396 4556
rect 18436 4516 18457 4556
rect 18543 4516 18560 4556
rect 18600 4516 18609 4556
rect 18223 4493 18289 4516
rect 18375 4493 18457 4516
rect 18543 4493 18609 4516
rect 18223 4474 18609 4493
rect 33343 4579 33729 4598
rect 33343 4556 33409 4579
rect 33495 4556 33577 4579
rect 33663 4556 33729 4579
rect 33343 4516 33352 4556
rect 33392 4516 33409 4556
rect 33495 4516 33516 4556
rect 33556 4516 33577 4556
rect 33663 4516 33680 4556
rect 33720 4516 33729 4556
rect 33343 4493 33409 4516
rect 33495 4493 33577 4516
rect 33663 4493 33729 4516
rect 33343 4474 33729 4493
rect 48463 4579 48849 4598
rect 48463 4556 48529 4579
rect 48615 4556 48697 4579
rect 48783 4556 48849 4579
rect 48463 4516 48472 4556
rect 48512 4516 48529 4556
rect 48615 4516 48636 4556
rect 48676 4516 48697 4556
rect 48783 4516 48800 4556
rect 48840 4516 48849 4556
rect 48463 4493 48529 4516
rect 48615 4493 48697 4516
rect 48783 4493 48849 4516
rect 48463 4474 48849 4493
rect 63583 4579 63969 4598
rect 63583 4556 63649 4579
rect 63735 4556 63817 4579
rect 63903 4556 63969 4579
rect 63583 4516 63592 4556
rect 63632 4516 63649 4556
rect 63735 4516 63756 4556
rect 63796 4516 63817 4556
rect 63903 4516 63920 4556
rect 63960 4516 63969 4556
rect 63583 4493 63649 4516
rect 63735 4493 63817 4516
rect 63903 4493 63969 4516
rect 63583 4474 63969 4493
rect 78703 4579 79089 4598
rect 78703 4556 78769 4579
rect 78855 4556 78937 4579
rect 79023 4556 79089 4579
rect 78703 4516 78712 4556
rect 78752 4516 78769 4556
rect 78855 4516 78876 4556
rect 78916 4516 78937 4556
rect 79023 4516 79040 4556
rect 79080 4516 79089 4556
rect 78703 4493 78769 4516
rect 78855 4493 78937 4516
rect 79023 4493 79089 4516
rect 78703 4474 79089 4493
rect 93823 4579 94209 4598
rect 93823 4556 93889 4579
rect 93975 4556 94057 4579
rect 94143 4556 94209 4579
rect 93823 4516 93832 4556
rect 93872 4516 93889 4556
rect 93975 4516 93996 4556
rect 94036 4516 94057 4556
rect 94143 4516 94160 4556
rect 94200 4516 94209 4556
rect 93823 4493 93889 4516
rect 93975 4493 94057 4516
rect 94143 4493 94209 4516
rect 93823 4474 94209 4493
rect 4343 3823 4729 3842
rect 4343 3800 4409 3823
rect 4495 3800 4577 3823
rect 4663 3800 4729 3823
rect 4343 3760 4352 3800
rect 4392 3760 4409 3800
rect 4495 3760 4516 3800
rect 4556 3760 4577 3800
rect 4663 3760 4680 3800
rect 4720 3760 4729 3800
rect 4343 3737 4409 3760
rect 4495 3737 4577 3760
rect 4663 3737 4729 3760
rect 4343 3718 4729 3737
rect 19463 3823 19849 3842
rect 19463 3800 19529 3823
rect 19615 3800 19697 3823
rect 19783 3800 19849 3823
rect 19463 3760 19472 3800
rect 19512 3760 19529 3800
rect 19615 3760 19636 3800
rect 19676 3760 19697 3800
rect 19783 3760 19800 3800
rect 19840 3760 19849 3800
rect 19463 3737 19529 3760
rect 19615 3737 19697 3760
rect 19783 3737 19849 3760
rect 19463 3718 19849 3737
rect 34583 3823 34969 3842
rect 34583 3800 34649 3823
rect 34735 3800 34817 3823
rect 34903 3800 34969 3823
rect 34583 3760 34592 3800
rect 34632 3760 34649 3800
rect 34735 3760 34756 3800
rect 34796 3760 34817 3800
rect 34903 3760 34920 3800
rect 34960 3760 34969 3800
rect 34583 3737 34649 3760
rect 34735 3737 34817 3760
rect 34903 3737 34969 3760
rect 34583 3718 34969 3737
rect 49703 3823 50089 3842
rect 49703 3800 49769 3823
rect 49855 3800 49937 3823
rect 50023 3800 50089 3823
rect 49703 3760 49712 3800
rect 49752 3760 49769 3800
rect 49855 3760 49876 3800
rect 49916 3760 49937 3800
rect 50023 3760 50040 3800
rect 50080 3760 50089 3800
rect 49703 3737 49769 3760
rect 49855 3737 49937 3760
rect 50023 3737 50089 3760
rect 49703 3718 50089 3737
rect 64823 3823 65209 3842
rect 64823 3800 64889 3823
rect 64975 3800 65057 3823
rect 65143 3800 65209 3823
rect 64823 3760 64832 3800
rect 64872 3760 64889 3800
rect 64975 3760 64996 3800
rect 65036 3760 65057 3800
rect 65143 3760 65160 3800
rect 65200 3760 65209 3800
rect 64823 3737 64889 3760
rect 64975 3737 65057 3760
rect 65143 3737 65209 3760
rect 64823 3718 65209 3737
rect 79943 3823 80329 3842
rect 79943 3800 80009 3823
rect 80095 3800 80177 3823
rect 80263 3800 80329 3823
rect 79943 3760 79952 3800
rect 79992 3760 80009 3800
rect 80095 3760 80116 3800
rect 80156 3760 80177 3800
rect 80263 3760 80280 3800
rect 80320 3760 80329 3800
rect 79943 3737 80009 3760
rect 80095 3737 80177 3760
rect 80263 3737 80329 3760
rect 79943 3718 80329 3737
rect 95063 3823 95449 3842
rect 95063 3800 95129 3823
rect 95215 3800 95297 3823
rect 95383 3800 95449 3823
rect 95063 3760 95072 3800
rect 95112 3760 95129 3800
rect 95215 3760 95236 3800
rect 95276 3760 95297 3800
rect 95383 3760 95400 3800
rect 95440 3760 95449 3800
rect 95063 3737 95129 3760
rect 95215 3737 95297 3760
rect 95383 3737 95449 3760
rect 95063 3718 95449 3737
rect 3103 3067 3489 3086
rect 3103 3044 3169 3067
rect 3255 3044 3337 3067
rect 3423 3044 3489 3067
rect 3103 3004 3112 3044
rect 3152 3004 3169 3044
rect 3255 3004 3276 3044
rect 3316 3004 3337 3044
rect 3423 3004 3440 3044
rect 3480 3004 3489 3044
rect 3103 2981 3169 3004
rect 3255 2981 3337 3004
rect 3423 2981 3489 3004
rect 3103 2962 3489 2981
rect 18223 3067 18609 3086
rect 18223 3044 18289 3067
rect 18375 3044 18457 3067
rect 18543 3044 18609 3067
rect 18223 3004 18232 3044
rect 18272 3004 18289 3044
rect 18375 3004 18396 3044
rect 18436 3004 18457 3044
rect 18543 3004 18560 3044
rect 18600 3004 18609 3044
rect 18223 2981 18289 3004
rect 18375 2981 18457 3004
rect 18543 2981 18609 3004
rect 18223 2962 18609 2981
rect 33343 3067 33729 3086
rect 33343 3044 33409 3067
rect 33495 3044 33577 3067
rect 33663 3044 33729 3067
rect 33343 3004 33352 3044
rect 33392 3004 33409 3044
rect 33495 3004 33516 3044
rect 33556 3004 33577 3044
rect 33663 3004 33680 3044
rect 33720 3004 33729 3044
rect 33343 2981 33409 3004
rect 33495 2981 33577 3004
rect 33663 2981 33729 3004
rect 33343 2962 33729 2981
rect 48463 3067 48849 3086
rect 48463 3044 48529 3067
rect 48615 3044 48697 3067
rect 48783 3044 48849 3067
rect 48463 3004 48472 3044
rect 48512 3004 48529 3044
rect 48615 3004 48636 3044
rect 48676 3004 48697 3044
rect 48783 3004 48800 3044
rect 48840 3004 48849 3044
rect 48463 2981 48529 3004
rect 48615 2981 48697 3004
rect 48783 2981 48849 3004
rect 48463 2962 48849 2981
rect 63583 3067 63969 3086
rect 63583 3044 63649 3067
rect 63735 3044 63817 3067
rect 63903 3044 63969 3067
rect 63583 3004 63592 3044
rect 63632 3004 63649 3044
rect 63735 3004 63756 3044
rect 63796 3004 63817 3044
rect 63903 3004 63920 3044
rect 63960 3004 63969 3044
rect 63583 2981 63649 3004
rect 63735 2981 63817 3004
rect 63903 2981 63969 3004
rect 63583 2962 63969 2981
rect 78703 3067 79089 3086
rect 78703 3044 78769 3067
rect 78855 3044 78937 3067
rect 79023 3044 79089 3067
rect 78703 3004 78712 3044
rect 78752 3004 78769 3044
rect 78855 3004 78876 3044
rect 78916 3004 78937 3044
rect 79023 3004 79040 3044
rect 79080 3004 79089 3044
rect 78703 2981 78769 3004
rect 78855 2981 78937 3004
rect 79023 2981 79089 3004
rect 78703 2962 79089 2981
rect 93823 3067 94209 3086
rect 93823 3044 93889 3067
rect 93975 3044 94057 3067
rect 94143 3044 94209 3067
rect 93823 3004 93832 3044
rect 93872 3004 93889 3044
rect 93975 3004 93996 3044
rect 94036 3004 94057 3044
rect 94143 3004 94160 3044
rect 94200 3004 94209 3044
rect 93823 2981 93889 3004
rect 93975 2981 94057 3004
rect 94143 2981 94209 3004
rect 93823 2962 94209 2981
rect 4343 2311 4729 2330
rect 4343 2288 4409 2311
rect 4495 2288 4577 2311
rect 4663 2288 4729 2311
rect 4343 2248 4352 2288
rect 4392 2248 4409 2288
rect 4495 2248 4516 2288
rect 4556 2248 4577 2288
rect 4663 2248 4680 2288
rect 4720 2248 4729 2288
rect 4343 2225 4409 2248
rect 4495 2225 4577 2248
rect 4663 2225 4729 2248
rect 4343 2206 4729 2225
rect 19463 2311 19849 2330
rect 19463 2288 19529 2311
rect 19615 2288 19697 2311
rect 19783 2288 19849 2311
rect 19463 2248 19472 2288
rect 19512 2248 19529 2288
rect 19615 2248 19636 2288
rect 19676 2248 19697 2288
rect 19783 2248 19800 2288
rect 19840 2248 19849 2288
rect 19463 2225 19529 2248
rect 19615 2225 19697 2248
rect 19783 2225 19849 2248
rect 19463 2206 19849 2225
rect 34583 2311 34969 2330
rect 34583 2288 34649 2311
rect 34735 2288 34817 2311
rect 34903 2288 34969 2311
rect 34583 2248 34592 2288
rect 34632 2248 34649 2288
rect 34735 2248 34756 2288
rect 34796 2248 34817 2288
rect 34903 2248 34920 2288
rect 34960 2248 34969 2288
rect 34583 2225 34649 2248
rect 34735 2225 34817 2248
rect 34903 2225 34969 2248
rect 34583 2206 34969 2225
rect 49703 2311 50089 2330
rect 49703 2288 49769 2311
rect 49855 2288 49937 2311
rect 50023 2288 50089 2311
rect 49703 2248 49712 2288
rect 49752 2248 49769 2288
rect 49855 2248 49876 2288
rect 49916 2248 49937 2288
rect 50023 2248 50040 2288
rect 50080 2248 50089 2288
rect 49703 2225 49769 2248
rect 49855 2225 49937 2248
rect 50023 2225 50089 2248
rect 49703 2206 50089 2225
rect 64823 2311 65209 2330
rect 64823 2288 64889 2311
rect 64975 2288 65057 2311
rect 65143 2288 65209 2311
rect 64823 2248 64832 2288
rect 64872 2248 64889 2288
rect 64975 2248 64996 2288
rect 65036 2248 65057 2288
rect 65143 2248 65160 2288
rect 65200 2248 65209 2288
rect 64823 2225 64889 2248
rect 64975 2225 65057 2248
rect 65143 2225 65209 2248
rect 64823 2206 65209 2225
rect 79943 2311 80329 2330
rect 79943 2288 80009 2311
rect 80095 2288 80177 2311
rect 80263 2288 80329 2311
rect 79943 2248 79952 2288
rect 79992 2248 80009 2288
rect 80095 2248 80116 2288
rect 80156 2248 80177 2288
rect 80263 2248 80280 2288
rect 80320 2248 80329 2288
rect 79943 2225 80009 2248
rect 80095 2225 80177 2248
rect 80263 2225 80329 2248
rect 79943 2206 80329 2225
rect 95063 2311 95449 2330
rect 95063 2288 95129 2311
rect 95215 2288 95297 2311
rect 95383 2288 95449 2311
rect 95063 2248 95072 2288
rect 95112 2248 95129 2288
rect 95215 2248 95236 2288
rect 95276 2248 95297 2288
rect 95383 2248 95400 2288
rect 95440 2248 95449 2288
rect 95063 2225 95129 2248
rect 95215 2225 95297 2248
rect 95383 2225 95449 2248
rect 95063 2206 95449 2225
rect 3103 1555 3489 1574
rect 3103 1532 3169 1555
rect 3255 1532 3337 1555
rect 3423 1532 3489 1555
rect 3103 1492 3112 1532
rect 3152 1492 3169 1532
rect 3255 1492 3276 1532
rect 3316 1492 3337 1532
rect 3423 1492 3440 1532
rect 3480 1492 3489 1532
rect 3103 1469 3169 1492
rect 3255 1469 3337 1492
rect 3423 1469 3489 1492
rect 3103 1450 3489 1469
rect 18223 1555 18609 1574
rect 18223 1532 18289 1555
rect 18375 1532 18457 1555
rect 18543 1532 18609 1555
rect 18223 1492 18232 1532
rect 18272 1492 18289 1532
rect 18375 1492 18396 1532
rect 18436 1492 18457 1532
rect 18543 1492 18560 1532
rect 18600 1492 18609 1532
rect 18223 1469 18289 1492
rect 18375 1469 18457 1492
rect 18543 1469 18609 1492
rect 18223 1450 18609 1469
rect 33343 1555 33729 1574
rect 33343 1532 33409 1555
rect 33495 1532 33577 1555
rect 33663 1532 33729 1555
rect 33343 1492 33352 1532
rect 33392 1492 33409 1532
rect 33495 1492 33516 1532
rect 33556 1492 33577 1532
rect 33663 1492 33680 1532
rect 33720 1492 33729 1532
rect 33343 1469 33409 1492
rect 33495 1469 33577 1492
rect 33663 1469 33729 1492
rect 33343 1450 33729 1469
rect 48463 1555 48849 1574
rect 48463 1532 48529 1555
rect 48615 1532 48697 1555
rect 48783 1532 48849 1555
rect 48463 1492 48472 1532
rect 48512 1492 48529 1532
rect 48615 1492 48636 1532
rect 48676 1492 48697 1532
rect 48783 1492 48800 1532
rect 48840 1492 48849 1532
rect 48463 1469 48529 1492
rect 48615 1469 48697 1492
rect 48783 1469 48849 1492
rect 48463 1450 48849 1469
rect 63583 1555 63969 1574
rect 63583 1532 63649 1555
rect 63735 1532 63817 1555
rect 63903 1532 63969 1555
rect 63583 1492 63592 1532
rect 63632 1492 63649 1532
rect 63735 1492 63756 1532
rect 63796 1492 63817 1532
rect 63903 1492 63920 1532
rect 63960 1492 63969 1532
rect 63583 1469 63649 1492
rect 63735 1469 63817 1492
rect 63903 1469 63969 1492
rect 63583 1450 63969 1469
rect 78703 1555 79089 1574
rect 78703 1532 78769 1555
rect 78855 1532 78937 1555
rect 79023 1532 79089 1555
rect 78703 1492 78712 1532
rect 78752 1492 78769 1532
rect 78855 1492 78876 1532
rect 78916 1492 78937 1532
rect 79023 1492 79040 1532
rect 79080 1492 79089 1532
rect 78703 1469 78769 1492
rect 78855 1469 78937 1492
rect 79023 1469 79089 1492
rect 78703 1450 79089 1469
rect 93823 1555 94209 1574
rect 93823 1532 93889 1555
rect 93975 1532 94057 1555
rect 94143 1532 94209 1555
rect 93823 1492 93832 1532
rect 93872 1492 93889 1532
rect 93975 1492 93996 1532
rect 94036 1492 94057 1532
rect 94143 1492 94160 1532
rect 94200 1492 94209 1532
rect 93823 1469 93889 1492
rect 93975 1469 94057 1492
rect 94143 1469 94209 1492
rect 93823 1450 94209 1469
rect 4343 799 4729 818
rect 4343 776 4409 799
rect 4495 776 4577 799
rect 4663 776 4729 799
rect 4343 736 4352 776
rect 4392 736 4409 776
rect 4495 736 4516 776
rect 4556 736 4577 776
rect 4663 736 4680 776
rect 4720 736 4729 776
rect 4343 713 4409 736
rect 4495 713 4577 736
rect 4663 713 4729 736
rect 4343 694 4729 713
rect 19463 799 19849 818
rect 19463 776 19529 799
rect 19615 776 19697 799
rect 19783 776 19849 799
rect 19463 736 19472 776
rect 19512 736 19529 776
rect 19615 736 19636 776
rect 19676 736 19697 776
rect 19783 736 19800 776
rect 19840 736 19849 776
rect 19463 713 19529 736
rect 19615 713 19697 736
rect 19783 713 19849 736
rect 19463 694 19849 713
rect 34583 799 34969 818
rect 34583 776 34649 799
rect 34735 776 34817 799
rect 34903 776 34969 799
rect 34583 736 34592 776
rect 34632 736 34649 776
rect 34735 736 34756 776
rect 34796 736 34817 776
rect 34903 736 34920 776
rect 34960 736 34969 776
rect 34583 713 34649 736
rect 34735 713 34817 736
rect 34903 713 34969 736
rect 34583 694 34969 713
rect 49703 799 50089 818
rect 49703 776 49769 799
rect 49855 776 49937 799
rect 50023 776 50089 799
rect 49703 736 49712 776
rect 49752 736 49769 776
rect 49855 736 49876 776
rect 49916 736 49937 776
rect 50023 736 50040 776
rect 50080 736 50089 776
rect 49703 713 49769 736
rect 49855 713 49937 736
rect 50023 713 50089 736
rect 49703 694 50089 713
rect 64823 799 65209 818
rect 64823 776 64889 799
rect 64975 776 65057 799
rect 65143 776 65209 799
rect 64823 736 64832 776
rect 64872 736 64889 776
rect 64975 736 64996 776
rect 65036 736 65057 776
rect 65143 736 65160 776
rect 65200 736 65209 776
rect 64823 713 64889 736
rect 64975 713 65057 736
rect 65143 713 65209 736
rect 64823 694 65209 713
rect 79943 799 80329 818
rect 79943 776 80009 799
rect 80095 776 80177 799
rect 80263 776 80329 799
rect 79943 736 79952 776
rect 79992 736 80009 776
rect 80095 736 80116 776
rect 80156 736 80177 776
rect 80263 736 80280 776
rect 80320 736 80329 776
rect 79943 713 80009 736
rect 80095 713 80177 736
rect 80263 713 80329 736
rect 79943 694 80329 713
rect 95063 799 95449 818
rect 95063 776 95129 799
rect 95215 776 95297 799
rect 95383 776 95449 799
rect 95063 736 95072 776
rect 95112 736 95129 776
rect 95215 736 95236 776
rect 95276 736 95297 776
rect 95383 736 95400 776
rect 95440 736 95449 776
rect 95063 713 95129 736
rect 95215 713 95297 736
rect 95383 713 95449 736
rect 95063 694 95449 713
<< via5 >>
rect 4409 38576 4495 38599
rect 4577 38576 4663 38599
rect 4409 38536 4434 38576
rect 4434 38536 4474 38576
rect 4474 38536 4495 38576
rect 4577 38536 4598 38576
rect 4598 38536 4638 38576
rect 4638 38536 4663 38576
rect 4409 38513 4495 38536
rect 4577 38513 4663 38536
rect 19529 38576 19615 38599
rect 19697 38576 19783 38599
rect 19529 38536 19554 38576
rect 19554 38536 19594 38576
rect 19594 38536 19615 38576
rect 19697 38536 19718 38576
rect 19718 38536 19758 38576
rect 19758 38536 19783 38576
rect 19529 38513 19615 38536
rect 19697 38513 19783 38536
rect 34649 38576 34735 38599
rect 34817 38576 34903 38599
rect 34649 38536 34674 38576
rect 34674 38536 34714 38576
rect 34714 38536 34735 38576
rect 34817 38536 34838 38576
rect 34838 38536 34878 38576
rect 34878 38536 34903 38576
rect 34649 38513 34735 38536
rect 34817 38513 34903 38536
rect 49769 38576 49855 38599
rect 49937 38576 50023 38599
rect 49769 38536 49794 38576
rect 49794 38536 49834 38576
rect 49834 38536 49855 38576
rect 49937 38536 49958 38576
rect 49958 38536 49998 38576
rect 49998 38536 50023 38576
rect 49769 38513 49855 38536
rect 49937 38513 50023 38536
rect 64889 38576 64975 38599
rect 65057 38576 65143 38599
rect 64889 38536 64914 38576
rect 64914 38536 64954 38576
rect 64954 38536 64975 38576
rect 65057 38536 65078 38576
rect 65078 38536 65118 38576
rect 65118 38536 65143 38576
rect 64889 38513 64975 38536
rect 65057 38513 65143 38536
rect 80009 38576 80095 38599
rect 80177 38576 80263 38599
rect 80009 38536 80034 38576
rect 80034 38536 80074 38576
rect 80074 38536 80095 38576
rect 80177 38536 80198 38576
rect 80198 38536 80238 38576
rect 80238 38536 80263 38576
rect 80009 38513 80095 38536
rect 80177 38513 80263 38536
rect 95129 38576 95215 38599
rect 95297 38576 95383 38599
rect 95129 38536 95154 38576
rect 95154 38536 95194 38576
rect 95194 38536 95215 38576
rect 95297 38536 95318 38576
rect 95318 38536 95358 38576
rect 95358 38536 95383 38576
rect 95129 38513 95215 38536
rect 95297 38513 95383 38536
rect 3169 37820 3255 37843
rect 3337 37820 3423 37843
rect 3169 37780 3194 37820
rect 3194 37780 3234 37820
rect 3234 37780 3255 37820
rect 3337 37780 3358 37820
rect 3358 37780 3398 37820
rect 3398 37780 3423 37820
rect 3169 37757 3255 37780
rect 3337 37757 3423 37780
rect 18289 37820 18375 37843
rect 18457 37820 18543 37843
rect 18289 37780 18314 37820
rect 18314 37780 18354 37820
rect 18354 37780 18375 37820
rect 18457 37780 18478 37820
rect 18478 37780 18518 37820
rect 18518 37780 18543 37820
rect 18289 37757 18375 37780
rect 18457 37757 18543 37780
rect 33409 37820 33495 37843
rect 33577 37820 33663 37843
rect 33409 37780 33434 37820
rect 33434 37780 33474 37820
rect 33474 37780 33495 37820
rect 33577 37780 33598 37820
rect 33598 37780 33638 37820
rect 33638 37780 33663 37820
rect 33409 37757 33495 37780
rect 33577 37757 33663 37780
rect 48529 37820 48615 37843
rect 48697 37820 48783 37843
rect 48529 37780 48554 37820
rect 48554 37780 48594 37820
rect 48594 37780 48615 37820
rect 48697 37780 48718 37820
rect 48718 37780 48758 37820
rect 48758 37780 48783 37820
rect 48529 37757 48615 37780
rect 48697 37757 48783 37780
rect 63649 37820 63735 37843
rect 63817 37820 63903 37843
rect 63649 37780 63674 37820
rect 63674 37780 63714 37820
rect 63714 37780 63735 37820
rect 63817 37780 63838 37820
rect 63838 37780 63878 37820
rect 63878 37780 63903 37820
rect 63649 37757 63735 37780
rect 63817 37757 63903 37780
rect 78769 37820 78855 37843
rect 78937 37820 79023 37843
rect 78769 37780 78794 37820
rect 78794 37780 78834 37820
rect 78834 37780 78855 37820
rect 78937 37780 78958 37820
rect 78958 37780 78998 37820
rect 78998 37780 79023 37820
rect 78769 37757 78855 37780
rect 78937 37757 79023 37780
rect 93889 37820 93975 37843
rect 94057 37820 94143 37843
rect 93889 37780 93914 37820
rect 93914 37780 93954 37820
rect 93954 37780 93975 37820
rect 94057 37780 94078 37820
rect 94078 37780 94118 37820
rect 94118 37780 94143 37820
rect 93889 37757 93975 37780
rect 94057 37757 94143 37780
rect 4409 37064 4495 37087
rect 4577 37064 4663 37087
rect 4409 37024 4434 37064
rect 4434 37024 4474 37064
rect 4474 37024 4495 37064
rect 4577 37024 4598 37064
rect 4598 37024 4638 37064
rect 4638 37024 4663 37064
rect 4409 37001 4495 37024
rect 4577 37001 4663 37024
rect 19529 37064 19615 37087
rect 19697 37064 19783 37087
rect 19529 37024 19554 37064
rect 19554 37024 19594 37064
rect 19594 37024 19615 37064
rect 19697 37024 19718 37064
rect 19718 37024 19758 37064
rect 19758 37024 19783 37064
rect 19529 37001 19615 37024
rect 19697 37001 19783 37024
rect 34649 37064 34735 37087
rect 34817 37064 34903 37087
rect 34649 37024 34674 37064
rect 34674 37024 34714 37064
rect 34714 37024 34735 37064
rect 34817 37024 34838 37064
rect 34838 37024 34878 37064
rect 34878 37024 34903 37064
rect 34649 37001 34735 37024
rect 34817 37001 34903 37024
rect 49769 37064 49855 37087
rect 49937 37064 50023 37087
rect 49769 37024 49794 37064
rect 49794 37024 49834 37064
rect 49834 37024 49855 37064
rect 49937 37024 49958 37064
rect 49958 37024 49998 37064
rect 49998 37024 50023 37064
rect 49769 37001 49855 37024
rect 49937 37001 50023 37024
rect 64889 37064 64975 37087
rect 65057 37064 65143 37087
rect 64889 37024 64914 37064
rect 64914 37024 64954 37064
rect 64954 37024 64975 37064
rect 65057 37024 65078 37064
rect 65078 37024 65118 37064
rect 65118 37024 65143 37064
rect 64889 37001 64975 37024
rect 65057 37001 65143 37024
rect 80009 37064 80095 37087
rect 80177 37064 80263 37087
rect 80009 37024 80034 37064
rect 80034 37024 80074 37064
rect 80074 37024 80095 37064
rect 80177 37024 80198 37064
rect 80198 37024 80238 37064
rect 80238 37024 80263 37064
rect 80009 37001 80095 37024
rect 80177 37001 80263 37024
rect 95129 37064 95215 37087
rect 95297 37064 95383 37087
rect 95129 37024 95154 37064
rect 95154 37024 95194 37064
rect 95194 37024 95215 37064
rect 95297 37024 95318 37064
rect 95318 37024 95358 37064
rect 95358 37024 95383 37064
rect 95129 37001 95215 37024
rect 95297 37001 95383 37024
rect 3169 36308 3255 36331
rect 3337 36308 3423 36331
rect 3169 36268 3194 36308
rect 3194 36268 3234 36308
rect 3234 36268 3255 36308
rect 3337 36268 3358 36308
rect 3358 36268 3398 36308
rect 3398 36268 3423 36308
rect 3169 36245 3255 36268
rect 3337 36245 3423 36268
rect 18289 36308 18375 36331
rect 18457 36308 18543 36331
rect 18289 36268 18314 36308
rect 18314 36268 18354 36308
rect 18354 36268 18375 36308
rect 18457 36268 18478 36308
rect 18478 36268 18518 36308
rect 18518 36268 18543 36308
rect 18289 36245 18375 36268
rect 18457 36245 18543 36268
rect 33409 36308 33495 36331
rect 33577 36308 33663 36331
rect 33409 36268 33434 36308
rect 33434 36268 33474 36308
rect 33474 36268 33495 36308
rect 33577 36268 33598 36308
rect 33598 36268 33638 36308
rect 33638 36268 33663 36308
rect 33409 36245 33495 36268
rect 33577 36245 33663 36268
rect 48529 36308 48615 36331
rect 48697 36308 48783 36331
rect 48529 36268 48554 36308
rect 48554 36268 48594 36308
rect 48594 36268 48615 36308
rect 48697 36268 48718 36308
rect 48718 36268 48758 36308
rect 48758 36268 48783 36308
rect 48529 36245 48615 36268
rect 48697 36245 48783 36268
rect 63649 36308 63735 36331
rect 63817 36308 63903 36331
rect 63649 36268 63674 36308
rect 63674 36268 63714 36308
rect 63714 36268 63735 36308
rect 63817 36268 63838 36308
rect 63838 36268 63878 36308
rect 63878 36268 63903 36308
rect 63649 36245 63735 36268
rect 63817 36245 63903 36268
rect 78769 36308 78855 36331
rect 78937 36308 79023 36331
rect 78769 36268 78794 36308
rect 78794 36268 78834 36308
rect 78834 36268 78855 36308
rect 78937 36268 78958 36308
rect 78958 36268 78998 36308
rect 78998 36268 79023 36308
rect 78769 36245 78855 36268
rect 78937 36245 79023 36268
rect 93889 36308 93975 36331
rect 94057 36308 94143 36331
rect 93889 36268 93914 36308
rect 93914 36268 93954 36308
rect 93954 36268 93975 36308
rect 94057 36268 94078 36308
rect 94078 36268 94118 36308
rect 94118 36268 94143 36308
rect 93889 36245 93975 36268
rect 94057 36245 94143 36268
rect 4409 35552 4495 35575
rect 4577 35552 4663 35575
rect 4409 35512 4434 35552
rect 4434 35512 4474 35552
rect 4474 35512 4495 35552
rect 4577 35512 4598 35552
rect 4598 35512 4638 35552
rect 4638 35512 4663 35552
rect 4409 35489 4495 35512
rect 4577 35489 4663 35512
rect 19529 35552 19615 35575
rect 19697 35552 19783 35575
rect 19529 35512 19554 35552
rect 19554 35512 19594 35552
rect 19594 35512 19615 35552
rect 19697 35512 19718 35552
rect 19718 35512 19758 35552
rect 19758 35512 19783 35552
rect 19529 35489 19615 35512
rect 19697 35489 19783 35512
rect 34649 35552 34735 35575
rect 34817 35552 34903 35575
rect 34649 35512 34674 35552
rect 34674 35512 34714 35552
rect 34714 35512 34735 35552
rect 34817 35512 34838 35552
rect 34838 35512 34878 35552
rect 34878 35512 34903 35552
rect 34649 35489 34735 35512
rect 34817 35489 34903 35512
rect 49769 35552 49855 35575
rect 49937 35552 50023 35575
rect 49769 35512 49794 35552
rect 49794 35512 49834 35552
rect 49834 35512 49855 35552
rect 49937 35512 49958 35552
rect 49958 35512 49998 35552
rect 49998 35512 50023 35552
rect 49769 35489 49855 35512
rect 49937 35489 50023 35512
rect 64889 35552 64975 35575
rect 65057 35552 65143 35575
rect 64889 35512 64914 35552
rect 64914 35512 64954 35552
rect 64954 35512 64975 35552
rect 65057 35512 65078 35552
rect 65078 35512 65118 35552
rect 65118 35512 65143 35552
rect 64889 35489 64975 35512
rect 65057 35489 65143 35512
rect 80009 35552 80095 35575
rect 80177 35552 80263 35575
rect 80009 35512 80034 35552
rect 80034 35512 80074 35552
rect 80074 35512 80095 35552
rect 80177 35512 80198 35552
rect 80198 35512 80238 35552
rect 80238 35512 80263 35552
rect 80009 35489 80095 35512
rect 80177 35489 80263 35512
rect 95129 35552 95215 35575
rect 95297 35552 95383 35575
rect 95129 35512 95154 35552
rect 95154 35512 95194 35552
rect 95194 35512 95215 35552
rect 95297 35512 95318 35552
rect 95318 35512 95358 35552
rect 95358 35512 95383 35552
rect 95129 35489 95215 35512
rect 95297 35489 95383 35512
rect 3169 34796 3255 34819
rect 3337 34796 3423 34819
rect 3169 34756 3194 34796
rect 3194 34756 3234 34796
rect 3234 34756 3255 34796
rect 3337 34756 3358 34796
rect 3358 34756 3398 34796
rect 3398 34756 3423 34796
rect 3169 34733 3255 34756
rect 3337 34733 3423 34756
rect 18289 34796 18375 34819
rect 18457 34796 18543 34819
rect 18289 34756 18314 34796
rect 18314 34756 18354 34796
rect 18354 34756 18375 34796
rect 18457 34756 18478 34796
rect 18478 34756 18518 34796
rect 18518 34756 18543 34796
rect 18289 34733 18375 34756
rect 18457 34733 18543 34756
rect 33409 34796 33495 34819
rect 33577 34796 33663 34819
rect 33409 34756 33434 34796
rect 33434 34756 33474 34796
rect 33474 34756 33495 34796
rect 33577 34756 33598 34796
rect 33598 34756 33638 34796
rect 33638 34756 33663 34796
rect 33409 34733 33495 34756
rect 33577 34733 33663 34756
rect 48529 34796 48615 34819
rect 48697 34796 48783 34819
rect 48529 34756 48554 34796
rect 48554 34756 48594 34796
rect 48594 34756 48615 34796
rect 48697 34756 48718 34796
rect 48718 34756 48758 34796
rect 48758 34756 48783 34796
rect 48529 34733 48615 34756
rect 48697 34733 48783 34756
rect 63649 34796 63735 34819
rect 63817 34796 63903 34819
rect 63649 34756 63674 34796
rect 63674 34756 63714 34796
rect 63714 34756 63735 34796
rect 63817 34756 63838 34796
rect 63838 34756 63878 34796
rect 63878 34756 63903 34796
rect 63649 34733 63735 34756
rect 63817 34733 63903 34756
rect 78769 34796 78855 34819
rect 78937 34796 79023 34819
rect 78769 34756 78794 34796
rect 78794 34756 78834 34796
rect 78834 34756 78855 34796
rect 78937 34756 78958 34796
rect 78958 34756 78998 34796
rect 78998 34756 79023 34796
rect 78769 34733 78855 34756
rect 78937 34733 79023 34756
rect 93889 34796 93975 34819
rect 94057 34796 94143 34819
rect 93889 34756 93914 34796
rect 93914 34756 93954 34796
rect 93954 34756 93975 34796
rect 94057 34756 94078 34796
rect 94078 34756 94118 34796
rect 94118 34756 94143 34796
rect 93889 34733 93975 34756
rect 94057 34733 94143 34756
rect 4409 34040 4495 34063
rect 4577 34040 4663 34063
rect 4409 34000 4434 34040
rect 4434 34000 4474 34040
rect 4474 34000 4495 34040
rect 4577 34000 4598 34040
rect 4598 34000 4638 34040
rect 4638 34000 4663 34040
rect 4409 33977 4495 34000
rect 4577 33977 4663 34000
rect 19529 34040 19615 34063
rect 19697 34040 19783 34063
rect 19529 34000 19554 34040
rect 19554 34000 19594 34040
rect 19594 34000 19615 34040
rect 19697 34000 19718 34040
rect 19718 34000 19758 34040
rect 19758 34000 19783 34040
rect 19529 33977 19615 34000
rect 19697 33977 19783 34000
rect 34649 34040 34735 34063
rect 34817 34040 34903 34063
rect 34649 34000 34674 34040
rect 34674 34000 34714 34040
rect 34714 34000 34735 34040
rect 34817 34000 34838 34040
rect 34838 34000 34878 34040
rect 34878 34000 34903 34040
rect 34649 33977 34735 34000
rect 34817 33977 34903 34000
rect 49769 34040 49855 34063
rect 49937 34040 50023 34063
rect 49769 34000 49794 34040
rect 49794 34000 49834 34040
rect 49834 34000 49855 34040
rect 49937 34000 49958 34040
rect 49958 34000 49998 34040
rect 49998 34000 50023 34040
rect 49769 33977 49855 34000
rect 49937 33977 50023 34000
rect 64889 34040 64975 34063
rect 65057 34040 65143 34063
rect 64889 34000 64914 34040
rect 64914 34000 64954 34040
rect 64954 34000 64975 34040
rect 65057 34000 65078 34040
rect 65078 34000 65118 34040
rect 65118 34000 65143 34040
rect 64889 33977 64975 34000
rect 65057 33977 65143 34000
rect 80009 34040 80095 34063
rect 80177 34040 80263 34063
rect 80009 34000 80034 34040
rect 80034 34000 80074 34040
rect 80074 34000 80095 34040
rect 80177 34000 80198 34040
rect 80198 34000 80238 34040
rect 80238 34000 80263 34040
rect 80009 33977 80095 34000
rect 80177 33977 80263 34000
rect 95129 34040 95215 34063
rect 95297 34040 95383 34063
rect 95129 34000 95154 34040
rect 95154 34000 95194 34040
rect 95194 34000 95215 34040
rect 95297 34000 95318 34040
rect 95318 34000 95358 34040
rect 95358 34000 95383 34040
rect 95129 33977 95215 34000
rect 95297 33977 95383 34000
rect 3169 33284 3255 33307
rect 3337 33284 3423 33307
rect 3169 33244 3194 33284
rect 3194 33244 3234 33284
rect 3234 33244 3255 33284
rect 3337 33244 3358 33284
rect 3358 33244 3398 33284
rect 3398 33244 3423 33284
rect 3169 33221 3255 33244
rect 3337 33221 3423 33244
rect 18289 33284 18375 33307
rect 18457 33284 18543 33307
rect 18289 33244 18314 33284
rect 18314 33244 18354 33284
rect 18354 33244 18375 33284
rect 18457 33244 18478 33284
rect 18478 33244 18518 33284
rect 18518 33244 18543 33284
rect 18289 33221 18375 33244
rect 18457 33221 18543 33244
rect 33409 33284 33495 33307
rect 33577 33284 33663 33307
rect 33409 33244 33434 33284
rect 33434 33244 33474 33284
rect 33474 33244 33495 33284
rect 33577 33244 33598 33284
rect 33598 33244 33638 33284
rect 33638 33244 33663 33284
rect 33409 33221 33495 33244
rect 33577 33221 33663 33244
rect 48529 33284 48615 33307
rect 48697 33284 48783 33307
rect 48529 33244 48554 33284
rect 48554 33244 48594 33284
rect 48594 33244 48615 33284
rect 48697 33244 48718 33284
rect 48718 33244 48758 33284
rect 48758 33244 48783 33284
rect 48529 33221 48615 33244
rect 48697 33221 48783 33244
rect 63649 33284 63735 33307
rect 63817 33284 63903 33307
rect 63649 33244 63674 33284
rect 63674 33244 63714 33284
rect 63714 33244 63735 33284
rect 63817 33244 63838 33284
rect 63838 33244 63878 33284
rect 63878 33244 63903 33284
rect 63649 33221 63735 33244
rect 63817 33221 63903 33244
rect 78769 33284 78855 33307
rect 78937 33284 79023 33307
rect 78769 33244 78794 33284
rect 78794 33244 78834 33284
rect 78834 33244 78855 33284
rect 78937 33244 78958 33284
rect 78958 33244 78998 33284
rect 78998 33244 79023 33284
rect 78769 33221 78855 33244
rect 78937 33221 79023 33244
rect 93889 33284 93975 33307
rect 94057 33284 94143 33307
rect 93889 33244 93914 33284
rect 93914 33244 93954 33284
rect 93954 33244 93975 33284
rect 94057 33244 94078 33284
rect 94078 33244 94118 33284
rect 94118 33244 94143 33284
rect 93889 33221 93975 33244
rect 94057 33221 94143 33244
rect 4409 32528 4495 32551
rect 4577 32528 4663 32551
rect 4409 32488 4434 32528
rect 4434 32488 4474 32528
rect 4474 32488 4495 32528
rect 4577 32488 4598 32528
rect 4598 32488 4638 32528
rect 4638 32488 4663 32528
rect 4409 32465 4495 32488
rect 4577 32465 4663 32488
rect 19529 32528 19615 32551
rect 19697 32528 19783 32551
rect 19529 32488 19554 32528
rect 19554 32488 19594 32528
rect 19594 32488 19615 32528
rect 19697 32488 19718 32528
rect 19718 32488 19758 32528
rect 19758 32488 19783 32528
rect 19529 32465 19615 32488
rect 19697 32465 19783 32488
rect 34649 32528 34735 32551
rect 34817 32528 34903 32551
rect 34649 32488 34674 32528
rect 34674 32488 34714 32528
rect 34714 32488 34735 32528
rect 34817 32488 34838 32528
rect 34838 32488 34878 32528
rect 34878 32488 34903 32528
rect 34649 32465 34735 32488
rect 34817 32465 34903 32488
rect 49769 32528 49855 32551
rect 49937 32528 50023 32551
rect 49769 32488 49794 32528
rect 49794 32488 49834 32528
rect 49834 32488 49855 32528
rect 49937 32488 49958 32528
rect 49958 32488 49998 32528
rect 49998 32488 50023 32528
rect 49769 32465 49855 32488
rect 49937 32465 50023 32488
rect 64889 32528 64975 32551
rect 65057 32528 65143 32551
rect 64889 32488 64914 32528
rect 64914 32488 64954 32528
rect 64954 32488 64975 32528
rect 65057 32488 65078 32528
rect 65078 32488 65118 32528
rect 65118 32488 65143 32528
rect 64889 32465 64975 32488
rect 65057 32465 65143 32488
rect 80009 32528 80095 32551
rect 80177 32528 80263 32551
rect 80009 32488 80034 32528
rect 80034 32488 80074 32528
rect 80074 32488 80095 32528
rect 80177 32488 80198 32528
rect 80198 32488 80238 32528
rect 80238 32488 80263 32528
rect 80009 32465 80095 32488
rect 80177 32465 80263 32488
rect 95129 32528 95215 32551
rect 95297 32528 95383 32551
rect 95129 32488 95154 32528
rect 95154 32488 95194 32528
rect 95194 32488 95215 32528
rect 95297 32488 95318 32528
rect 95318 32488 95358 32528
rect 95358 32488 95383 32528
rect 95129 32465 95215 32488
rect 95297 32465 95383 32488
rect 3169 31772 3255 31795
rect 3337 31772 3423 31795
rect 3169 31732 3194 31772
rect 3194 31732 3234 31772
rect 3234 31732 3255 31772
rect 3337 31732 3358 31772
rect 3358 31732 3398 31772
rect 3398 31732 3423 31772
rect 3169 31709 3255 31732
rect 3337 31709 3423 31732
rect 18289 31772 18375 31795
rect 18457 31772 18543 31795
rect 18289 31732 18314 31772
rect 18314 31732 18354 31772
rect 18354 31732 18375 31772
rect 18457 31732 18478 31772
rect 18478 31732 18518 31772
rect 18518 31732 18543 31772
rect 18289 31709 18375 31732
rect 18457 31709 18543 31732
rect 33409 31772 33495 31795
rect 33577 31772 33663 31795
rect 33409 31732 33434 31772
rect 33434 31732 33474 31772
rect 33474 31732 33495 31772
rect 33577 31732 33598 31772
rect 33598 31732 33638 31772
rect 33638 31732 33663 31772
rect 33409 31709 33495 31732
rect 33577 31709 33663 31732
rect 48529 31772 48615 31795
rect 48697 31772 48783 31795
rect 48529 31732 48554 31772
rect 48554 31732 48594 31772
rect 48594 31732 48615 31772
rect 48697 31732 48718 31772
rect 48718 31732 48758 31772
rect 48758 31732 48783 31772
rect 48529 31709 48615 31732
rect 48697 31709 48783 31732
rect 63649 31772 63735 31795
rect 63817 31772 63903 31795
rect 63649 31732 63674 31772
rect 63674 31732 63714 31772
rect 63714 31732 63735 31772
rect 63817 31732 63838 31772
rect 63838 31732 63878 31772
rect 63878 31732 63903 31772
rect 63649 31709 63735 31732
rect 63817 31709 63903 31732
rect 78769 31772 78855 31795
rect 78937 31772 79023 31795
rect 78769 31732 78794 31772
rect 78794 31732 78834 31772
rect 78834 31732 78855 31772
rect 78937 31732 78958 31772
rect 78958 31732 78998 31772
rect 78998 31732 79023 31772
rect 78769 31709 78855 31732
rect 78937 31709 79023 31732
rect 93889 31772 93975 31795
rect 94057 31772 94143 31795
rect 93889 31732 93914 31772
rect 93914 31732 93954 31772
rect 93954 31732 93975 31772
rect 94057 31732 94078 31772
rect 94078 31732 94118 31772
rect 94118 31732 94143 31772
rect 93889 31709 93975 31732
rect 94057 31709 94143 31732
rect 4409 31016 4495 31039
rect 4577 31016 4663 31039
rect 4409 30976 4434 31016
rect 4434 30976 4474 31016
rect 4474 30976 4495 31016
rect 4577 30976 4598 31016
rect 4598 30976 4638 31016
rect 4638 30976 4663 31016
rect 4409 30953 4495 30976
rect 4577 30953 4663 30976
rect 19529 31016 19615 31039
rect 19697 31016 19783 31039
rect 19529 30976 19554 31016
rect 19554 30976 19594 31016
rect 19594 30976 19615 31016
rect 19697 30976 19718 31016
rect 19718 30976 19758 31016
rect 19758 30976 19783 31016
rect 19529 30953 19615 30976
rect 19697 30953 19783 30976
rect 34649 31016 34735 31039
rect 34817 31016 34903 31039
rect 34649 30976 34674 31016
rect 34674 30976 34714 31016
rect 34714 30976 34735 31016
rect 34817 30976 34838 31016
rect 34838 30976 34878 31016
rect 34878 30976 34903 31016
rect 34649 30953 34735 30976
rect 34817 30953 34903 30976
rect 49769 31016 49855 31039
rect 49937 31016 50023 31039
rect 49769 30976 49794 31016
rect 49794 30976 49834 31016
rect 49834 30976 49855 31016
rect 49937 30976 49958 31016
rect 49958 30976 49998 31016
rect 49998 30976 50023 31016
rect 49769 30953 49855 30976
rect 49937 30953 50023 30976
rect 64889 31016 64975 31039
rect 65057 31016 65143 31039
rect 64889 30976 64914 31016
rect 64914 30976 64954 31016
rect 64954 30976 64975 31016
rect 65057 30976 65078 31016
rect 65078 30976 65118 31016
rect 65118 30976 65143 31016
rect 64889 30953 64975 30976
rect 65057 30953 65143 30976
rect 80009 31016 80095 31039
rect 80177 31016 80263 31039
rect 80009 30976 80034 31016
rect 80034 30976 80074 31016
rect 80074 30976 80095 31016
rect 80177 30976 80198 31016
rect 80198 30976 80238 31016
rect 80238 30976 80263 31016
rect 80009 30953 80095 30976
rect 80177 30953 80263 30976
rect 95129 31016 95215 31039
rect 95297 31016 95383 31039
rect 95129 30976 95154 31016
rect 95154 30976 95194 31016
rect 95194 30976 95215 31016
rect 95297 30976 95318 31016
rect 95318 30976 95358 31016
rect 95358 30976 95383 31016
rect 95129 30953 95215 30976
rect 95297 30953 95383 30976
rect 3169 30260 3255 30283
rect 3337 30260 3423 30283
rect 3169 30220 3194 30260
rect 3194 30220 3234 30260
rect 3234 30220 3255 30260
rect 3337 30220 3358 30260
rect 3358 30220 3398 30260
rect 3398 30220 3423 30260
rect 3169 30197 3255 30220
rect 3337 30197 3423 30220
rect 18289 30260 18375 30283
rect 18457 30260 18543 30283
rect 18289 30220 18314 30260
rect 18314 30220 18354 30260
rect 18354 30220 18375 30260
rect 18457 30220 18478 30260
rect 18478 30220 18518 30260
rect 18518 30220 18543 30260
rect 18289 30197 18375 30220
rect 18457 30197 18543 30220
rect 33409 30260 33495 30283
rect 33577 30260 33663 30283
rect 33409 30220 33434 30260
rect 33434 30220 33474 30260
rect 33474 30220 33495 30260
rect 33577 30220 33598 30260
rect 33598 30220 33638 30260
rect 33638 30220 33663 30260
rect 33409 30197 33495 30220
rect 33577 30197 33663 30220
rect 48529 30260 48615 30283
rect 48697 30260 48783 30283
rect 48529 30220 48554 30260
rect 48554 30220 48594 30260
rect 48594 30220 48615 30260
rect 48697 30220 48718 30260
rect 48718 30220 48758 30260
rect 48758 30220 48783 30260
rect 48529 30197 48615 30220
rect 48697 30197 48783 30220
rect 63649 30260 63735 30283
rect 63817 30260 63903 30283
rect 63649 30220 63674 30260
rect 63674 30220 63714 30260
rect 63714 30220 63735 30260
rect 63817 30220 63838 30260
rect 63838 30220 63878 30260
rect 63878 30220 63903 30260
rect 63649 30197 63735 30220
rect 63817 30197 63903 30220
rect 78769 30260 78855 30283
rect 78937 30260 79023 30283
rect 78769 30220 78794 30260
rect 78794 30220 78834 30260
rect 78834 30220 78855 30260
rect 78937 30220 78958 30260
rect 78958 30220 78998 30260
rect 78998 30220 79023 30260
rect 78769 30197 78855 30220
rect 78937 30197 79023 30220
rect 93889 30260 93975 30283
rect 94057 30260 94143 30283
rect 93889 30220 93914 30260
rect 93914 30220 93954 30260
rect 93954 30220 93975 30260
rect 94057 30220 94078 30260
rect 94078 30220 94118 30260
rect 94118 30220 94143 30260
rect 93889 30197 93975 30220
rect 94057 30197 94143 30220
rect 4409 29504 4495 29527
rect 4577 29504 4663 29527
rect 4409 29464 4434 29504
rect 4434 29464 4474 29504
rect 4474 29464 4495 29504
rect 4577 29464 4598 29504
rect 4598 29464 4638 29504
rect 4638 29464 4663 29504
rect 4409 29441 4495 29464
rect 4577 29441 4663 29464
rect 19529 29504 19615 29527
rect 19697 29504 19783 29527
rect 19529 29464 19554 29504
rect 19554 29464 19594 29504
rect 19594 29464 19615 29504
rect 19697 29464 19718 29504
rect 19718 29464 19758 29504
rect 19758 29464 19783 29504
rect 19529 29441 19615 29464
rect 19697 29441 19783 29464
rect 34649 29504 34735 29527
rect 34817 29504 34903 29527
rect 34649 29464 34674 29504
rect 34674 29464 34714 29504
rect 34714 29464 34735 29504
rect 34817 29464 34838 29504
rect 34838 29464 34878 29504
rect 34878 29464 34903 29504
rect 34649 29441 34735 29464
rect 34817 29441 34903 29464
rect 49769 29504 49855 29527
rect 49937 29504 50023 29527
rect 49769 29464 49794 29504
rect 49794 29464 49834 29504
rect 49834 29464 49855 29504
rect 49937 29464 49958 29504
rect 49958 29464 49998 29504
rect 49998 29464 50023 29504
rect 49769 29441 49855 29464
rect 49937 29441 50023 29464
rect 64889 29504 64975 29527
rect 65057 29504 65143 29527
rect 64889 29464 64914 29504
rect 64914 29464 64954 29504
rect 64954 29464 64975 29504
rect 65057 29464 65078 29504
rect 65078 29464 65118 29504
rect 65118 29464 65143 29504
rect 64889 29441 64975 29464
rect 65057 29441 65143 29464
rect 80009 29504 80095 29527
rect 80177 29504 80263 29527
rect 80009 29464 80034 29504
rect 80034 29464 80074 29504
rect 80074 29464 80095 29504
rect 80177 29464 80198 29504
rect 80198 29464 80238 29504
rect 80238 29464 80263 29504
rect 80009 29441 80095 29464
rect 80177 29441 80263 29464
rect 95129 29504 95215 29527
rect 95297 29504 95383 29527
rect 95129 29464 95154 29504
rect 95154 29464 95194 29504
rect 95194 29464 95215 29504
rect 95297 29464 95318 29504
rect 95318 29464 95358 29504
rect 95358 29464 95383 29504
rect 95129 29441 95215 29464
rect 95297 29441 95383 29464
rect 3169 28748 3255 28771
rect 3337 28748 3423 28771
rect 3169 28708 3194 28748
rect 3194 28708 3234 28748
rect 3234 28708 3255 28748
rect 3337 28708 3358 28748
rect 3358 28708 3398 28748
rect 3398 28708 3423 28748
rect 3169 28685 3255 28708
rect 3337 28685 3423 28708
rect 18289 28748 18375 28771
rect 18457 28748 18543 28771
rect 18289 28708 18314 28748
rect 18314 28708 18354 28748
rect 18354 28708 18375 28748
rect 18457 28708 18478 28748
rect 18478 28708 18518 28748
rect 18518 28708 18543 28748
rect 18289 28685 18375 28708
rect 18457 28685 18543 28708
rect 33409 28748 33495 28771
rect 33577 28748 33663 28771
rect 33409 28708 33434 28748
rect 33434 28708 33474 28748
rect 33474 28708 33495 28748
rect 33577 28708 33598 28748
rect 33598 28708 33638 28748
rect 33638 28708 33663 28748
rect 33409 28685 33495 28708
rect 33577 28685 33663 28708
rect 48529 28748 48615 28771
rect 48697 28748 48783 28771
rect 48529 28708 48554 28748
rect 48554 28708 48594 28748
rect 48594 28708 48615 28748
rect 48697 28708 48718 28748
rect 48718 28708 48758 28748
rect 48758 28708 48783 28748
rect 48529 28685 48615 28708
rect 48697 28685 48783 28708
rect 63649 28748 63735 28771
rect 63817 28748 63903 28771
rect 63649 28708 63674 28748
rect 63674 28708 63714 28748
rect 63714 28708 63735 28748
rect 63817 28708 63838 28748
rect 63838 28708 63878 28748
rect 63878 28708 63903 28748
rect 63649 28685 63735 28708
rect 63817 28685 63903 28708
rect 78769 28748 78855 28771
rect 78937 28748 79023 28771
rect 78769 28708 78794 28748
rect 78794 28708 78834 28748
rect 78834 28708 78855 28748
rect 78937 28708 78958 28748
rect 78958 28708 78998 28748
rect 78998 28708 79023 28748
rect 78769 28685 78855 28708
rect 78937 28685 79023 28708
rect 93889 28748 93975 28771
rect 94057 28748 94143 28771
rect 93889 28708 93914 28748
rect 93914 28708 93954 28748
rect 93954 28708 93975 28748
rect 94057 28708 94078 28748
rect 94078 28708 94118 28748
rect 94118 28708 94143 28748
rect 93889 28685 93975 28708
rect 94057 28685 94143 28708
rect 4409 27992 4495 28015
rect 4577 27992 4663 28015
rect 4409 27952 4434 27992
rect 4434 27952 4474 27992
rect 4474 27952 4495 27992
rect 4577 27952 4598 27992
rect 4598 27952 4638 27992
rect 4638 27952 4663 27992
rect 4409 27929 4495 27952
rect 4577 27929 4663 27952
rect 19529 27992 19615 28015
rect 19697 27992 19783 28015
rect 19529 27952 19554 27992
rect 19554 27952 19594 27992
rect 19594 27952 19615 27992
rect 19697 27952 19718 27992
rect 19718 27952 19758 27992
rect 19758 27952 19783 27992
rect 19529 27929 19615 27952
rect 19697 27929 19783 27952
rect 34649 27992 34735 28015
rect 34817 27992 34903 28015
rect 34649 27952 34674 27992
rect 34674 27952 34714 27992
rect 34714 27952 34735 27992
rect 34817 27952 34838 27992
rect 34838 27952 34878 27992
rect 34878 27952 34903 27992
rect 34649 27929 34735 27952
rect 34817 27929 34903 27952
rect 49769 27992 49855 28015
rect 49937 27992 50023 28015
rect 49769 27952 49794 27992
rect 49794 27952 49834 27992
rect 49834 27952 49855 27992
rect 49937 27952 49958 27992
rect 49958 27952 49998 27992
rect 49998 27952 50023 27992
rect 49769 27929 49855 27952
rect 49937 27929 50023 27952
rect 64889 27992 64975 28015
rect 65057 27992 65143 28015
rect 64889 27952 64914 27992
rect 64914 27952 64954 27992
rect 64954 27952 64975 27992
rect 65057 27952 65078 27992
rect 65078 27952 65118 27992
rect 65118 27952 65143 27992
rect 64889 27929 64975 27952
rect 65057 27929 65143 27952
rect 80009 27992 80095 28015
rect 80177 27992 80263 28015
rect 80009 27952 80034 27992
rect 80034 27952 80074 27992
rect 80074 27952 80095 27992
rect 80177 27952 80198 27992
rect 80198 27952 80238 27992
rect 80238 27952 80263 27992
rect 80009 27929 80095 27952
rect 80177 27929 80263 27952
rect 95129 27992 95215 28015
rect 95297 27992 95383 28015
rect 95129 27952 95154 27992
rect 95154 27952 95194 27992
rect 95194 27952 95215 27992
rect 95297 27952 95318 27992
rect 95318 27952 95358 27992
rect 95358 27952 95383 27992
rect 95129 27929 95215 27952
rect 95297 27929 95383 27952
rect 3169 27236 3255 27259
rect 3337 27236 3423 27259
rect 3169 27196 3194 27236
rect 3194 27196 3234 27236
rect 3234 27196 3255 27236
rect 3337 27196 3358 27236
rect 3358 27196 3398 27236
rect 3398 27196 3423 27236
rect 3169 27173 3255 27196
rect 3337 27173 3423 27196
rect 18289 27236 18375 27259
rect 18457 27236 18543 27259
rect 18289 27196 18314 27236
rect 18314 27196 18354 27236
rect 18354 27196 18375 27236
rect 18457 27196 18478 27236
rect 18478 27196 18518 27236
rect 18518 27196 18543 27236
rect 18289 27173 18375 27196
rect 18457 27173 18543 27196
rect 33409 27236 33495 27259
rect 33577 27236 33663 27259
rect 33409 27196 33434 27236
rect 33434 27196 33474 27236
rect 33474 27196 33495 27236
rect 33577 27196 33598 27236
rect 33598 27196 33638 27236
rect 33638 27196 33663 27236
rect 33409 27173 33495 27196
rect 33577 27173 33663 27196
rect 48529 27236 48615 27259
rect 48697 27236 48783 27259
rect 48529 27196 48554 27236
rect 48554 27196 48594 27236
rect 48594 27196 48615 27236
rect 48697 27196 48718 27236
rect 48718 27196 48758 27236
rect 48758 27196 48783 27236
rect 48529 27173 48615 27196
rect 48697 27173 48783 27196
rect 63649 27236 63735 27259
rect 63817 27236 63903 27259
rect 63649 27196 63674 27236
rect 63674 27196 63714 27236
rect 63714 27196 63735 27236
rect 63817 27196 63838 27236
rect 63838 27196 63878 27236
rect 63878 27196 63903 27236
rect 63649 27173 63735 27196
rect 63817 27173 63903 27196
rect 78769 27236 78855 27259
rect 78937 27236 79023 27259
rect 78769 27196 78794 27236
rect 78794 27196 78834 27236
rect 78834 27196 78855 27236
rect 78937 27196 78958 27236
rect 78958 27196 78998 27236
rect 78998 27196 79023 27236
rect 78769 27173 78855 27196
rect 78937 27173 79023 27196
rect 93889 27236 93975 27259
rect 94057 27236 94143 27259
rect 93889 27196 93914 27236
rect 93914 27196 93954 27236
rect 93954 27196 93975 27236
rect 94057 27196 94078 27236
rect 94078 27196 94118 27236
rect 94118 27196 94143 27236
rect 93889 27173 93975 27196
rect 94057 27173 94143 27196
rect 4409 26480 4495 26503
rect 4577 26480 4663 26503
rect 4409 26440 4434 26480
rect 4434 26440 4474 26480
rect 4474 26440 4495 26480
rect 4577 26440 4598 26480
rect 4598 26440 4638 26480
rect 4638 26440 4663 26480
rect 4409 26417 4495 26440
rect 4577 26417 4663 26440
rect 19529 26480 19615 26503
rect 19697 26480 19783 26503
rect 19529 26440 19554 26480
rect 19554 26440 19594 26480
rect 19594 26440 19615 26480
rect 19697 26440 19718 26480
rect 19718 26440 19758 26480
rect 19758 26440 19783 26480
rect 19529 26417 19615 26440
rect 19697 26417 19783 26440
rect 34649 26480 34735 26503
rect 34817 26480 34903 26503
rect 34649 26440 34674 26480
rect 34674 26440 34714 26480
rect 34714 26440 34735 26480
rect 34817 26440 34838 26480
rect 34838 26440 34878 26480
rect 34878 26440 34903 26480
rect 34649 26417 34735 26440
rect 34817 26417 34903 26440
rect 49769 26480 49855 26503
rect 49937 26480 50023 26503
rect 49769 26440 49794 26480
rect 49794 26440 49834 26480
rect 49834 26440 49855 26480
rect 49937 26440 49958 26480
rect 49958 26440 49998 26480
rect 49998 26440 50023 26480
rect 49769 26417 49855 26440
rect 49937 26417 50023 26440
rect 64889 26480 64975 26503
rect 65057 26480 65143 26503
rect 64889 26440 64914 26480
rect 64914 26440 64954 26480
rect 64954 26440 64975 26480
rect 65057 26440 65078 26480
rect 65078 26440 65118 26480
rect 65118 26440 65143 26480
rect 64889 26417 64975 26440
rect 65057 26417 65143 26440
rect 80009 26480 80095 26503
rect 80177 26480 80263 26503
rect 80009 26440 80034 26480
rect 80034 26440 80074 26480
rect 80074 26440 80095 26480
rect 80177 26440 80198 26480
rect 80198 26440 80238 26480
rect 80238 26440 80263 26480
rect 80009 26417 80095 26440
rect 80177 26417 80263 26440
rect 95129 26480 95215 26503
rect 95297 26480 95383 26503
rect 95129 26440 95154 26480
rect 95154 26440 95194 26480
rect 95194 26440 95215 26480
rect 95297 26440 95318 26480
rect 95318 26440 95358 26480
rect 95358 26440 95383 26480
rect 95129 26417 95215 26440
rect 95297 26417 95383 26440
rect 3169 25724 3255 25747
rect 3337 25724 3423 25747
rect 3169 25684 3194 25724
rect 3194 25684 3234 25724
rect 3234 25684 3255 25724
rect 3337 25684 3358 25724
rect 3358 25684 3398 25724
rect 3398 25684 3423 25724
rect 3169 25661 3255 25684
rect 3337 25661 3423 25684
rect 18289 25724 18375 25747
rect 18457 25724 18543 25747
rect 18289 25684 18314 25724
rect 18314 25684 18354 25724
rect 18354 25684 18375 25724
rect 18457 25684 18478 25724
rect 18478 25684 18518 25724
rect 18518 25684 18543 25724
rect 18289 25661 18375 25684
rect 18457 25661 18543 25684
rect 33409 25724 33495 25747
rect 33577 25724 33663 25747
rect 33409 25684 33434 25724
rect 33434 25684 33474 25724
rect 33474 25684 33495 25724
rect 33577 25684 33598 25724
rect 33598 25684 33638 25724
rect 33638 25684 33663 25724
rect 33409 25661 33495 25684
rect 33577 25661 33663 25684
rect 48529 25724 48615 25747
rect 48697 25724 48783 25747
rect 48529 25684 48554 25724
rect 48554 25684 48594 25724
rect 48594 25684 48615 25724
rect 48697 25684 48718 25724
rect 48718 25684 48758 25724
rect 48758 25684 48783 25724
rect 48529 25661 48615 25684
rect 48697 25661 48783 25684
rect 63649 25724 63735 25747
rect 63817 25724 63903 25747
rect 63649 25684 63674 25724
rect 63674 25684 63714 25724
rect 63714 25684 63735 25724
rect 63817 25684 63838 25724
rect 63838 25684 63878 25724
rect 63878 25684 63903 25724
rect 63649 25661 63735 25684
rect 63817 25661 63903 25684
rect 78769 25724 78855 25747
rect 78937 25724 79023 25747
rect 78769 25684 78794 25724
rect 78794 25684 78834 25724
rect 78834 25684 78855 25724
rect 78937 25684 78958 25724
rect 78958 25684 78998 25724
rect 78998 25684 79023 25724
rect 78769 25661 78855 25684
rect 78937 25661 79023 25684
rect 93889 25724 93975 25747
rect 94057 25724 94143 25747
rect 93889 25684 93914 25724
rect 93914 25684 93954 25724
rect 93954 25684 93975 25724
rect 94057 25684 94078 25724
rect 94078 25684 94118 25724
rect 94118 25684 94143 25724
rect 93889 25661 93975 25684
rect 94057 25661 94143 25684
rect 4409 24968 4495 24991
rect 4577 24968 4663 24991
rect 4409 24928 4434 24968
rect 4434 24928 4474 24968
rect 4474 24928 4495 24968
rect 4577 24928 4598 24968
rect 4598 24928 4638 24968
rect 4638 24928 4663 24968
rect 4409 24905 4495 24928
rect 4577 24905 4663 24928
rect 19529 24968 19615 24991
rect 19697 24968 19783 24991
rect 19529 24928 19554 24968
rect 19554 24928 19594 24968
rect 19594 24928 19615 24968
rect 19697 24928 19718 24968
rect 19718 24928 19758 24968
rect 19758 24928 19783 24968
rect 19529 24905 19615 24928
rect 19697 24905 19783 24928
rect 34649 24968 34735 24991
rect 34817 24968 34903 24991
rect 34649 24928 34674 24968
rect 34674 24928 34714 24968
rect 34714 24928 34735 24968
rect 34817 24928 34838 24968
rect 34838 24928 34878 24968
rect 34878 24928 34903 24968
rect 34649 24905 34735 24928
rect 34817 24905 34903 24928
rect 49769 24968 49855 24991
rect 49937 24968 50023 24991
rect 49769 24928 49794 24968
rect 49794 24928 49834 24968
rect 49834 24928 49855 24968
rect 49937 24928 49958 24968
rect 49958 24928 49998 24968
rect 49998 24928 50023 24968
rect 49769 24905 49855 24928
rect 49937 24905 50023 24928
rect 64889 24968 64975 24991
rect 65057 24968 65143 24991
rect 64889 24928 64914 24968
rect 64914 24928 64954 24968
rect 64954 24928 64975 24968
rect 65057 24928 65078 24968
rect 65078 24928 65118 24968
rect 65118 24928 65143 24968
rect 64889 24905 64975 24928
rect 65057 24905 65143 24928
rect 80009 24968 80095 24991
rect 80177 24968 80263 24991
rect 80009 24928 80034 24968
rect 80034 24928 80074 24968
rect 80074 24928 80095 24968
rect 80177 24928 80198 24968
rect 80198 24928 80238 24968
rect 80238 24928 80263 24968
rect 80009 24905 80095 24928
rect 80177 24905 80263 24928
rect 95129 24968 95215 24991
rect 95297 24968 95383 24991
rect 95129 24928 95154 24968
rect 95154 24928 95194 24968
rect 95194 24928 95215 24968
rect 95297 24928 95318 24968
rect 95318 24928 95358 24968
rect 95358 24928 95383 24968
rect 95129 24905 95215 24928
rect 95297 24905 95383 24928
rect 3169 24212 3255 24235
rect 3337 24212 3423 24235
rect 3169 24172 3194 24212
rect 3194 24172 3234 24212
rect 3234 24172 3255 24212
rect 3337 24172 3358 24212
rect 3358 24172 3398 24212
rect 3398 24172 3423 24212
rect 3169 24149 3255 24172
rect 3337 24149 3423 24172
rect 18289 24212 18375 24235
rect 18457 24212 18543 24235
rect 18289 24172 18314 24212
rect 18314 24172 18354 24212
rect 18354 24172 18375 24212
rect 18457 24172 18478 24212
rect 18478 24172 18518 24212
rect 18518 24172 18543 24212
rect 18289 24149 18375 24172
rect 18457 24149 18543 24172
rect 33409 24212 33495 24235
rect 33577 24212 33663 24235
rect 33409 24172 33434 24212
rect 33434 24172 33474 24212
rect 33474 24172 33495 24212
rect 33577 24172 33598 24212
rect 33598 24172 33638 24212
rect 33638 24172 33663 24212
rect 33409 24149 33495 24172
rect 33577 24149 33663 24172
rect 48529 24212 48615 24235
rect 48697 24212 48783 24235
rect 48529 24172 48554 24212
rect 48554 24172 48594 24212
rect 48594 24172 48615 24212
rect 48697 24172 48718 24212
rect 48718 24172 48758 24212
rect 48758 24172 48783 24212
rect 48529 24149 48615 24172
rect 48697 24149 48783 24172
rect 63649 24212 63735 24235
rect 63817 24212 63903 24235
rect 63649 24172 63674 24212
rect 63674 24172 63714 24212
rect 63714 24172 63735 24212
rect 63817 24172 63838 24212
rect 63838 24172 63878 24212
rect 63878 24172 63903 24212
rect 63649 24149 63735 24172
rect 63817 24149 63903 24172
rect 78769 24212 78855 24235
rect 78937 24212 79023 24235
rect 78769 24172 78794 24212
rect 78794 24172 78834 24212
rect 78834 24172 78855 24212
rect 78937 24172 78958 24212
rect 78958 24172 78998 24212
rect 78998 24172 79023 24212
rect 78769 24149 78855 24172
rect 78937 24149 79023 24172
rect 93889 24212 93975 24235
rect 94057 24212 94143 24235
rect 93889 24172 93914 24212
rect 93914 24172 93954 24212
rect 93954 24172 93975 24212
rect 94057 24172 94078 24212
rect 94078 24172 94118 24212
rect 94118 24172 94143 24212
rect 93889 24149 93975 24172
rect 94057 24149 94143 24172
rect 4409 23456 4495 23479
rect 4577 23456 4663 23479
rect 4409 23416 4434 23456
rect 4434 23416 4474 23456
rect 4474 23416 4495 23456
rect 4577 23416 4598 23456
rect 4598 23416 4638 23456
rect 4638 23416 4663 23456
rect 4409 23393 4495 23416
rect 4577 23393 4663 23416
rect 19529 23456 19615 23479
rect 19697 23456 19783 23479
rect 19529 23416 19554 23456
rect 19554 23416 19594 23456
rect 19594 23416 19615 23456
rect 19697 23416 19718 23456
rect 19718 23416 19758 23456
rect 19758 23416 19783 23456
rect 19529 23393 19615 23416
rect 19697 23393 19783 23416
rect 34649 23456 34735 23479
rect 34817 23456 34903 23479
rect 34649 23416 34674 23456
rect 34674 23416 34714 23456
rect 34714 23416 34735 23456
rect 34817 23416 34838 23456
rect 34838 23416 34878 23456
rect 34878 23416 34903 23456
rect 34649 23393 34735 23416
rect 34817 23393 34903 23416
rect 49769 23456 49855 23479
rect 49937 23456 50023 23479
rect 49769 23416 49794 23456
rect 49794 23416 49834 23456
rect 49834 23416 49855 23456
rect 49937 23416 49958 23456
rect 49958 23416 49998 23456
rect 49998 23416 50023 23456
rect 49769 23393 49855 23416
rect 49937 23393 50023 23416
rect 64889 23456 64975 23479
rect 65057 23456 65143 23479
rect 64889 23416 64914 23456
rect 64914 23416 64954 23456
rect 64954 23416 64975 23456
rect 65057 23416 65078 23456
rect 65078 23416 65118 23456
rect 65118 23416 65143 23456
rect 64889 23393 64975 23416
rect 65057 23393 65143 23416
rect 80009 23456 80095 23479
rect 80177 23456 80263 23479
rect 80009 23416 80034 23456
rect 80034 23416 80074 23456
rect 80074 23416 80095 23456
rect 80177 23416 80198 23456
rect 80198 23416 80238 23456
rect 80238 23416 80263 23456
rect 80009 23393 80095 23416
rect 80177 23393 80263 23416
rect 95129 23456 95215 23479
rect 95297 23456 95383 23479
rect 95129 23416 95154 23456
rect 95154 23416 95194 23456
rect 95194 23416 95215 23456
rect 95297 23416 95318 23456
rect 95318 23416 95358 23456
rect 95358 23416 95383 23456
rect 95129 23393 95215 23416
rect 95297 23393 95383 23416
rect 3169 22700 3255 22723
rect 3337 22700 3423 22723
rect 3169 22660 3194 22700
rect 3194 22660 3234 22700
rect 3234 22660 3255 22700
rect 3337 22660 3358 22700
rect 3358 22660 3398 22700
rect 3398 22660 3423 22700
rect 3169 22637 3255 22660
rect 3337 22637 3423 22660
rect 18289 22700 18375 22723
rect 18457 22700 18543 22723
rect 18289 22660 18314 22700
rect 18314 22660 18354 22700
rect 18354 22660 18375 22700
rect 18457 22660 18478 22700
rect 18478 22660 18518 22700
rect 18518 22660 18543 22700
rect 18289 22637 18375 22660
rect 18457 22637 18543 22660
rect 33409 22700 33495 22723
rect 33577 22700 33663 22723
rect 33409 22660 33434 22700
rect 33434 22660 33474 22700
rect 33474 22660 33495 22700
rect 33577 22660 33598 22700
rect 33598 22660 33638 22700
rect 33638 22660 33663 22700
rect 33409 22637 33495 22660
rect 33577 22637 33663 22660
rect 48529 22700 48615 22723
rect 48697 22700 48783 22723
rect 48529 22660 48554 22700
rect 48554 22660 48594 22700
rect 48594 22660 48615 22700
rect 48697 22660 48718 22700
rect 48718 22660 48758 22700
rect 48758 22660 48783 22700
rect 48529 22637 48615 22660
rect 48697 22637 48783 22660
rect 63649 22700 63735 22723
rect 63817 22700 63903 22723
rect 63649 22660 63674 22700
rect 63674 22660 63714 22700
rect 63714 22660 63735 22700
rect 63817 22660 63838 22700
rect 63838 22660 63878 22700
rect 63878 22660 63903 22700
rect 63649 22637 63735 22660
rect 63817 22637 63903 22660
rect 78769 22700 78855 22723
rect 78937 22700 79023 22723
rect 78769 22660 78794 22700
rect 78794 22660 78834 22700
rect 78834 22660 78855 22700
rect 78937 22660 78958 22700
rect 78958 22660 78998 22700
rect 78998 22660 79023 22700
rect 78769 22637 78855 22660
rect 78937 22637 79023 22660
rect 93889 22700 93975 22723
rect 94057 22700 94143 22723
rect 93889 22660 93914 22700
rect 93914 22660 93954 22700
rect 93954 22660 93975 22700
rect 94057 22660 94078 22700
rect 94078 22660 94118 22700
rect 94118 22660 94143 22700
rect 93889 22637 93975 22660
rect 94057 22637 94143 22660
rect 4409 21944 4495 21967
rect 4577 21944 4663 21967
rect 4409 21904 4434 21944
rect 4434 21904 4474 21944
rect 4474 21904 4495 21944
rect 4577 21904 4598 21944
rect 4598 21904 4638 21944
rect 4638 21904 4663 21944
rect 4409 21881 4495 21904
rect 4577 21881 4663 21904
rect 19529 21944 19615 21967
rect 19697 21944 19783 21967
rect 19529 21904 19554 21944
rect 19554 21904 19594 21944
rect 19594 21904 19615 21944
rect 19697 21904 19718 21944
rect 19718 21904 19758 21944
rect 19758 21904 19783 21944
rect 19529 21881 19615 21904
rect 19697 21881 19783 21904
rect 34649 21944 34735 21967
rect 34817 21944 34903 21967
rect 34649 21904 34674 21944
rect 34674 21904 34714 21944
rect 34714 21904 34735 21944
rect 34817 21904 34838 21944
rect 34838 21904 34878 21944
rect 34878 21904 34903 21944
rect 34649 21881 34735 21904
rect 34817 21881 34903 21904
rect 49769 21944 49855 21967
rect 49937 21944 50023 21967
rect 49769 21904 49794 21944
rect 49794 21904 49834 21944
rect 49834 21904 49855 21944
rect 49937 21904 49958 21944
rect 49958 21904 49998 21944
rect 49998 21904 50023 21944
rect 49769 21881 49855 21904
rect 49937 21881 50023 21904
rect 64889 21944 64975 21967
rect 65057 21944 65143 21967
rect 64889 21904 64914 21944
rect 64914 21904 64954 21944
rect 64954 21904 64975 21944
rect 65057 21904 65078 21944
rect 65078 21904 65118 21944
rect 65118 21904 65143 21944
rect 64889 21881 64975 21904
rect 65057 21881 65143 21904
rect 80009 21944 80095 21967
rect 80177 21944 80263 21967
rect 80009 21904 80034 21944
rect 80034 21904 80074 21944
rect 80074 21904 80095 21944
rect 80177 21904 80198 21944
rect 80198 21904 80238 21944
rect 80238 21904 80263 21944
rect 80009 21881 80095 21904
rect 80177 21881 80263 21904
rect 95129 21944 95215 21967
rect 95297 21944 95383 21967
rect 95129 21904 95154 21944
rect 95154 21904 95194 21944
rect 95194 21904 95215 21944
rect 95297 21904 95318 21944
rect 95318 21904 95358 21944
rect 95358 21904 95383 21944
rect 95129 21881 95215 21904
rect 95297 21881 95383 21904
rect 3169 21188 3255 21211
rect 3337 21188 3423 21211
rect 3169 21148 3194 21188
rect 3194 21148 3234 21188
rect 3234 21148 3255 21188
rect 3337 21148 3358 21188
rect 3358 21148 3398 21188
rect 3398 21148 3423 21188
rect 3169 21125 3255 21148
rect 3337 21125 3423 21148
rect 18289 21188 18375 21211
rect 18457 21188 18543 21211
rect 18289 21148 18314 21188
rect 18314 21148 18354 21188
rect 18354 21148 18375 21188
rect 18457 21148 18478 21188
rect 18478 21148 18518 21188
rect 18518 21148 18543 21188
rect 18289 21125 18375 21148
rect 18457 21125 18543 21148
rect 33409 21188 33495 21211
rect 33577 21188 33663 21211
rect 33409 21148 33434 21188
rect 33434 21148 33474 21188
rect 33474 21148 33495 21188
rect 33577 21148 33598 21188
rect 33598 21148 33638 21188
rect 33638 21148 33663 21188
rect 33409 21125 33495 21148
rect 33577 21125 33663 21148
rect 48529 21188 48615 21211
rect 48697 21188 48783 21211
rect 48529 21148 48554 21188
rect 48554 21148 48594 21188
rect 48594 21148 48615 21188
rect 48697 21148 48718 21188
rect 48718 21148 48758 21188
rect 48758 21148 48783 21188
rect 48529 21125 48615 21148
rect 48697 21125 48783 21148
rect 63649 21188 63735 21211
rect 63817 21188 63903 21211
rect 63649 21148 63674 21188
rect 63674 21148 63714 21188
rect 63714 21148 63735 21188
rect 63817 21148 63838 21188
rect 63838 21148 63878 21188
rect 63878 21148 63903 21188
rect 63649 21125 63735 21148
rect 63817 21125 63903 21148
rect 78769 21188 78855 21211
rect 78937 21188 79023 21211
rect 78769 21148 78794 21188
rect 78794 21148 78834 21188
rect 78834 21148 78855 21188
rect 78937 21148 78958 21188
rect 78958 21148 78998 21188
rect 78998 21148 79023 21188
rect 78769 21125 78855 21148
rect 78937 21125 79023 21148
rect 93889 21188 93975 21211
rect 94057 21188 94143 21211
rect 93889 21148 93914 21188
rect 93914 21148 93954 21188
rect 93954 21148 93975 21188
rect 94057 21148 94078 21188
rect 94078 21148 94118 21188
rect 94118 21148 94143 21188
rect 93889 21125 93975 21148
rect 94057 21125 94143 21148
rect 4409 20432 4495 20455
rect 4577 20432 4663 20455
rect 4409 20392 4434 20432
rect 4434 20392 4474 20432
rect 4474 20392 4495 20432
rect 4577 20392 4598 20432
rect 4598 20392 4638 20432
rect 4638 20392 4663 20432
rect 4409 20369 4495 20392
rect 4577 20369 4663 20392
rect 19529 20432 19615 20455
rect 19697 20432 19783 20455
rect 19529 20392 19554 20432
rect 19554 20392 19594 20432
rect 19594 20392 19615 20432
rect 19697 20392 19718 20432
rect 19718 20392 19758 20432
rect 19758 20392 19783 20432
rect 19529 20369 19615 20392
rect 19697 20369 19783 20392
rect 34649 20432 34735 20455
rect 34817 20432 34903 20455
rect 34649 20392 34674 20432
rect 34674 20392 34714 20432
rect 34714 20392 34735 20432
rect 34817 20392 34838 20432
rect 34838 20392 34878 20432
rect 34878 20392 34903 20432
rect 34649 20369 34735 20392
rect 34817 20369 34903 20392
rect 49769 20432 49855 20455
rect 49937 20432 50023 20455
rect 49769 20392 49794 20432
rect 49794 20392 49834 20432
rect 49834 20392 49855 20432
rect 49937 20392 49958 20432
rect 49958 20392 49998 20432
rect 49998 20392 50023 20432
rect 49769 20369 49855 20392
rect 49937 20369 50023 20392
rect 64889 20432 64975 20455
rect 65057 20432 65143 20455
rect 64889 20392 64914 20432
rect 64914 20392 64954 20432
rect 64954 20392 64975 20432
rect 65057 20392 65078 20432
rect 65078 20392 65118 20432
rect 65118 20392 65143 20432
rect 64889 20369 64975 20392
rect 65057 20369 65143 20392
rect 80009 20432 80095 20455
rect 80177 20432 80263 20455
rect 80009 20392 80034 20432
rect 80034 20392 80074 20432
rect 80074 20392 80095 20432
rect 80177 20392 80198 20432
rect 80198 20392 80238 20432
rect 80238 20392 80263 20432
rect 80009 20369 80095 20392
rect 80177 20369 80263 20392
rect 95129 20432 95215 20455
rect 95297 20432 95383 20455
rect 95129 20392 95154 20432
rect 95154 20392 95194 20432
rect 95194 20392 95215 20432
rect 95297 20392 95318 20432
rect 95318 20392 95358 20432
rect 95358 20392 95383 20432
rect 95129 20369 95215 20392
rect 95297 20369 95383 20392
rect 3169 19676 3255 19699
rect 3337 19676 3423 19699
rect 3169 19636 3194 19676
rect 3194 19636 3234 19676
rect 3234 19636 3255 19676
rect 3337 19636 3358 19676
rect 3358 19636 3398 19676
rect 3398 19636 3423 19676
rect 3169 19613 3255 19636
rect 3337 19613 3423 19636
rect 18289 19676 18375 19699
rect 18457 19676 18543 19699
rect 18289 19636 18314 19676
rect 18314 19636 18354 19676
rect 18354 19636 18375 19676
rect 18457 19636 18478 19676
rect 18478 19636 18518 19676
rect 18518 19636 18543 19676
rect 18289 19613 18375 19636
rect 18457 19613 18543 19636
rect 33409 19676 33495 19699
rect 33577 19676 33663 19699
rect 33409 19636 33434 19676
rect 33434 19636 33474 19676
rect 33474 19636 33495 19676
rect 33577 19636 33598 19676
rect 33598 19636 33638 19676
rect 33638 19636 33663 19676
rect 33409 19613 33495 19636
rect 33577 19613 33663 19636
rect 48529 19676 48615 19699
rect 48697 19676 48783 19699
rect 48529 19636 48554 19676
rect 48554 19636 48594 19676
rect 48594 19636 48615 19676
rect 48697 19636 48718 19676
rect 48718 19636 48758 19676
rect 48758 19636 48783 19676
rect 48529 19613 48615 19636
rect 48697 19613 48783 19636
rect 63649 19676 63735 19699
rect 63817 19676 63903 19699
rect 63649 19636 63674 19676
rect 63674 19636 63714 19676
rect 63714 19636 63735 19676
rect 63817 19636 63838 19676
rect 63838 19636 63878 19676
rect 63878 19636 63903 19676
rect 63649 19613 63735 19636
rect 63817 19613 63903 19636
rect 78769 19676 78855 19699
rect 78937 19676 79023 19699
rect 78769 19636 78794 19676
rect 78794 19636 78834 19676
rect 78834 19636 78855 19676
rect 78937 19636 78958 19676
rect 78958 19636 78998 19676
rect 78998 19636 79023 19676
rect 78769 19613 78855 19636
rect 78937 19613 79023 19636
rect 93889 19676 93975 19699
rect 94057 19676 94143 19699
rect 93889 19636 93914 19676
rect 93914 19636 93954 19676
rect 93954 19636 93975 19676
rect 94057 19636 94078 19676
rect 94078 19636 94118 19676
rect 94118 19636 94143 19676
rect 93889 19613 93975 19636
rect 94057 19613 94143 19636
rect 4409 18920 4495 18943
rect 4577 18920 4663 18943
rect 4409 18880 4434 18920
rect 4434 18880 4474 18920
rect 4474 18880 4495 18920
rect 4577 18880 4598 18920
rect 4598 18880 4638 18920
rect 4638 18880 4663 18920
rect 4409 18857 4495 18880
rect 4577 18857 4663 18880
rect 19529 18920 19615 18943
rect 19697 18920 19783 18943
rect 19529 18880 19554 18920
rect 19554 18880 19594 18920
rect 19594 18880 19615 18920
rect 19697 18880 19718 18920
rect 19718 18880 19758 18920
rect 19758 18880 19783 18920
rect 19529 18857 19615 18880
rect 19697 18857 19783 18880
rect 34649 18920 34735 18943
rect 34817 18920 34903 18943
rect 34649 18880 34674 18920
rect 34674 18880 34714 18920
rect 34714 18880 34735 18920
rect 34817 18880 34838 18920
rect 34838 18880 34878 18920
rect 34878 18880 34903 18920
rect 34649 18857 34735 18880
rect 34817 18857 34903 18880
rect 49769 18920 49855 18943
rect 49937 18920 50023 18943
rect 49769 18880 49794 18920
rect 49794 18880 49834 18920
rect 49834 18880 49855 18920
rect 49937 18880 49958 18920
rect 49958 18880 49998 18920
rect 49998 18880 50023 18920
rect 49769 18857 49855 18880
rect 49937 18857 50023 18880
rect 64889 18920 64975 18943
rect 65057 18920 65143 18943
rect 64889 18880 64914 18920
rect 64914 18880 64954 18920
rect 64954 18880 64975 18920
rect 65057 18880 65078 18920
rect 65078 18880 65118 18920
rect 65118 18880 65143 18920
rect 64889 18857 64975 18880
rect 65057 18857 65143 18880
rect 80009 18920 80095 18943
rect 80177 18920 80263 18943
rect 80009 18880 80034 18920
rect 80034 18880 80074 18920
rect 80074 18880 80095 18920
rect 80177 18880 80198 18920
rect 80198 18880 80238 18920
rect 80238 18880 80263 18920
rect 80009 18857 80095 18880
rect 80177 18857 80263 18880
rect 95129 18920 95215 18943
rect 95297 18920 95383 18943
rect 95129 18880 95154 18920
rect 95154 18880 95194 18920
rect 95194 18880 95215 18920
rect 95297 18880 95318 18920
rect 95318 18880 95358 18920
rect 95358 18880 95383 18920
rect 95129 18857 95215 18880
rect 95297 18857 95383 18880
rect 3169 18164 3255 18187
rect 3337 18164 3423 18187
rect 3169 18124 3194 18164
rect 3194 18124 3234 18164
rect 3234 18124 3255 18164
rect 3337 18124 3358 18164
rect 3358 18124 3398 18164
rect 3398 18124 3423 18164
rect 3169 18101 3255 18124
rect 3337 18101 3423 18124
rect 18289 18164 18375 18187
rect 18457 18164 18543 18187
rect 18289 18124 18314 18164
rect 18314 18124 18354 18164
rect 18354 18124 18375 18164
rect 18457 18124 18478 18164
rect 18478 18124 18518 18164
rect 18518 18124 18543 18164
rect 18289 18101 18375 18124
rect 18457 18101 18543 18124
rect 33409 18164 33495 18187
rect 33577 18164 33663 18187
rect 33409 18124 33434 18164
rect 33434 18124 33474 18164
rect 33474 18124 33495 18164
rect 33577 18124 33598 18164
rect 33598 18124 33638 18164
rect 33638 18124 33663 18164
rect 33409 18101 33495 18124
rect 33577 18101 33663 18124
rect 48529 18164 48615 18187
rect 48697 18164 48783 18187
rect 48529 18124 48554 18164
rect 48554 18124 48594 18164
rect 48594 18124 48615 18164
rect 48697 18124 48718 18164
rect 48718 18124 48758 18164
rect 48758 18124 48783 18164
rect 48529 18101 48615 18124
rect 48697 18101 48783 18124
rect 63649 18164 63735 18187
rect 63817 18164 63903 18187
rect 63649 18124 63674 18164
rect 63674 18124 63714 18164
rect 63714 18124 63735 18164
rect 63817 18124 63838 18164
rect 63838 18124 63878 18164
rect 63878 18124 63903 18164
rect 63649 18101 63735 18124
rect 63817 18101 63903 18124
rect 78769 18164 78855 18187
rect 78937 18164 79023 18187
rect 78769 18124 78794 18164
rect 78794 18124 78834 18164
rect 78834 18124 78855 18164
rect 78937 18124 78958 18164
rect 78958 18124 78998 18164
rect 78998 18124 79023 18164
rect 78769 18101 78855 18124
rect 78937 18101 79023 18124
rect 93889 18164 93975 18187
rect 94057 18164 94143 18187
rect 93889 18124 93914 18164
rect 93914 18124 93954 18164
rect 93954 18124 93975 18164
rect 94057 18124 94078 18164
rect 94078 18124 94118 18164
rect 94118 18124 94143 18164
rect 93889 18101 93975 18124
rect 94057 18101 94143 18124
rect 4409 17408 4495 17431
rect 4577 17408 4663 17431
rect 4409 17368 4434 17408
rect 4434 17368 4474 17408
rect 4474 17368 4495 17408
rect 4577 17368 4598 17408
rect 4598 17368 4638 17408
rect 4638 17368 4663 17408
rect 4409 17345 4495 17368
rect 4577 17345 4663 17368
rect 19529 17408 19615 17431
rect 19697 17408 19783 17431
rect 19529 17368 19554 17408
rect 19554 17368 19594 17408
rect 19594 17368 19615 17408
rect 19697 17368 19718 17408
rect 19718 17368 19758 17408
rect 19758 17368 19783 17408
rect 19529 17345 19615 17368
rect 19697 17345 19783 17368
rect 34649 17408 34735 17431
rect 34817 17408 34903 17431
rect 34649 17368 34674 17408
rect 34674 17368 34714 17408
rect 34714 17368 34735 17408
rect 34817 17368 34838 17408
rect 34838 17368 34878 17408
rect 34878 17368 34903 17408
rect 34649 17345 34735 17368
rect 34817 17345 34903 17368
rect 49769 17408 49855 17431
rect 49937 17408 50023 17431
rect 49769 17368 49794 17408
rect 49794 17368 49834 17408
rect 49834 17368 49855 17408
rect 49937 17368 49958 17408
rect 49958 17368 49998 17408
rect 49998 17368 50023 17408
rect 49769 17345 49855 17368
rect 49937 17345 50023 17368
rect 64889 17408 64975 17431
rect 65057 17408 65143 17431
rect 64889 17368 64914 17408
rect 64914 17368 64954 17408
rect 64954 17368 64975 17408
rect 65057 17368 65078 17408
rect 65078 17368 65118 17408
rect 65118 17368 65143 17408
rect 64889 17345 64975 17368
rect 65057 17345 65143 17368
rect 80009 17408 80095 17431
rect 80177 17408 80263 17431
rect 80009 17368 80034 17408
rect 80034 17368 80074 17408
rect 80074 17368 80095 17408
rect 80177 17368 80198 17408
rect 80198 17368 80238 17408
rect 80238 17368 80263 17408
rect 80009 17345 80095 17368
rect 80177 17345 80263 17368
rect 95129 17408 95215 17431
rect 95297 17408 95383 17431
rect 95129 17368 95154 17408
rect 95154 17368 95194 17408
rect 95194 17368 95215 17408
rect 95297 17368 95318 17408
rect 95318 17368 95358 17408
rect 95358 17368 95383 17408
rect 95129 17345 95215 17368
rect 95297 17345 95383 17368
rect 3169 16652 3255 16675
rect 3337 16652 3423 16675
rect 3169 16612 3194 16652
rect 3194 16612 3234 16652
rect 3234 16612 3255 16652
rect 3337 16612 3358 16652
rect 3358 16612 3398 16652
rect 3398 16612 3423 16652
rect 3169 16589 3255 16612
rect 3337 16589 3423 16612
rect 18289 16652 18375 16675
rect 18457 16652 18543 16675
rect 18289 16612 18314 16652
rect 18314 16612 18354 16652
rect 18354 16612 18375 16652
rect 18457 16612 18478 16652
rect 18478 16612 18518 16652
rect 18518 16612 18543 16652
rect 18289 16589 18375 16612
rect 18457 16589 18543 16612
rect 33409 16652 33495 16675
rect 33577 16652 33663 16675
rect 33409 16612 33434 16652
rect 33434 16612 33474 16652
rect 33474 16612 33495 16652
rect 33577 16612 33598 16652
rect 33598 16612 33638 16652
rect 33638 16612 33663 16652
rect 33409 16589 33495 16612
rect 33577 16589 33663 16612
rect 48529 16652 48615 16675
rect 48697 16652 48783 16675
rect 48529 16612 48554 16652
rect 48554 16612 48594 16652
rect 48594 16612 48615 16652
rect 48697 16612 48718 16652
rect 48718 16612 48758 16652
rect 48758 16612 48783 16652
rect 48529 16589 48615 16612
rect 48697 16589 48783 16612
rect 63649 16652 63735 16675
rect 63817 16652 63903 16675
rect 63649 16612 63674 16652
rect 63674 16612 63714 16652
rect 63714 16612 63735 16652
rect 63817 16612 63838 16652
rect 63838 16612 63878 16652
rect 63878 16612 63903 16652
rect 63649 16589 63735 16612
rect 63817 16589 63903 16612
rect 78769 16652 78855 16675
rect 78937 16652 79023 16675
rect 78769 16612 78794 16652
rect 78794 16612 78834 16652
rect 78834 16612 78855 16652
rect 78937 16612 78958 16652
rect 78958 16612 78998 16652
rect 78998 16612 79023 16652
rect 78769 16589 78855 16612
rect 78937 16589 79023 16612
rect 93889 16652 93975 16675
rect 94057 16652 94143 16675
rect 93889 16612 93914 16652
rect 93914 16612 93954 16652
rect 93954 16612 93975 16652
rect 94057 16612 94078 16652
rect 94078 16612 94118 16652
rect 94118 16612 94143 16652
rect 93889 16589 93975 16612
rect 94057 16589 94143 16612
rect 4409 15896 4495 15919
rect 4577 15896 4663 15919
rect 4409 15856 4434 15896
rect 4434 15856 4474 15896
rect 4474 15856 4495 15896
rect 4577 15856 4598 15896
rect 4598 15856 4638 15896
rect 4638 15856 4663 15896
rect 4409 15833 4495 15856
rect 4577 15833 4663 15856
rect 19529 15896 19615 15919
rect 19697 15896 19783 15919
rect 19529 15856 19554 15896
rect 19554 15856 19594 15896
rect 19594 15856 19615 15896
rect 19697 15856 19718 15896
rect 19718 15856 19758 15896
rect 19758 15856 19783 15896
rect 19529 15833 19615 15856
rect 19697 15833 19783 15856
rect 34649 15896 34735 15919
rect 34817 15896 34903 15919
rect 34649 15856 34674 15896
rect 34674 15856 34714 15896
rect 34714 15856 34735 15896
rect 34817 15856 34838 15896
rect 34838 15856 34878 15896
rect 34878 15856 34903 15896
rect 34649 15833 34735 15856
rect 34817 15833 34903 15856
rect 49769 15896 49855 15919
rect 49937 15896 50023 15919
rect 49769 15856 49794 15896
rect 49794 15856 49834 15896
rect 49834 15856 49855 15896
rect 49937 15856 49958 15896
rect 49958 15856 49998 15896
rect 49998 15856 50023 15896
rect 49769 15833 49855 15856
rect 49937 15833 50023 15856
rect 64889 15896 64975 15919
rect 65057 15896 65143 15919
rect 64889 15856 64914 15896
rect 64914 15856 64954 15896
rect 64954 15856 64975 15896
rect 65057 15856 65078 15896
rect 65078 15856 65118 15896
rect 65118 15856 65143 15896
rect 64889 15833 64975 15856
rect 65057 15833 65143 15856
rect 80009 15896 80095 15919
rect 80177 15896 80263 15919
rect 80009 15856 80034 15896
rect 80034 15856 80074 15896
rect 80074 15856 80095 15896
rect 80177 15856 80198 15896
rect 80198 15856 80238 15896
rect 80238 15856 80263 15896
rect 80009 15833 80095 15856
rect 80177 15833 80263 15856
rect 95129 15896 95215 15919
rect 95297 15896 95383 15919
rect 95129 15856 95154 15896
rect 95154 15856 95194 15896
rect 95194 15856 95215 15896
rect 95297 15856 95318 15896
rect 95318 15856 95358 15896
rect 95358 15856 95383 15896
rect 95129 15833 95215 15856
rect 95297 15833 95383 15856
rect 3169 15140 3255 15163
rect 3337 15140 3423 15163
rect 3169 15100 3194 15140
rect 3194 15100 3234 15140
rect 3234 15100 3255 15140
rect 3337 15100 3358 15140
rect 3358 15100 3398 15140
rect 3398 15100 3423 15140
rect 3169 15077 3255 15100
rect 3337 15077 3423 15100
rect 18289 15140 18375 15163
rect 18457 15140 18543 15163
rect 18289 15100 18314 15140
rect 18314 15100 18354 15140
rect 18354 15100 18375 15140
rect 18457 15100 18478 15140
rect 18478 15100 18518 15140
rect 18518 15100 18543 15140
rect 18289 15077 18375 15100
rect 18457 15077 18543 15100
rect 33409 15140 33495 15163
rect 33577 15140 33663 15163
rect 33409 15100 33434 15140
rect 33434 15100 33474 15140
rect 33474 15100 33495 15140
rect 33577 15100 33598 15140
rect 33598 15100 33638 15140
rect 33638 15100 33663 15140
rect 33409 15077 33495 15100
rect 33577 15077 33663 15100
rect 48529 15140 48615 15163
rect 48697 15140 48783 15163
rect 48529 15100 48554 15140
rect 48554 15100 48594 15140
rect 48594 15100 48615 15140
rect 48697 15100 48718 15140
rect 48718 15100 48758 15140
rect 48758 15100 48783 15140
rect 48529 15077 48615 15100
rect 48697 15077 48783 15100
rect 63649 15140 63735 15163
rect 63817 15140 63903 15163
rect 63649 15100 63674 15140
rect 63674 15100 63714 15140
rect 63714 15100 63735 15140
rect 63817 15100 63838 15140
rect 63838 15100 63878 15140
rect 63878 15100 63903 15140
rect 63649 15077 63735 15100
rect 63817 15077 63903 15100
rect 78769 15140 78855 15163
rect 78937 15140 79023 15163
rect 78769 15100 78794 15140
rect 78794 15100 78834 15140
rect 78834 15100 78855 15140
rect 78937 15100 78958 15140
rect 78958 15100 78998 15140
rect 78998 15100 79023 15140
rect 78769 15077 78855 15100
rect 78937 15077 79023 15100
rect 93889 15140 93975 15163
rect 94057 15140 94143 15163
rect 93889 15100 93914 15140
rect 93914 15100 93954 15140
rect 93954 15100 93975 15140
rect 94057 15100 94078 15140
rect 94078 15100 94118 15140
rect 94118 15100 94143 15140
rect 93889 15077 93975 15100
rect 94057 15077 94143 15100
rect 4409 14384 4495 14407
rect 4577 14384 4663 14407
rect 4409 14344 4434 14384
rect 4434 14344 4474 14384
rect 4474 14344 4495 14384
rect 4577 14344 4598 14384
rect 4598 14344 4638 14384
rect 4638 14344 4663 14384
rect 4409 14321 4495 14344
rect 4577 14321 4663 14344
rect 19529 14384 19615 14407
rect 19697 14384 19783 14407
rect 19529 14344 19554 14384
rect 19554 14344 19594 14384
rect 19594 14344 19615 14384
rect 19697 14344 19718 14384
rect 19718 14344 19758 14384
rect 19758 14344 19783 14384
rect 19529 14321 19615 14344
rect 19697 14321 19783 14344
rect 34649 14384 34735 14407
rect 34817 14384 34903 14407
rect 34649 14344 34674 14384
rect 34674 14344 34714 14384
rect 34714 14344 34735 14384
rect 34817 14344 34838 14384
rect 34838 14344 34878 14384
rect 34878 14344 34903 14384
rect 34649 14321 34735 14344
rect 34817 14321 34903 14344
rect 49769 14384 49855 14407
rect 49937 14384 50023 14407
rect 49769 14344 49794 14384
rect 49794 14344 49834 14384
rect 49834 14344 49855 14384
rect 49937 14344 49958 14384
rect 49958 14344 49998 14384
rect 49998 14344 50023 14384
rect 49769 14321 49855 14344
rect 49937 14321 50023 14344
rect 64889 14384 64975 14407
rect 65057 14384 65143 14407
rect 64889 14344 64914 14384
rect 64914 14344 64954 14384
rect 64954 14344 64975 14384
rect 65057 14344 65078 14384
rect 65078 14344 65118 14384
rect 65118 14344 65143 14384
rect 64889 14321 64975 14344
rect 65057 14321 65143 14344
rect 80009 14384 80095 14407
rect 80177 14384 80263 14407
rect 80009 14344 80034 14384
rect 80034 14344 80074 14384
rect 80074 14344 80095 14384
rect 80177 14344 80198 14384
rect 80198 14344 80238 14384
rect 80238 14344 80263 14384
rect 80009 14321 80095 14344
rect 80177 14321 80263 14344
rect 95129 14384 95215 14407
rect 95297 14384 95383 14407
rect 95129 14344 95154 14384
rect 95154 14344 95194 14384
rect 95194 14344 95215 14384
rect 95297 14344 95318 14384
rect 95318 14344 95358 14384
rect 95358 14344 95383 14384
rect 95129 14321 95215 14344
rect 95297 14321 95383 14344
rect 3169 13628 3255 13651
rect 3337 13628 3423 13651
rect 3169 13588 3194 13628
rect 3194 13588 3234 13628
rect 3234 13588 3255 13628
rect 3337 13588 3358 13628
rect 3358 13588 3398 13628
rect 3398 13588 3423 13628
rect 3169 13565 3255 13588
rect 3337 13565 3423 13588
rect 18289 13628 18375 13651
rect 18457 13628 18543 13651
rect 18289 13588 18314 13628
rect 18314 13588 18354 13628
rect 18354 13588 18375 13628
rect 18457 13588 18478 13628
rect 18478 13588 18518 13628
rect 18518 13588 18543 13628
rect 18289 13565 18375 13588
rect 18457 13565 18543 13588
rect 33409 13628 33495 13651
rect 33577 13628 33663 13651
rect 33409 13588 33434 13628
rect 33434 13588 33474 13628
rect 33474 13588 33495 13628
rect 33577 13588 33598 13628
rect 33598 13588 33638 13628
rect 33638 13588 33663 13628
rect 33409 13565 33495 13588
rect 33577 13565 33663 13588
rect 48529 13628 48615 13651
rect 48697 13628 48783 13651
rect 48529 13588 48554 13628
rect 48554 13588 48594 13628
rect 48594 13588 48615 13628
rect 48697 13588 48718 13628
rect 48718 13588 48758 13628
rect 48758 13588 48783 13628
rect 48529 13565 48615 13588
rect 48697 13565 48783 13588
rect 63649 13628 63735 13651
rect 63817 13628 63903 13651
rect 63649 13588 63674 13628
rect 63674 13588 63714 13628
rect 63714 13588 63735 13628
rect 63817 13588 63838 13628
rect 63838 13588 63878 13628
rect 63878 13588 63903 13628
rect 63649 13565 63735 13588
rect 63817 13565 63903 13588
rect 78769 13628 78855 13651
rect 78937 13628 79023 13651
rect 78769 13588 78794 13628
rect 78794 13588 78834 13628
rect 78834 13588 78855 13628
rect 78937 13588 78958 13628
rect 78958 13588 78998 13628
rect 78998 13588 79023 13628
rect 78769 13565 78855 13588
rect 78937 13565 79023 13588
rect 93889 13628 93975 13651
rect 94057 13628 94143 13651
rect 93889 13588 93914 13628
rect 93914 13588 93954 13628
rect 93954 13588 93975 13628
rect 94057 13588 94078 13628
rect 94078 13588 94118 13628
rect 94118 13588 94143 13628
rect 93889 13565 93975 13588
rect 94057 13565 94143 13588
rect 4409 12872 4495 12895
rect 4577 12872 4663 12895
rect 4409 12832 4434 12872
rect 4434 12832 4474 12872
rect 4474 12832 4495 12872
rect 4577 12832 4598 12872
rect 4598 12832 4638 12872
rect 4638 12832 4663 12872
rect 4409 12809 4495 12832
rect 4577 12809 4663 12832
rect 19529 12872 19615 12895
rect 19697 12872 19783 12895
rect 19529 12832 19554 12872
rect 19554 12832 19594 12872
rect 19594 12832 19615 12872
rect 19697 12832 19718 12872
rect 19718 12832 19758 12872
rect 19758 12832 19783 12872
rect 19529 12809 19615 12832
rect 19697 12809 19783 12832
rect 34649 12872 34735 12895
rect 34817 12872 34903 12895
rect 34649 12832 34674 12872
rect 34674 12832 34714 12872
rect 34714 12832 34735 12872
rect 34817 12832 34838 12872
rect 34838 12832 34878 12872
rect 34878 12832 34903 12872
rect 34649 12809 34735 12832
rect 34817 12809 34903 12832
rect 49769 12872 49855 12895
rect 49937 12872 50023 12895
rect 49769 12832 49794 12872
rect 49794 12832 49834 12872
rect 49834 12832 49855 12872
rect 49937 12832 49958 12872
rect 49958 12832 49998 12872
rect 49998 12832 50023 12872
rect 49769 12809 49855 12832
rect 49937 12809 50023 12832
rect 64889 12872 64975 12895
rect 65057 12872 65143 12895
rect 64889 12832 64914 12872
rect 64914 12832 64954 12872
rect 64954 12832 64975 12872
rect 65057 12832 65078 12872
rect 65078 12832 65118 12872
rect 65118 12832 65143 12872
rect 64889 12809 64975 12832
rect 65057 12809 65143 12832
rect 80009 12872 80095 12895
rect 80177 12872 80263 12895
rect 80009 12832 80034 12872
rect 80034 12832 80074 12872
rect 80074 12832 80095 12872
rect 80177 12832 80198 12872
rect 80198 12832 80238 12872
rect 80238 12832 80263 12872
rect 80009 12809 80095 12832
rect 80177 12809 80263 12832
rect 95129 12872 95215 12895
rect 95297 12872 95383 12895
rect 95129 12832 95154 12872
rect 95154 12832 95194 12872
rect 95194 12832 95215 12872
rect 95297 12832 95318 12872
rect 95318 12832 95358 12872
rect 95358 12832 95383 12872
rect 95129 12809 95215 12832
rect 95297 12809 95383 12832
rect 3169 12116 3255 12139
rect 3337 12116 3423 12139
rect 3169 12076 3194 12116
rect 3194 12076 3234 12116
rect 3234 12076 3255 12116
rect 3337 12076 3358 12116
rect 3358 12076 3398 12116
rect 3398 12076 3423 12116
rect 3169 12053 3255 12076
rect 3337 12053 3423 12076
rect 18289 12116 18375 12139
rect 18457 12116 18543 12139
rect 18289 12076 18314 12116
rect 18314 12076 18354 12116
rect 18354 12076 18375 12116
rect 18457 12076 18478 12116
rect 18478 12076 18518 12116
rect 18518 12076 18543 12116
rect 18289 12053 18375 12076
rect 18457 12053 18543 12076
rect 33409 12116 33495 12139
rect 33577 12116 33663 12139
rect 33409 12076 33434 12116
rect 33434 12076 33474 12116
rect 33474 12076 33495 12116
rect 33577 12076 33598 12116
rect 33598 12076 33638 12116
rect 33638 12076 33663 12116
rect 33409 12053 33495 12076
rect 33577 12053 33663 12076
rect 48529 12116 48615 12139
rect 48697 12116 48783 12139
rect 48529 12076 48554 12116
rect 48554 12076 48594 12116
rect 48594 12076 48615 12116
rect 48697 12076 48718 12116
rect 48718 12076 48758 12116
rect 48758 12076 48783 12116
rect 48529 12053 48615 12076
rect 48697 12053 48783 12076
rect 63649 12116 63735 12139
rect 63817 12116 63903 12139
rect 63649 12076 63674 12116
rect 63674 12076 63714 12116
rect 63714 12076 63735 12116
rect 63817 12076 63838 12116
rect 63838 12076 63878 12116
rect 63878 12076 63903 12116
rect 63649 12053 63735 12076
rect 63817 12053 63903 12076
rect 78769 12116 78855 12139
rect 78937 12116 79023 12139
rect 78769 12076 78794 12116
rect 78794 12076 78834 12116
rect 78834 12076 78855 12116
rect 78937 12076 78958 12116
rect 78958 12076 78998 12116
rect 78998 12076 79023 12116
rect 78769 12053 78855 12076
rect 78937 12053 79023 12076
rect 93889 12116 93975 12139
rect 94057 12116 94143 12139
rect 93889 12076 93914 12116
rect 93914 12076 93954 12116
rect 93954 12076 93975 12116
rect 94057 12076 94078 12116
rect 94078 12076 94118 12116
rect 94118 12076 94143 12116
rect 93889 12053 93975 12076
rect 94057 12053 94143 12076
rect 4409 11360 4495 11383
rect 4577 11360 4663 11383
rect 4409 11320 4434 11360
rect 4434 11320 4474 11360
rect 4474 11320 4495 11360
rect 4577 11320 4598 11360
rect 4598 11320 4638 11360
rect 4638 11320 4663 11360
rect 4409 11297 4495 11320
rect 4577 11297 4663 11320
rect 19529 11360 19615 11383
rect 19697 11360 19783 11383
rect 19529 11320 19554 11360
rect 19554 11320 19594 11360
rect 19594 11320 19615 11360
rect 19697 11320 19718 11360
rect 19718 11320 19758 11360
rect 19758 11320 19783 11360
rect 19529 11297 19615 11320
rect 19697 11297 19783 11320
rect 34649 11360 34735 11383
rect 34817 11360 34903 11383
rect 34649 11320 34674 11360
rect 34674 11320 34714 11360
rect 34714 11320 34735 11360
rect 34817 11320 34838 11360
rect 34838 11320 34878 11360
rect 34878 11320 34903 11360
rect 34649 11297 34735 11320
rect 34817 11297 34903 11320
rect 49769 11360 49855 11383
rect 49937 11360 50023 11383
rect 49769 11320 49794 11360
rect 49794 11320 49834 11360
rect 49834 11320 49855 11360
rect 49937 11320 49958 11360
rect 49958 11320 49998 11360
rect 49998 11320 50023 11360
rect 49769 11297 49855 11320
rect 49937 11297 50023 11320
rect 64889 11360 64975 11383
rect 65057 11360 65143 11383
rect 64889 11320 64914 11360
rect 64914 11320 64954 11360
rect 64954 11320 64975 11360
rect 65057 11320 65078 11360
rect 65078 11320 65118 11360
rect 65118 11320 65143 11360
rect 64889 11297 64975 11320
rect 65057 11297 65143 11320
rect 80009 11360 80095 11383
rect 80177 11360 80263 11383
rect 80009 11320 80034 11360
rect 80034 11320 80074 11360
rect 80074 11320 80095 11360
rect 80177 11320 80198 11360
rect 80198 11320 80238 11360
rect 80238 11320 80263 11360
rect 80009 11297 80095 11320
rect 80177 11297 80263 11320
rect 95129 11360 95215 11383
rect 95297 11360 95383 11383
rect 95129 11320 95154 11360
rect 95154 11320 95194 11360
rect 95194 11320 95215 11360
rect 95297 11320 95318 11360
rect 95318 11320 95358 11360
rect 95358 11320 95383 11360
rect 95129 11297 95215 11320
rect 95297 11297 95383 11320
rect 3169 10604 3255 10627
rect 3337 10604 3423 10627
rect 3169 10564 3194 10604
rect 3194 10564 3234 10604
rect 3234 10564 3255 10604
rect 3337 10564 3358 10604
rect 3358 10564 3398 10604
rect 3398 10564 3423 10604
rect 3169 10541 3255 10564
rect 3337 10541 3423 10564
rect 18289 10604 18375 10627
rect 18457 10604 18543 10627
rect 18289 10564 18314 10604
rect 18314 10564 18354 10604
rect 18354 10564 18375 10604
rect 18457 10564 18478 10604
rect 18478 10564 18518 10604
rect 18518 10564 18543 10604
rect 18289 10541 18375 10564
rect 18457 10541 18543 10564
rect 33409 10604 33495 10627
rect 33577 10604 33663 10627
rect 33409 10564 33434 10604
rect 33434 10564 33474 10604
rect 33474 10564 33495 10604
rect 33577 10564 33598 10604
rect 33598 10564 33638 10604
rect 33638 10564 33663 10604
rect 33409 10541 33495 10564
rect 33577 10541 33663 10564
rect 48529 10604 48615 10627
rect 48697 10604 48783 10627
rect 48529 10564 48554 10604
rect 48554 10564 48594 10604
rect 48594 10564 48615 10604
rect 48697 10564 48718 10604
rect 48718 10564 48758 10604
rect 48758 10564 48783 10604
rect 48529 10541 48615 10564
rect 48697 10541 48783 10564
rect 63649 10604 63735 10627
rect 63817 10604 63903 10627
rect 63649 10564 63674 10604
rect 63674 10564 63714 10604
rect 63714 10564 63735 10604
rect 63817 10564 63838 10604
rect 63838 10564 63878 10604
rect 63878 10564 63903 10604
rect 63649 10541 63735 10564
rect 63817 10541 63903 10564
rect 78769 10604 78855 10627
rect 78937 10604 79023 10627
rect 78769 10564 78794 10604
rect 78794 10564 78834 10604
rect 78834 10564 78855 10604
rect 78937 10564 78958 10604
rect 78958 10564 78998 10604
rect 78998 10564 79023 10604
rect 78769 10541 78855 10564
rect 78937 10541 79023 10564
rect 93889 10604 93975 10627
rect 94057 10604 94143 10627
rect 93889 10564 93914 10604
rect 93914 10564 93954 10604
rect 93954 10564 93975 10604
rect 94057 10564 94078 10604
rect 94078 10564 94118 10604
rect 94118 10564 94143 10604
rect 93889 10541 93975 10564
rect 94057 10541 94143 10564
rect 4409 9848 4495 9871
rect 4577 9848 4663 9871
rect 4409 9808 4434 9848
rect 4434 9808 4474 9848
rect 4474 9808 4495 9848
rect 4577 9808 4598 9848
rect 4598 9808 4638 9848
rect 4638 9808 4663 9848
rect 4409 9785 4495 9808
rect 4577 9785 4663 9808
rect 19529 9848 19615 9871
rect 19697 9848 19783 9871
rect 19529 9808 19554 9848
rect 19554 9808 19594 9848
rect 19594 9808 19615 9848
rect 19697 9808 19718 9848
rect 19718 9808 19758 9848
rect 19758 9808 19783 9848
rect 19529 9785 19615 9808
rect 19697 9785 19783 9808
rect 34649 9848 34735 9871
rect 34817 9848 34903 9871
rect 34649 9808 34674 9848
rect 34674 9808 34714 9848
rect 34714 9808 34735 9848
rect 34817 9808 34838 9848
rect 34838 9808 34878 9848
rect 34878 9808 34903 9848
rect 34649 9785 34735 9808
rect 34817 9785 34903 9808
rect 49769 9848 49855 9871
rect 49937 9848 50023 9871
rect 49769 9808 49794 9848
rect 49794 9808 49834 9848
rect 49834 9808 49855 9848
rect 49937 9808 49958 9848
rect 49958 9808 49998 9848
rect 49998 9808 50023 9848
rect 49769 9785 49855 9808
rect 49937 9785 50023 9808
rect 64889 9848 64975 9871
rect 65057 9848 65143 9871
rect 64889 9808 64914 9848
rect 64914 9808 64954 9848
rect 64954 9808 64975 9848
rect 65057 9808 65078 9848
rect 65078 9808 65118 9848
rect 65118 9808 65143 9848
rect 64889 9785 64975 9808
rect 65057 9785 65143 9808
rect 80009 9848 80095 9871
rect 80177 9848 80263 9871
rect 80009 9808 80034 9848
rect 80034 9808 80074 9848
rect 80074 9808 80095 9848
rect 80177 9808 80198 9848
rect 80198 9808 80238 9848
rect 80238 9808 80263 9848
rect 80009 9785 80095 9808
rect 80177 9785 80263 9808
rect 95129 9848 95215 9871
rect 95297 9848 95383 9871
rect 95129 9808 95154 9848
rect 95154 9808 95194 9848
rect 95194 9808 95215 9848
rect 95297 9808 95318 9848
rect 95318 9808 95358 9848
rect 95358 9808 95383 9848
rect 95129 9785 95215 9808
rect 95297 9785 95383 9808
rect 3169 9092 3255 9115
rect 3337 9092 3423 9115
rect 3169 9052 3194 9092
rect 3194 9052 3234 9092
rect 3234 9052 3255 9092
rect 3337 9052 3358 9092
rect 3358 9052 3398 9092
rect 3398 9052 3423 9092
rect 3169 9029 3255 9052
rect 3337 9029 3423 9052
rect 18289 9092 18375 9115
rect 18457 9092 18543 9115
rect 18289 9052 18314 9092
rect 18314 9052 18354 9092
rect 18354 9052 18375 9092
rect 18457 9052 18478 9092
rect 18478 9052 18518 9092
rect 18518 9052 18543 9092
rect 18289 9029 18375 9052
rect 18457 9029 18543 9052
rect 33409 9092 33495 9115
rect 33577 9092 33663 9115
rect 33409 9052 33434 9092
rect 33434 9052 33474 9092
rect 33474 9052 33495 9092
rect 33577 9052 33598 9092
rect 33598 9052 33638 9092
rect 33638 9052 33663 9092
rect 33409 9029 33495 9052
rect 33577 9029 33663 9052
rect 48529 9092 48615 9115
rect 48697 9092 48783 9115
rect 48529 9052 48554 9092
rect 48554 9052 48594 9092
rect 48594 9052 48615 9092
rect 48697 9052 48718 9092
rect 48718 9052 48758 9092
rect 48758 9052 48783 9092
rect 48529 9029 48615 9052
rect 48697 9029 48783 9052
rect 63649 9092 63735 9115
rect 63817 9092 63903 9115
rect 63649 9052 63674 9092
rect 63674 9052 63714 9092
rect 63714 9052 63735 9092
rect 63817 9052 63838 9092
rect 63838 9052 63878 9092
rect 63878 9052 63903 9092
rect 63649 9029 63735 9052
rect 63817 9029 63903 9052
rect 78769 9092 78855 9115
rect 78937 9092 79023 9115
rect 78769 9052 78794 9092
rect 78794 9052 78834 9092
rect 78834 9052 78855 9092
rect 78937 9052 78958 9092
rect 78958 9052 78998 9092
rect 78998 9052 79023 9092
rect 78769 9029 78855 9052
rect 78937 9029 79023 9052
rect 93889 9092 93975 9115
rect 94057 9092 94143 9115
rect 93889 9052 93914 9092
rect 93914 9052 93954 9092
rect 93954 9052 93975 9092
rect 94057 9052 94078 9092
rect 94078 9052 94118 9092
rect 94118 9052 94143 9092
rect 93889 9029 93975 9052
rect 94057 9029 94143 9052
rect 4409 8336 4495 8359
rect 4577 8336 4663 8359
rect 4409 8296 4434 8336
rect 4434 8296 4474 8336
rect 4474 8296 4495 8336
rect 4577 8296 4598 8336
rect 4598 8296 4638 8336
rect 4638 8296 4663 8336
rect 4409 8273 4495 8296
rect 4577 8273 4663 8296
rect 19529 8336 19615 8359
rect 19697 8336 19783 8359
rect 19529 8296 19554 8336
rect 19554 8296 19594 8336
rect 19594 8296 19615 8336
rect 19697 8296 19718 8336
rect 19718 8296 19758 8336
rect 19758 8296 19783 8336
rect 19529 8273 19615 8296
rect 19697 8273 19783 8296
rect 34649 8336 34735 8359
rect 34817 8336 34903 8359
rect 34649 8296 34674 8336
rect 34674 8296 34714 8336
rect 34714 8296 34735 8336
rect 34817 8296 34838 8336
rect 34838 8296 34878 8336
rect 34878 8296 34903 8336
rect 34649 8273 34735 8296
rect 34817 8273 34903 8296
rect 49769 8336 49855 8359
rect 49937 8336 50023 8359
rect 49769 8296 49794 8336
rect 49794 8296 49834 8336
rect 49834 8296 49855 8336
rect 49937 8296 49958 8336
rect 49958 8296 49998 8336
rect 49998 8296 50023 8336
rect 49769 8273 49855 8296
rect 49937 8273 50023 8296
rect 64889 8336 64975 8359
rect 65057 8336 65143 8359
rect 64889 8296 64914 8336
rect 64914 8296 64954 8336
rect 64954 8296 64975 8336
rect 65057 8296 65078 8336
rect 65078 8296 65118 8336
rect 65118 8296 65143 8336
rect 64889 8273 64975 8296
rect 65057 8273 65143 8296
rect 80009 8336 80095 8359
rect 80177 8336 80263 8359
rect 80009 8296 80034 8336
rect 80034 8296 80074 8336
rect 80074 8296 80095 8336
rect 80177 8296 80198 8336
rect 80198 8296 80238 8336
rect 80238 8296 80263 8336
rect 80009 8273 80095 8296
rect 80177 8273 80263 8296
rect 95129 8336 95215 8359
rect 95297 8336 95383 8359
rect 95129 8296 95154 8336
rect 95154 8296 95194 8336
rect 95194 8296 95215 8336
rect 95297 8296 95318 8336
rect 95318 8296 95358 8336
rect 95358 8296 95383 8336
rect 95129 8273 95215 8296
rect 95297 8273 95383 8296
rect 3169 7580 3255 7603
rect 3337 7580 3423 7603
rect 3169 7540 3194 7580
rect 3194 7540 3234 7580
rect 3234 7540 3255 7580
rect 3337 7540 3358 7580
rect 3358 7540 3398 7580
rect 3398 7540 3423 7580
rect 3169 7517 3255 7540
rect 3337 7517 3423 7540
rect 18289 7580 18375 7603
rect 18457 7580 18543 7603
rect 18289 7540 18314 7580
rect 18314 7540 18354 7580
rect 18354 7540 18375 7580
rect 18457 7540 18478 7580
rect 18478 7540 18518 7580
rect 18518 7540 18543 7580
rect 18289 7517 18375 7540
rect 18457 7517 18543 7540
rect 33409 7580 33495 7603
rect 33577 7580 33663 7603
rect 33409 7540 33434 7580
rect 33434 7540 33474 7580
rect 33474 7540 33495 7580
rect 33577 7540 33598 7580
rect 33598 7540 33638 7580
rect 33638 7540 33663 7580
rect 33409 7517 33495 7540
rect 33577 7517 33663 7540
rect 48529 7580 48615 7603
rect 48697 7580 48783 7603
rect 48529 7540 48554 7580
rect 48554 7540 48594 7580
rect 48594 7540 48615 7580
rect 48697 7540 48718 7580
rect 48718 7540 48758 7580
rect 48758 7540 48783 7580
rect 48529 7517 48615 7540
rect 48697 7517 48783 7540
rect 63649 7580 63735 7603
rect 63817 7580 63903 7603
rect 63649 7540 63674 7580
rect 63674 7540 63714 7580
rect 63714 7540 63735 7580
rect 63817 7540 63838 7580
rect 63838 7540 63878 7580
rect 63878 7540 63903 7580
rect 63649 7517 63735 7540
rect 63817 7517 63903 7540
rect 78769 7580 78855 7603
rect 78937 7580 79023 7603
rect 78769 7540 78794 7580
rect 78794 7540 78834 7580
rect 78834 7540 78855 7580
rect 78937 7540 78958 7580
rect 78958 7540 78998 7580
rect 78998 7540 79023 7580
rect 78769 7517 78855 7540
rect 78937 7517 79023 7540
rect 93889 7580 93975 7603
rect 94057 7580 94143 7603
rect 93889 7540 93914 7580
rect 93914 7540 93954 7580
rect 93954 7540 93975 7580
rect 94057 7540 94078 7580
rect 94078 7540 94118 7580
rect 94118 7540 94143 7580
rect 93889 7517 93975 7540
rect 94057 7517 94143 7540
rect 4409 6824 4495 6847
rect 4577 6824 4663 6847
rect 4409 6784 4434 6824
rect 4434 6784 4474 6824
rect 4474 6784 4495 6824
rect 4577 6784 4598 6824
rect 4598 6784 4638 6824
rect 4638 6784 4663 6824
rect 4409 6761 4495 6784
rect 4577 6761 4663 6784
rect 19529 6824 19615 6847
rect 19697 6824 19783 6847
rect 19529 6784 19554 6824
rect 19554 6784 19594 6824
rect 19594 6784 19615 6824
rect 19697 6784 19718 6824
rect 19718 6784 19758 6824
rect 19758 6784 19783 6824
rect 19529 6761 19615 6784
rect 19697 6761 19783 6784
rect 34649 6824 34735 6847
rect 34817 6824 34903 6847
rect 34649 6784 34674 6824
rect 34674 6784 34714 6824
rect 34714 6784 34735 6824
rect 34817 6784 34838 6824
rect 34838 6784 34878 6824
rect 34878 6784 34903 6824
rect 34649 6761 34735 6784
rect 34817 6761 34903 6784
rect 49769 6824 49855 6847
rect 49937 6824 50023 6847
rect 49769 6784 49794 6824
rect 49794 6784 49834 6824
rect 49834 6784 49855 6824
rect 49937 6784 49958 6824
rect 49958 6784 49998 6824
rect 49998 6784 50023 6824
rect 49769 6761 49855 6784
rect 49937 6761 50023 6784
rect 64889 6824 64975 6847
rect 65057 6824 65143 6847
rect 64889 6784 64914 6824
rect 64914 6784 64954 6824
rect 64954 6784 64975 6824
rect 65057 6784 65078 6824
rect 65078 6784 65118 6824
rect 65118 6784 65143 6824
rect 64889 6761 64975 6784
rect 65057 6761 65143 6784
rect 80009 6824 80095 6847
rect 80177 6824 80263 6847
rect 80009 6784 80034 6824
rect 80034 6784 80074 6824
rect 80074 6784 80095 6824
rect 80177 6784 80198 6824
rect 80198 6784 80238 6824
rect 80238 6784 80263 6824
rect 80009 6761 80095 6784
rect 80177 6761 80263 6784
rect 95129 6824 95215 6847
rect 95297 6824 95383 6847
rect 95129 6784 95154 6824
rect 95154 6784 95194 6824
rect 95194 6784 95215 6824
rect 95297 6784 95318 6824
rect 95318 6784 95358 6824
rect 95358 6784 95383 6824
rect 95129 6761 95215 6784
rect 95297 6761 95383 6784
rect 3169 6068 3255 6091
rect 3337 6068 3423 6091
rect 3169 6028 3194 6068
rect 3194 6028 3234 6068
rect 3234 6028 3255 6068
rect 3337 6028 3358 6068
rect 3358 6028 3398 6068
rect 3398 6028 3423 6068
rect 3169 6005 3255 6028
rect 3337 6005 3423 6028
rect 18289 6068 18375 6091
rect 18457 6068 18543 6091
rect 18289 6028 18314 6068
rect 18314 6028 18354 6068
rect 18354 6028 18375 6068
rect 18457 6028 18478 6068
rect 18478 6028 18518 6068
rect 18518 6028 18543 6068
rect 18289 6005 18375 6028
rect 18457 6005 18543 6028
rect 33409 6068 33495 6091
rect 33577 6068 33663 6091
rect 33409 6028 33434 6068
rect 33434 6028 33474 6068
rect 33474 6028 33495 6068
rect 33577 6028 33598 6068
rect 33598 6028 33638 6068
rect 33638 6028 33663 6068
rect 33409 6005 33495 6028
rect 33577 6005 33663 6028
rect 48529 6068 48615 6091
rect 48697 6068 48783 6091
rect 48529 6028 48554 6068
rect 48554 6028 48594 6068
rect 48594 6028 48615 6068
rect 48697 6028 48718 6068
rect 48718 6028 48758 6068
rect 48758 6028 48783 6068
rect 48529 6005 48615 6028
rect 48697 6005 48783 6028
rect 63649 6068 63735 6091
rect 63817 6068 63903 6091
rect 63649 6028 63674 6068
rect 63674 6028 63714 6068
rect 63714 6028 63735 6068
rect 63817 6028 63838 6068
rect 63838 6028 63878 6068
rect 63878 6028 63903 6068
rect 63649 6005 63735 6028
rect 63817 6005 63903 6028
rect 78769 6068 78855 6091
rect 78937 6068 79023 6091
rect 78769 6028 78794 6068
rect 78794 6028 78834 6068
rect 78834 6028 78855 6068
rect 78937 6028 78958 6068
rect 78958 6028 78998 6068
rect 78998 6028 79023 6068
rect 78769 6005 78855 6028
rect 78937 6005 79023 6028
rect 93889 6068 93975 6091
rect 94057 6068 94143 6091
rect 93889 6028 93914 6068
rect 93914 6028 93954 6068
rect 93954 6028 93975 6068
rect 94057 6028 94078 6068
rect 94078 6028 94118 6068
rect 94118 6028 94143 6068
rect 93889 6005 93975 6028
rect 94057 6005 94143 6028
rect 4409 5312 4495 5335
rect 4577 5312 4663 5335
rect 4409 5272 4434 5312
rect 4434 5272 4474 5312
rect 4474 5272 4495 5312
rect 4577 5272 4598 5312
rect 4598 5272 4638 5312
rect 4638 5272 4663 5312
rect 4409 5249 4495 5272
rect 4577 5249 4663 5272
rect 19529 5312 19615 5335
rect 19697 5312 19783 5335
rect 19529 5272 19554 5312
rect 19554 5272 19594 5312
rect 19594 5272 19615 5312
rect 19697 5272 19718 5312
rect 19718 5272 19758 5312
rect 19758 5272 19783 5312
rect 19529 5249 19615 5272
rect 19697 5249 19783 5272
rect 34649 5312 34735 5335
rect 34817 5312 34903 5335
rect 34649 5272 34674 5312
rect 34674 5272 34714 5312
rect 34714 5272 34735 5312
rect 34817 5272 34838 5312
rect 34838 5272 34878 5312
rect 34878 5272 34903 5312
rect 34649 5249 34735 5272
rect 34817 5249 34903 5272
rect 49769 5312 49855 5335
rect 49937 5312 50023 5335
rect 49769 5272 49794 5312
rect 49794 5272 49834 5312
rect 49834 5272 49855 5312
rect 49937 5272 49958 5312
rect 49958 5272 49998 5312
rect 49998 5272 50023 5312
rect 49769 5249 49855 5272
rect 49937 5249 50023 5272
rect 64889 5312 64975 5335
rect 65057 5312 65143 5335
rect 64889 5272 64914 5312
rect 64914 5272 64954 5312
rect 64954 5272 64975 5312
rect 65057 5272 65078 5312
rect 65078 5272 65118 5312
rect 65118 5272 65143 5312
rect 64889 5249 64975 5272
rect 65057 5249 65143 5272
rect 80009 5312 80095 5335
rect 80177 5312 80263 5335
rect 80009 5272 80034 5312
rect 80034 5272 80074 5312
rect 80074 5272 80095 5312
rect 80177 5272 80198 5312
rect 80198 5272 80238 5312
rect 80238 5272 80263 5312
rect 80009 5249 80095 5272
rect 80177 5249 80263 5272
rect 95129 5312 95215 5335
rect 95297 5312 95383 5335
rect 95129 5272 95154 5312
rect 95154 5272 95194 5312
rect 95194 5272 95215 5312
rect 95297 5272 95318 5312
rect 95318 5272 95358 5312
rect 95358 5272 95383 5312
rect 95129 5249 95215 5272
rect 95297 5249 95383 5272
rect 3169 4556 3255 4579
rect 3337 4556 3423 4579
rect 3169 4516 3194 4556
rect 3194 4516 3234 4556
rect 3234 4516 3255 4556
rect 3337 4516 3358 4556
rect 3358 4516 3398 4556
rect 3398 4516 3423 4556
rect 3169 4493 3255 4516
rect 3337 4493 3423 4516
rect 18289 4556 18375 4579
rect 18457 4556 18543 4579
rect 18289 4516 18314 4556
rect 18314 4516 18354 4556
rect 18354 4516 18375 4556
rect 18457 4516 18478 4556
rect 18478 4516 18518 4556
rect 18518 4516 18543 4556
rect 18289 4493 18375 4516
rect 18457 4493 18543 4516
rect 33409 4556 33495 4579
rect 33577 4556 33663 4579
rect 33409 4516 33434 4556
rect 33434 4516 33474 4556
rect 33474 4516 33495 4556
rect 33577 4516 33598 4556
rect 33598 4516 33638 4556
rect 33638 4516 33663 4556
rect 33409 4493 33495 4516
rect 33577 4493 33663 4516
rect 48529 4556 48615 4579
rect 48697 4556 48783 4579
rect 48529 4516 48554 4556
rect 48554 4516 48594 4556
rect 48594 4516 48615 4556
rect 48697 4516 48718 4556
rect 48718 4516 48758 4556
rect 48758 4516 48783 4556
rect 48529 4493 48615 4516
rect 48697 4493 48783 4516
rect 63649 4556 63735 4579
rect 63817 4556 63903 4579
rect 63649 4516 63674 4556
rect 63674 4516 63714 4556
rect 63714 4516 63735 4556
rect 63817 4516 63838 4556
rect 63838 4516 63878 4556
rect 63878 4516 63903 4556
rect 63649 4493 63735 4516
rect 63817 4493 63903 4516
rect 78769 4556 78855 4579
rect 78937 4556 79023 4579
rect 78769 4516 78794 4556
rect 78794 4516 78834 4556
rect 78834 4516 78855 4556
rect 78937 4516 78958 4556
rect 78958 4516 78998 4556
rect 78998 4516 79023 4556
rect 78769 4493 78855 4516
rect 78937 4493 79023 4516
rect 93889 4556 93975 4579
rect 94057 4556 94143 4579
rect 93889 4516 93914 4556
rect 93914 4516 93954 4556
rect 93954 4516 93975 4556
rect 94057 4516 94078 4556
rect 94078 4516 94118 4556
rect 94118 4516 94143 4556
rect 93889 4493 93975 4516
rect 94057 4493 94143 4516
rect 4409 3800 4495 3823
rect 4577 3800 4663 3823
rect 4409 3760 4434 3800
rect 4434 3760 4474 3800
rect 4474 3760 4495 3800
rect 4577 3760 4598 3800
rect 4598 3760 4638 3800
rect 4638 3760 4663 3800
rect 4409 3737 4495 3760
rect 4577 3737 4663 3760
rect 19529 3800 19615 3823
rect 19697 3800 19783 3823
rect 19529 3760 19554 3800
rect 19554 3760 19594 3800
rect 19594 3760 19615 3800
rect 19697 3760 19718 3800
rect 19718 3760 19758 3800
rect 19758 3760 19783 3800
rect 19529 3737 19615 3760
rect 19697 3737 19783 3760
rect 34649 3800 34735 3823
rect 34817 3800 34903 3823
rect 34649 3760 34674 3800
rect 34674 3760 34714 3800
rect 34714 3760 34735 3800
rect 34817 3760 34838 3800
rect 34838 3760 34878 3800
rect 34878 3760 34903 3800
rect 34649 3737 34735 3760
rect 34817 3737 34903 3760
rect 49769 3800 49855 3823
rect 49937 3800 50023 3823
rect 49769 3760 49794 3800
rect 49794 3760 49834 3800
rect 49834 3760 49855 3800
rect 49937 3760 49958 3800
rect 49958 3760 49998 3800
rect 49998 3760 50023 3800
rect 49769 3737 49855 3760
rect 49937 3737 50023 3760
rect 64889 3800 64975 3823
rect 65057 3800 65143 3823
rect 64889 3760 64914 3800
rect 64914 3760 64954 3800
rect 64954 3760 64975 3800
rect 65057 3760 65078 3800
rect 65078 3760 65118 3800
rect 65118 3760 65143 3800
rect 64889 3737 64975 3760
rect 65057 3737 65143 3760
rect 80009 3800 80095 3823
rect 80177 3800 80263 3823
rect 80009 3760 80034 3800
rect 80034 3760 80074 3800
rect 80074 3760 80095 3800
rect 80177 3760 80198 3800
rect 80198 3760 80238 3800
rect 80238 3760 80263 3800
rect 80009 3737 80095 3760
rect 80177 3737 80263 3760
rect 95129 3800 95215 3823
rect 95297 3800 95383 3823
rect 95129 3760 95154 3800
rect 95154 3760 95194 3800
rect 95194 3760 95215 3800
rect 95297 3760 95318 3800
rect 95318 3760 95358 3800
rect 95358 3760 95383 3800
rect 95129 3737 95215 3760
rect 95297 3737 95383 3760
rect 3169 3044 3255 3067
rect 3337 3044 3423 3067
rect 3169 3004 3194 3044
rect 3194 3004 3234 3044
rect 3234 3004 3255 3044
rect 3337 3004 3358 3044
rect 3358 3004 3398 3044
rect 3398 3004 3423 3044
rect 3169 2981 3255 3004
rect 3337 2981 3423 3004
rect 18289 3044 18375 3067
rect 18457 3044 18543 3067
rect 18289 3004 18314 3044
rect 18314 3004 18354 3044
rect 18354 3004 18375 3044
rect 18457 3004 18478 3044
rect 18478 3004 18518 3044
rect 18518 3004 18543 3044
rect 18289 2981 18375 3004
rect 18457 2981 18543 3004
rect 33409 3044 33495 3067
rect 33577 3044 33663 3067
rect 33409 3004 33434 3044
rect 33434 3004 33474 3044
rect 33474 3004 33495 3044
rect 33577 3004 33598 3044
rect 33598 3004 33638 3044
rect 33638 3004 33663 3044
rect 33409 2981 33495 3004
rect 33577 2981 33663 3004
rect 48529 3044 48615 3067
rect 48697 3044 48783 3067
rect 48529 3004 48554 3044
rect 48554 3004 48594 3044
rect 48594 3004 48615 3044
rect 48697 3004 48718 3044
rect 48718 3004 48758 3044
rect 48758 3004 48783 3044
rect 48529 2981 48615 3004
rect 48697 2981 48783 3004
rect 63649 3044 63735 3067
rect 63817 3044 63903 3067
rect 63649 3004 63674 3044
rect 63674 3004 63714 3044
rect 63714 3004 63735 3044
rect 63817 3004 63838 3044
rect 63838 3004 63878 3044
rect 63878 3004 63903 3044
rect 63649 2981 63735 3004
rect 63817 2981 63903 3004
rect 78769 3044 78855 3067
rect 78937 3044 79023 3067
rect 78769 3004 78794 3044
rect 78794 3004 78834 3044
rect 78834 3004 78855 3044
rect 78937 3004 78958 3044
rect 78958 3004 78998 3044
rect 78998 3004 79023 3044
rect 78769 2981 78855 3004
rect 78937 2981 79023 3004
rect 93889 3044 93975 3067
rect 94057 3044 94143 3067
rect 93889 3004 93914 3044
rect 93914 3004 93954 3044
rect 93954 3004 93975 3044
rect 94057 3004 94078 3044
rect 94078 3004 94118 3044
rect 94118 3004 94143 3044
rect 93889 2981 93975 3004
rect 94057 2981 94143 3004
rect 4409 2288 4495 2311
rect 4577 2288 4663 2311
rect 4409 2248 4434 2288
rect 4434 2248 4474 2288
rect 4474 2248 4495 2288
rect 4577 2248 4598 2288
rect 4598 2248 4638 2288
rect 4638 2248 4663 2288
rect 4409 2225 4495 2248
rect 4577 2225 4663 2248
rect 19529 2288 19615 2311
rect 19697 2288 19783 2311
rect 19529 2248 19554 2288
rect 19554 2248 19594 2288
rect 19594 2248 19615 2288
rect 19697 2248 19718 2288
rect 19718 2248 19758 2288
rect 19758 2248 19783 2288
rect 19529 2225 19615 2248
rect 19697 2225 19783 2248
rect 34649 2288 34735 2311
rect 34817 2288 34903 2311
rect 34649 2248 34674 2288
rect 34674 2248 34714 2288
rect 34714 2248 34735 2288
rect 34817 2248 34838 2288
rect 34838 2248 34878 2288
rect 34878 2248 34903 2288
rect 34649 2225 34735 2248
rect 34817 2225 34903 2248
rect 49769 2288 49855 2311
rect 49937 2288 50023 2311
rect 49769 2248 49794 2288
rect 49794 2248 49834 2288
rect 49834 2248 49855 2288
rect 49937 2248 49958 2288
rect 49958 2248 49998 2288
rect 49998 2248 50023 2288
rect 49769 2225 49855 2248
rect 49937 2225 50023 2248
rect 64889 2288 64975 2311
rect 65057 2288 65143 2311
rect 64889 2248 64914 2288
rect 64914 2248 64954 2288
rect 64954 2248 64975 2288
rect 65057 2248 65078 2288
rect 65078 2248 65118 2288
rect 65118 2248 65143 2288
rect 64889 2225 64975 2248
rect 65057 2225 65143 2248
rect 80009 2288 80095 2311
rect 80177 2288 80263 2311
rect 80009 2248 80034 2288
rect 80034 2248 80074 2288
rect 80074 2248 80095 2288
rect 80177 2248 80198 2288
rect 80198 2248 80238 2288
rect 80238 2248 80263 2288
rect 80009 2225 80095 2248
rect 80177 2225 80263 2248
rect 95129 2288 95215 2311
rect 95297 2288 95383 2311
rect 95129 2248 95154 2288
rect 95154 2248 95194 2288
rect 95194 2248 95215 2288
rect 95297 2248 95318 2288
rect 95318 2248 95358 2288
rect 95358 2248 95383 2288
rect 95129 2225 95215 2248
rect 95297 2225 95383 2248
rect 3169 1532 3255 1555
rect 3337 1532 3423 1555
rect 3169 1492 3194 1532
rect 3194 1492 3234 1532
rect 3234 1492 3255 1532
rect 3337 1492 3358 1532
rect 3358 1492 3398 1532
rect 3398 1492 3423 1532
rect 3169 1469 3255 1492
rect 3337 1469 3423 1492
rect 18289 1532 18375 1555
rect 18457 1532 18543 1555
rect 18289 1492 18314 1532
rect 18314 1492 18354 1532
rect 18354 1492 18375 1532
rect 18457 1492 18478 1532
rect 18478 1492 18518 1532
rect 18518 1492 18543 1532
rect 18289 1469 18375 1492
rect 18457 1469 18543 1492
rect 33409 1532 33495 1555
rect 33577 1532 33663 1555
rect 33409 1492 33434 1532
rect 33434 1492 33474 1532
rect 33474 1492 33495 1532
rect 33577 1492 33598 1532
rect 33598 1492 33638 1532
rect 33638 1492 33663 1532
rect 33409 1469 33495 1492
rect 33577 1469 33663 1492
rect 48529 1532 48615 1555
rect 48697 1532 48783 1555
rect 48529 1492 48554 1532
rect 48554 1492 48594 1532
rect 48594 1492 48615 1532
rect 48697 1492 48718 1532
rect 48718 1492 48758 1532
rect 48758 1492 48783 1532
rect 48529 1469 48615 1492
rect 48697 1469 48783 1492
rect 63649 1532 63735 1555
rect 63817 1532 63903 1555
rect 63649 1492 63674 1532
rect 63674 1492 63714 1532
rect 63714 1492 63735 1532
rect 63817 1492 63838 1532
rect 63838 1492 63878 1532
rect 63878 1492 63903 1532
rect 63649 1469 63735 1492
rect 63817 1469 63903 1492
rect 78769 1532 78855 1555
rect 78937 1532 79023 1555
rect 78769 1492 78794 1532
rect 78794 1492 78834 1532
rect 78834 1492 78855 1532
rect 78937 1492 78958 1532
rect 78958 1492 78998 1532
rect 78998 1492 79023 1532
rect 78769 1469 78855 1492
rect 78937 1469 79023 1492
rect 93889 1532 93975 1555
rect 94057 1532 94143 1555
rect 93889 1492 93914 1532
rect 93914 1492 93954 1532
rect 93954 1492 93975 1532
rect 94057 1492 94078 1532
rect 94078 1492 94118 1532
rect 94118 1492 94143 1532
rect 93889 1469 93975 1492
rect 94057 1469 94143 1492
rect 4409 776 4495 799
rect 4577 776 4663 799
rect 4409 736 4434 776
rect 4434 736 4474 776
rect 4474 736 4495 776
rect 4577 736 4598 776
rect 4598 736 4638 776
rect 4638 736 4663 776
rect 4409 713 4495 736
rect 4577 713 4663 736
rect 19529 776 19615 799
rect 19697 776 19783 799
rect 19529 736 19554 776
rect 19554 736 19594 776
rect 19594 736 19615 776
rect 19697 736 19718 776
rect 19718 736 19758 776
rect 19758 736 19783 776
rect 19529 713 19615 736
rect 19697 713 19783 736
rect 34649 776 34735 799
rect 34817 776 34903 799
rect 34649 736 34674 776
rect 34674 736 34714 776
rect 34714 736 34735 776
rect 34817 736 34838 776
rect 34838 736 34878 776
rect 34878 736 34903 776
rect 34649 713 34735 736
rect 34817 713 34903 736
rect 49769 776 49855 799
rect 49937 776 50023 799
rect 49769 736 49794 776
rect 49794 736 49834 776
rect 49834 736 49855 776
rect 49937 736 49958 776
rect 49958 736 49998 776
rect 49998 736 50023 776
rect 49769 713 49855 736
rect 49937 713 50023 736
rect 64889 776 64975 799
rect 65057 776 65143 799
rect 64889 736 64914 776
rect 64914 736 64954 776
rect 64954 736 64975 776
rect 65057 736 65078 776
rect 65078 736 65118 776
rect 65118 736 65143 776
rect 64889 713 64975 736
rect 65057 713 65143 736
rect 80009 776 80095 799
rect 80177 776 80263 799
rect 80009 736 80034 776
rect 80034 736 80074 776
rect 80074 736 80095 776
rect 80177 736 80198 776
rect 80198 736 80238 776
rect 80238 736 80263 776
rect 80009 713 80095 736
rect 80177 713 80263 736
rect 95129 776 95215 799
rect 95297 776 95383 799
rect 95129 736 95154 776
rect 95154 736 95194 776
rect 95194 736 95215 776
rect 95297 736 95318 776
rect 95318 736 95358 776
rect 95358 736 95383 776
rect 95129 713 95215 736
rect 95297 713 95383 736
<< metal6 >>
rect 3076 37843 3516 38600
rect 3076 37757 3169 37843
rect 3255 37757 3337 37843
rect 3423 37757 3516 37843
rect 3076 36331 3516 37757
rect 3076 36245 3169 36331
rect 3255 36245 3337 36331
rect 3423 36245 3516 36331
rect 3076 34819 3516 36245
rect 3076 34733 3169 34819
rect 3255 34733 3337 34819
rect 3423 34733 3516 34819
rect 3076 33307 3516 34733
rect 3076 33221 3169 33307
rect 3255 33221 3337 33307
rect 3423 33221 3516 33307
rect 3076 31795 3516 33221
rect 3076 31709 3169 31795
rect 3255 31709 3337 31795
rect 3423 31709 3516 31795
rect 3076 30283 3516 31709
rect 3076 30197 3169 30283
rect 3255 30197 3337 30283
rect 3423 30197 3516 30283
rect 3076 28771 3516 30197
rect 3076 28685 3169 28771
rect 3255 28685 3337 28771
rect 3423 28685 3516 28771
rect 3076 27259 3516 28685
rect 3076 27173 3169 27259
rect 3255 27173 3337 27259
rect 3423 27173 3516 27259
rect 3076 25747 3516 27173
rect 3076 25661 3169 25747
rect 3255 25661 3337 25747
rect 3423 25661 3516 25747
rect 3076 24235 3516 25661
rect 3076 24149 3169 24235
rect 3255 24149 3337 24235
rect 3423 24149 3516 24235
rect 3076 22723 3516 24149
rect 3076 22637 3169 22723
rect 3255 22637 3337 22723
rect 3423 22637 3516 22723
rect 3076 21211 3516 22637
rect 3076 21125 3169 21211
rect 3255 21125 3337 21211
rect 3423 21125 3516 21211
rect 3076 19699 3516 21125
rect 3076 19613 3169 19699
rect 3255 19613 3337 19699
rect 3423 19613 3516 19699
rect 3076 18187 3516 19613
rect 3076 18101 3169 18187
rect 3255 18101 3337 18187
rect 3423 18101 3516 18187
rect 3076 16675 3516 18101
rect 3076 16589 3169 16675
rect 3255 16589 3337 16675
rect 3423 16589 3516 16675
rect 3076 15163 3516 16589
rect 3076 15077 3169 15163
rect 3255 15077 3337 15163
rect 3423 15077 3516 15163
rect 3076 13651 3516 15077
rect 3076 13565 3169 13651
rect 3255 13565 3337 13651
rect 3423 13565 3516 13651
rect 3076 12139 3516 13565
rect 3076 12053 3169 12139
rect 3255 12053 3337 12139
rect 3423 12053 3516 12139
rect 3076 10627 3516 12053
rect 3076 10541 3169 10627
rect 3255 10541 3337 10627
rect 3423 10541 3516 10627
rect 3076 9115 3516 10541
rect 3076 9029 3169 9115
rect 3255 9029 3337 9115
rect 3423 9029 3516 9115
rect 3076 7603 3516 9029
rect 3076 7517 3169 7603
rect 3255 7517 3337 7603
rect 3423 7517 3516 7603
rect 3076 6091 3516 7517
rect 3076 6005 3169 6091
rect 3255 6005 3337 6091
rect 3423 6005 3516 6091
rect 3076 4579 3516 6005
rect 3076 4493 3169 4579
rect 3255 4493 3337 4579
rect 3423 4493 3516 4579
rect 3076 3067 3516 4493
rect 3076 2981 3169 3067
rect 3255 2981 3337 3067
rect 3423 2981 3516 3067
rect 3076 1555 3516 2981
rect 3076 1469 3169 1555
rect 3255 1469 3337 1555
rect 3423 1469 3516 1555
rect 3076 712 3516 1469
rect 4316 38599 4756 38682
rect 4316 38513 4409 38599
rect 4495 38513 4577 38599
rect 4663 38513 4756 38599
rect 4316 37087 4756 38513
rect 4316 37001 4409 37087
rect 4495 37001 4577 37087
rect 4663 37001 4756 37087
rect 4316 35575 4756 37001
rect 4316 35489 4409 35575
rect 4495 35489 4577 35575
rect 4663 35489 4756 35575
rect 4316 34063 4756 35489
rect 4316 33977 4409 34063
rect 4495 33977 4577 34063
rect 4663 33977 4756 34063
rect 4316 32551 4756 33977
rect 4316 32465 4409 32551
rect 4495 32465 4577 32551
rect 4663 32465 4756 32551
rect 4316 31039 4756 32465
rect 4316 30953 4409 31039
rect 4495 30953 4577 31039
rect 4663 30953 4756 31039
rect 4316 29527 4756 30953
rect 4316 29441 4409 29527
rect 4495 29441 4577 29527
rect 4663 29441 4756 29527
rect 4316 28015 4756 29441
rect 4316 27929 4409 28015
rect 4495 27929 4577 28015
rect 4663 27929 4756 28015
rect 4316 26503 4756 27929
rect 4316 26417 4409 26503
rect 4495 26417 4577 26503
rect 4663 26417 4756 26503
rect 4316 24991 4756 26417
rect 4316 24905 4409 24991
rect 4495 24905 4577 24991
rect 4663 24905 4756 24991
rect 4316 23479 4756 24905
rect 4316 23393 4409 23479
rect 4495 23393 4577 23479
rect 4663 23393 4756 23479
rect 4316 21967 4756 23393
rect 4316 21881 4409 21967
rect 4495 21881 4577 21967
rect 4663 21881 4756 21967
rect 4316 20455 4756 21881
rect 4316 20369 4409 20455
rect 4495 20369 4577 20455
rect 4663 20369 4756 20455
rect 4316 18943 4756 20369
rect 4316 18857 4409 18943
rect 4495 18857 4577 18943
rect 4663 18857 4756 18943
rect 4316 17431 4756 18857
rect 4316 17345 4409 17431
rect 4495 17345 4577 17431
rect 4663 17345 4756 17431
rect 4316 15919 4756 17345
rect 4316 15833 4409 15919
rect 4495 15833 4577 15919
rect 4663 15833 4756 15919
rect 4316 14407 4756 15833
rect 4316 14321 4409 14407
rect 4495 14321 4577 14407
rect 4663 14321 4756 14407
rect 4316 12895 4756 14321
rect 4316 12809 4409 12895
rect 4495 12809 4577 12895
rect 4663 12809 4756 12895
rect 4316 11383 4756 12809
rect 4316 11297 4409 11383
rect 4495 11297 4577 11383
rect 4663 11297 4756 11383
rect 4316 9871 4756 11297
rect 4316 9785 4409 9871
rect 4495 9785 4577 9871
rect 4663 9785 4756 9871
rect 4316 8359 4756 9785
rect 4316 8273 4409 8359
rect 4495 8273 4577 8359
rect 4663 8273 4756 8359
rect 4316 6847 4756 8273
rect 4316 6761 4409 6847
rect 4495 6761 4577 6847
rect 4663 6761 4756 6847
rect 4316 5335 4756 6761
rect 4316 5249 4409 5335
rect 4495 5249 4577 5335
rect 4663 5249 4756 5335
rect 4316 3823 4756 5249
rect 4316 3737 4409 3823
rect 4495 3737 4577 3823
rect 4663 3737 4756 3823
rect 4316 2311 4756 3737
rect 4316 2225 4409 2311
rect 4495 2225 4577 2311
rect 4663 2225 4756 2311
rect 4316 799 4756 2225
rect 4316 713 4409 799
rect 4495 713 4577 799
rect 4663 713 4756 799
rect 4316 630 4756 713
rect 18196 37843 18636 38600
rect 18196 37757 18289 37843
rect 18375 37757 18457 37843
rect 18543 37757 18636 37843
rect 18196 36331 18636 37757
rect 18196 36245 18289 36331
rect 18375 36245 18457 36331
rect 18543 36245 18636 36331
rect 18196 34819 18636 36245
rect 18196 34733 18289 34819
rect 18375 34733 18457 34819
rect 18543 34733 18636 34819
rect 18196 33307 18636 34733
rect 18196 33221 18289 33307
rect 18375 33221 18457 33307
rect 18543 33221 18636 33307
rect 18196 31795 18636 33221
rect 18196 31709 18289 31795
rect 18375 31709 18457 31795
rect 18543 31709 18636 31795
rect 18196 30283 18636 31709
rect 18196 30197 18289 30283
rect 18375 30197 18457 30283
rect 18543 30197 18636 30283
rect 18196 28771 18636 30197
rect 18196 28685 18289 28771
rect 18375 28685 18457 28771
rect 18543 28685 18636 28771
rect 18196 27259 18636 28685
rect 18196 27173 18289 27259
rect 18375 27173 18457 27259
rect 18543 27173 18636 27259
rect 18196 25747 18636 27173
rect 18196 25661 18289 25747
rect 18375 25661 18457 25747
rect 18543 25661 18636 25747
rect 18196 24235 18636 25661
rect 18196 24149 18289 24235
rect 18375 24149 18457 24235
rect 18543 24149 18636 24235
rect 18196 22723 18636 24149
rect 18196 22637 18289 22723
rect 18375 22637 18457 22723
rect 18543 22637 18636 22723
rect 18196 21211 18636 22637
rect 18196 21125 18289 21211
rect 18375 21125 18457 21211
rect 18543 21125 18636 21211
rect 18196 19699 18636 21125
rect 18196 19613 18289 19699
rect 18375 19613 18457 19699
rect 18543 19613 18636 19699
rect 18196 18187 18636 19613
rect 18196 18101 18289 18187
rect 18375 18101 18457 18187
rect 18543 18101 18636 18187
rect 18196 16675 18636 18101
rect 18196 16589 18289 16675
rect 18375 16589 18457 16675
rect 18543 16589 18636 16675
rect 18196 15163 18636 16589
rect 18196 15077 18289 15163
rect 18375 15077 18457 15163
rect 18543 15077 18636 15163
rect 18196 13651 18636 15077
rect 18196 13565 18289 13651
rect 18375 13565 18457 13651
rect 18543 13565 18636 13651
rect 18196 12139 18636 13565
rect 18196 12053 18289 12139
rect 18375 12053 18457 12139
rect 18543 12053 18636 12139
rect 18196 10627 18636 12053
rect 18196 10541 18289 10627
rect 18375 10541 18457 10627
rect 18543 10541 18636 10627
rect 18196 9115 18636 10541
rect 18196 9029 18289 9115
rect 18375 9029 18457 9115
rect 18543 9029 18636 9115
rect 18196 7603 18636 9029
rect 18196 7517 18289 7603
rect 18375 7517 18457 7603
rect 18543 7517 18636 7603
rect 18196 6091 18636 7517
rect 18196 6005 18289 6091
rect 18375 6005 18457 6091
rect 18543 6005 18636 6091
rect 18196 4579 18636 6005
rect 18196 4493 18289 4579
rect 18375 4493 18457 4579
rect 18543 4493 18636 4579
rect 18196 3067 18636 4493
rect 18196 2981 18289 3067
rect 18375 2981 18457 3067
rect 18543 2981 18636 3067
rect 18196 1555 18636 2981
rect 18196 1469 18289 1555
rect 18375 1469 18457 1555
rect 18543 1469 18636 1555
rect 18196 712 18636 1469
rect 19436 38599 19876 38682
rect 19436 38513 19529 38599
rect 19615 38513 19697 38599
rect 19783 38513 19876 38599
rect 19436 37087 19876 38513
rect 19436 37001 19529 37087
rect 19615 37001 19697 37087
rect 19783 37001 19876 37087
rect 19436 35575 19876 37001
rect 19436 35489 19529 35575
rect 19615 35489 19697 35575
rect 19783 35489 19876 35575
rect 19436 34063 19876 35489
rect 19436 33977 19529 34063
rect 19615 33977 19697 34063
rect 19783 33977 19876 34063
rect 19436 32551 19876 33977
rect 19436 32465 19529 32551
rect 19615 32465 19697 32551
rect 19783 32465 19876 32551
rect 19436 31039 19876 32465
rect 19436 30953 19529 31039
rect 19615 30953 19697 31039
rect 19783 30953 19876 31039
rect 19436 29527 19876 30953
rect 19436 29441 19529 29527
rect 19615 29441 19697 29527
rect 19783 29441 19876 29527
rect 19436 28015 19876 29441
rect 19436 27929 19529 28015
rect 19615 27929 19697 28015
rect 19783 27929 19876 28015
rect 19436 26503 19876 27929
rect 19436 26417 19529 26503
rect 19615 26417 19697 26503
rect 19783 26417 19876 26503
rect 19436 24991 19876 26417
rect 19436 24905 19529 24991
rect 19615 24905 19697 24991
rect 19783 24905 19876 24991
rect 19436 23479 19876 24905
rect 19436 23393 19529 23479
rect 19615 23393 19697 23479
rect 19783 23393 19876 23479
rect 19436 21967 19876 23393
rect 19436 21881 19529 21967
rect 19615 21881 19697 21967
rect 19783 21881 19876 21967
rect 19436 20455 19876 21881
rect 19436 20369 19529 20455
rect 19615 20369 19697 20455
rect 19783 20369 19876 20455
rect 19436 18943 19876 20369
rect 19436 18857 19529 18943
rect 19615 18857 19697 18943
rect 19783 18857 19876 18943
rect 19436 17431 19876 18857
rect 19436 17345 19529 17431
rect 19615 17345 19697 17431
rect 19783 17345 19876 17431
rect 19436 15919 19876 17345
rect 19436 15833 19529 15919
rect 19615 15833 19697 15919
rect 19783 15833 19876 15919
rect 19436 14407 19876 15833
rect 19436 14321 19529 14407
rect 19615 14321 19697 14407
rect 19783 14321 19876 14407
rect 19436 12895 19876 14321
rect 19436 12809 19529 12895
rect 19615 12809 19697 12895
rect 19783 12809 19876 12895
rect 19436 11383 19876 12809
rect 19436 11297 19529 11383
rect 19615 11297 19697 11383
rect 19783 11297 19876 11383
rect 19436 9871 19876 11297
rect 19436 9785 19529 9871
rect 19615 9785 19697 9871
rect 19783 9785 19876 9871
rect 19436 8359 19876 9785
rect 19436 8273 19529 8359
rect 19615 8273 19697 8359
rect 19783 8273 19876 8359
rect 19436 6847 19876 8273
rect 19436 6761 19529 6847
rect 19615 6761 19697 6847
rect 19783 6761 19876 6847
rect 19436 5335 19876 6761
rect 19436 5249 19529 5335
rect 19615 5249 19697 5335
rect 19783 5249 19876 5335
rect 19436 3823 19876 5249
rect 19436 3737 19529 3823
rect 19615 3737 19697 3823
rect 19783 3737 19876 3823
rect 19436 2311 19876 3737
rect 19436 2225 19529 2311
rect 19615 2225 19697 2311
rect 19783 2225 19876 2311
rect 19436 799 19876 2225
rect 19436 713 19529 799
rect 19615 713 19697 799
rect 19783 713 19876 799
rect 19436 630 19876 713
rect 33316 37843 33756 38600
rect 33316 37757 33409 37843
rect 33495 37757 33577 37843
rect 33663 37757 33756 37843
rect 33316 36331 33756 37757
rect 33316 36245 33409 36331
rect 33495 36245 33577 36331
rect 33663 36245 33756 36331
rect 33316 34819 33756 36245
rect 33316 34733 33409 34819
rect 33495 34733 33577 34819
rect 33663 34733 33756 34819
rect 33316 33307 33756 34733
rect 33316 33221 33409 33307
rect 33495 33221 33577 33307
rect 33663 33221 33756 33307
rect 33316 31795 33756 33221
rect 33316 31709 33409 31795
rect 33495 31709 33577 31795
rect 33663 31709 33756 31795
rect 33316 30283 33756 31709
rect 33316 30197 33409 30283
rect 33495 30197 33577 30283
rect 33663 30197 33756 30283
rect 33316 28771 33756 30197
rect 33316 28685 33409 28771
rect 33495 28685 33577 28771
rect 33663 28685 33756 28771
rect 33316 27259 33756 28685
rect 33316 27173 33409 27259
rect 33495 27173 33577 27259
rect 33663 27173 33756 27259
rect 33316 25747 33756 27173
rect 33316 25661 33409 25747
rect 33495 25661 33577 25747
rect 33663 25661 33756 25747
rect 33316 24235 33756 25661
rect 33316 24149 33409 24235
rect 33495 24149 33577 24235
rect 33663 24149 33756 24235
rect 33316 22723 33756 24149
rect 33316 22637 33409 22723
rect 33495 22637 33577 22723
rect 33663 22637 33756 22723
rect 33316 21211 33756 22637
rect 33316 21125 33409 21211
rect 33495 21125 33577 21211
rect 33663 21125 33756 21211
rect 33316 19699 33756 21125
rect 33316 19613 33409 19699
rect 33495 19613 33577 19699
rect 33663 19613 33756 19699
rect 33316 18187 33756 19613
rect 33316 18101 33409 18187
rect 33495 18101 33577 18187
rect 33663 18101 33756 18187
rect 33316 16675 33756 18101
rect 33316 16589 33409 16675
rect 33495 16589 33577 16675
rect 33663 16589 33756 16675
rect 33316 15163 33756 16589
rect 33316 15077 33409 15163
rect 33495 15077 33577 15163
rect 33663 15077 33756 15163
rect 33316 13651 33756 15077
rect 33316 13565 33409 13651
rect 33495 13565 33577 13651
rect 33663 13565 33756 13651
rect 33316 12139 33756 13565
rect 33316 12053 33409 12139
rect 33495 12053 33577 12139
rect 33663 12053 33756 12139
rect 33316 10627 33756 12053
rect 33316 10541 33409 10627
rect 33495 10541 33577 10627
rect 33663 10541 33756 10627
rect 33316 9115 33756 10541
rect 33316 9029 33409 9115
rect 33495 9029 33577 9115
rect 33663 9029 33756 9115
rect 33316 7603 33756 9029
rect 33316 7517 33409 7603
rect 33495 7517 33577 7603
rect 33663 7517 33756 7603
rect 33316 6091 33756 7517
rect 33316 6005 33409 6091
rect 33495 6005 33577 6091
rect 33663 6005 33756 6091
rect 33316 4579 33756 6005
rect 33316 4493 33409 4579
rect 33495 4493 33577 4579
rect 33663 4493 33756 4579
rect 33316 3067 33756 4493
rect 33316 2981 33409 3067
rect 33495 2981 33577 3067
rect 33663 2981 33756 3067
rect 33316 1555 33756 2981
rect 33316 1469 33409 1555
rect 33495 1469 33577 1555
rect 33663 1469 33756 1555
rect 33316 712 33756 1469
rect 34556 38599 34996 38682
rect 34556 38513 34649 38599
rect 34735 38513 34817 38599
rect 34903 38513 34996 38599
rect 34556 37087 34996 38513
rect 34556 37001 34649 37087
rect 34735 37001 34817 37087
rect 34903 37001 34996 37087
rect 34556 35575 34996 37001
rect 34556 35489 34649 35575
rect 34735 35489 34817 35575
rect 34903 35489 34996 35575
rect 34556 34063 34996 35489
rect 34556 33977 34649 34063
rect 34735 33977 34817 34063
rect 34903 33977 34996 34063
rect 34556 32551 34996 33977
rect 34556 32465 34649 32551
rect 34735 32465 34817 32551
rect 34903 32465 34996 32551
rect 34556 31039 34996 32465
rect 34556 30953 34649 31039
rect 34735 30953 34817 31039
rect 34903 30953 34996 31039
rect 34556 29527 34996 30953
rect 34556 29441 34649 29527
rect 34735 29441 34817 29527
rect 34903 29441 34996 29527
rect 34556 28015 34996 29441
rect 34556 27929 34649 28015
rect 34735 27929 34817 28015
rect 34903 27929 34996 28015
rect 34556 26503 34996 27929
rect 34556 26417 34649 26503
rect 34735 26417 34817 26503
rect 34903 26417 34996 26503
rect 34556 24991 34996 26417
rect 34556 24905 34649 24991
rect 34735 24905 34817 24991
rect 34903 24905 34996 24991
rect 34556 23479 34996 24905
rect 34556 23393 34649 23479
rect 34735 23393 34817 23479
rect 34903 23393 34996 23479
rect 34556 21967 34996 23393
rect 34556 21881 34649 21967
rect 34735 21881 34817 21967
rect 34903 21881 34996 21967
rect 34556 20455 34996 21881
rect 34556 20369 34649 20455
rect 34735 20369 34817 20455
rect 34903 20369 34996 20455
rect 34556 18943 34996 20369
rect 34556 18857 34649 18943
rect 34735 18857 34817 18943
rect 34903 18857 34996 18943
rect 34556 17431 34996 18857
rect 34556 17345 34649 17431
rect 34735 17345 34817 17431
rect 34903 17345 34996 17431
rect 34556 15919 34996 17345
rect 34556 15833 34649 15919
rect 34735 15833 34817 15919
rect 34903 15833 34996 15919
rect 34556 14407 34996 15833
rect 34556 14321 34649 14407
rect 34735 14321 34817 14407
rect 34903 14321 34996 14407
rect 34556 12895 34996 14321
rect 34556 12809 34649 12895
rect 34735 12809 34817 12895
rect 34903 12809 34996 12895
rect 34556 11383 34996 12809
rect 34556 11297 34649 11383
rect 34735 11297 34817 11383
rect 34903 11297 34996 11383
rect 34556 9871 34996 11297
rect 34556 9785 34649 9871
rect 34735 9785 34817 9871
rect 34903 9785 34996 9871
rect 34556 8359 34996 9785
rect 34556 8273 34649 8359
rect 34735 8273 34817 8359
rect 34903 8273 34996 8359
rect 34556 6847 34996 8273
rect 34556 6761 34649 6847
rect 34735 6761 34817 6847
rect 34903 6761 34996 6847
rect 34556 5335 34996 6761
rect 34556 5249 34649 5335
rect 34735 5249 34817 5335
rect 34903 5249 34996 5335
rect 34556 3823 34996 5249
rect 34556 3737 34649 3823
rect 34735 3737 34817 3823
rect 34903 3737 34996 3823
rect 34556 2311 34996 3737
rect 34556 2225 34649 2311
rect 34735 2225 34817 2311
rect 34903 2225 34996 2311
rect 34556 799 34996 2225
rect 34556 713 34649 799
rect 34735 713 34817 799
rect 34903 713 34996 799
rect 34556 630 34996 713
rect 48436 37843 48876 38600
rect 48436 37757 48529 37843
rect 48615 37757 48697 37843
rect 48783 37757 48876 37843
rect 48436 36331 48876 37757
rect 48436 36245 48529 36331
rect 48615 36245 48697 36331
rect 48783 36245 48876 36331
rect 48436 34819 48876 36245
rect 48436 34733 48529 34819
rect 48615 34733 48697 34819
rect 48783 34733 48876 34819
rect 48436 33307 48876 34733
rect 48436 33221 48529 33307
rect 48615 33221 48697 33307
rect 48783 33221 48876 33307
rect 48436 31795 48876 33221
rect 48436 31709 48529 31795
rect 48615 31709 48697 31795
rect 48783 31709 48876 31795
rect 48436 30283 48876 31709
rect 48436 30197 48529 30283
rect 48615 30197 48697 30283
rect 48783 30197 48876 30283
rect 48436 28771 48876 30197
rect 48436 28685 48529 28771
rect 48615 28685 48697 28771
rect 48783 28685 48876 28771
rect 48436 27259 48876 28685
rect 48436 27173 48529 27259
rect 48615 27173 48697 27259
rect 48783 27173 48876 27259
rect 48436 25747 48876 27173
rect 48436 25661 48529 25747
rect 48615 25661 48697 25747
rect 48783 25661 48876 25747
rect 48436 24235 48876 25661
rect 48436 24149 48529 24235
rect 48615 24149 48697 24235
rect 48783 24149 48876 24235
rect 48436 22723 48876 24149
rect 48436 22637 48529 22723
rect 48615 22637 48697 22723
rect 48783 22637 48876 22723
rect 48436 21211 48876 22637
rect 48436 21125 48529 21211
rect 48615 21125 48697 21211
rect 48783 21125 48876 21211
rect 48436 19699 48876 21125
rect 48436 19613 48529 19699
rect 48615 19613 48697 19699
rect 48783 19613 48876 19699
rect 48436 18187 48876 19613
rect 48436 18101 48529 18187
rect 48615 18101 48697 18187
rect 48783 18101 48876 18187
rect 48436 16675 48876 18101
rect 48436 16589 48529 16675
rect 48615 16589 48697 16675
rect 48783 16589 48876 16675
rect 48436 15163 48876 16589
rect 48436 15077 48529 15163
rect 48615 15077 48697 15163
rect 48783 15077 48876 15163
rect 48436 13651 48876 15077
rect 48436 13565 48529 13651
rect 48615 13565 48697 13651
rect 48783 13565 48876 13651
rect 48436 12139 48876 13565
rect 48436 12053 48529 12139
rect 48615 12053 48697 12139
rect 48783 12053 48876 12139
rect 48436 10627 48876 12053
rect 48436 10541 48529 10627
rect 48615 10541 48697 10627
rect 48783 10541 48876 10627
rect 48436 9115 48876 10541
rect 48436 9029 48529 9115
rect 48615 9029 48697 9115
rect 48783 9029 48876 9115
rect 48436 7603 48876 9029
rect 48436 7517 48529 7603
rect 48615 7517 48697 7603
rect 48783 7517 48876 7603
rect 48436 6091 48876 7517
rect 48436 6005 48529 6091
rect 48615 6005 48697 6091
rect 48783 6005 48876 6091
rect 48436 4579 48876 6005
rect 48436 4493 48529 4579
rect 48615 4493 48697 4579
rect 48783 4493 48876 4579
rect 48436 3067 48876 4493
rect 48436 2981 48529 3067
rect 48615 2981 48697 3067
rect 48783 2981 48876 3067
rect 48436 1555 48876 2981
rect 48436 1469 48529 1555
rect 48615 1469 48697 1555
rect 48783 1469 48876 1555
rect 48436 712 48876 1469
rect 49676 38599 50116 38682
rect 49676 38513 49769 38599
rect 49855 38513 49937 38599
rect 50023 38513 50116 38599
rect 49676 37087 50116 38513
rect 49676 37001 49769 37087
rect 49855 37001 49937 37087
rect 50023 37001 50116 37087
rect 49676 35575 50116 37001
rect 49676 35489 49769 35575
rect 49855 35489 49937 35575
rect 50023 35489 50116 35575
rect 49676 34063 50116 35489
rect 49676 33977 49769 34063
rect 49855 33977 49937 34063
rect 50023 33977 50116 34063
rect 49676 32551 50116 33977
rect 49676 32465 49769 32551
rect 49855 32465 49937 32551
rect 50023 32465 50116 32551
rect 49676 31039 50116 32465
rect 49676 30953 49769 31039
rect 49855 30953 49937 31039
rect 50023 30953 50116 31039
rect 49676 29527 50116 30953
rect 49676 29441 49769 29527
rect 49855 29441 49937 29527
rect 50023 29441 50116 29527
rect 49676 28015 50116 29441
rect 49676 27929 49769 28015
rect 49855 27929 49937 28015
rect 50023 27929 50116 28015
rect 49676 26503 50116 27929
rect 49676 26417 49769 26503
rect 49855 26417 49937 26503
rect 50023 26417 50116 26503
rect 49676 24991 50116 26417
rect 49676 24905 49769 24991
rect 49855 24905 49937 24991
rect 50023 24905 50116 24991
rect 49676 23479 50116 24905
rect 49676 23393 49769 23479
rect 49855 23393 49937 23479
rect 50023 23393 50116 23479
rect 49676 21967 50116 23393
rect 49676 21881 49769 21967
rect 49855 21881 49937 21967
rect 50023 21881 50116 21967
rect 49676 20455 50116 21881
rect 49676 20369 49769 20455
rect 49855 20369 49937 20455
rect 50023 20369 50116 20455
rect 49676 18943 50116 20369
rect 49676 18857 49769 18943
rect 49855 18857 49937 18943
rect 50023 18857 50116 18943
rect 49676 17431 50116 18857
rect 49676 17345 49769 17431
rect 49855 17345 49937 17431
rect 50023 17345 50116 17431
rect 49676 15919 50116 17345
rect 49676 15833 49769 15919
rect 49855 15833 49937 15919
rect 50023 15833 50116 15919
rect 49676 14407 50116 15833
rect 49676 14321 49769 14407
rect 49855 14321 49937 14407
rect 50023 14321 50116 14407
rect 49676 12895 50116 14321
rect 49676 12809 49769 12895
rect 49855 12809 49937 12895
rect 50023 12809 50116 12895
rect 49676 11383 50116 12809
rect 49676 11297 49769 11383
rect 49855 11297 49937 11383
rect 50023 11297 50116 11383
rect 49676 9871 50116 11297
rect 49676 9785 49769 9871
rect 49855 9785 49937 9871
rect 50023 9785 50116 9871
rect 49676 8359 50116 9785
rect 49676 8273 49769 8359
rect 49855 8273 49937 8359
rect 50023 8273 50116 8359
rect 49676 6847 50116 8273
rect 49676 6761 49769 6847
rect 49855 6761 49937 6847
rect 50023 6761 50116 6847
rect 49676 5335 50116 6761
rect 49676 5249 49769 5335
rect 49855 5249 49937 5335
rect 50023 5249 50116 5335
rect 49676 3823 50116 5249
rect 49676 3737 49769 3823
rect 49855 3737 49937 3823
rect 50023 3737 50116 3823
rect 49676 2311 50116 3737
rect 49676 2225 49769 2311
rect 49855 2225 49937 2311
rect 50023 2225 50116 2311
rect 49676 799 50116 2225
rect 49676 713 49769 799
rect 49855 713 49937 799
rect 50023 713 50116 799
rect 49676 630 50116 713
rect 63556 37843 63996 38600
rect 63556 37757 63649 37843
rect 63735 37757 63817 37843
rect 63903 37757 63996 37843
rect 63556 36331 63996 37757
rect 63556 36245 63649 36331
rect 63735 36245 63817 36331
rect 63903 36245 63996 36331
rect 63556 34819 63996 36245
rect 63556 34733 63649 34819
rect 63735 34733 63817 34819
rect 63903 34733 63996 34819
rect 63556 33307 63996 34733
rect 63556 33221 63649 33307
rect 63735 33221 63817 33307
rect 63903 33221 63996 33307
rect 63556 31795 63996 33221
rect 63556 31709 63649 31795
rect 63735 31709 63817 31795
rect 63903 31709 63996 31795
rect 63556 30283 63996 31709
rect 63556 30197 63649 30283
rect 63735 30197 63817 30283
rect 63903 30197 63996 30283
rect 63556 28771 63996 30197
rect 63556 28685 63649 28771
rect 63735 28685 63817 28771
rect 63903 28685 63996 28771
rect 63556 27259 63996 28685
rect 63556 27173 63649 27259
rect 63735 27173 63817 27259
rect 63903 27173 63996 27259
rect 63556 25747 63996 27173
rect 63556 25661 63649 25747
rect 63735 25661 63817 25747
rect 63903 25661 63996 25747
rect 63556 24235 63996 25661
rect 63556 24149 63649 24235
rect 63735 24149 63817 24235
rect 63903 24149 63996 24235
rect 63556 22723 63996 24149
rect 63556 22637 63649 22723
rect 63735 22637 63817 22723
rect 63903 22637 63996 22723
rect 63556 21211 63996 22637
rect 63556 21125 63649 21211
rect 63735 21125 63817 21211
rect 63903 21125 63996 21211
rect 63556 19699 63996 21125
rect 63556 19613 63649 19699
rect 63735 19613 63817 19699
rect 63903 19613 63996 19699
rect 63556 18187 63996 19613
rect 63556 18101 63649 18187
rect 63735 18101 63817 18187
rect 63903 18101 63996 18187
rect 63556 16675 63996 18101
rect 63556 16589 63649 16675
rect 63735 16589 63817 16675
rect 63903 16589 63996 16675
rect 63556 15163 63996 16589
rect 63556 15077 63649 15163
rect 63735 15077 63817 15163
rect 63903 15077 63996 15163
rect 63556 13651 63996 15077
rect 63556 13565 63649 13651
rect 63735 13565 63817 13651
rect 63903 13565 63996 13651
rect 63556 12139 63996 13565
rect 63556 12053 63649 12139
rect 63735 12053 63817 12139
rect 63903 12053 63996 12139
rect 63556 10627 63996 12053
rect 63556 10541 63649 10627
rect 63735 10541 63817 10627
rect 63903 10541 63996 10627
rect 63556 9115 63996 10541
rect 63556 9029 63649 9115
rect 63735 9029 63817 9115
rect 63903 9029 63996 9115
rect 63556 7603 63996 9029
rect 63556 7517 63649 7603
rect 63735 7517 63817 7603
rect 63903 7517 63996 7603
rect 63556 6091 63996 7517
rect 63556 6005 63649 6091
rect 63735 6005 63817 6091
rect 63903 6005 63996 6091
rect 63556 4579 63996 6005
rect 63556 4493 63649 4579
rect 63735 4493 63817 4579
rect 63903 4493 63996 4579
rect 63556 3067 63996 4493
rect 63556 2981 63649 3067
rect 63735 2981 63817 3067
rect 63903 2981 63996 3067
rect 63556 1555 63996 2981
rect 63556 1469 63649 1555
rect 63735 1469 63817 1555
rect 63903 1469 63996 1555
rect 63556 712 63996 1469
rect 64796 38599 65236 38682
rect 64796 38513 64889 38599
rect 64975 38513 65057 38599
rect 65143 38513 65236 38599
rect 64796 37087 65236 38513
rect 64796 37001 64889 37087
rect 64975 37001 65057 37087
rect 65143 37001 65236 37087
rect 64796 35575 65236 37001
rect 64796 35489 64889 35575
rect 64975 35489 65057 35575
rect 65143 35489 65236 35575
rect 64796 34063 65236 35489
rect 64796 33977 64889 34063
rect 64975 33977 65057 34063
rect 65143 33977 65236 34063
rect 64796 32551 65236 33977
rect 64796 32465 64889 32551
rect 64975 32465 65057 32551
rect 65143 32465 65236 32551
rect 64796 31039 65236 32465
rect 64796 30953 64889 31039
rect 64975 30953 65057 31039
rect 65143 30953 65236 31039
rect 64796 29527 65236 30953
rect 64796 29441 64889 29527
rect 64975 29441 65057 29527
rect 65143 29441 65236 29527
rect 64796 28015 65236 29441
rect 64796 27929 64889 28015
rect 64975 27929 65057 28015
rect 65143 27929 65236 28015
rect 64796 26503 65236 27929
rect 64796 26417 64889 26503
rect 64975 26417 65057 26503
rect 65143 26417 65236 26503
rect 64796 24991 65236 26417
rect 64796 24905 64889 24991
rect 64975 24905 65057 24991
rect 65143 24905 65236 24991
rect 64796 23479 65236 24905
rect 64796 23393 64889 23479
rect 64975 23393 65057 23479
rect 65143 23393 65236 23479
rect 64796 21967 65236 23393
rect 64796 21881 64889 21967
rect 64975 21881 65057 21967
rect 65143 21881 65236 21967
rect 64796 20455 65236 21881
rect 64796 20369 64889 20455
rect 64975 20369 65057 20455
rect 65143 20369 65236 20455
rect 64796 18943 65236 20369
rect 64796 18857 64889 18943
rect 64975 18857 65057 18943
rect 65143 18857 65236 18943
rect 64796 17431 65236 18857
rect 64796 17345 64889 17431
rect 64975 17345 65057 17431
rect 65143 17345 65236 17431
rect 64796 15919 65236 17345
rect 64796 15833 64889 15919
rect 64975 15833 65057 15919
rect 65143 15833 65236 15919
rect 64796 14407 65236 15833
rect 64796 14321 64889 14407
rect 64975 14321 65057 14407
rect 65143 14321 65236 14407
rect 64796 12895 65236 14321
rect 64796 12809 64889 12895
rect 64975 12809 65057 12895
rect 65143 12809 65236 12895
rect 64796 11383 65236 12809
rect 64796 11297 64889 11383
rect 64975 11297 65057 11383
rect 65143 11297 65236 11383
rect 64796 9871 65236 11297
rect 64796 9785 64889 9871
rect 64975 9785 65057 9871
rect 65143 9785 65236 9871
rect 64796 8359 65236 9785
rect 64796 8273 64889 8359
rect 64975 8273 65057 8359
rect 65143 8273 65236 8359
rect 64796 6847 65236 8273
rect 64796 6761 64889 6847
rect 64975 6761 65057 6847
rect 65143 6761 65236 6847
rect 64796 5335 65236 6761
rect 64796 5249 64889 5335
rect 64975 5249 65057 5335
rect 65143 5249 65236 5335
rect 64796 3823 65236 5249
rect 64796 3737 64889 3823
rect 64975 3737 65057 3823
rect 65143 3737 65236 3823
rect 64796 2311 65236 3737
rect 64796 2225 64889 2311
rect 64975 2225 65057 2311
rect 65143 2225 65236 2311
rect 64796 799 65236 2225
rect 64796 713 64889 799
rect 64975 713 65057 799
rect 65143 713 65236 799
rect 64796 630 65236 713
rect 78676 37843 79116 38600
rect 78676 37757 78769 37843
rect 78855 37757 78937 37843
rect 79023 37757 79116 37843
rect 78676 36331 79116 37757
rect 78676 36245 78769 36331
rect 78855 36245 78937 36331
rect 79023 36245 79116 36331
rect 78676 34819 79116 36245
rect 78676 34733 78769 34819
rect 78855 34733 78937 34819
rect 79023 34733 79116 34819
rect 78676 33307 79116 34733
rect 78676 33221 78769 33307
rect 78855 33221 78937 33307
rect 79023 33221 79116 33307
rect 78676 31795 79116 33221
rect 78676 31709 78769 31795
rect 78855 31709 78937 31795
rect 79023 31709 79116 31795
rect 78676 30283 79116 31709
rect 78676 30197 78769 30283
rect 78855 30197 78937 30283
rect 79023 30197 79116 30283
rect 78676 28771 79116 30197
rect 78676 28685 78769 28771
rect 78855 28685 78937 28771
rect 79023 28685 79116 28771
rect 78676 27259 79116 28685
rect 78676 27173 78769 27259
rect 78855 27173 78937 27259
rect 79023 27173 79116 27259
rect 78676 25747 79116 27173
rect 78676 25661 78769 25747
rect 78855 25661 78937 25747
rect 79023 25661 79116 25747
rect 78676 24235 79116 25661
rect 78676 24149 78769 24235
rect 78855 24149 78937 24235
rect 79023 24149 79116 24235
rect 78676 22723 79116 24149
rect 78676 22637 78769 22723
rect 78855 22637 78937 22723
rect 79023 22637 79116 22723
rect 78676 21211 79116 22637
rect 78676 21125 78769 21211
rect 78855 21125 78937 21211
rect 79023 21125 79116 21211
rect 78676 19699 79116 21125
rect 78676 19613 78769 19699
rect 78855 19613 78937 19699
rect 79023 19613 79116 19699
rect 78676 18187 79116 19613
rect 78676 18101 78769 18187
rect 78855 18101 78937 18187
rect 79023 18101 79116 18187
rect 78676 16675 79116 18101
rect 78676 16589 78769 16675
rect 78855 16589 78937 16675
rect 79023 16589 79116 16675
rect 78676 15163 79116 16589
rect 78676 15077 78769 15163
rect 78855 15077 78937 15163
rect 79023 15077 79116 15163
rect 78676 13651 79116 15077
rect 78676 13565 78769 13651
rect 78855 13565 78937 13651
rect 79023 13565 79116 13651
rect 78676 12139 79116 13565
rect 78676 12053 78769 12139
rect 78855 12053 78937 12139
rect 79023 12053 79116 12139
rect 78676 10627 79116 12053
rect 78676 10541 78769 10627
rect 78855 10541 78937 10627
rect 79023 10541 79116 10627
rect 78676 9115 79116 10541
rect 78676 9029 78769 9115
rect 78855 9029 78937 9115
rect 79023 9029 79116 9115
rect 78676 7603 79116 9029
rect 78676 7517 78769 7603
rect 78855 7517 78937 7603
rect 79023 7517 79116 7603
rect 78676 6091 79116 7517
rect 78676 6005 78769 6091
rect 78855 6005 78937 6091
rect 79023 6005 79116 6091
rect 78676 4579 79116 6005
rect 78676 4493 78769 4579
rect 78855 4493 78937 4579
rect 79023 4493 79116 4579
rect 78676 3067 79116 4493
rect 78676 2981 78769 3067
rect 78855 2981 78937 3067
rect 79023 2981 79116 3067
rect 78676 1555 79116 2981
rect 78676 1469 78769 1555
rect 78855 1469 78937 1555
rect 79023 1469 79116 1555
rect 78676 712 79116 1469
rect 79916 38599 80356 38682
rect 79916 38513 80009 38599
rect 80095 38513 80177 38599
rect 80263 38513 80356 38599
rect 79916 37087 80356 38513
rect 79916 37001 80009 37087
rect 80095 37001 80177 37087
rect 80263 37001 80356 37087
rect 79916 35575 80356 37001
rect 79916 35489 80009 35575
rect 80095 35489 80177 35575
rect 80263 35489 80356 35575
rect 79916 34063 80356 35489
rect 79916 33977 80009 34063
rect 80095 33977 80177 34063
rect 80263 33977 80356 34063
rect 79916 32551 80356 33977
rect 79916 32465 80009 32551
rect 80095 32465 80177 32551
rect 80263 32465 80356 32551
rect 79916 31039 80356 32465
rect 79916 30953 80009 31039
rect 80095 30953 80177 31039
rect 80263 30953 80356 31039
rect 79916 29527 80356 30953
rect 79916 29441 80009 29527
rect 80095 29441 80177 29527
rect 80263 29441 80356 29527
rect 79916 28015 80356 29441
rect 79916 27929 80009 28015
rect 80095 27929 80177 28015
rect 80263 27929 80356 28015
rect 79916 26503 80356 27929
rect 79916 26417 80009 26503
rect 80095 26417 80177 26503
rect 80263 26417 80356 26503
rect 79916 24991 80356 26417
rect 79916 24905 80009 24991
rect 80095 24905 80177 24991
rect 80263 24905 80356 24991
rect 79916 23479 80356 24905
rect 79916 23393 80009 23479
rect 80095 23393 80177 23479
rect 80263 23393 80356 23479
rect 79916 21967 80356 23393
rect 79916 21881 80009 21967
rect 80095 21881 80177 21967
rect 80263 21881 80356 21967
rect 79916 20455 80356 21881
rect 79916 20369 80009 20455
rect 80095 20369 80177 20455
rect 80263 20369 80356 20455
rect 79916 18943 80356 20369
rect 79916 18857 80009 18943
rect 80095 18857 80177 18943
rect 80263 18857 80356 18943
rect 79916 17431 80356 18857
rect 79916 17345 80009 17431
rect 80095 17345 80177 17431
rect 80263 17345 80356 17431
rect 79916 15919 80356 17345
rect 79916 15833 80009 15919
rect 80095 15833 80177 15919
rect 80263 15833 80356 15919
rect 79916 14407 80356 15833
rect 79916 14321 80009 14407
rect 80095 14321 80177 14407
rect 80263 14321 80356 14407
rect 79916 12895 80356 14321
rect 79916 12809 80009 12895
rect 80095 12809 80177 12895
rect 80263 12809 80356 12895
rect 79916 11383 80356 12809
rect 79916 11297 80009 11383
rect 80095 11297 80177 11383
rect 80263 11297 80356 11383
rect 79916 9871 80356 11297
rect 79916 9785 80009 9871
rect 80095 9785 80177 9871
rect 80263 9785 80356 9871
rect 79916 8359 80356 9785
rect 79916 8273 80009 8359
rect 80095 8273 80177 8359
rect 80263 8273 80356 8359
rect 79916 6847 80356 8273
rect 79916 6761 80009 6847
rect 80095 6761 80177 6847
rect 80263 6761 80356 6847
rect 79916 5335 80356 6761
rect 79916 5249 80009 5335
rect 80095 5249 80177 5335
rect 80263 5249 80356 5335
rect 79916 3823 80356 5249
rect 79916 3737 80009 3823
rect 80095 3737 80177 3823
rect 80263 3737 80356 3823
rect 79916 2311 80356 3737
rect 79916 2225 80009 2311
rect 80095 2225 80177 2311
rect 80263 2225 80356 2311
rect 79916 799 80356 2225
rect 79916 713 80009 799
rect 80095 713 80177 799
rect 80263 713 80356 799
rect 79916 630 80356 713
rect 93796 37843 94236 38600
rect 93796 37757 93889 37843
rect 93975 37757 94057 37843
rect 94143 37757 94236 37843
rect 93796 36331 94236 37757
rect 93796 36245 93889 36331
rect 93975 36245 94057 36331
rect 94143 36245 94236 36331
rect 93796 34819 94236 36245
rect 93796 34733 93889 34819
rect 93975 34733 94057 34819
rect 94143 34733 94236 34819
rect 93796 33307 94236 34733
rect 93796 33221 93889 33307
rect 93975 33221 94057 33307
rect 94143 33221 94236 33307
rect 93796 31795 94236 33221
rect 93796 31709 93889 31795
rect 93975 31709 94057 31795
rect 94143 31709 94236 31795
rect 93796 30283 94236 31709
rect 93796 30197 93889 30283
rect 93975 30197 94057 30283
rect 94143 30197 94236 30283
rect 93796 28771 94236 30197
rect 93796 28685 93889 28771
rect 93975 28685 94057 28771
rect 94143 28685 94236 28771
rect 93796 27259 94236 28685
rect 93796 27173 93889 27259
rect 93975 27173 94057 27259
rect 94143 27173 94236 27259
rect 93796 25747 94236 27173
rect 93796 25661 93889 25747
rect 93975 25661 94057 25747
rect 94143 25661 94236 25747
rect 93796 24235 94236 25661
rect 93796 24149 93889 24235
rect 93975 24149 94057 24235
rect 94143 24149 94236 24235
rect 93796 22723 94236 24149
rect 93796 22637 93889 22723
rect 93975 22637 94057 22723
rect 94143 22637 94236 22723
rect 93796 21211 94236 22637
rect 93796 21125 93889 21211
rect 93975 21125 94057 21211
rect 94143 21125 94236 21211
rect 93796 19699 94236 21125
rect 93796 19613 93889 19699
rect 93975 19613 94057 19699
rect 94143 19613 94236 19699
rect 93796 18187 94236 19613
rect 93796 18101 93889 18187
rect 93975 18101 94057 18187
rect 94143 18101 94236 18187
rect 93796 16675 94236 18101
rect 93796 16589 93889 16675
rect 93975 16589 94057 16675
rect 94143 16589 94236 16675
rect 93796 15163 94236 16589
rect 93796 15077 93889 15163
rect 93975 15077 94057 15163
rect 94143 15077 94236 15163
rect 93796 13651 94236 15077
rect 93796 13565 93889 13651
rect 93975 13565 94057 13651
rect 94143 13565 94236 13651
rect 93796 12139 94236 13565
rect 93796 12053 93889 12139
rect 93975 12053 94057 12139
rect 94143 12053 94236 12139
rect 93796 10627 94236 12053
rect 93796 10541 93889 10627
rect 93975 10541 94057 10627
rect 94143 10541 94236 10627
rect 93796 9115 94236 10541
rect 93796 9029 93889 9115
rect 93975 9029 94057 9115
rect 94143 9029 94236 9115
rect 93796 7603 94236 9029
rect 93796 7517 93889 7603
rect 93975 7517 94057 7603
rect 94143 7517 94236 7603
rect 93796 6091 94236 7517
rect 93796 6005 93889 6091
rect 93975 6005 94057 6091
rect 94143 6005 94236 6091
rect 93796 4579 94236 6005
rect 93796 4493 93889 4579
rect 93975 4493 94057 4579
rect 94143 4493 94236 4579
rect 93796 3067 94236 4493
rect 93796 2981 93889 3067
rect 93975 2981 94057 3067
rect 94143 2981 94236 3067
rect 93796 1555 94236 2981
rect 93796 1469 93889 1555
rect 93975 1469 94057 1555
rect 94143 1469 94236 1555
rect 93796 712 94236 1469
rect 95036 38599 95476 38682
rect 95036 38513 95129 38599
rect 95215 38513 95297 38599
rect 95383 38513 95476 38599
rect 95036 37087 95476 38513
rect 95036 37001 95129 37087
rect 95215 37001 95297 37087
rect 95383 37001 95476 37087
rect 95036 35575 95476 37001
rect 95036 35489 95129 35575
rect 95215 35489 95297 35575
rect 95383 35489 95476 35575
rect 95036 34063 95476 35489
rect 95036 33977 95129 34063
rect 95215 33977 95297 34063
rect 95383 33977 95476 34063
rect 95036 32551 95476 33977
rect 95036 32465 95129 32551
rect 95215 32465 95297 32551
rect 95383 32465 95476 32551
rect 95036 31039 95476 32465
rect 95036 30953 95129 31039
rect 95215 30953 95297 31039
rect 95383 30953 95476 31039
rect 95036 29527 95476 30953
rect 95036 29441 95129 29527
rect 95215 29441 95297 29527
rect 95383 29441 95476 29527
rect 95036 28015 95476 29441
rect 95036 27929 95129 28015
rect 95215 27929 95297 28015
rect 95383 27929 95476 28015
rect 95036 26503 95476 27929
rect 95036 26417 95129 26503
rect 95215 26417 95297 26503
rect 95383 26417 95476 26503
rect 95036 24991 95476 26417
rect 95036 24905 95129 24991
rect 95215 24905 95297 24991
rect 95383 24905 95476 24991
rect 95036 23479 95476 24905
rect 95036 23393 95129 23479
rect 95215 23393 95297 23479
rect 95383 23393 95476 23479
rect 95036 21967 95476 23393
rect 95036 21881 95129 21967
rect 95215 21881 95297 21967
rect 95383 21881 95476 21967
rect 95036 20455 95476 21881
rect 95036 20369 95129 20455
rect 95215 20369 95297 20455
rect 95383 20369 95476 20455
rect 95036 18943 95476 20369
rect 95036 18857 95129 18943
rect 95215 18857 95297 18943
rect 95383 18857 95476 18943
rect 95036 17431 95476 18857
rect 95036 17345 95129 17431
rect 95215 17345 95297 17431
rect 95383 17345 95476 17431
rect 95036 15919 95476 17345
rect 95036 15833 95129 15919
rect 95215 15833 95297 15919
rect 95383 15833 95476 15919
rect 95036 14407 95476 15833
rect 95036 14321 95129 14407
rect 95215 14321 95297 14407
rect 95383 14321 95476 14407
rect 95036 12895 95476 14321
rect 95036 12809 95129 12895
rect 95215 12809 95297 12895
rect 95383 12809 95476 12895
rect 95036 11383 95476 12809
rect 95036 11297 95129 11383
rect 95215 11297 95297 11383
rect 95383 11297 95476 11383
rect 95036 9871 95476 11297
rect 95036 9785 95129 9871
rect 95215 9785 95297 9871
rect 95383 9785 95476 9871
rect 95036 8359 95476 9785
rect 95036 8273 95129 8359
rect 95215 8273 95297 8359
rect 95383 8273 95476 8359
rect 95036 6847 95476 8273
rect 95036 6761 95129 6847
rect 95215 6761 95297 6847
rect 95383 6761 95476 6847
rect 95036 5335 95476 6761
rect 95036 5249 95129 5335
rect 95215 5249 95297 5335
rect 95383 5249 95476 5335
rect 95036 3823 95476 5249
rect 95036 3737 95129 3823
rect 95215 3737 95297 3823
rect 95383 3737 95476 3823
rect 95036 2311 95476 3737
rect 95036 2225 95129 2311
rect 95215 2225 95297 2311
rect 95383 2225 95476 2311
rect 95036 799 95476 2225
rect 95036 713 95129 799
rect 95215 713 95297 799
rect 95383 713 95476 799
rect 95036 630 95476 713
use sg13g2_and2_1  _222_
timestamp 1676905363
transform 1 0 10368 0 1 34020
box -48 -56 528 834
use sg13g2_and2_1  _223_
timestamp 1676905363
transform 1 0 12480 0 -1 3780
box -48 -56 528 834
use sg13g2_nand2_1  _224_
timestamp 1676560849
transform 1 0 29568 0 -1 6804
box -48 -56 432 834
use sg13g2_xor2_1  _225_
timestamp 1677581577
transform -1 0 28992 0 1 6804
box -48 -56 816 834
use sg13g2_and2_1  _226_
timestamp 1676905363
transform -1 0 37056 0 -1 35532
box -48 -56 528 834
use sg13g2_and2_1  _227_
timestamp 1676905363
transform 1 0 19968 0 1 30996
box -48 -56 528 834
use sg13g2_and2_1  _228_
timestamp 1676905363
transform 1 0 5184 0 -1 9828
box -48 -56 528 834
use sg13g2_nand2_1  _229_
timestamp 1676560849
transform 1 0 30528 0 1 6804
box -48 -56 432 834
use sg13g2_nor2_1  _230_
timestamp 1676630787
transform -1 0 30336 0 1 8316
box -48 -56 432 834
use sg13g2_xor2_1  _231_
timestamp 1677581577
transform -1 0 30528 0 1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _232_
timestamp 1677520200
transform -1 0 29760 0 1 6804
box -48 -56 816 834
use sg13g2_and2_1  _233_
timestamp 1676905363
transform 1 0 11712 0 -1 18900
box -48 -56 528 834
use sg13g2_and2_1  _234_
timestamp 1676905363
transform -1 0 39168 0 -1 23436
box -48 -56 528 834
use sg13g2_and2_1  _235_
timestamp 1676905363
transform 1 0 33696 0 -1 21924
box -48 -56 528 834
use sg13g2_and2_1  _236_
timestamp 1676905363
transform 1 0 32160 0 1 12852
box -48 -56 528 834
use sg13g2_and2_1  _237_
timestamp 1676905363
transform 1 0 26976 0 1 17388
box -48 -56 528 834
use sg13g2_and2_1  _238_
timestamp 1676905363
transform -1 0 55296 0 -1 12852
box -48 -56 528 834
use sg13g2_and2_1  _239_
timestamp 1676905363
transform 1 0 48000 0 1 17388
box -48 -56 528 834
use sg13g2_and2_1  _240_
timestamp 1676905363
transform 1 0 40320 0 1 3780
box -48 -56 528 834
use sg13g2_and2_1  _241_
timestamp 1676905363
transform -1 0 52320 0 -1 5292
box -48 -56 528 834
use sg13g2_and2_1  _242_
timestamp 1676905363
transform 1 0 6336 0 1 27972
box -48 -56 528 834
use sg13g2_and2_1  _243_
timestamp 1676905363
transform -1 0 25920 0 -1 35532
box -48 -56 528 834
use sg13g2_and2_1  _244_
timestamp 1676905363
transform -1 0 46080 0 1 29484
box -48 -56 528 834
use sg13g2_and2_1  _245_
timestamp 1676905363
transform 1 0 5952 0 -1 23436
box -48 -56 528 834
use sg13g2_nand2_1  _246_
timestamp 1676560849
transform -1 0 41664 0 -1 9828
box -48 -56 432 834
use sg13g2_xor2_1  _247_
timestamp 1677581577
transform -1 0 40512 0 -1 8316
box -48 -56 816 834
use sg13g2_xor2_1  _248_
timestamp 1677581577
transform -1 0 44256 0 -1 11340
box -48 -56 816 834
use sg13g2_xnor2_1  _249_
timestamp 1677520200
transform -1 0 41280 0 1 8316
box -48 -56 816 834
use sg13g2_nand2_1  _250_
timestamp 1676560849
transform -1 0 18720 0 -1 24948
box -48 -56 432 834
use sg13g2_xor2_1  _251_
timestamp 1677581577
transform 1 0 16704 0 1 24948
box -48 -56 816 834
use sg13g2_xnor2_1  _252_
timestamp 1677520200
transform 1 0 17568 0 1 24948
box -48 -56 816 834
use sg13g2_xor2_1  _253_
timestamp 1677581577
transform 1 0 18528 0 -1 23436
box -48 -56 816 834
use sg13g2_nand2_1  _254_
timestamp 1676560849
transform 1 0 22560 0 -1 21924
box -48 -56 432 834
use sg13g2_xor2_1  _255_
timestamp 1677581577
transform 1 0 22752 0 1 24948
box -48 -56 816 834
use sg13g2_xnor2_1  _256_
timestamp 1677520200
transform -1 0 22272 0 -1 23436
box -48 -56 816 834
use sg13g2_xor2_1  _257_
timestamp 1677581577
transform -1 0 22560 0 -1 21924
box -48 -56 816 834
use sg13g2_nand2_1  _258_
timestamp 1676560849
transform 1 0 19680 0 1 8316
box -48 -56 432 834
use sg13g2_nand2_1  _259_
timestamp 1676560849
transform 1 0 21984 0 1 8316
box -48 -56 432 834
use sg13g2_nor2_1  _260_
timestamp 1676630787
transform 1 0 20832 0 1 8316
box -48 -56 432 834
use sg13g2_xor2_1  _261_
timestamp 1677581577
transform -1 0 22464 0 -1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _262_
timestamp 1677520200
transform -1 0 21984 0 1 8316
box -48 -56 816 834
use sg13g2_o21ai_1  _263_
timestamp 1685179043
transform 1 0 22848 0 -1 8316
box -48 -56 538 834
use sg13g2_and2_1  _264_
timestamp 1676905363
transform -1 0 26592 0 -1 9828
box -48 -56 528 834
use sg13g2_or2_1  _265_
timestamp 1684239771
transform -1 0 27072 0 -1 9828
box -48 -56 528 834
use sg13g2_nand2b_1  _266_
timestamp 1676570795
transform -1 0 26208 0 1 8316
box -48 -56 528 834
use sg13g2_xnor2_1  _267_
timestamp 1677520200
transform -1 0 26112 0 1 9828
box -48 -56 816 834
use sg13g2_xor2_1  _268_
timestamp 1677581577
transform -1 0 19296 0 -1 8316
box -48 -56 816 834
use sg13g2_nand2_1  _269_
timestamp 1676560849
transform 1 0 39648 0 -1 20412
box -48 -56 432 834
use sg13g2_xor2_1  _270_
timestamp 1677581577
transform 1 0 40224 0 1 24948
box -48 -56 816 834
use sg13g2_xnor2_1  _271_
timestamp 1677520200
transform 1 0 40224 0 -1 20412
box -48 -56 816 834
use sg13g2_xor2_1  _272_
timestamp 1677581577
transform 1 0 39264 0 1 18900
box -48 -56 816 834
use sg13g2_nand2_1  _273_
timestamp 1676560849
transform 1 0 35616 0 -1 15876
box -48 -56 432 834
use sg13g2_xor2_1  _274_
timestamp 1677581577
transform 1 0 33504 0 -1 17388
box -48 -56 816 834
use sg13g2_xnor2_1  _275_
timestamp 1677520200
transform 1 0 35712 0 1 15876
box -48 -56 816 834
use sg13g2_xor2_1  _276_
timestamp 1677581577
transform 1 0 35904 0 1 14364
box -48 -56 816 834
use sg13g2_nand2_1  _277_
timestamp 1676560849
transform 1 0 51168 0 1 14364
box -48 -56 432 834
use sg13g2_xor2_1  _278_
timestamp 1677581577
transform 1 0 54432 0 -1 17388
box -48 -56 816 834
use sg13g2_xnor2_1  _279_
timestamp 1677520200
transform -1 0 53280 0 1 14364
box -48 -56 816 834
use sg13g2_xor2_1  _280_
timestamp 1677581577
transform -1 0 53568 0 -1 14364
box -48 -56 816 834
use sg13g2_nand2_1  _281_
timestamp 1676560849
transform 1 0 46368 0 1 5292
box -48 -56 432 834
use sg13g2_xor2_1  _282_
timestamp 1677581577
transform -1 0 48192 0 -1 3780
box -48 -56 816 834
use sg13g2_xnor2_1  _283_
timestamp 1677520200
transform 1 0 46848 0 1 5292
box -48 -56 816 834
use sg13g2_xor2_1  _284_
timestamp 1677581577
transform 1 0 44736 0 -1 6804
box -48 -56 816 834
use sg13g2_nand2_1  _285_
timestamp 1676560849
transform 1 0 40704 0 1 14364
box -48 -56 432 834
use sg13g2_xor2_1  _286_
timestamp 1677581577
transform 1 0 41376 0 1 17388
box -48 -56 816 834
use sg13g2_xnor2_1  _287_
timestamp 1677520200
transform -1 0 41952 0 1 14364
box -48 -56 816 834
use sg13g2_xor2_1  _288_
timestamp 1677581577
transform 1 0 39744 0 1 12852
box -48 -56 816 834
use sg13g2_nand2_1  _289_
timestamp 1676560849
transform 1 0 46848 0 1 9828
box -48 -56 432 834
use sg13g2_xor2_1  _290_
timestamp 1677581577
transform -1 0 50400 0 1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _291_
timestamp 1677520200
transform -1 0 48864 0 1 9828
box -48 -56 816 834
use sg13g2_xor2_1  _292_
timestamp 1677581577
transform -1 0 47808 0 -1 9828
box -48 -56 816 834
use sg13g2_nand2_1  _293_
timestamp 1676560849
transform 1 0 17088 0 1 11340
box -48 -56 432 834
use sg13g2_nand2_1  _294_
timestamp 1676560849
transform -1 0 20544 0 1 12852
box -48 -56 432 834
use sg13g2_nor2_1  _295_
timestamp 1676630787
transform 1 0 18528 0 -1 14364
box -48 -56 432 834
use sg13g2_xor2_1  _296_
timestamp 1677581577
transform -1 0 19200 0 1 12852
box -48 -56 816 834
use sg13g2_xnor2_1  _297_
timestamp 1677520200
transform 1 0 18144 0 -1 12852
box -48 -56 816 834
use sg13g2_xor2_1  _298_
timestamp 1677581577
transform 1 0 15936 0 1 9828
box -48 -56 816 834
use sg13g2_nand2_1  _299_
timestamp 1676560849
transform -1 0 13248 0 1 27972
box -48 -56 432 834
use sg13g2_xor2_1  _300_
timestamp 1677581577
transform 1 0 11040 0 1 29484
box -48 -56 816 834
use sg13g2_xnor2_1  _301_
timestamp 1677520200
transform 1 0 12096 0 -1 29484
box -48 -56 816 834
use sg13g2_xor2_1  _302_
timestamp 1677581577
transform 1 0 13632 0 -1 27972
box -48 -56 816 834
use sg13g2_nand2_1  _303_
timestamp 1676560849
transform -1 0 26496 0 1 30996
box -48 -56 432 834
use sg13g2_xor2_1  _304_
timestamp 1677581577
transform 1 0 24096 0 1 34020
box -48 -56 816 834
use sg13g2_xnor2_1  _305_
timestamp 1677520200
transform 1 0 25920 0 -1 32508
box -48 -56 816 834
use sg13g2_xor2_1  _306_
timestamp 1677581577
transform -1 0 27552 0 -1 30996
box -48 -56 816 834
use sg13g2_nand2_1  _307_
timestamp 1676560849
transform 1 0 37824 0 1 29484
box -48 -56 432 834
use sg13g2_xor2_1  _308_
timestamp 1677581577
transform -1 0 43488 0 -1 32508
box -48 -56 816 834
use sg13g2_xnor2_1  _309_
timestamp 1677520200
transform -1 0 38784 0 -1 32508
box -48 -56 816 834
use sg13g2_xor2_1  _310_
timestamp 1677581577
transform -1 0 37824 0 1 29484
box -48 -56 816 834
use sg13g2_nand2_1  _311_
timestamp 1676560849
transform 1 0 28416 0 -1 29484
box -48 -56 432 834
use sg13g2_xor2_1  _312_
timestamp 1677581577
transform 1 0 30528 0 -1 30996
box -48 -56 816 834
use sg13g2_xnor2_1  _313_
timestamp 1677520200
transform 1 0 28416 0 1 27972
box -48 -56 816 834
use sg13g2_xor2_1  _314_
timestamp 1677581577
transform -1 0 28416 0 1 27972
box -48 -56 816 834
use sg13g2_nand2_1  _315_
timestamp 1676560849
transform -1 0 14208 0 1 21924
box -48 -56 432 834
use sg13g2_xor2_1  _316_
timestamp 1677581577
transform 1 0 11040 0 1 21924
box -48 -56 816 834
use sg13g2_xnor2_1  _317_
timestamp 1677520200
transform -1 0 14400 0 -1 23436
box -48 -56 816 834
use sg13g2_xor2_1  _318_
timestamp 1677581577
transform 1 0 14400 0 1 21924
box -48 -56 816 834
use sg13g2_o21ai_1  _319_
timestamp 1685179043
transform -1 0 29952 0 -1 8316
box -48 -56 538 834
use sg13g2_nand2_1  _320_
timestamp 1676560849
transform 1 0 8832 0 -1 35532
box -48 -56 432 834
use sg13g2_nand2_1  _321_
timestamp 1676560849
transform -1 0 10752 0 1 35532
box -48 -56 432 834
use sg13g2_xor2_1  _322_
timestamp 1677581577
transform 1 0 9216 0 1 34020
box -48 -56 816 834
use sg13g2_nand2_1  _323_
timestamp 1676560849
transform 1 0 10848 0 -1 3780
box -48 -56 432 834
use sg13g2_nand2_1  _324_
timestamp 1676560849
transform 1 0 11232 0 -1 3780
box -48 -56 432 834
use sg13g2_xor2_1  _325_
timestamp 1677581577
transform 1 0 11616 0 1 2268
box -48 -56 816 834
use sg13g2_nand2_1  _326_
timestamp 1676560849
transform 1 0 37056 0 -1 35532
box -48 -56 432 834
use sg13g2_nand2_1  _327_
timestamp 1676560849
transform -1 0 39936 0 1 35532
box -48 -56 432 834
use sg13g2_xor2_1  _328_
timestamp 1677581577
transform 1 0 38976 0 -1 35532
box -48 -56 816 834
use sg13g2_nand2_1  _329_
timestamp 1676560849
transform 1 0 18240 0 -1 34020
box -48 -56 432 834
use sg13g2_nand2_1  _330_
timestamp 1676560849
transform 1 0 17952 0 1 32508
box -48 -56 432 834
use sg13g2_xor2_1  _331_
timestamp 1677581577
transform 1 0 18624 0 -1 34020
box -48 -56 816 834
use sg13g2_a21o_2  _332_
timestamp 1683999997
transform 1 0 25344 0 -1 9828
box -48 -56 816 834
use sg13g2_nand2_1  _333_
timestamp 1676560849
transform 1 0 3840 0 1 11340
box -48 -56 432 834
use sg13g2_nand2_1  _334_
timestamp 1676560849
transform 1 0 3072 0 -1 9828
box -48 -56 432 834
use sg13g2_xor2_1  _335_
timestamp 1677581577
transform 1 0 5088 0 1 11340
box -48 -56 816 834
use sg13g2_nand2_1  _336_
timestamp 1676560849
transform 1 0 8160 0 -1 17388
box -48 -56 432 834
use sg13g2_nand2_1  _337_
timestamp 1676560849
transform 1 0 8736 0 1 17388
box -48 -56 432 834
use sg13g2_xor2_1  _338_
timestamp 1677581577
transform 1 0 8160 0 -1 18900
box -48 -56 816 834
use sg13g2_nand2_1  _339_
timestamp 1676560849
transform -1 0 39840 0 1 24948
box -48 -56 432 834
use sg13g2_nand2_1  _340_
timestamp 1676560849
transform -1 0 43104 0 1 23436
box -48 -56 432 834
use sg13g2_xor2_1  _341_
timestamp 1677581577
transform 1 0 41184 0 1 24948
box -48 -56 816 834
use sg13g2_nand2_1  _342_
timestamp 1676560849
transform 1 0 31584 0 -1 23436
box -48 -56 432 834
use sg13g2_nand2_1  _343_
timestamp 1676560849
transform 1 0 31776 0 -1 24948
box -48 -56 432 834
use sg13g2_xor2_1  _344_
timestamp 1677581577
transform 1 0 32160 0 -1 24948
box -48 -56 816 834
use sg13g2_nand2_1  _345_
timestamp 1676560849
transform -1 0 31488 0 1 11340
box -48 -56 432 834
use sg13g2_nand2_1  _346_
timestamp 1676560849
transform 1 0 28800 0 1 12852
box -48 -56 432 834
use sg13g2_xor2_1  _347_
timestamp 1677581577
transform -1 0 31008 0 1 12852
box -48 -56 816 834
use sg13g2_nand2_1  _348_
timestamp 1676560849
transform 1 0 26496 0 1 18900
box -48 -56 432 834
use sg13g2_nand2_1  _349_
timestamp 1676560849
transform 1 0 26400 0 1 17388
box -48 -56 432 834
use sg13g2_xor2_1  _350_
timestamp 1677581577
transform 1 0 27456 0 1 17388
box -48 -56 816 834
use sg13g2_nand2_1  _351_
timestamp 1676560849
transform -1 0 56928 0 -1 12852
box -48 -56 432 834
use sg13g2_nand2_1  _352_
timestamp 1676560849
transform -1 0 56064 0 -1 11340
box -48 -56 432 834
use sg13g2_xor2_1  _353_
timestamp 1677581577
transform 1 0 55392 0 -1 14364
box -48 -56 816 834
use sg13g2_nand2_1  _354_
timestamp 1676560849
transform -1 0 49632 0 -1 20412
box -48 -56 432 834
use sg13g2_nand2_1  _355_
timestamp 1676560849
transform -1 0 50016 0 -1 20412
box -48 -56 432 834
use sg13g2_xor2_1  _356_
timestamp 1677581577
transform 1 0 50112 0 1 18900
box -48 -56 816 834
use sg13g2_nand2_1  _357_
timestamp 1676560849
transform 1 0 40128 0 -1 3780
box -48 -56 432 834
use sg13g2_nand2_1  _358_
timestamp 1676560849
transform 1 0 39936 0 1 3780
box -48 -56 432 834
use sg13g2_xor2_1  _359_
timestamp 1677581577
transform 1 0 40992 0 1 3780
box -48 -56 816 834
use sg13g2_nand2_1  _360_
timestamp 1676560849
transform -1 0 52224 0 -1 3780
box -48 -56 432 834
use sg13g2_nand2_1  _361_
timestamp 1676560849
transform -1 0 54336 0 1 3780
box -48 -56 432 834
use sg13g2_xor2_1  _362_
timestamp 1677581577
transform 1 0 53088 0 -1 3780
box -48 -56 816 834
use sg13g2_o21ai_1  _363_
timestamp 1685179043
transform 1 0 19776 0 -1 12852
box -48 -56 538 834
use sg13g2_nand2_1  _364_
timestamp 1676560849
transform 1 0 3936 0 -1 30996
box -48 -56 432 834
use sg13g2_nand2_1  _365_
timestamp 1676560849
transform 1 0 4992 0 -1 29484
box -48 -56 432 834
use sg13g2_xor2_1  _366_
timestamp 1677581577
transform 1 0 5088 0 1 29484
box -48 -56 816 834
use sg13g2_nand2_1  _367_
timestamp 1676560849
transform 1 0 21696 0 1 35532
box -48 -56 432 834
use sg13g2_nand2_1  _368_
timestamp 1676560849
transform -1 0 26496 0 1 35532
box -48 -56 432 834
use sg13g2_xor2_1  _369_
timestamp 1677581577
transform 1 0 22080 0 1 37044
box -48 -56 816 834
use sg13g2_nand2_1  _370_
timestamp 1676560849
transform -1 0 47136 0 -1 29484
box -48 -56 432 834
use sg13g2_nand2_1  _371_
timestamp 1676560849
transform -1 0 48672 0 -1 30996
box -48 -56 432 834
use sg13g2_xor2_1  _372_
timestamp 1677581577
transform 1 0 47328 0 1 29484
box -48 -56 816 834
use sg13g2_nand2_1  _373_
timestamp 1676560849
transform 1 0 4032 0 1 23436
box -48 -56 432 834
use sg13g2_nand2_1  _374_
timestamp 1676560849
transform 1 0 4032 0 1 21924
box -48 -56 432 834
use sg13g2_xor2_1  _375_
timestamp 1677581577
transform 1 0 5184 0 -1 23436
box -48 -56 816 834
use sg13g2_buf_1  _376_
timestamp 1676385511
transform 1 0 42144 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  _377_
timestamp 1676385511
transform -1 0 38496 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  _378_
timestamp 1676385511
transform -1 0 32640 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  _379_
timestamp 1676385511
transform 1 0 29568 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  _380_
timestamp 1676385511
transform -1 0 28704 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  _381_
timestamp 1676385511
transform -1 0 31968 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  _382_
timestamp 1676385511
transform -1 0 26208 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  _383_
timestamp 1676385511
transform -1 0 26208 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  _384_
timestamp 1676385511
transform -1 0 54144 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  _385_
timestamp 1676385511
transform -1 0 57120 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  _386_
timestamp 1676385511
transform -1 0 47904 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  _387_
timestamp 1676385511
transform -1 0 48384 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  _388_
timestamp 1676385511
transform -1 0 34560 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _389_
timestamp 1676385511
transform -1 0 38496 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _390_
timestamp 1676385511
transform 1 0 52128 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _391_
timestamp 1676385511
transform -1 0 54816 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _392_
timestamp 1676385511
transform -1 0 12096 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _393_
timestamp 1676385511
transform -1 0 8544 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _394_
timestamp 1676385511
transform -1 0 38016 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  _395_
timestamp 1676385511
transform 1 0 43104 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  _396_
timestamp 1676385511
transform -1 0 31200 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  _397_
timestamp 1676385511
transform -1 0 32160 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  _398_
timestamp 1676385511
transform -1 0 32352 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _399_
timestamp 1676385511
transform -1 0 25440 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  _400_
timestamp 1676385511
transform -1 0 22080 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  _401_
timestamp 1676385511
transform -1 0 24096 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  _402_
timestamp 1676385511
transform -1 0 56544 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _403_
timestamp 1676385511
transform -1 0 55872 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  _404_
timestamp 1676385511
transform -1 0 47520 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  _405_
timestamp 1676385511
transform -1 0 49344 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  _406_
timestamp 1676385511
transform -1 0 40128 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _407_
timestamp 1676385511
transform -1 0 38880 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _408_
timestamp 1676385511
transform -1 0 51552 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _409_
timestamp 1676385511
transform 1 0 54336 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _410_
timestamp 1676385511
transform 1 0 10752 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _411_
timestamp 1676385511
transform -1 0 8160 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _412_
timestamp 1676385511
transform -1 0 3744 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  _413_
timestamp 1676385511
transform -1 0 3552 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  _414_
timestamp 1676385511
transform -1 0 11136 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  _415_
timestamp 1676385511
transform -1 0 5568 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  _416_
timestamp 1676385511
transform -1 0 7488 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _417_
timestamp 1676385511
transform 1 0 10464 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _418_
timestamp 1676385511
transform -1 0 4800 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  _419_
timestamp 1676385511
transform -1 0 2496 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  _420_
timestamp 1676385511
transform -1 0 18240 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  _421_
timestamp 1676385511
transform -1 0 17184 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _422_
timestamp 1676385511
transform -1 0 25824 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _423_
timestamp 1676385511
transform -1 0 18240 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _424_
timestamp 1676385511
transform 1 0 46656 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  _425_
timestamp 1676385511
transform -1 0 47136 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  _426_
timestamp 1676385511
transform -1 0 37728 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _427_
timestamp 1676385511
transform -1 0 34464 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _428_
timestamp 1676385511
transform -1 0 3072 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _429_
timestamp 1676385511
transform -1 0 2496 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _430_
timestamp 1676385511
transform -1 0 3744 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  _431_
timestamp 1676385511
transform -1 0 2976 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  _432_
timestamp 1676385511
transform 1 0 10272 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  _433_
timestamp 1676385511
transform -1 0 6912 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  _434_
timestamp 1676385511
transform -1 0 11136 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _435_
timestamp 1676385511
transform -1 0 6240 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _436_
timestamp 1676385511
transform -1 0 3648 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  _437_
timestamp 1676385511
transform -1 0 3552 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  _438_
timestamp 1676385511
transform -1 0 18336 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  _439_
timestamp 1676385511
transform -1 0 15840 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  _440_
timestamp 1676385511
transform -1 0 23904 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  _441_
timestamp 1676385511
transform 1 0 27360 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _442_
timestamp 1676385511
transform -1 0 45024 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  _443_
timestamp 1676385511
transform 1 0 48672 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  _444_
timestamp 1676385511
transform -1 0 34464 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _445_
timestamp 1676385511
transform -1 0 39936 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _446_
timestamp 1676385511
transform -1 0 3552 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _447_
timestamp 1676385511
transform -1 0 2592 0 -1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _448_
timestamp 1746538728
transform 1 0 37344 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _449_
timestamp 1746538728
transform 1 0 41280 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _450_
timestamp 1746538728
transform 1 0 36000 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _451_
timestamp 1746538728
transform 1 0 34464 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _452_
timestamp 1746538728
transform 1 0 33600 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _453_
timestamp 1746538728
transform 1 0 30528 0 -1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _454_
timestamp 1746538728
transform 1 0 30912 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _455_
timestamp 1746538728
transform 1 0 29856 0 1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _456_
timestamp 1746538728
transform -1 0 54336 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _457_
timestamp 1746538728
transform -1 0 57792 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _458_
timestamp 1746538728
transform 1 0 49152 0 -1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _459_
timestamp 1746538728
transform 1 0 51936 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _460_
timestamp 1746538728
transform 1 0 41184 0 -1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _461_
timestamp 1746538728
transform 1 0 43968 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _462_
timestamp 1746538728
transform -1 0 47808 0 -1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _463_
timestamp 1746538728
transform -1 0 49632 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _464_
timestamp 1746538728
transform 1 0 14016 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _465_
timestamp 1746538728
transform 1 0 17568 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _466_
timestamp 1746538728
transform 1 0 39936 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _467_
timestamp 1746538728
transform 1 0 40992 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _468_
timestamp 1746538728
transform 1 0 37152 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _469_
timestamp 1746538728
transform 1 0 37152 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _470_
timestamp 1746538728
transform -1 0 48480 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _471_
timestamp 1746538728
transform -1 0 50496 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _472_
timestamp 1746538728
transform 1 0 45408 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _473_
timestamp 1746538728
transform 1 0 48288 0 1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _474_
timestamp 1746538728
transform 1 0 17376 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _475_
timestamp 1746538728
transform 1 0 21312 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _476_
timestamp 1746538728
transform -1 0 40896 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _477_
timestamp 1746538728
transform 1 0 41376 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _478_
timestamp 1746538728
transform -1 0 41280 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _479_
timestamp 1746538728
transform -1 0 46656 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _480_
timestamp 1746538728
transform 1 0 22080 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _481_
timestamp 1746538728
transform 1 0 24672 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _482_
timestamp 1746538728
transform -1 0 36000 0 1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_2  _483_
timestamp 1746538784
transform -1 0 36096 0 -1 8316
box -48 -56 2736 834
use sg13g2_dfrbpq_1  _484_
timestamp 1746538728
transform 1 0 26400 0 -1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _485_
timestamp 1746538728
transform 1 0 27840 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _486_
timestamp 1746538728
transform 1 0 16128 0 1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _487_
timestamp 1746538728
transform -1 0 22848 0 1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _488_
timestamp 1746538728
transform -1 0 27456 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _489_
timestamp 1746538728
transform 1 0 9024 0 1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _490_
timestamp 1746538728
transform 1 0 7488 0 -1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _491_
timestamp 1746538728
transform 1 0 12960 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _492_
timestamp 1746538728
transform 1 0 8640 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _493_
timestamp 1746538728
transform 1 0 10944 0 -1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _494_
timestamp 1746538728
transform 1 0 9216 0 1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _495_
timestamp 1746538728
transform 1 0 8544 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _496_
timestamp 1746538728
transform 1 0 7200 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _497_
timestamp 1746538728
transform 1 0 21888 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _498_
timestamp 1746538728
transform 1 0 20832 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _499_
timestamp 1746538728
transform 1 0 25632 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _500_
timestamp 1746538728
transform 1 0 21792 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _501_
timestamp 1746538728
transform -1 0 39552 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _502_
timestamp 1746538728
transform -1 0 44832 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _503_
timestamp 1746538728
transform 1 0 35424 0 -1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _504_
timestamp 1746538728
transform 1 0 40224 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _505_
timestamp 1746538728
transform 1 0 4704 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _506_
timestamp 1746538728
transform 1 0 6144 0 -1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _507_
timestamp 1746538728
transform 1 0 16032 0 1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _508_
timestamp 1746538728
transform 1 0 14304 0 1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _509_
timestamp 1746538728
transform 1 0 15264 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _510_
timestamp 1746538728
transform 1 0 12672 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _511_
timestamp 1746538728
transform 1 0 25632 0 1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _512_
timestamp 1746538728
transform 1 0 28032 0 -1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _513_
timestamp 1746538728
transform -1 0 34656 0 -1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _514_
timestamp 1746538728
transform -1 0 34848 0 1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _515_
timestamp 1746538728
transform 1 0 7296 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _516_
timestamp 1746538728
transform 1 0 9408 0 -1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _517_
timestamp 1746538728
transform 1 0 19680 0 1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _518_
timestamp 1746538728
transform 1 0 19776 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _519_
timestamp 1746538728
transform -1 0 23424 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _520_
timestamp 1746538728
transform -1 0 30336 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _521_
timestamp 1746538728
transform 1 0 9888 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _522_
timestamp 1746538728
transform 1 0 12192 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _523_
timestamp 1746538728
transform -1 0 19008 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _524_
timestamp 1746538728
transform -1 0 19872 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _525_
timestamp 1746538728
transform 1 0 11808 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _526_
timestamp 1746538728
transform 1 0 15936 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _527_
timestamp 1746538728
transform 1 0 15840 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _528_
timestamp 1746538728
transform 1 0 18912 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _529_
timestamp 1746538728
transform 1 0 22944 0 -1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _530_
timestamp 1746538728
transform 1 0 42528 0 1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _531_
timestamp 1746538728
transform 1 0 37056 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _532_
timestamp 1746538728
transform 1 0 32064 0 1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _533_
timestamp 1746538728
transform -1 0 30720 0 1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _534_
timestamp 1746538728
transform 1 0 27552 0 -1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _535_
timestamp 1746538728
transform 1 0 31008 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _536_
timestamp 1746538728
transform 1 0 25056 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _537_
timestamp 1746538728
transform 1 0 24864 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _538_
timestamp 1746538728
transform 1 0 52704 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _539_
timestamp 1746538728
transform 1 0 56256 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _540_
timestamp 1746538728
transform 1 0 46656 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _541_
timestamp 1746538728
transform 1 0 47808 0 -1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _542_
timestamp 1746538728
transform 1 0 33312 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _543_
timestamp 1746538728
transform 1 0 36672 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _544_
timestamp 1746538728
transform 1 0 52512 0 1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _545_
timestamp 1746538728
transform 1 0 54336 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _546_
timestamp 1746538728
transform 1 0 11424 0 -1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _547_
timestamp 1746538728
transform 1 0 7200 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _548_
timestamp 1746538728
transform 1 0 36768 0 1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _549_
timestamp 1746538728
transform -1 0 46080 0 -1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _550_
timestamp 1746538728
transform 1 0 30240 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _551_
timestamp 1746538728
transform 1 0 30816 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _552_
timestamp 1746538728
transform 1 0 31488 0 1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _553_
timestamp 1746538728
transform 1 0 23808 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _554_
timestamp 1746538728
transform 1 0 20928 0 1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _555_
timestamp 1746538728
transform 1 0 22656 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _556_
timestamp 1746538728
transform 1 0 56160 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _557_
timestamp 1746538728
transform 1 0 54816 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _558_
timestamp 1746538728
transform 1 0 46272 0 1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _559_
timestamp 1746538728
transform 1 0 48384 0 1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _560_
timestamp 1746538728
transform 1 0 39264 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _561_
timestamp 1746538728
transform 1 0 37632 0 1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _562_
timestamp 1746538728
transform 1 0 50400 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _563_
timestamp 1746538728
transform 1 0 54720 0 -1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _564_
timestamp 1746538728
transform 1 0 11136 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _565_
timestamp 1746538728
transform 1 0 7008 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _566_
timestamp 1746538728
transform 1 0 2592 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _567_
timestamp 1746538728
transform 1 0 2304 0 1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _568_
timestamp 1746538728
transform 1 0 10848 0 1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _569_
timestamp 1746538728
transform 1 0 4032 0 1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _570_
timestamp 1746538728
transform 1 0 6240 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _571_
timestamp 1746538728
transform 1 0 10848 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _572_
timestamp 1746538728
transform 1 0 3840 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _573_
timestamp 1746538728
transform 1 0 1824 0 -1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _574_
timestamp 1746538728
transform 1 0 17472 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _575_
timestamp 1746538728
transform 1 0 15744 0 1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _576_
timestamp 1746538728
transform 1 0 25056 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _577_
timestamp 1746538728
transform 1 0 16704 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _578_
timestamp 1746538728
transform 1 0 47040 0 1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _579_
timestamp 1746538728
transform 1 0 46944 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _580_
timestamp 1746538728
transform 1 0 37056 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _581_
timestamp 1746538728
transform 1 0 33120 0 1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _582_
timestamp 1746538728
transform 1 0 2592 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _583_
timestamp 1746538728
transform 1 0 2016 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _584_
timestamp 1746538728
transform 1 0 2592 0 -1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _585_
timestamp 1746538728
transform 1 0 1632 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _586_
timestamp 1746538728
transform 1 0 10656 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _587_
timestamp 1746538728
transform 1 0 5568 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _588_
timestamp 1746538728
transform 1 0 10848 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _589_
timestamp 1746538728
transform 1 0 5664 0 1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _590_
timestamp 1746538728
transform 1 0 2496 0 1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _591_
timestamp 1746538728
transform 1 0 2208 0 1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _592_
timestamp 1746538728
transform 1 0 17376 0 1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _593_
timestamp 1746538728
transform 1 0 14400 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_2  _594_
timestamp 1746538784
transform 1 0 23520 0 1 24948
box -48 -56 2736 834
use sg13g2_dfrbpq_1  _595_
timestamp 1746538728
transform 1 0 27744 0 1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _596_
timestamp 1746538728
transform 1 0 43680 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _597_
timestamp 1746538728
transform 1 0 49056 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _598_
timestamp 1746538728
transform 1 0 33120 0 -1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _599_
timestamp 1746538728
transform 1 0 39648 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _600_
timestamp 1746538728
transform 1 0 2496 0 -1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _601_
timestamp 1746538728
transform 1 0 1920 0 1 8316
box -48 -56 2640 834
use sg13g2_buf_8  clkbuf_0_clk
timestamp 1676454965
transform 1 0 30336 0 -1 20412
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_0_0_clk
timestamp 1676454965
transform -1 0 8256 0 1 12852
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_1_0_clk
timestamp 1676454965
transform -1 0 9984 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_2_0_clk
timestamp 1676454965
transform -1 0 19968 0 -1 9828
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_3_0_clk
timestamp 1676454965
transform 1 0 18720 0 1 11340
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_4_0_clk
timestamp 1676454965
transform -1 0 9984 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_5_0_clk
timestamp 1676454965
transform -1 0 10752 0 -1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_6_0_clk
timestamp 1676454965
transform -1 0 23328 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_7_0_clk
timestamp 1676454965
transform -1 0 23616 0 1 30996
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_8_0_clk
timestamp 1676454965
transform -1 0 37440 0 -1 8316
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_9_0_clk
timestamp 1676454965
transform -1 0 37248 0 -1 11340
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_10_0_clk
timestamp 1676454965
transform 1 0 50688 0 -1 8316
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_11_0_clk
timestamp 1676454965
transform 1 0 51456 0 1 9828
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_12_0_clk
timestamp 1676454965
transform -1 0 33888 0 -1 23436
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_13_0_clk
timestamp 1676454965
transform -1 0 35232 0 1 24948
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_14_0_clk
timestamp 1676454965
transform -1 0 46848 0 -1 26460
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_15_0_clk
timestamp 1676454965
transform -1 0 43680 0 -1 27972
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_0__f_clk
timestamp 1676454965
transform -1 0 4512 0 1 9828
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_1__f_clk
timestamp 1676454965
transform 1 0 8448 0 -1 8316
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_2__f_clk
timestamp 1676454965
transform -1 0 8160 0 -1 18900
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_3__f_clk
timestamp 1676454965
transform 1 0 12480 0 1 15876
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_4__f_clk
timestamp 1676454965
transform -1 0 18336 0 1 5292
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_5__f_clk
timestamp 1676454965
transform 1 0 21408 0 -1 6804
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_6__f_clk
timestamp 1676454965
transform -1 0 19680 0 1 8316
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_7__f_clk
timestamp 1676454965
transform 1 0 19008 0 -1 17388
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_8__f_clk
timestamp 1676454965
transform -1 0 6336 0 1 27972
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_9__f_clk
timestamp 1676454965
transform 1 0 11136 0 -1 26460
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_10__f_clk
timestamp 1676454965
transform -1 0 7392 0 -1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_11__f_clk
timestamp 1676454965
transform 1 0 12000 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_12__f_clk
timestamp 1676454965
transform -1 0 20736 0 1 26460
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_13__f_clk
timestamp 1676454965
transform 1 0 24960 0 1 27972
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_14__f_clk
timestamp 1676454965
transform -1 0 21696 0 -1 35532
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_15__f_clk
timestamp 1676454965
transform 1 0 25152 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_16__f_clk
timestamp 1676454965
transform -1 0 34080 0 1 5292
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_17__f_clk
timestamp 1676454965
transform 1 0 39168 0 -1 6804
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_18__f_clk
timestamp 1676454965
transform -1 0 33696 0 -1 12852
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_19__f_clk
timestamp 1676454965
transform 1 0 38784 0 -1 14364
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_20__f_clk
timestamp 1676454965
transform -1 0 48864 0 1 5292
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_21__f_clk
timestamp 1676454965
transform 1 0 53856 0 -1 6804
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_22__f_clk
timestamp 1676454965
transform -1 0 50496 0 1 12852
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_23__f_clk
timestamp 1676454965
transform 1 0 54432 0 1 12852
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_24__f_clk
timestamp 1676454965
transform -1 0 30336 0 -1 20412
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_25__f_clk
timestamp 1676454965
transform 1 0 34752 0 1 18900
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_26__f_clk
timestamp 1676454965
transform -1 0 34176 0 -1 24948
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_27__f_clk
timestamp 1676454965
transform 1 0 34368 0 -1 30996
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_28__f_clk
timestamp 1676454965
transform -1 0 43488 0 -1 24948
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_29__f_clk
timestamp 1676454965
transform 1 0 47136 0 1 21924
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_30__f_clk
timestamp 1676454965
transform -1 0 42624 0 1 30996
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_31__f_clk
timestamp 1676454965
transform 1 0 46080 0 1 29484
box -48 -56 1296 834
use sg13g2_inv_1  clkload0
timestamp 1676386529
transform 1 0 18912 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  clkload1
timestamp 1676386529
transform -1 0 12000 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  clkload2
timestamp 1676385511
transform 1 0 19392 0 1 24948
box -48 -56 432 834
use sg13g2_inv_1  clkload3
timestamp 1676386529
transform -1 0 25440 0 -1 34020
box -48 -56 336 834
use sg13g2_buf_1  clkload4
timestamp 1676385511
transform 1 0 39168 0 -1 5292
box -48 -56 432 834
use sg13g2_inv_1  clkload5
timestamp 1676386529
transform -1 0 54720 0 -1 14364
box -48 -56 336 834
use sg13g2_inv_1  clkload6
timestamp 1676386529
transform 1 0 34080 0 -1 30996
box -48 -56 336 834
use sg13g2_inv_1  clkload7
timestamp 1676386529
transform 1 0 46080 0 -1 30996
box -48 -56 336 834
use sg13g2_buf_8  fanout60
timestamp 1676454965
transform 1 0 14976 0 1 5292
box -48 -56 1296 834
use sg13g2_buf_8  fanout61
timestamp 1676454965
transform -1 0 12096 0 1 6804
box -48 -56 1296 834
use sg13g2_buf_8  fanout62
timestamp 1676454965
transform -1 0 11904 0 1 12852
box -48 -56 1296 834
use sg13g2_buf_8  fanout63
timestamp 1676454965
transform -1 0 14304 0 -1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout64
timestamp 1676454965
transform -1 0 23808 0 1 12852
box -48 -56 1296 834
use sg13g2_buf_8  fanout65
timestamp 1676454965
transform 1 0 21408 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout66
timestamp 1676454965
transform 1 0 22656 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout67
timestamp 1676454965
transform 1 0 9696 0 1 20412
box -48 -56 1296 834
use sg13g2_buf_8  fanout68
timestamp 1676454965
transform -1 0 10368 0 1 26460
box -48 -56 1296 834
use sg13g2_buf_8  fanout69
timestamp 1676454965
transform -1 0 14880 0 1 20412
box -48 -56 1296 834
use sg13g2_buf_8  fanout70
timestamp 1676454965
transform 1 0 15648 0 1 29484
box -48 -56 1296 834
use sg13g2_buf_8  fanout71
timestamp 1676454965
transform -1 0 23520 0 1 21924
box -48 -56 1296 834
use sg13g2_buf_8  fanout72
timestamp 1676454965
transform -1 0 26016 0 -1 23436
box -48 -56 1296 834
use sg13g2_buf_8  fanout73
timestamp 1676454965
transform 1 0 37632 0 -1 8316
box -48 -56 1296 834
use sg13g2_buf_8  fanout74
timestamp 1676454965
transform -1 0 42912 0 -1 15876
box -48 -56 1296 834
use sg13g2_buf_8  fanout75
timestamp 1676454965
transform -1 0 52512 0 -1 9828
box -48 -56 1296 834
use sg13g2_buf_2  fanout76
timestamp 1676385467
transform -1 0 53280 0 -1 9828
box -48 -56 528 834
use sg13g2_buf_8  fanout77
timestamp 1676454965
transform 1 0 46464 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout78
timestamp 1676454965
transform 1 0 44928 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout79
timestamp 1676454965
transform 1 0 29568 0 -1 26460
box -48 -56 1296 834
use sg13g2_buf_8  fanout80
timestamp 1676454965
transform -1 0 30336 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  fanout81
timestamp 1676454965
transform -1 0 42912 0 1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout82
timestamp 1676454965
transform -1 0 42240 0 -1 30996
box -48 -56 1296 834
use sg13g2_buf_8  fanout83
timestamp 1676454965
transform 1 0 42624 0 1 29484
box -48 -56 1296 834
use sg13g2_buf_8  fanout84
timestamp 1676454965
transform -1 0 44736 0 1 26460
box -48 -56 1296 834
use sg13g2_buf_8  fanout85
timestamp 1676454965
transform 1 0 26016 0 -1 23436
box -48 -56 1296 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679585382
transform 1 0 576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679585382
transform 1 0 1248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679585382
transform 1 0 1920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679585382
transform 1 0 2592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679585382
transform 1 0 3264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679585382
transform 1 0 3936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679585382
transform 1 0 4608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679585382
transform 1 0 5280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679585382
transform 1 0 5952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679585382
transform 1 0 6624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679585382
transform 1 0 7296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679585382
transform 1 0 7968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679585382
transform 1 0 8640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679585382
transform 1 0 9312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679585382
transform 1 0 9984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679585382
transform 1 0 10656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679585382
transform 1 0 11328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679585382
transform 1 0 12000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679585382
transform 1 0 12672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679585382
transform 1 0 13344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679585382
transform 1 0 14016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679585382
transform 1 0 14688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679585382
transform 1 0 15360 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679585382
transform 1 0 16032 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679585382
transform 1 0 16704 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679585382
transform 1 0 17376 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679585382
transform 1 0 18048 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679585382
transform 1 0 18720 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1679585382
transform 1 0 19392 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1679585382
transform 1 0 20064 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1679585382
transform 1 0 20736 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1679585382
transform 1 0 21408 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_224
timestamp 1679585382
transform 1 0 22080 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_231
timestamp 1679585382
transform 1 0 22752 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_238
timestamp 1679585382
transform 1 0 23424 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_245
timestamp 1679585382
transform 1 0 24096 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_252
timestamp 1679585382
transform 1 0 24768 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_259
timestamp 1679585382
transform 1 0 25440 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_266
timestamp 1679585382
transform 1 0 26112 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_273
timestamp 1679585382
transform 1 0 26784 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_280
timestamp 1679585382
transform 1 0 27456 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_287
timestamp 1679585382
transform 1 0 28128 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_294
timestamp 1679585382
transform 1 0 28800 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_301
timestamp 1679585382
transform 1 0 29472 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_308
timestamp 1679585382
transform 1 0 30144 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_315
timestamp 1679585382
transform 1 0 30816 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_322
timestamp 1679585382
transform 1 0 31488 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_329
timestamp 1679585382
transform 1 0 32160 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_336
timestamp 1679585382
transform 1 0 32832 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_343
timestamp 1679585382
transform 1 0 33504 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_350
timestamp 1679585382
transform 1 0 34176 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_357
timestamp 1679585382
transform 1 0 34848 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_364
timestamp 1679585382
transform 1 0 35520 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_371
timestamp 1679585382
transform 1 0 36192 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_378
timestamp 1679585382
transform 1 0 36864 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_385
timestamp 1679585382
transform 1 0 37536 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_392
timestamp 1679585382
transform 1 0 38208 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_399
timestamp 1679585382
transform 1 0 38880 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_406
timestamp 1679585382
transform 1 0 39552 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_413
timestamp 1679585382
transform 1 0 40224 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_420
timestamp 1679585382
transform 1 0 40896 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_427
timestamp 1679585382
transform 1 0 41568 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_434
timestamp 1679585382
transform 1 0 42240 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_441
timestamp 1679585382
transform 1 0 42912 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_448
timestamp 1679585382
transform 1 0 43584 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_455
timestamp 1679585382
transform 1 0 44256 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_462
timestamp 1679585382
transform 1 0 44928 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_469
timestamp 1679585382
transform 1 0 45600 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_476
timestamp 1679585382
transform 1 0 46272 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_483
timestamp 1679585382
transform 1 0 46944 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_490
timestamp 1679585382
transform 1 0 47616 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_497
timestamp 1679585382
transform 1 0 48288 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_504
timestamp 1679585382
transform 1 0 48960 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_511
timestamp 1679585382
transform 1 0 49632 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_518
timestamp 1679585382
transform 1 0 50304 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_525
timestamp 1679585382
transform 1 0 50976 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_532
timestamp 1679585382
transform 1 0 51648 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_539
timestamp 1679585382
transform 1 0 52320 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_546
timestamp 1679585382
transform 1 0 52992 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_553
timestamp 1679585382
transform 1 0 53664 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_560
timestamp 1679585382
transform 1 0 54336 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_567
timestamp 1679585382
transform 1 0 55008 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_574
timestamp 1679585382
transform 1 0 55680 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_581
timestamp 1679585382
transform 1 0 56352 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_588
timestamp 1679585382
transform 1 0 57024 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_595
timestamp 1679585382
transform 1 0 57696 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_602
timestamp 1679585382
transform 1 0 58368 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_609
timestamp 1679585382
transform 1 0 59040 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_616
timestamp 1679585382
transform 1 0 59712 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_623
timestamp 1679585382
transform 1 0 60384 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_630
timestamp 1679585382
transform 1 0 61056 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_637
timestamp 1679585382
transform 1 0 61728 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_644
timestamp 1679585382
transform 1 0 62400 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_651
timestamp 1679585382
transform 1 0 63072 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_658
timestamp 1679585382
transform 1 0 63744 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_665
timestamp 1679585382
transform 1 0 64416 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_672
timestamp 1679585382
transform 1 0 65088 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_679
timestamp 1679585382
transform 1 0 65760 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_686
timestamp 1679585382
transform 1 0 66432 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_693
timestamp 1679585382
transform 1 0 67104 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_700
timestamp 1679585382
transform 1 0 67776 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_707
timestamp 1679585382
transform 1 0 68448 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_714
timestamp 1679585382
transform 1 0 69120 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_721
timestamp 1679585382
transform 1 0 69792 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_728
timestamp 1679585382
transform 1 0 70464 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_735
timestamp 1679585382
transform 1 0 71136 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_742
timestamp 1679585382
transform 1 0 71808 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_749
timestamp 1679585382
transform 1 0 72480 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_756
timestamp 1679585382
transform 1 0 73152 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_763
timestamp 1679585382
transform 1 0 73824 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_770
timestamp 1679585382
transform 1 0 74496 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_777
timestamp 1679585382
transform 1 0 75168 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_784
timestamp 1679585382
transform 1 0 75840 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_791
timestamp 1679585382
transform 1 0 76512 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_798
timestamp 1679585382
transform 1 0 77184 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_805
timestamp 1679585382
transform 1 0 77856 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_812
timestamp 1679585382
transform 1 0 78528 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_819
timestamp 1679585382
transform 1 0 79200 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_826
timestamp 1679585382
transform 1 0 79872 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_833
timestamp 1679585382
transform 1 0 80544 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_840
timestamp 1679585382
transform 1 0 81216 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_847
timestamp 1679585382
transform 1 0 81888 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_854
timestamp 1679585382
transform 1 0 82560 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_861
timestamp 1679585382
transform 1 0 83232 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_868
timestamp 1679585382
transform 1 0 83904 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_875
timestamp 1679585382
transform 1 0 84576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_882
timestamp 1679585382
transform 1 0 85248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_889
timestamp 1679585382
transform 1 0 85920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_896
timestamp 1679585382
transform 1 0 86592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_903
timestamp 1679585382
transform 1 0 87264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_910
timestamp 1679585382
transform 1 0 87936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_917
timestamp 1679585382
transform 1 0 88608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_924
timestamp 1679585382
transform 1 0 89280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_931
timestamp 1679585382
transform 1 0 89952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_938
timestamp 1679585382
transform 1 0 90624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_945
timestamp 1679585382
transform 1 0 91296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_952
timestamp 1679585382
transform 1 0 91968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_959
timestamp 1679585382
transform 1 0 92640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_966
timestamp 1679585382
transform 1 0 93312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_973
timestamp 1679585382
transform 1 0 93984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_980
timestamp 1679585382
transform 1 0 94656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_987
timestamp 1679585382
transform 1 0 95328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_994
timestamp 1679585382
transform 1 0 96000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1001
timestamp 1679585382
transform 1 0 96672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1008
timestamp 1679585382
transform 1 0 97344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1015
timestamp 1679585382
transform 1 0 98016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1022
timestamp 1679585382
transform 1 0 98688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679585382
transform 1 0 576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679585382
transform 1 0 1248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679585382
transform 1 0 1920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679585382
transform 1 0 2592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679585382
transform 1 0 3264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679585382
transform 1 0 3936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679585382
transform 1 0 4608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679585382
transform 1 0 5280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679585382
transform 1 0 5952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679585382
transform 1 0 6624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_70
timestamp 1679581501
transform 1 0 7296 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_74
timestamp 1677583258
transform 1 0 7680 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_83
timestamp 1677583704
transform 1 0 8544 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_85
timestamp 1677583258
transform 1 0 8736 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_95
timestamp 1679585382
transform 1 0 9696 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_102
timestamp 1679585382
transform 1 0 10368 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_109
timestamp 1679585382
transform 1 0 11040 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_116
timestamp 1679585382
transform 1 0 11712 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_123
timestamp 1679585382
transform 1 0 12384 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_130
timestamp 1679585382
transform 1 0 13056 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_137
timestamp 1679585382
transform 1 0 13728 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_144
timestamp 1679585382
transform 1 0 14400 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_151
timestamp 1679585382
transform 1 0 15072 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_158
timestamp 1679585382
transform 1 0 15744 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_165
timestamp 1679581501
transform 1 0 16416 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_169
timestamp 1677583704
transform 1 0 16800 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_180
timestamp 1679585382
transform 1 0 17856 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_187
timestamp 1679585382
transform 1 0 18528 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_194
timestamp 1679585382
transform 1 0 19200 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_201
timestamp 1679585382
transform 1 0 19872 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_208
timestamp 1679585382
transform 1 0 20544 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_215
timestamp 1679585382
transform 1 0 21216 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_222
timestamp 1679585382
transform 1 0 21888 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_229
timestamp 1679585382
transform 1 0 22560 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_236
timestamp 1679585382
transform 1 0 23232 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_243
timestamp 1679585382
transform 1 0 23904 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_250
timestamp 1679585382
transform 1 0 24576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_257
timestamp 1679585382
transform 1 0 25248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_264
timestamp 1679585382
transform 1 0 25920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_271
timestamp 1679585382
transform 1 0 26592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_278
timestamp 1679585382
transform 1 0 27264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_285
timestamp 1679585382
transform 1 0 27936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_292
timestamp 1679585382
transform 1 0 28608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_299
timestamp 1679585382
transform 1 0 29280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_306
timestamp 1679585382
transform 1 0 29952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_313
timestamp 1679585382
transform 1 0 30624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_320
timestamp 1679585382
transform 1 0 31296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_327
timestamp 1679585382
transform 1 0 31968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_334
timestamp 1679585382
transform 1 0 32640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_341
timestamp 1679585382
transform 1 0 33312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_348
timestamp 1679585382
transform 1 0 33984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_355
timestamp 1679585382
transform 1 0 34656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_362
timestamp 1679585382
transform 1 0 35328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_369
timestamp 1679585382
transform 1 0 36000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_376
timestamp 1679585382
transform 1 0 36672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_383
timestamp 1679585382
transform 1 0 37344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_390
timestamp 1679585382
transform 1 0 38016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_397
timestamp 1679585382
transform 1 0 38688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_404
timestamp 1679585382
transform 1 0 39360 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_411
timestamp 1679585382
transform 1 0 40032 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_418
timestamp 1679585382
transform 1 0 40704 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_425
timestamp 1679585382
transform 1 0 41376 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_432
timestamp 1679585382
transform 1 0 42048 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_439
timestamp 1679585382
transform 1 0 42720 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_446
timestamp 1679585382
transform 1 0 43392 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_453
timestamp 1679585382
transform 1 0 44064 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_460
timestamp 1679585382
transform 1 0 44736 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_467
timestamp 1679585382
transform 1 0 45408 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_474
timestamp 1679585382
transform 1 0 46080 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_481
timestamp 1679585382
transform 1 0 46752 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_488
timestamp 1679585382
transform 1 0 47424 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_495
timestamp 1679585382
transform 1 0 48096 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_502
timestamp 1679585382
transform 1 0 48768 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_509
timestamp 1679585382
transform 1 0 49440 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_516
timestamp 1679585382
transform 1 0 50112 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_523
timestamp 1679585382
transform 1 0 50784 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_530
timestamp 1679585382
transform 1 0 51456 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_537
timestamp 1679585382
transform 1 0 52128 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_544
timestamp 1679585382
transform 1 0 52800 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_551
timestamp 1679585382
transform 1 0 53472 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_558
timestamp 1679585382
transform 1 0 54144 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_565
timestamp 1679585382
transform 1 0 54816 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_572
timestamp 1679585382
transform 1 0 55488 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_579
timestamp 1679585382
transform 1 0 56160 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_586
timestamp 1679585382
transform 1 0 56832 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_593
timestamp 1679585382
transform 1 0 57504 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_600
timestamp 1679585382
transform 1 0 58176 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_607
timestamp 1679585382
transform 1 0 58848 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_614
timestamp 1679585382
transform 1 0 59520 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_621
timestamp 1679585382
transform 1 0 60192 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_628
timestamp 1679585382
transform 1 0 60864 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_635
timestamp 1679585382
transform 1 0 61536 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_642
timestamp 1679585382
transform 1 0 62208 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_649
timestamp 1679585382
transform 1 0 62880 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_656
timestamp 1679585382
transform 1 0 63552 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_663
timestamp 1679585382
transform 1 0 64224 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_670
timestamp 1679585382
transform 1 0 64896 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_677
timestamp 1679585382
transform 1 0 65568 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_684
timestamp 1679585382
transform 1 0 66240 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_691
timestamp 1679585382
transform 1 0 66912 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_698
timestamp 1679585382
transform 1 0 67584 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_705
timestamp 1679585382
transform 1 0 68256 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_712
timestamp 1679585382
transform 1 0 68928 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_719
timestamp 1679585382
transform 1 0 69600 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_726
timestamp 1679585382
transform 1 0 70272 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_733
timestamp 1679585382
transform 1 0 70944 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_740
timestamp 1679585382
transform 1 0 71616 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_747
timestamp 1679585382
transform 1 0 72288 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_754
timestamp 1679585382
transform 1 0 72960 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_761
timestamp 1679585382
transform 1 0 73632 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_768
timestamp 1679585382
transform 1 0 74304 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_775
timestamp 1679585382
transform 1 0 74976 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_782
timestamp 1679585382
transform 1 0 75648 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_789
timestamp 1679585382
transform 1 0 76320 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_796
timestamp 1679585382
transform 1 0 76992 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_803
timestamp 1679585382
transform 1 0 77664 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_810
timestamp 1679585382
transform 1 0 78336 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_817
timestamp 1679585382
transform 1 0 79008 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_824
timestamp 1679585382
transform 1 0 79680 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_831
timestamp 1679585382
transform 1 0 80352 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_838
timestamp 1679585382
transform 1 0 81024 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_845
timestamp 1679585382
transform 1 0 81696 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_852
timestamp 1679585382
transform 1 0 82368 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_859
timestamp 1679585382
transform 1 0 83040 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_866
timestamp 1679585382
transform 1 0 83712 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_873
timestamp 1679585382
transform 1 0 84384 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_880
timestamp 1679585382
transform 1 0 85056 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_887
timestamp 1679585382
transform 1 0 85728 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_894
timestamp 1679585382
transform 1 0 86400 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_901
timestamp 1679585382
transform 1 0 87072 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_908
timestamp 1679585382
transform 1 0 87744 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_915
timestamp 1679585382
transform 1 0 88416 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_922
timestamp 1679585382
transform 1 0 89088 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_929
timestamp 1679585382
transform 1 0 89760 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_936
timestamp 1679585382
transform 1 0 90432 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_943
timestamp 1679585382
transform 1 0 91104 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_950
timestamp 1679585382
transform 1 0 91776 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_957
timestamp 1679585382
transform 1 0 92448 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_964
timestamp 1679585382
transform 1 0 93120 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_971
timestamp 1679585382
transform 1 0 93792 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_978
timestamp 1679585382
transform 1 0 94464 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_985
timestamp 1679585382
transform 1 0 95136 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_992
timestamp 1679585382
transform 1 0 95808 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_999
timestamp 1679585382
transform 1 0 96480 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1006
timestamp 1679585382
transform 1 0 97152 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1013
timestamp 1679585382
transform 1 0 97824 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1020
timestamp 1679585382
transform 1 0 98496 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_1027
timestamp 1677583704
transform 1 0 99168 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_4
timestamp 1679585382
transform 1 0 960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_11
timestamp 1679585382
transform 1 0 1632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_18
timestamp 1679585382
transform 1 0 2304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_25
timestamp 1679585382
transform 1 0 2976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_32
timestamp 1679585382
transform 1 0 3648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_39
timestamp 1679585382
transform 1 0 4320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_46
timestamp 1679585382
transform 1 0 4992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_53
timestamp 1679585382
transform 1 0 5664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_60
timestamp 1679585382
transform 1 0 6336 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_67
timestamp 1677583704
transform 1 0 7008 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_105
timestamp 1679585382
transform 1 0 10656 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_112
timestamp 1677583704
transform 1 0 11328 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_114
timestamp 1677583258
transform 1 0 11520 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_123
timestamp 1679585382
transform 1 0 12384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_130
timestamp 1679585382
transform 1 0 13056 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_137
timestamp 1677583704
transform 1 0 13728 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_139
timestamp 1677583258
transform 1 0 13920 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_167
timestamp 1679585382
transform 1 0 16608 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_174
timestamp 1677583258
transform 1 0 17280 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_202
timestamp 1679585382
transform 1 0 19968 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_209
timestamp 1679585382
transform 1 0 20640 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_216
timestamp 1679585382
transform 1 0 21312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_223
timestamp 1679585382
transform 1 0 21984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_230
timestamp 1679585382
transform 1 0 22656 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_237
timestamp 1679585382
transform 1 0 23328 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_244
timestamp 1679585382
transform 1 0 24000 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_251
timestamp 1679585382
transform 1 0 24672 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_258
timestamp 1679585382
transform 1 0 25344 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_265
timestamp 1679585382
transform 1 0 26016 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_272
timestamp 1679585382
transform 1 0 26688 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_279
timestamp 1679585382
transform 1 0 27360 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_286
timestamp 1679585382
transform 1 0 28032 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_293
timestamp 1679585382
transform 1 0 28704 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_300
timestamp 1679585382
transform 1 0 29376 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_307
timestamp 1679585382
transform 1 0 30048 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_314
timestamp 1679585382
transform 1 0 30720 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_321
timestamp 1679585382
transform 1 0 31392 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_328
timestamp 1679585382
transform 1 0 32064 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_335
timestamp 1679585382
transform 1 0 32736 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_342
timestamp 1679585382
transform 1 0 33408 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_349
timestamp 1679585382
transform 1 0 34080 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_356
timestamp 1679585382
transform 1 0 34752 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_363
timestamp 1679585382
transform 1 0 35424 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_370
timestamp 1679581501
transform 1 0 36096 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_374
timestamp 1677583704
transform 1 0 36480 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_430
timestamp 1679585382
transform 1 0 41856 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_437
timestamp 1679585382
transform 1 0 42528 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_444
timestamp 1679585382
transform 1 0 43200 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_451
timestamp 1677583258
transform 1 0 43872 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_479
timestamp 1679581501
transform 1 0 46560 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_483
timestamp 1677583258
transform 1 0 46944 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_511
timestamp 1679585382
transform 1 0 49632 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_518
timestamp 1677583258
transform 1 0 50304 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_546
timestamp 1679585382
transform 1 0 52992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_553
timestamp 1679585382
transform 1 0 53664 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_560
timestamp 1677583258
transform 1 0 54336 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_565
timestamp 1679585382
transform 1 0 54816 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_572
timestamp 1679585382
transform 1 0 55488 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_579
timestamp 1679585382
transform 1 0 56160 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_586
timestamp 1679585382
transform 1 0 56832 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_593
timestamp 1679585382
transform 1 0 57504 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_600
timestamp 1679585382
transform 1 0 58176 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_607
timestamp 1679585382
transform 1 0 58848 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_614
timestamp 1679585382
transform 1 0 59520 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_621
timestamp 1679585382
transform 1 0 60192 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_628
timestamp 1679585382
transform 1 0 60864 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_635
timestamp 1679585382
transform 1 0 61536 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_642
timestamp 1679585382
transform 1 0 62208 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_649
timestamp 1679585382
transform 1 0 62880 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_656
timestamp 1679585382
transform 1 0 63552 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_663
timestamp 1679585382
transform 1 0 64224 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_670
timestamp 1679585382
transform 1 0 64896 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_677
timestamp 1679585382
transform 1 0 65568 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_684
timestamp 1679585382
transform 1 0 66240 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_691
timestamp 1679585382
transform 1 0 66912 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_698
timestamp 1679585382
transform 1 0 67584 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_705
timestamp 1679585382
transform 1 0 68256 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_712
timestamp 1679585382
transform 1 0 68928 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_719
timestamp 1679585382
transform 1 0 69600 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_726
timestamp 1679585382
transform 1 0 70272 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_733
timestamp 1679585382
transform 1 0 70944 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_740
timestamp 1679585382
transform 1 0 71616 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_747
timestamp 1679585382
transform 1 0 72288 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_754
timestamp 1679585382
transform 1 0 72960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_761
timestamp 1679585382
transform 1 0 73632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_768
timestamp 1679585382
transform 1 0 74304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_775
timestamp 1679585382
transform 1 0 74976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_782
timestamp 1679585382
transform 1 0 75648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_789
timestamp 1679585382
transform 1 0 76320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_796
timestamp 1679585382
transform 1 0 76992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_803
timestamp 1679585382
transform 1 0 77664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_810
timestamp 1679585382
transform 1 0 78336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_817
timestamp 1679585382
transform 1 0 79008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_824
timestamp 1679585382
transform 1 0 79680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_831
timestamp 1679585382
transform 1 0 80352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_838
timestamp 1679585382
transform 1 0 81024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_845
timestamp 1679585382
transform 1 0 81696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_852
timestamp 1679585382
transform 1 0 82368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_859
timestamp 1679585382
transform 1 0 83040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_866
timestamp 1679585382
transform 1 0 83712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_873
timestamp 1679585382
transform 1 0 84384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_880
timestamp 1679585382
transform 1 0 85056 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_887
timestamp 1679585382
transform 1 0 85728 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_894
timestamp 1679585382
transform 1 0 86400 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_901
timestamp 1679585382
transform 1 0 87072 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_908
timestamp 1679585382
transform 1 0 87744 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_915
timestamp 1679585382
transform 1 0 88416 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_922
timestamp 1679585382
transform 1 0 89088 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_929
timestamp 1679585382
transform 1 0 89760 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_936
timestamp 1679585382
transform 1 0 90432 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_943
timestamp 1679585382
transform 1 0 91104 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_950
timestamp 1679585382
transform 1 0 91776 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_957
timestamp 1679585382
transform 1 0 92448 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_964
timestamp 1679585382
transform 1 0 93120 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_971
timestamp 1679585382
transform 1 0 93792 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_978
timestamp 1679585382
transform 1 0 94464 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_985
timestamp 1679585382
transform 1 0 95136 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_992
timestamp 1679585382
transform 1 0 95808 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_999
timestamp 1679585382
transform 1 0 96480 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1006
timestamp 1679585382
transform 1 0 97152 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1013
timestamp 1679585382
transform 1 0 97824 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1020
timestamp 1679585382
transform 1 0 98496 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_1027
timestamp 1677583704
transform 1 0 99168 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_4
timestamp 1679585382
transform 1 0 960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_11
timestamp 1679585382
transform 1 0 1632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_18
timestamp 1679585382
transform 1 0 2304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_25
timestamp 1679585382
transform 1 0 2976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_32
timestamp 1679585382
transform 1 0 3648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_39
timestamp 1679585382
transform 1 0 4320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_46
timestamp 1679585382
transform 1 0 4992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_53
timestamp 1679585382
transform 1 0 5664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_60
timestamp 1679585382
transform 1 0 6336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_94
timestamp 1679585382
transform 1 0 9600 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_101
timestamp 1679581501
transform 1 0 10272 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_105
timestamp 1677583704
transform 1 0 10656 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_115
timestamp 1677583258
transform 1 0 11616 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_120
timestamp 1679581501
transform 1 0 12096 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_138
timestamp 1679585382
transform 1 0 13824 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_145
timestamp 1679585382
transform 1 0 14496 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_152
timestamp 1679585382
transform 1 0 15168 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_159
timestamp 1679585382
transform 1 0 15840 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_166
timestamp 1679585382
transform 1 0 16512 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_173
timestamp 1679581501
transform 1 0 17184 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_204
timestamp 1679585382
transform 1 0 20160 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_211
timestamp 1677583704
transform 1 0 20832 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_222
timestamp 1677583704
transform 1 0 21888 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_278
timestamp 1679585382
transform 1 0 27264 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_285
timestamp 1679585382
transform 1 0 27936 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_292
timestamp 1679585382
transform 1 0 28608 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_299
timestamp 1679585382
transform 1 0 29280 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_306
timestamp 1679585382
transform 1 0 29952 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_313
timestamp 1679585382
transform 1 0 30624 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_320
timestamp 1679585382
transform 1 0 31296 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_327
timestamp 1679585382
transform 1 0 31968 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_334
timestamp 1679585382
transform 1 0 32640 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_368
timestamp 1679585382
transform 1 0 35904 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_375
timestamp 1679585382
transform 1 0 36576 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_382
timestamp 1679585382
transform 1 0 37248 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_389
timestamp 1677583704
transform 1 0 37920 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_395
timestamp 1677583704
transform 1 0 38496 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_397
timestamp 1677583258
transform 1 0 38688 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_407
timestamp 1677583258
transform 1 0 39648 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_416
timestamp 1679581501
transform 1 0 40512 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_429
timestamp 1679585382
transform 1 0 41760 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_436
timestamp 1679585382
transform 1 0 42432 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_443
timestamp 1679585382
transform 1 0 43104 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_450
timestamp 1679585382
transform 1 0 43776 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_457
timestamp 1679585382
transform 1 0 44448 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_464
timestamp 1679585382
transform 1 0 45120 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_471
timestamp 1679585382
transform 1 0 45792 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_478
timestamp 1679585382
transform 1 0 46464 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_485
timestamp 1677583704
transform 1 0 47136 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_487
timestamp 1677583258
transform 1 0 47328 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_496
timestamp 1679585382
transform 1 0 48192 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_503
timestamp 1679585382
transform 1 0 48864 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_510
timestamp 1679585382
transform 1 0 49536 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_517
timestamp 1679585382
transform 1 0 50208 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_524
timestamp 1677583704
transform 1 0 50880 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_526
timestamp 1677583258
transform 1 0 51072 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_531
timestamp 1677583704
transform 1 0 51552 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_533
timestamp 1677583258
transform 1 0 51744 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_555
timestamp 1679581501
transform 1 0 53856 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_559
timestamp 1677583258
transform 1 0 54240 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_587
timestamp 1679585382
transform 1 0 56928 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_594
timestamp 1679585382
transform 1 0 57600 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_601
timestamp 1679585382
transform 1 0 58272 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_608
timestamp 1679585382
transform 1 0 58944 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_615
timestamp 1679585382
transform 1 0 59616 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_622
timestamp 1679585382
transform 1 0 60288 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_629
timestamp 1679585382
transform 1 0 60960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_636
timestamp 1679585382
transform 1 0 61632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_643
timestamp 1679585382
transform 1 0 62304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_650
timestamp 1679585382
transform 1 0 62976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_657
timestamp 1679585382
transform 1 0 63648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_664
timestamp 1679585382
transform 1 0 64320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_671
timestamp 1679585382
transform 1 0 64992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_678
timestamp 1679585382
transform 1 0 65664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_685
timestamp 1679585382
transform 1 0 66336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_692
timestamp 1679585382
transform 1 0 67008 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_699
timestamp 1679585382
transform 1 0 67680 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_706
timestamp 1679585382
transform 1 0 68352 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_713
timestamp 1679585382
transform 1 0 69024 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_720
timestamp 1679585382
transform 1 0 69696 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_727
timestamp 1679585382
transform 1 0 70368 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_734
timestamp 1679585382
transform 1 0 71040 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_741
timestamp 1679585382
transform 1 0 71712 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_748
timestamp 1679585382
transform 1 0 72384 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_755
timestamp 1679585382
transform 1 0 73056 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_762
timestamp 1679585382
transform 1 0 73728 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_769
timestamp 1679585382
transform 1 0 74400 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_776
timestamp 1679585382
transform 1 0 75072 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_783
timestamp 1679585382
transform 1 0 75744 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_790
timestamp 1679585382
transform 1 0 76416 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_797
timestamp 1679585382
transform 1 0 77088 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_804
timestamp 1679585382
transform 1 0 77760 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_811
timestamp 1679585382
transform 1 0 78432 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_818
timestamp 1679585382
transform 1 0 79104 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_825
timestamp 1679585382
transform 1 0 79776 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_832
timestamp 1679585382
transform 1 0 80448 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_839
timestamp 1679585382
transform 1 0 81120 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_846
timestamp 1679585382
transform 1 0 81792 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_853
timestamp 1679585382
transform 1 0 82464 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_860
timestamp 1679585382
transform 1 0 83136 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_867
timestamp 1679585382
transform 1 0 83808 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_874
timestamp 1679585382
transform 1 0 84480 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_881
timestamp 1679585382
transform 1 0 85152 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_888
timestamp 1679585382
transform 1 0 85824 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_895
timestamp 1679585382
transform 1 0 86496 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_902
timestamp 1679585382
transform 1 0 87168 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_909
timestamp 1679585382
transform 1 0 87840 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_916
timestamp 1679585382
transform 1 0 88512 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_923
timestamp 1679585382
transform 1 0 89184 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_930
timestamp 1679585382
transform 1 0 89856 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_937
timestamp 1679585382
transform 1 0 90528 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_944
timestamp 1679585382
transform 1 0 91200 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_951
timestamp 1679585382
transform 1 0 91872 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_958
timestamp 1679585382
transform 1 0 92544 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_965
timestamp 1679585382
transform 1 0 93216 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_972
timestamp 1679585382
transform 1 0 93888 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_979
timestamp 1679585382
transform 1 0 94560 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_986
timestamp 1679585382
transform 1 0 95232 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_993
timestamp 1679585382
transform 1 0 95904 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1000
timestamp 1679585382
transform 1 0 96576 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1007
timestamp 1679585382
transform 1 0 97248 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1014
timestamp 1679585382
transform 1 0 97920 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1021
timestamp 1679585382
transform 1 0 98592 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_1028
timestamp 1677583258
transform 1 0 99264 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_4
timestamp 1679585382
transform 1 0 960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_11
timestamp 1679585382
transform 1 0 1632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_18
timestamp 1679585382
transform 1 0 2304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_25
timestamp 1679585382
transform 1 0 2976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_32
timestamp 1679585382
transform 1 0 3648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_39
timestamp 1679585382
transform 1 0 4320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_46
timestamp 1679585382
transform 1 0 4992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_53
timestamp 1679585382
transform 1 0 5664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_60
timestamp 1679585382
transform 1 0 6336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_67
timestamp 1679585382
transform 1 0 7008 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_74
timestamp 1679585382
transform 1 0 7680 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_81
timestamp 1679585382
transform 1 0 8352 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_88
timestamp 1679585382
transform 1 0 9024 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_95
timestamp 1679585382
transform 1 0 9696 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_102
timestamp 1679581501
transform 1 0 10368 0 1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_137
timestamp 1679585382
transform 1 0 13728 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_144
timestamp 1679585382
transform 1 0 14400 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_151
timestamp 1679585382
transform 1 0 15072 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_158
timestamp 1679585382
transform 1 0 15744 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_165
timestamp 1679585382
transform 1 0 16416 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_172
timestamp 1679585382
transform 1 0 17088 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_179
timestamp 1679585382
transform 1 0 17760 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_186
timestamp 1679585382
transform 1 0 18432 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_193
timestamp 1679585382
transform 1 0 19104 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_200
timestamp 1679585382
transform 1 0 19776 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_243
timestamp 1679581501
transform 1 0 23904 0 1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_256
timestamp 1679585382
transform 1 0 25152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_263
timestamp 1679585382
transform 1 0 25824 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_270
timestamp 1679581501
transform 1 0 26496 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_274
timestamp 1677583258
transform 1 0 26880 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_311
timestamp 1679585382
transform 1 0 30432 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_318
timestamp 1679585382
transform 1 0 31104 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_325
timestamp 1679585382
transform 1 0 31776 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_332
timestamp 1679585382
transform 1 0 32448 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_339
timestamp 1679585382
transform 1 0 33120 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_346
timestamp 1679581501
transform 1 0 33792 0 1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_354
timestamp 1679585382
transform 1 0 34560 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_361
timestamp 1679585382
transform 1 0 35232 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_368
timestamp 1679585382
transform 1 0 35904 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_375
timestamp 1679585382
transform 1 0 36576 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_382
timestamp 1679585382
transform 1 0 37248 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_389
timestamp 1677583704
transform 1 0 37920 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_391
timestamp 1677583258
transform 1 0 38112 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_401
timestamp 1679585382
transform 1 0 39072 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_408
timestamp 1677583704
transform 1 0 39744 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_419
timestamp 1677583704
transform 1 0 40800 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_429
timestamp 1679585382
transform 1 0 41760 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_436
timestamp 1679585382
transform 1 0 42432 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_443
timestamp 1679585382
transform 1 0 43104 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_450
timestamp 1679585382
transform 1 0 43776 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_457
timestamp 1679585382
transform 1 0 44448 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_464
timestamp 1679585382
transform 1 0 45120 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_471
timestamp 1679585382
transform 1 0 45792 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_478
timestamp 1679585382
transform 1 0 46464 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_485
timestamp 1679585382
transform 1 0 47136 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_492
timestamp 1679585382
transform 1 0 47808 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_499
timestamp 1679585382
transform 1 0 48480 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_506
timestamp 1679585382
transform 1 0 49152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_513
timestamp 1679585382
transform 1 0 49824 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_520
timestamp 1679585382
transform 1 0 50496 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_527
timestamp 1679585382
transform 1 0 51168 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_534
timestamp 1679585382
transform 1 0 51840 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_541
timestamp 1679585382
transform 1 0 52512 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_548
timestamp 1679585382
transform 1 0 53184 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_555
timestamp 1677583258
transform 1 0 53856 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_560
timestamp 1679585382
transform 1 0 54336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_567
timestamp 1679585382
transform 1 0 55008 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_574
timestamp 1677583258
transform 1 0 55680 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_584
timestamp 1679585382
transform 1 0 56640 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_591
timestamp 1679585382
transform 1 0 57312 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_598
timestamp 1679585382
transform 1 0 57984 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_605
timestamp 1679585382
transform 1 0 58656 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_612
timestamp 1679585382
transform 1 0 59328 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_619
timestamp 1679585382
transform 1 0 60000 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_626
timestamp 1679585382
transform 1 0 60672 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_633
timestamp 1679585382
transform 1 0 61344 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_640
timestamp 1679585382
transform 1 0 62016 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_647
timestamp 1679585382
transform 1 0 62688 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_654
timestamp 1679585382
transform 1 0 63360 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_661
timestamp 1679585382
transform 1 0 64032 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_668
timestamp 1679585382
transform 1 0 64704 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_675
timestamp 1679585382
transform 1 0 65376 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_682
timestamp 1679585382
transform 1 0 66048 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_689
timestamp 1679585382
transform 1 0 66720 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_696
timestamp 1679585382
transform 1 0 67392 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_703
timestamp 1679585382
transform 1 0 68064 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_710
timestamp 1679585382
transform 1 0 68736 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_717
timestamp 1679585382
transform 1 0 69408 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_724
timestamp 1679585382
transform 1 0 70080 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_731
timestamp 1679585382
transform 1 0 70752 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_738
timestamp 1679585382
transform 1 0 71424 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_745
timestamp 1679585382
transform 1 0 72096 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_752
timestamp 1679585382
transform 1 0 72768 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_759
timestamp 1679585382
transform 1 0 73440 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_766
timestamp 1679585382
transform 1 0 74112 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_773
timestamp 1679585382
transform 1 0 74784 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_780
timestamp 1679585382
transform 1 0 75456 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_787
timestamp 1679585382
transform 1 0 76128 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_794
timestamp 1679585382
transform 1 0 76800 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_801
timestamp 1679585382
transform 1 0 77472 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_808
timestamp 1679585382
transform 1 0 78144 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_815
timestamp 1679585382
transform 1 0 78816 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_822
timestamp 1679585382
transform 1 0 79488 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_829
timestamp 1679585382
transform 1 0 80160 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_836
timestamp 1679585382
transform 1 0 80832 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_843
timestamp 1679585382
transform 1 0 81504 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_850
timestamp 1679585382
transform 1 0 82176 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_857
timestamp 1679585382
transform 1 0 82848 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_864
timestamp 1679585382
transform 1 0 83520 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_871
timestamp 1679585382
transform 1 0 84192 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_878
timestamp 1679585382
transform 1 0 84864 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_885
timestamp 1679585382
transform 1 0 85536 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_892
timestamp 1679585382
transform 1 0 86208 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_899
timestamp 1679585382
transform 1 0 86880 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_906
timestamp 1679585382
transform 1 0 87552 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_913
timestamp 1679585382
transform 1 0 88224 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_920
timestamp 1679585382
transform 1 0 88896 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_927
timestamp 1679585382
transform 1 0 89568 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_934
timestamp 1679585382
transform 1 0 90240 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_941
timestamp 1679585382
transform 1 0 90912 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_948
timestamp 1679585382
transform 1 0 91584 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_955
timestamp 1679585382
transform 1 0 92256 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_962
timestamp 1679585382
transform 1 0 92928 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_969
timestamp 1679585382
transform 1 0 93600 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_976
timestamp 1679585382
transform 1 0 94272 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_983
timestamp 1679585382
transform 1 0 94944 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_990
timestamp 1679585382
transform 1 0 95616 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_997
timestamp 1679585382
transform 1 0 96288 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1004
timestamp 1679585382
transform 1 0 96960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1011
timestamp 1679585382
transform 1 0 97632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1018
timestamp 1679585382
transform 1 0 98304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_1025
timestamp 1679581501
transform 1 0 98976 0 1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_4
timestamp 1679585382
transform 1 0 960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_11
timestamp 1679585382
transform 1 0 1632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_18
timestamp 1679585382
transform 1 0 2304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_25
timestamp 1679585382
transform 1 0 2976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_32
timestamp 1679585382
transform 1 0 3648 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_39
timestamp 1679585382
transform 1 0 4320 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_46
timestamp 1679585382
transform 1 0 4992 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_53
timestamp 1679585382
transform 1 0 5664 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_60
timestamp 1679585382
transform 1 0 6336 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_67
timestamp 1679585382
transform 1 0 7008 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_74
timestamp 1679585382
transform 1 0 7680 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_81
timestamp 1679585382
transform 1 0 8352 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_88
timestamp 1679585382
transform 1 0 9024 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_95
timestamp 1679585382
transform 1 0 9696 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_102
timestamp 1679585382
transform 1 0 10368 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_109
timestamp 1679581501
transform 1 0 11040 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_140
timestamp 1679585382
transform 1 0 14016 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_147
timestamp 1679585382
transform 1 0 14688 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_154
timestamp 1679585382
transform 1 0 15360 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_161
timestamp 1679585382
transform 1 0 16032 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_168
timestamp 1679585382
transform 1 0 16704 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_175
timestamp 1679585382
transform 1 0 17376 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_182
timestamp 1679585382
transform 1 0 18048 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_189
timestamp 1679585382
transform 1 0 18720 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_196
timestamp 1679585382
transform 1 0 19392 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_203
timestamp 1679585382
transform 1 0 20064 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_210
timestamp 1679585382
transform 1 0 20736 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_217
timestamp 1679585382
transform 1 0 21408 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_224
timestamp 1679585382
transform 1 0 22080 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_231
timestamp 1679585382
transform 1 0 22752 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_238
timestamp 1679585382
transform 1 0 23424 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_245
timestamp 1679585382
transform 1 0 24096 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_252
timestamp 1679585382
transform 1 0 24768 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_259
timestamp 1677583258
transform 1 0 25440 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_296
timestamp 1679585382
transform 1 0 28992 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_303
timestamp 1679585382
transform 1 0 29664 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_310
timestamp 1679585382
transform 1 0 30336 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_317
timestamp 1679585382
transform 1 0 31008 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_324
timestamp 1679585382
transform 1 0 31680 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_331
timestamp 1679585382
transform 1 0 32352 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_338
timestamp 1679585382
transform 1 0 33024 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_345
timestamp 1679585382
transform 1 0 33696 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_352
timestamp 1679585382
transform 1 0 34368 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_359
timestamp 1679585382
transform 1 0 35040 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_366
timestamp 1679585382
transform 1 0 35712 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_373
timestamp 1679585382
transform 1 0 36384 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_380
timestamp 1679585382
transform 1 0 37056 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_387
timestamp 1679585382
transform 1 0 37728 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_394
timestamp 1679585382
transform 1 0 38400 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_401
timestamp 1677583258
transform 1 0 39072 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_406
timestamp 1679585382
transform 1 0 39552 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_413
timestamp 1679585382
transform 1 0 40224 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_420
timestamp 1677583704
transform 1 0 40896 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_422
timestamp 1677583258
transform 1 0 41088 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_450
timestamp 1679585382
transform 1 0 43776 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_457
timestamp 1679585382
transform 1 0 44448 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_464
timestamp 1677583258
transform 1 0 45120 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_492
timestamp 1679585382
transform 1 0 47808 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_499
timestamp 1679585382
transform 1 0 48480 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_506
timestamp 1679585382
transform 1 0 49152 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_513
timestamp 1679585382
transform 1 0 49824 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_520
timestamp 1679585382
transform 1 0 50496 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_527
timestamp 1679585382
transform 1 0 51168 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_539
timestamp 1679585382
transform 1 0 52320 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_546
timestamp 1679585382
transform 1 0 52992 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_553
timestamp 1679585382
transform 1 0 53664 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_591
timestamp 1679585382
transform 1 0 57312 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_598
timestamp 1679585382
transform 1 0 57984 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_605
timestamp 1679585382
transform 1 0 58656 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_612
timestamp 1679585382
transform 1 0 59328 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_619
timestamp 1679585382
transform 1 0 60000 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_626
timestamp 1679585382
transform 1 0 60672 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_633
timestamp 1679585382
transform 1 0 61344 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_640
timestamp 1679585382
transform 1 0 62016 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_647
timestamp 1679585382
transform 1 0 62688 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_654
timestamp 1679585382
transform 1 0 63360 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_661
timestamp 1679585382
transform 1 0 64032 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_668
timestamp 1679585382
transform 1 0 64704 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_675
timestamp 1679585382
transform 1 0 65376 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_682
timestamp 1679585382
transform 1 0 66048 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_689
timestamp 1679585382
transform 1 0 66720 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_696
timestamp 1679585382
transform 1 0 67392 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_703
timestamp 1679585382
transform 1 0 68064 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_710
timestamp 1679585382
transform 1 0 68736 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_717
timestamp 1679585382
transform 1 0 69408 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_724
timestamp 1679585382
transform 1 0 70080 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_731
timestamp 1679585382
transform 1 0 70752 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_738
timestamp 1679585382
transform 1 0 71424 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_745
timestamp 1679585382
transform 1 0 72096 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_752
timestamp 1679585382
transform 1 0 72768 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_759
timestamp 1679585382
transform 1 0 73440 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_766
timestamp 1679585382
transform 1 0 74112 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_773
timestamp 1679585382
transform 1 0 74784 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_780
timestamp 1679585382
transform 1 0 75456 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_787
timestamp 1679585382
transform 1 0 76128 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_794
timestamp 1679585382
transform 1 0 76800 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_801
timestamp 1679585382
transform 1 0 77472 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_808
timestamp 1679585382
transform 1 0 78144 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_815
timestamp 1679585382
transform 1 0 78816 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_822
timestamp 1679585382
transform 1 0 79488 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_829
timestamp 1679585382
transform 1 0 80160 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_836
timestamp 1679585382
transform 1 0 80832 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_843
timestamp 1679585382
transform 1 0 81504 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_850
timestamp 1679585382
transform 1 0 82176 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_857
timestamp 1679585382
transform 1 0 82848 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_864
timestamp 1679585382
transform 1 0 83520 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_871
timestamp 1679585382
transform 1 0 84192 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_878
timestamp 1679585382
transform 1 0 84864 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_885
timestamp 1679585382
transform 1 0 85536 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_892
timestamp 1679585382
transform 1 0 86208 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_899
timestamp 1679585382
transform 1 0 86880 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_906
timestamp 1679585382
transform 1 0 87552 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_913
timestamp 1679585382
transform 1 0 88224 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_920
timestamp 1679585382
transform 1 0 88896 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_927
timestamp 1679585382
transform 1 0 89568 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_934
timestamp 1679585382
transform 1 0 90240 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_941
timestamp 1679585382
transform 1 0 90912 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_948
timestamp 1679585382
transform 1 0 91584 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_955
timestamp 1679585382
transform 1 0 92256 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_962
timestamp 1679585382
transform 1 0 92928 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_969
timestamp 1679585382
transform 1 0 93600 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_976
timestamp 1679585382
transform 1 0 94272 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_983
timestamp 1679585382
transform 1 0 94944 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_990
timestamp 1679585382
transform 1 0 95616 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_997
timestamp 1679585382
transform 1 0 96288 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1004
timestamp 1679585382
transform 1 0 96960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1011
timestamp 1679585382
transform 1 0 97632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1018
timestamp 1679585382
transform 1 0 98304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_1025
timestamp 1679581501
transform 1 0 98976 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_4
timestamp 1679585382
transform 1 0 960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_11
timestamp 1679585382
transform 1 0 1632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_18
timestamp 1679585382
transform 1 0 2304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_25
timestamp 1679585382
transform 1 0 2976 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_32
timestamp 1679585382
transform 1 0 3648 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_39
timestamp 1679585382
transform 1 0 4320 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_46
timestamp 1679585382
transform 1 0 4992 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_53
timestamp 1679585382
transform 1 0 5664 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_60
timestamp 1679585382
transform 1 0 6336 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_67
timestamp 1679585382
transform 1 0 7008 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_74
timestamp 1679585382
transform 1 0 7680 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_81
timestamp 1679585382
transform 1 0 8352 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_88
timestamp 1679585382
transform 1 0 9024 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_95
timestamp 1679585382
transform 1 0 9696 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_102
timestamp 1679585382
transform 1 0 10368 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_109
timestamp 1679585382
transform 1 0 11040 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_116
timestamp 1679581501
transform 1 0 11712 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_120
timestamp 1677583704
transform 1 0 12096 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_131
timestamp 1679585382
transform 1 0 13152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_138
timestamp 1679585382
transform 1 0 13824 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_145
timestamp 1679581501
transform 1 0 14496 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_149
timestamp 1677583258
transform 1 0 14880 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_163
timestamp 1679585382
transform 1 0 16224 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_170
timestamp 1677583704
transform 1 0 16896 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_185
timestamp 1679585382
transform 1 0 18336 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_192
timestamp 1679585382
transform 1 0 19008 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_199
timestamp 1679585382
transform 1 0 19680 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_206
timestamp 1679585382
transform 1 0 20352 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_213
timestamp 1679585382
transform 1 0 21024 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_220
timestamp 1679585382
transform 1 0 21696 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_227
timestamp 1679585382
transform 1 0 22368 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_234
timestamp 1679585382
transform 1 0 23040 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_241
timestamp 1679585382
transform 1 0 23712 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_248
timestamp 1679585382
transform 1 0 24384 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_255
timestamp 1679585382
transform 1 0 25056 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_262
timestamp 1679585382
transform 1 0 25728 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_269
timestamp 1679585382
transform 1 0 26400 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_276
timestamp 1679585382
transform 1 0 27072 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_283
timestamp 1679585382
transform 1 0 27744 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_290
timestamp 1679585382
transform 1 0 28416 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_297
timestamp 1679585382
transform 1 0 29088 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_304
timestamp 1679585382
transform 1 0 29760 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_311
timestamp 1679585382
transform 1 0 30432 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_318
timestamp 1679585382
transform 1 0 31104 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_325
timestamp 1679585382
transform 1 0 31776 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_332
timestamp 1679581501
transform 1 0 32448 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_349
timestamp 1679585382
transform 1 0 34080 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_356
timestamp 1679585382
transform 1 0 34752 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_363
timestamp 1679585382
transform 1 0 35424 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_370
timestamp 1679585382
transform 1 0 36096 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_377
timestamp 1679585382
transform 1 0 36768 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_384
timestamp 1677583704
transform 1 0 37440 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_413
timestamp 1679585382
transform 1 0 40224 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_420
timestamp 1679585382
transform 1 0 40896 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_427
timestamp 1679585382
transform 1 0 41568 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_434
timestamp 1679585382
transform 1 0 42240 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_441
timestamp 1679585382
transform 1 0 42912 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_448
timestamp 1679585382
transform 1 0 43584 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_455
timestamp 1679585382
transform 1 0 44256 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_462
timestamp 1677583704
transform 1 0 44928 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_464
timestamp 1677583258
transform 1 0 45120 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_474
timestamp 1677583704
transform 1 0 46080 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_476
timestamp 1677583258
transform 1 0 46272 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_481
timestamp 1677583258
transform 1 0 46752 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_503
timestamp 1679585382
transform 1 0 48864 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_510
timestamp 1679585382
transform 1 0 49536 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_517
timestamp 1679585382
transform 1 0 50208 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_524
timestamp 1679585382
transform 1 0 50880 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_531
timestamp 1679581501
transform 1 0 51552 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_535
timestamp 1677583704
transform 1 0 51936 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_568
timestamp 1679585382
transform 1 0 55104 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_575
timestamp 1677583258
transform 1 0 55776 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_585
timestamp 1679585382
transform 1 0 56736 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_592
timestamp 1679585382
transform 1 0 57408 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_599
timestamp 1679585382
transform 1 0 58080 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_606
timestamp 1679585382
transform 1 0 58752 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_613
timestamp 1679585382
transform 1 0 59424 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_620
timestamp 1679585382
transform 1 0 60096 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_627
timestamp 1679585382
transform 1 0 60768 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_634
timestamp 1679585382
transform 1 0 61440 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_641
timestamp 1679585382
transform 1 0 62112 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_648
timestamp 1679585382
transform 1 0 62784 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_655
timestamp 1679585382
transform 1 0 63456 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_662
timestamp 1679585382
transform 1 0 64128 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_669
timestamp 1679585382
transform 1 0 64800 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_676
timestamp 1679585382
transform 1 0 65472 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_683
timestamp 1679585382
transform 1 0 66144 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_690
timestamp 1679585382
transform 1 0 66816 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_697
timestamp 1679585382
transform 1 0 67488 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_704
timestamp 1679585382
transform 1 0 68160 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_711
timestamp 1679585382
transform 1 0 68832 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_718
timestamp 1679585382
transform 1 0 69504 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_725
timestamp 1679585382
transform 1 0 70176 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_732
timestamp 1679585382
transform 1 0 70848 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_739
timestamp 1679585382
transform 1 0 71520 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_746
timestamp 1679585382
transform 1 0 72192 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_753
timestamp 1679585382
transform 1 0 72864 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_760
timestamp 1679585382
transform 1 0 73536 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_767
timestamp 1679585382
transform 1 0 74208 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_774
timestamp 1679585382
transform 1 0 74880 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_781
timestamp 1679585382
transform 1 0 75552 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_788
timestamp 1679585382
transform 1 0 76224 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_795
timestamp 1679585382
transform 1 0 76896 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_802
timestamp 1679585382
transform 1 0 77568 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_809
timestamp 1679585382
transform 1 0 78240 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_816
timestamp 1679585382
transform 1 0 78912 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_823
timestamp 1679585382
transform 1 0 79584 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_830
timestamp 1679585382
transform 1 0 80256 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_837
timestamp 1679585382
transform 1 0 80928 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_844
timestamp 1679585382
transform 1 0 81600 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_851
timestamp 1679585382
transform 1 0 82272 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_858
timestamp 1679585382
transform 1 0 82944 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_865
timestamp 1679585382
transform 1 0 83616 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_872
timestamp 1679585382
transform 1 0 84288 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_879
timestamp 1679585382
transform 1 0 84960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_886
timestamp 1679585382
transform 1 0 85632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_893
timestamp 1679585382
transform 1 0 86304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_900
timestamp 1679585382
transform 1 0 86976 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_907
timestamp 1679585382
transform 1 0 87648 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_914
timestamp 1679585382
transform 1 0 88320 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_921
timestamp 1679585382
transform 1 0 88992 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_928
timestamp 1679585382
transform 1 0 89664 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_935
timestamp 1679585382
transform 1 0 90336 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_942
timestamp 1679585382
transform 1 0 91008 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_949
timestamp 1679585382
transform 1 0 91680 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_956
timestamp 1679585382
transform 1 0 92352 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_963
timestamp 1679585382
transform 1 0 93024 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_970
timestamp 1679585382
transform 1 0 93696 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_977
timestamp 1679585382
transform 1 0 94368 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_984
timestamp 1679585382
transform 1 0 95040 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_991
timestamp 1679585382
transform 1 0 95712 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_998
timestamp 1679585382
transform 1 0 96384 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1005
timestamp 1679585382
transform 1 0 97056 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1012
timestamp 1679585382
transform 1 0 97728 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1019
timestamp 1679585382
transform 1 0 98400 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_1026
timestamp 1677583704
transform 1 0 99072 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_1028
timestamp 1677583258
transform 1 0 99264 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679585382
transform 1 0 576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679585382
transform 1 0 1248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679585382
transform 1 0 1920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_21
timestamp 1679585382
transform 1 0 2592 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_28
timestamp 1679585382
transform 1 0 3264 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_35
timestamp 1679585382
transform 1 0 3936 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_42
timestamp 1679585382
transform 1 0 4608 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_49
timestamp 1679585382
transform 1 0 5280 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_56
timestamp 1679585382
transform 1 0 5952 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_63
timestamp 1679585382
transform 1 0 6624 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_70
timestamp 1679585382
transform 1 0 7296 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_77
timestamp 1679585382
transform 1 0 7968 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_84
timestamp 1679585382
transform 1 0 8640 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_91
timestamp 1679585382
transform 1 0 9312 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_98
timestamp 1679585382
transform 1 0 9984 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_105
timestamp 1679585382
transform 1 0 10656 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_112
timestamp 1679585382
transform 1 0 11328 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_119
timestamp 1679585382
transform 1 0 12000 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_126
timestamp 1679585382
transform 1 0 12672 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_133
timestamp 1679585382
transform 1 0 13344 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_140
timestamp 1679585382
transform 1 0 14016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_147
timestamp 1679585382
transform 1 0 14688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_154
timestamp 1679585382
transform 1 0 15360 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_161
timestamp 1679585382
transform 1 0 16032 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_168
timestamp 1679585382
transform 1 0 16704 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_175
timestamp 1679585382
transform 1 0 17376 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_182
timestamp 1679585382
transform 1 0 18048 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_189
timestamp 1679585382
transform 1 0 18720 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_196
timestamp 1679585382
transform 1 0 19392 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_203
timestamp 1679585382
transform 1 0 20064 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_210
timestamp 1679585382
transform 1 0 20736 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_230
timestamp 1679585382
transform 1 0 22656 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_237
timestamp 1679585382
transform 1 0 23328 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_244
timestamp 1679585382
transform 1 0 24000 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_251
timestamp 1679585382
transform 1 0 24672 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_258
timestamp 1679585382
transform 1 0 25344 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_265
timestamp 1679585382
transform 1 0 26016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_272
timestamp 1679585382
transform 1 0 26688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_279
timestamp 1679585382
transform 1 0 27360 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_286
timestamp 1679585382
transform 1 0 28032 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_306
timestamp 1679585382
transform 1 0 29952 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_313
timestamp 1679585382
transform 1 0 30624 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_320
timestamp 1679585382
transform 1 0 31296 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_327
timestamp 1679585382
transform 1 0 31968 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_334
timestamp 1679585382
transform 1 0 32640 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_341
timestamp 1679585382
transform 1 0 33312 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_348
timestamp 1679585382
transform 1 0 33984 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_355
timestamp 1679585382
transform 1 0 34656 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_362
timestamp 1679585382
transform 1 0 35328 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_369
timestamp 1679585382
transform 1 0 36000 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_376
timestamp 1679585382
transform 1 0 36672 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_383
timestamp 1679585382
transform 1 0 37344 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_390
timestamp 1679581501
transform 1 0 38016 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_394
timestamp 1677583258
transform 1 0 38400 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_399
timestamp 1677583704
transform 1 0 38880 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_401
timestamp 1677583258
transform 1 0 39072 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_415
timestamp 1679585382
transform 1 0 40416 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_422
timestamp 1679585382
transform 1 0 41088 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_429
timestamp 1679585382
transform 1 0 41760 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_436
timestamp 1679585382
transform 1 0 42432 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_443
timestamp 1679585382
transform 1 0 43104 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_450
timestamp 1679585382
transform 1 0 43776 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_457
timestamp 1677583704
transform 1 0 44448 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_459
timestamp 1677583258
transform 1 0 44640 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_477
timestamp 1679585382
transform 1 0 46368 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_484
timestamp 1679585382
transform 1 0 47040 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_491
timestamp 1677583704
transform 1 0 47712 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_502
timestamp 1679585382
transform 1 0 48768 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_509
timestamp 1679585382
transform 1 0 49440 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_516
timestamp 1679585382
transform 1 0 50112 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_523
timestamp 1679585382
transform 1 0 50784 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_530
timestamp 1679585382
transform 1 0 51456 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_537
timestamp 1679585382
transform 1 0 52128 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_544
timestamp 1677583704
transform 1 0 52800 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_568
timestamp 1679585382
transform 1 0 55104 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_575
timestamp 1679585382
transform 1 0 55776 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_582
timestamp 1679585382
transform 1 0 56448 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_589
timestamp 1679585382
transform 1 0 57120 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_596
timestamp 1679585382
transform 1 0 57792 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_603
timestamp 1679585382
transform 1 0 58464 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_610
timestamp 1679585382
transform 1 0 59136 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_617
timestamp 1679585382
transform 1 0 59808 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_624
timestamp 1679585382
transform 1 0 60480 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_631
timestamp 1679585382
transform 1 0 61152 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_638
timestamp 1679585382
transform 1 0 61824 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_645
timestamp 1679585382
transform 1 0 62496 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_652
timestamp 1679585382
transform 1 0 63168 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_659
timestamp 1679585382
transform 1 0 63840 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_666
timestamp 1679585382
transform 1 0 64512 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_673
timestamp 1679585382
transform 1 0 65184 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_680
timestamp 1679585382
transform 1 0 65856 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_687
timestamp 1679585382
transform 1 0 66528 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_694
timestamp 1679585382
transform 1 0 67200 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_701
timestamp 1679585382
transform 1 0 67872 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_708
timestamp 1679585382
transform 1 0 68544 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_715
timestamp 1679585382
transform 1 0 69216 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_722
timestamp 1679585382
transform 1 0 69888 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_729
timestamp 1679585382
transform 1 0 70560 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_736
timestamp 1679585382
transform 1 0 71232 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_743
timestamp 1679585382
transform 1 0 71904 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_750
timestamp 1679585382
transform 1 0 72576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_757
timestamp 1679585382
transform 1 0 73248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_764
timestamp 1679585382
transform 1 0 73920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_771
timestamp 1679585382
transform 1 0 74592 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_778
timestamp 1679585382
transform 1 0 75264 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_785
timestamp 1679585382
transform 1 0 75936 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_792
timestamp 1679585382
transform 1 0 76608 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_799
timestamp 1679585382
transform 1 0 77280 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_806
timestamp 1679585382
transform 1 0 77952 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_813
timestamp 1679585382
transform 1 0 78624 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_820
timestamp 1679585382
transform 1 0 79296 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_827
timestamp 1679585382
transform 1 0 79968 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_834
timestamp 1679585382
transform 1 0 80640 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_841
timestamp 1679585382
transform 1 0 81312 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_848
timestamp 1679585382
transform 1 0 81984 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_855
timestamp 1679585382
transform 1 0 82656 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_862
timestamp 1679585382
transform 1 0 83328 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_869
timestamp 1679585382
transform 1 0 84000 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_876
timestamp 1679585382
transform 1 0 84672 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_883
timestamp 1679585382
transform 1 0 85344 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_890
timestamp 1679585382
transform 1 0 86016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_897
timestamp 1679585382
transform 1 0 86688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_904
timestamp 1679585382
transform 1 0 87360 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_911
timestamp 1679585382
transform 1 0 88032 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_918
timestamp 1679585382
transform 1 0 88704 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_925
timestamp 1679585382
transform 1 0 89376 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_932
timestamp 1679585382
transform 1 0 90048 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_939
timestamp 1679585382
transform 1 0 90720 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_946
timestamp 1679585382
transform 1 0 91392 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_953
timestamp 1679585382
transform 1 0 92064 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_960
timestamp 1679585382
transform 1 0 92736 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_967
timestamp 1679585382
transform 1 0 93408 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_974
timestamp 1679585382
transform 1 0 94080 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_981
timestamp 1679585382
transform 1 0 94752 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_988
timestamp 1679585382
transform 1 0 95424 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_995
timestamp 1679585382
transform 1 0 96096 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1002
timestamp 1679585382
transform 1 0 96768 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1009
timestamp 1679585382
transform 1 0 97440 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1016
timestamp 1679585382
transform 1 0 98112 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_1023
timestamp 1679581501
transform 1 0 98784 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_1027
timestamp 1677583704
transform 1 0 99168 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_4
timestamp 1679585382
transform 1 0 960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_11
timestamp 1679585382
transform 1 0 1632 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_18
timestamp 1679585382
transform 1 0 2304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_25
timestamp 1679585382
transform 1 0 2976 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_32
timestamp 1679585382
transform 1 0 3648 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_39
timestamp 1679585382
transform 1 0 4320 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_46
timestamp 1679585382
transform 1 0 4992 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_53
timestamp 1679585382
transform 1 0 5664 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_60
timestamp 1679585382
transform 1 0 6336 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_67
timestamp 1679585382
transform 1 0 7008 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_74
timestamp 1679585382
transform 1 0 7680 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_81
timestamp 1679585382
transform 1 0 8352 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_88
timestamp 1679585382
transform 1 0 9024 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_95
timestamp 1679585382
transform 1 0 9696 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_102
timestamp 1679581501
transform 1 0 10368 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_106
timestamp 1677583258
transform 1 0 10752 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_120
timestamp 1679585382
transform 1 0 12096 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_127
timestamp 1679585382
transform 1 0 12768 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_134
timestamp 1679585382
transform 1 0 13440 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_141
timestamp 1679585382
transform 1 0 14112 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_148
timestamp 1679585382
transform 1 0 14784 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_155
timestamp 1679585382
transform 1 0 15456 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_189
timestamp 1679585382
transform 1 0 18720 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_196
timestamp 1679585382
transform 1 0 19392 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_203
timestamp 1677583704
transform 1 0 20064 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_241
timestamp 1679585382
transform 1 0 23712 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_248
timestamp 1679585382
transform 1 0 24384 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_255
timestamp 1679585382
transform 1 0 25056 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_262
timestamp 1677583704
transform 1 0 25728 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_273
timestamp 1679585382
transform 1 0 26784 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_280
timestamp 1679585382
transform 1 0 27456 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_287
timestamp 1677583258
transform 1 0 28128 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_316
timestamp 1679585382
transform 1 0 30912 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_332
timestamp 1679585382
transform 1 0 32448 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_339
timestamp 1677583704
transform 1 0 33120 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_341
timestamp 1677583258
transform 1 0 33312 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_369
timestamp 1679585382
transform 1 0 36000 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_376
timestamp 1679585382
transform 1 0 36672 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_383
timestamp 1679581501
transform 1 0 37344 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_387
timestamp 1677583704
transform 1 0 37728 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_398
timestamp 1679585382
transform 1 0 38784 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_414
timestamp 1679585382
transform 1 0 40320 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_421
timestamp 1679585382
transform 1 0 40992 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_428
timestamp 1679585382
transform 1 0 41664 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_435
timestamp 1679585382
transform 1 0 42336 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_442
timestamp 1679585382
transform 1 0 43008 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_449
timestamp 1679585382
transform 1 0 43680 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_456
timestamp 1679585382
transform 1 0 44352 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_463
timestamp 1679585382
transform 1 0 45024 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_470
timestamp 1679585382
transform 1 0 45696 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_477
timestamp 1679585382
transform 1 0 46368 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_484
timestamp 1679585382
transform 1 0 47040 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_491
timestamp 1679581501
transform 1 0 47712 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_495
timestamp 1677583704
transform 1 0 48096 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_524
timestamp 1679585382
transform 1 0 50880 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_531
timestamp 1679585382
transform 1 0 51552 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_538
timestamp 1679585382
transform 1 0 52224 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_545
timestamp 1679585382
transform 1 0 52896 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_552
timestamp 1679585382
transform 1 0 53568 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_559
timestamp 1679585382
transform 1 0 54240 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_566
timestamp 1679585382
transform 1 0 54912 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_573
timestamp 1679585382
transform 1 0 55584 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_580
timestamp 1679585382
transform 1 0 56256 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_587
timestamp 1679585382
transform 1 0 56928 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_594
timestamp 1679585382
transform 1 0 57600 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_601
timestamp 1679585382
transform 1 0 58272 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_608
timestamp 1679585382
transform 1 0 58944 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_615
timestamp 1679585382
transform 1 0 59616 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_622
timestamp 1679585382
transform 1 0 60288 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_629
timestamp 1679585382
transform 1 0 60960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_636
timestamp 1679585382
transform 1 0 61632 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_643
timestamp 1679585382
transform 1 0 62304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_650
timestamp 1679585382
transform 1 0 62976 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_657
timestamp 1679585382
transform 1 0 63648 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_664
timestamp 1679585382
transform 1 0 64320 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_671
timestamp 1679585382
transform 1 0 64992 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_678
timestamp 1679585382
transform 1 0 65664 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_685
timestamp 1679585382
transform 1 0 66336 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_692
timestamp 1679585382
transform 1 0 67008 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_699
timestamp 1679585382
transform 1 0 67680 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_706
timestamp 1679585382
transform 1 0 68352 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_713
timestamp 1679585382
transform 1 0 69024 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_720
timestamp 1679585382
transform 1 0 69696 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_727
timestamp 1679585382
transform 1 0 70368 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_734
timestamp 1679585382
transform 1 0 71040 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_741
timestamp 1679585382
transform 1 0 71712 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_748
timestamp 1679585382
transform 1 0 72384 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_755
timestamp 1679585382
transform 1 0 73056 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_762
timestamp 1679585382
transform 1 0 73728 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_769
timestamp 1679585382
transform 1 0 74400 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_776
timestamp 1679585382
transform 1 0 75072 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_783
timestamp 1679585382
transform 1 0 75744 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_790
timestamp 1679585382
transform 1 0 76416 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_797
timestamp 1679585382
transform 1 0 77088 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_804
timestamp 1679585382
transform 1 0 77760 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_811
timestamp 1679585382
transform 1 0 78432 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_818
timestamp 1679585382
transform 1 0 79104 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_825
timestamp 1679585382
transform 1 0 79776 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_832
timestamp 1679585382
transform 1 0 80448 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_839
timestamp 1679585382
transform 1 0 81120 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_846
timestamp 1679585382
transform 1 0 81792 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_853
timestamp 1679585382
transform 1 0 82464 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_860
timestamp 1679585382
transform 1 0 83136 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_867
timestamp 1679585382
transform 1 0 83808 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_874
timestamp 1679585382
transform 1 0 84480 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_881
timestamp 1679585382
transform 1 0 85152 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_888
timestamp 1679585382
transform 1 0 85824 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_895
timestamp 1679585382
transform 1 0 86496 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_902
timestamp 1679585382
transform 1 0 87168 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_909
timestamp 1679585382
transform 1 0 87840 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_916
timestamp 1679585382
transform 1 0 88512 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_923
timestamp 1679585382
transform 1 0 89184 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_930
timestamp 1679585382
transform 1 0 89856 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_937
timestamp 1679585382
transform 1 0 90528 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_944
timestamp 1679585382
transform 1 0 91200 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_951
timestamp 1679585382
transform 1 0 91872 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_958
timestamp 1679585382
transform 1 0 92544 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_965
timestamp 1679585382
transform 1 0 93216 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_972
timestamp 1679585382
transform 1 0 93888 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_979
timestamp 1679585382
transform 1 0 94560 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_986
timestamp 1679585382
transform 1 0 95232 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_993
timestamp 1679585382
transform 1 0 95904 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1000
timestamp 1679585382
transform 1 0 96576 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1007
timestamp 1679585382
transform 1 0 97248 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1014
timestamp 1679585382
transform 1 0 97920 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1021
timestamp 1679585382
transform 1 0 98592 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_1028
timestamp 1677583258
transform 1 0 99264 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_4
timestamp 1679585382
transform 1 0 960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_11
timestamp 1679581501
transform 1 0 1632 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_15
timestamp 1677583704
transform 1 0 2016 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_48
timestamp 1679585382
transform 1 0 5184 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_55
timestamp 1679585382
transform 1 0 5856 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_62
timestamp 1679585382
transform 1 0 6528 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_69
timestamp 1679585382
transform 1 0 7200 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_76
timestamp 1679581501
transform 1 0 7872 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_80
timestamp 1677583704
transform 1 0 8256 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_95
timestamp 1679585382
transform 1 0 9696 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_102
timestamp 1679585382
transform 1 0 10368 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_109
timestamp 1679585382
transform 1 0 11040 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_116
timestamp 1679585382
transform 1 0 11712 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_123
timestamp 1679585382
transform 1 0 12384 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_130
timestamp 1679585382
transform 1 0 13056 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_137
timestamp 1679585382
transform 1 0 13728 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_144
timestamp 1679585382
transform 1 0 14400 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_151
timestamp 1679585382
transform 1 0 15072 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_158
timestamp 1679585382
transform 1 0 15744 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_165
timestamp 1679585382
transform 1 0 16416 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_172
timestamp 1679585382
transform 1 0 17088 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_179
timestamp 1679585382
transform 1 0 17760 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_186
timestamp 1677583258
transform 1 0 18432 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_195
timestamp 1679585382
transform 1 0 19296 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_202
timestamp 1679585382
transform 1 0 19968 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_209
timestamp 1679585382
transform 1 0 20640 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_216
timestamp 1679581501
transform 1 0 21312 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_4  FILLER_9_228
timestamp 1679581501
transform 1 0 22464 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_237
timestamp 1679585382
transform 1 0 23328 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_244
timestamp 1679585382
transform 1 0 24000 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_251
timestamp 1677583704
transform 1 0 24672 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_280
timestamp 1679585382
transform 1 0 27456 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_287
timestamp 1679585382
transform 1 0 28128 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_294
timestamp 1679585382
transform 1 0 28800 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_306
timestamp 1677583704
transform 1 0 29952 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_308
timestamp 1677583258
transform 1 0 30144 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_318
timestamp 1679585382
transform 1 0 31104 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_325
timestamp 1679581501
transform 1 0 31776 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_4  FILLER_9_338
timestamp 1679581501
transform 1 0 33024 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_370
timestamp 1677583258
transform 1 0 36096 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_384
timestamp 1677583704
transform 1 0 37440 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_399
timestamp 1679585382
transform 1 0 38880 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_406
timestamp 1677583704
transform 1 0 39552 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_416
timestamp 1679585382
transform 1 0 40512 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_423
timestamp 1679585382
transform 1 0 41184 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_430
timestamp 1679585382
transform 1 0 41856 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_437
timestamp 1679585382
transform 1 0 42528 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_444
timestamp 1679585382
transform 1 0 43200 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_451
timestamp 1679585382
transform 1 0 43872 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_458
timestamp 1679585382
transform 1 0 44544 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_465
timestamp 1677583704
transform 1 0 45216 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_467
timestamp 1677583258
transform 1 0 45408 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_477
timestamp 1679585382
transform 1 0 46368 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_484
timestamp 1679585382
transform 1 0 47040 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_491
timestamp 1679585382
transform 1 0 47712 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_498
timestamp 1679585382
transform 1 0 48384 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_505
timestamp 1679585382
transform 1 0 49056 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_512
timestamp 1679585382
transform 1 0 49728 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_519
timestamp 1677583704
transform 1 0 50400 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_521
timestamp 1677583258
transform 1 0 50592 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_535
timestamp 1679585382
transform 1 0 51936 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_542
timestamp 1679585382
transform 1 0 52608 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_549
timestamp 1679585382
transform 1 0 53280 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_556
timestamp 1679585382
transform 1 0 53952 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_563
timestamp 1679585382
transform 1 0 54624 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_570
timestamp 1679585382
transform 1 0 55296 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_577
timestamp 1679585382
transform 1 0 55968 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_584
timestamp 1679585382
transform 1 0 56640 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_591
timestamp 1679585382
transform 1 0 57312 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_598
timestamp 1679585382
transform 1 0 57984 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_605
timestamp 1679585382
transform 1 0 58656 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_612
timestamp 1679585382
transform 1 0 59328 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_619
timestamp 1679585382
transform 1 0 60000 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_626
timestamp 1679585382
transform 1 0 60672 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_633
timestamp 1679585382
transform 1 0 61344 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_640
timestamp 1679585382
transform 1 0 62016 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_647
timestamp 1679585382
transform 1 0 62688 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_654
timestamp 1679585382
transform 1 0 63360 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_661
timestamp 1679585382
transform 1 0 64032 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_668
timestamp 1679585382
transform 1 0 64704 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_675
timestamp 1679585382
transform 1 0 65376 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_682
timestamp 1679585382
transform 1 0 66048 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_689
timestamp 1679585382
transform 1 0 66720 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_696
timestamp 1679585382
transform 1 0 67392 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_703
timestamp 1679585382
transform 1 0 68064 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_710
timestamp 1679585382
transform 1 0 68736 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_717
timestamp 1679585382
transform 1 0 69408 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_724
timestamp 1679585382
transform 1 0 70080 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_731
timestamp 1679585382
transform 1 0 70752 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_738
timestamp 1679585382
transform 1 0 71424 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_745
timestamp 1679585382
transform 1 0 72096 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_752
timestamp 1679585382
transform 1 0 72768 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_759
timestamp 1679585382
transform 1 0 73440 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_766
timestamp 1679585382
transform 1 0 74112 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_773
timestamp 1679585382
transform 1 0 74784 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_780
timestamp 1679585382
transform 1 0 75456 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_787
timestamp 1679585382
transform 1 0 76128 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_794
timestamp 1679585382
transform 1 0 76800 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_801
timestamp 1679585382
transform 1 0 77472 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_808
timestamp 1679585382
transform 1 0 78144 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_815
timestamp 1679585382
transform 1 0 78816 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_822
timestamp 1679585382
transform 1 0 79488 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_829
timestamp 1679585382
transform 1 0 80160 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_836
timestamp 1679585382
transform 1 0 80832 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_843
timestamp 1679585382
transform 1 0 81504 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_850
timestamp 1679585382
transform 1 0 82176 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_857
timestamp 1679585382
transform 1 0 82848 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_864
timestamp 1679585382
transform 1 0 83520 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_871
timestamp 1679585382
transform 1 0 84192 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_878
timestamp 1679585382
transform 1 0 84864 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_885
timestamp 1679585382
transform 1 0 85536 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_892
timestamp 1679585382
transform 1 0 86208 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_899
timestamp 1679585382
transform 1 0 86880 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_906
timestamp 1679585382
transform 1 0 87552 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_913
timestamp 1679585382
transform 1 0 88224 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_920
timestamp 1679585382
transform 1 0 88896 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_927
timestamp 1679585382
transform 1 0 89568 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_934
timestamp 1679585382
transform 1 0 90240 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_941
timestamp 1679585382
transform 1 0 90912 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_948
timestamp 1679585382
transform 1 0 91584 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_955
timestamp 1679585382
transform 1 0 92256 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_962
timestamp 1679585382
transform 1 0 92928 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_969
timestamp 1679585382
transform 1 0 93600 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_976
timestamp 1679585382
transform 1 0 94272 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_983
timestamp 1679585382
transform 1 0 94944 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_990
timestamp 1679585382
transform 1 0 95616 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_997
timestamp 1679585382
transform 1 0 96288 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1004
timestamp 1679585382
transform 1 0 96960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1011
timestamp 1679585382
transform 1 0 97632 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1018
timestamp 1679585382
transform 1 0 98304 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_1025
timestamp 1679581501
transform 1 0 98976 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_10_4
timestamp 1679585382
transform 1 0 960 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_11
timestamp 1677583704
transform 1 0 1632 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_13
timestamp 1677583258
transform 1 0 1824 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_41
timestamp 1677583704
transform 1 0 4512 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_124
timestamp 1679585382
transform 1 0 12480 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_131
timestamp 1679585382
transform 1 0 13152 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_138
timestamp 1679585382
transform 1 0 13824 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_145
timestamp 1679585382
transform 1 0 14496 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_152
timestamp 1679585382
transform 1 0 15168 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_159
timestamp 1679585382
transform 1 0 15840 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_166
timestamp 1679585382
transform 1 0 16512 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_173
timestamp 1679585382
transform 1 0 17184 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_180
timestamp 1679581501
transform 1 0 17856 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_184
timestamp 1677583704
transform 1 0 18240 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_203
timestamp 1679585382
transform 1 0 20064 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_210
timestamp 1677583258
transform 1 0 20736 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_227
timestamp 1679585382
transform 1 0 22368 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_234
timestamp 1679585382
transform 1 0 23040 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_241
timestamp 1679585382
transform 1 0 23712 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_248
timestamp 1679585382
transform 1 0 24384 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_255
timestamp 1679585382
transform 1 0 25056 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_267
timestamp 1679585382
transform 1 0 26208 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_274
timestamp 1679585382
transform 1 0 26880 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_281
timestamp 1679585382
transform 1 0 27552 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_288
timestamp 1679581501
transform 1 0 28224 0 1 8316
box -48 -56 432 834
use sg13g2_decap_4  FILLER_10_301
timestamp 1679581501
transform 1 0 29472 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_305
timestamp 1677583258
transform 1 0 29856 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_310
timestamp 1679585382
transform 1 0 30336 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_317
timestamp 1679585382
transform 1 0 31008 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_324
timestamp 1679585382
transform 1 0 31680 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_331
timestamp 1679585382
transform 1 0 32352 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_338
timestamp 1679585382
transform 1 0 33024 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_345
timestamp 1679585382
transform 1 0 33696 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_352
timestamp 1679585382
transform 1 0 34368 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_359
timestamp 1679585382
transform 1 0 35040 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_366
timestamp 1679585382
transform 1 0 35712 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_373
timestamp 1679585382
transform 1 0 36384 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_380
timestamp 1679585382
transform 1 0 37056 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_387
timestamp 1679581501
transform 1 0 37728 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_391
timestamp 1677583704
transform 1 0 38112 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_402
timestamp 1677583704
transform 1 0 39168 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_404
timestamp 1677583258
transform 1 0 39360 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_414
timestamp 1677583704
transform 1 0 40320 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_424
timestamp 1679585382
transform 1 0 41280 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_431
timestamp 1679585382
transform 1 0 41952 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_438
timestamp 1679585382
transform 1 0 42624 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_445
timestamp 1679585382
transform 1 0 43296 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_452
timestamp 1679585382
transform 1 0 43968 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_459
timestamp 1679585382
transform 1 0 44640 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_466
timestamp 1677583258
transform 1 0 45312 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_494
timestamp 1679585382
transform 1 0 48000 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_501
timestamp 1679585382
transform 1 0 48672 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_508
timestamp 1679585382
transform 1 0 49344 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_515
timestamp 1679585382
transform 1 0 50016 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_522
timestamp 1679585382
transform 1 0 50688 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_529
timestamp 1679585382
transform 1 0 51360 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_536
timestamp 1679585382
transform 1 0 52032 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_543
timestamp 1679585382
transform 1 0 52704 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_550
timestamp 1679585382
transform 1 0 53376 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_557
timestamp 1679585382
transform 1 0 54048 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_564
timestamp 1679585382
transform 1 0 54720 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_571
timestamp 1679585382
transform 1 0 55392 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_578
timestamp 1679585382
transform 1 0 56064 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_585
timestamp 1679585382
transform 1 0 56736 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_592
timestamp 1679585382
transform 1 0 57408 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_599
timestamp 1679585382
transform 1 0 58080 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_606
timestamp 1679585382
transform 1 0 58752 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_613
timestamp 1679585382
transform 1 0 59424 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_620
timestamp 1679585382
transform 1 0 60096 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_627
timestamp 1679585382
transform 1 0 60768 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_634
timestamp 1679585382
transform 1 0 61440 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_641
timestamp 1679585382
transform 1 0 62112 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_648
timestamp 1679585382
transform 1 0 62784 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_655
timestamp 1679585382
transform 1 0 63456 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_662
timestamp 1679585382
transform 1 0 64128 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_669
timestamp 1679585382
transform 1 0 64800 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_676
timestamp 1679585382
transform 1 0 65472 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_683
timestamp 1679585382
transform 1 0 66144 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_690
timestamp 1679585382
transform 1 0 66816 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_697
timestamp 1679585382
transform 1 0 67488 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_704
timestamp 1679585382
transform 1 0 68160 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_711
timestamp 1679585382
transform 1 0 68832 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_718
timestamp 1679585382
transform 1 0 69504 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_725
timestamp 1679585382
transform 1 0 70176 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_732
timestamp 1679585382
transform 1 0 70848 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_739
timestamp 1679585382
transform 1 0 71520 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_746
timestamp 1679585382
transform 1 0 72192 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_753
timestamp 1679585382
transform 1 0 72864 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_760
timestamp 1679585382
transform 1 0 73536 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_767
timestamp 1679585382
transform 1 0 74208 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_774
timestamp 1679585382
transform 1 0 74880 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_781
timestamp 1679585382
transform 1 0 75552 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_788
timestamp 1679585382
transform 1 0 76224 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_795
timestamp 1679585382
transform 1 0 76896 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_802
timestamp 1679585382
transform 1 0 77568 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_809
timestamp 1679585382
transform 1 0 78240 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_816
timestamp 1679585382
transform 1 0 78912 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_823
timestamp 1679585382
transform 1 0 79584 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_830
timestamp 1679585382
transform 1 0 80256 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_837
timestamp 1679585382
transform 1 0 80928 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_844
timestamp 1679585382
transform 1 0 81600 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_851
timestamp 1679585382
transform 1 0 82272 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_858
timestamp 1679585382
transform 1 0 82944 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_865
timestamp 1679585382
transform 1 0 83616 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_872
timestamp 1679585382
transform 1 0 84288 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_879
timestamp 1679585382
transform 1 0 84960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_886
timestamp 1679585382
transform 1 0 85632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_893
timestamp 1679585382
transform 1 0 86304 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_900
timestamp 1679585382
transform 1 0 86976 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_907
timestamp 1679585382
transform 1 0 87648 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_914
timestamp 1679585382
transform 1 0 88320 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_921
timestamp 1679585382
transform 1 0 88992 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_928
timestamp 1679585382
transform 1 0 89664 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_935
timestamp 1679585382
transform 1 0 90336 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_942
timestamp 1679585382
transform 1 0 91008 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_949
timestamp 1679585382
transform 1 0 91680 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_956
timestamp 1679585382
transform 1 0 92352 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_963
timestamp 1679585382
transform 1 0 93024 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_970
timestamp 1679585382
transform 1 0 93696 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_977
timestamp 1679585382
transform 1 0 94368 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_984
timestamp 1679585382
transform 1 0 95040 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_991
timestamp 1679585382
transform 1 0 95712 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_998
timestamp 1679585382
transform 1 0 96384 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1005
timestamp 1679585382
transform 1 0 97056 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1012
timestamp 1679585382
transform 1 0 97728 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1019
timestamp 1679585382
transform 1 0 98400 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_1026
timestamp 1677583704
transform 1 0 99072 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_1028
timestamp 1677583258
transform 1 0 99264 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_4
timestamp 1679585382
transform 1 0 960 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_11
timestamp 1679585382
transform 1 0 1632 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_18
timestamp 1679581501
transform 1 0 2304 0 -1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_53
timestamp 1679585382
transform 1 0 5664 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_60
timestamp 1679585382
transform 1 0 6336 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_67
timestamp 1677583704
transform 1 0 7008 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_69
timestamp 1677583258
transform 1 0 7200 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_79
timestamp 1679585382
transform 1 0 8160 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_86
timestamp 1679585382
transform 1 0 8832 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_93
timestamp 1679581501
transform 1 0 9504 0 -1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_106
timestamp 1679585382
transform 1 0 10752 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_113
timestamp 1679581501
transform 1 0 11424 0 -1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_144
timestamp 1679585382
transform 1 0 14400 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_151
timestamp 1679585382
transform 1 0 15072 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_158
timestamp 1677583258
transform 1 0 15744 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_186
timestamp 1677583704
transform 1 0 18432 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_188
timestamp 1677583258
transform 1 0 18624 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_202
timestamp 1679585382
transform 1 0 19968 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_209
timestamp 1679585382
transform 1 0 20640 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_216
timestamp 1679585382
transform 1 0 21312 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_223
timestamp 1679585382
transform 1 0 21984 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_230
timestamp 1679585382
transform 1 0 22656 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_237
timestamp 1679585382
transform 1 0 23328 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_244
timestamp 1679585382
transform 1 0 24000 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_251
timestamp 1679585382
transform 1 0 24672 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_276
timestamp 1679585382
transform 1 0 27072 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_283
timestamp 1679585382
transform 1 0 27744 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_290
timestamp 1679585382
transform 1 0 28416 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_297
timestamp 1679585382
transform 1 0 29088 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_304
timestamp 1679585382
transform 1 0 29760 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_311
timestamp 1679585382
transform 1 0 30432 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_318
timestamp 1679585382
transform 1 0 31104 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_325
timestamp 1679585382
transform 1 0 31776 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_332
timestamp 1679585382
transform 1 0 32448 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_339
timestamp 1679585382
transform 1 0 33120 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_346
timestamp 1679585382
transform 1 0 33792 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_353
timestamp 1679585382
transform 1 0 34464 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_360
timestamp 1679585382
transform 1 0 35136 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_367
timestamp 1679585382
transform 1 0 35808 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_374
timestamp 1679585382
transform 1 0 36480 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_381
timestamp 1679585382
transform 1 0 37152 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_388
timestamp 1679585382
transform 1 0 37824 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_395
timestamp 1677583704
transform 1 0 38496 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_428
timestamp 1679585382
transform 1 0 41664 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_435
timestamp 1679585382
transform 1 0 42336 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_442
timestamp 1679585382
transform 1 0 43008 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_449
timestamp 1679585382
transform 1 0 43680 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_456
timestamp 1679585382
transform 1 0 44352 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_463
timestamp 1679585382
transform 1 0 45024 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_470
timestamp 1679585382
transform 1 0 45696 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_477
timestamp 1679585382
transform 1 0 46368 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_501
timestamp 1679585382
transform 1 0 48672 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_508
timestamp 1679585382
transform 1 0 49344 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_515
timestamp 1679585382
transform 1 0 50016 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_522
timestamp 1679581501
transform 1 0 50688 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_526
timestamp 1677583704
transform 1 0 51072 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_541
timestamp 1677583704
transform 1 0 52512 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_543
timestamp 1677583258
transform 1 0 52704 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_549
timestamp 1679585382
transform 1 0 53280 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_556
timestamp 1679585382
transform 1 0 53952 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_563
timestamp 1677583704
transform 1 0 54624 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_592
timestamp 1679585382
transform 1 0 57408 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_599
timestamp 1679585382
transform 1 0 58080 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_606
timestamp 1679585382
transform 1 0 58752 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_613
timestamp 1679585382
transform 1 0 59424 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_620
timestamp 1679585382
transform 1 0 60096 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_627
timestamp 1679585382
transform 1 0 60768 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_634
timestamp 1679585382
transform 1 0 61440 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_641
timestamp 1679585382
transform 1 0 62112 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_648
timestamp 1679585382
transform 1 0 62784 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_655
timestamp 1679585382
transform 1 0 63456 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_662
timestamp 1679585382
transform 1 0 64128 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_669
timestamp 1679585382
transform 1 0 64800 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_676
timestamp 1679585382
transform 1 0 65472 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_683
timestamp 1679585382
transform 1 0 66144 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_690
timestamp 1679585382
transform 1 0 66816 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_697
timestamp 1679585382
transform 1 0 67488 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_704
timestamp 1679585382
transform 1 0 68160 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_711
timestamp 1679585382
transform 1 0 68832 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_718
timestamp 1679585382
transform 1 0 69504 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_725
timestamp 1679585382
transform 1 0 70176 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_732
timestamp 1679585382
transform 1 0 70848 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_739
timestamp 1679585382
transform 1 0 71520 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_746
timestamp 1679585382
transform 1 0 72192 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_753
timestamp 1679585382
transform 1 0 72864 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_760
timestamp 1679585382
transform 1 0 73536 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_767
timestamp 1679585382
transform 1 0 74208 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_774
timestamp 1679585382
transform 1 0 74880 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_781
timestamp 1679585382
transform 1 0 75552 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_788
timestamp 1679585382
transform 1 0 76224 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_795
timestamp 1679585382
transform 1 0 76896 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_802
timestamp 1679585382
transform 1 0 77568 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_809
timestamp 1679585382
transform 1 0 78240 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_816
timestamp 1679585382
transform 1 0 78912 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_823
timestamp 1679585382
transform 1 0 79584 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_830
timestamp 1679585382
transform 1 0 80256 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_837
timestamp 1679585382
transform 1 0 80928 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_844
timestamp 1679585382
transform 1 0 81600 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_851
timestamp 1679585382
transform 1 0 82272 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_858
timestamp 1679585382
transform 1 0 82944 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_865
timestamp 1679585382
transform 1 0 83616 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_872
timestamp 1679585382
transform 1 0 84288 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_879
timestamp 1679585382
transform 1 0 84960 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_886
timestamp 1679585382
transform 1 0 85632 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_893
timestamp 1679585382
transform 1 0 86304 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_900
timestamp 1679585382
transform 1 0 86976 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_907
timestamp 1679585382
transform 1 0 87648 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_914
timestamp 1679585382
transform 1 0 88320 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_921
timestamp 1679585382
transform 1 0 88992 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_928
timestamp 1679585382
transform 1 0 89664 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_935
timestamp 1679585382
transform 1 0 90336 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_942
timestamp 1679585382
transform 1 0 91008 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_949
timestamp 1679585382
transform 1 0 91680 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_956
timestamp 1679585382
transform 1 0 92352 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_963
timestamp 1679585382
transform 1 0 93024 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_970
timestamp 1679585382
transform 1 0 93696 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_977
timestamp 1679585382
transform 1 0 94368 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_984
timestamp 1679585382
transform 1 0 95040 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_991
timestamp 1679585382
transform 1 0 95712 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_998
timestamp 1679585382
transform 1 0 96384 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1005
timestamp 1679585382
transform 1 0 97056 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1012
timestamp 1679585382
transform 1 0 97728 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1019
timestamp 1679585382
transform 1 0 98400 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_1026
timestamp 1677583704
transform 1 0 99072 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_1028
timestamp 1677583258
transform 1 0 99264 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_4
timestamp 1679585382
transform 1 0 960 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_11
timestamp 1679585382
transform 1 0 1632 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_18
timestamp 1679585382
transform 1 0 2304 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_25
timestamp 1677583704
transform 1 0 2976 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_27
timestamp 1677583258
transform 1 0 3168 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_41
timestamp 1679585382
transform 1 0 4512 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_48
timestamp 1679585382
transform 1 0 5184 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_55
timestamp 1679585382
transform 1 0 5856 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_62
timestamp 1679585382
transform 1 0 6528 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_69
timestamp 1679585382
transform 1 0 7200 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_76
timestamp 1679585382
transform 1 0 7872 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_83
timestamp 1679585382
transform 1 0 8544 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_90
timestamp 1679585382
transform 1 0 9216 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_97
timestamp 1679585382
transform 1 0 9888 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_104
timestamp 1679585382
transform 1 0 10560 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_111
timestamp 1679585382
transform 1 0 11232 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_118
timestamp 1677583704
transform 1 0 11904 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_120
timestamp 1677583258
transform 1 0 12096 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_130
timestamp 1679585382
transform 1 0 13056 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_137
timestamp 1679585382
transform 1 0 13728 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_144
timestamp 1679585382
transform 1 0 14400 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_151
timestamp 1679585382
transform 1 0 15072 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_158
timestamp 1677583704
transform 1 0 15744 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_168
timestamp 1679585382
transform 1 0 16704 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_175
timestamp 1679585382
transform 1 0 17376 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_182
timestamp 1679585382
transform 1 0 18048 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_189
timestamp 1677583704
transform 1 0 18720 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_218
timestamp 1679585382
transform 1 0 21504 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_225
timestamp 1679585382
transform 1 0 22176 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_232
timestamp 1679585382
transform 1 0 22848 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_239
timestamp 1679585382
transform 1 0 23520 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_246
timestamp 1679585382
transform 1 0 24192 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_253
timestamp 1679581501
transform 1 0 24864 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_257
timestamp 1677583258
transform 1 0 25248 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_266
timestamp 1679585382
transform 1 0 26112 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_273
timestamp 1679585382
transform 1 0 26784 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_280
timestamp 1679585382
transform 1 0 27456 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_287
timestamp 1679585382
transform 1 0 28128 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_294
timestamp 1679585382
transform 1 0 28800 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_301
timestamp 1679585382
transform 1 0 29472 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_308
timestamp 1679585382
transform 1 0 30144 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_315
timestamp 1677583704
transform 1 0 30816 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_344
timestamp 1679585382
transform 1 0 33600 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_351
timestamp 1679585382
transform 1 0 34272 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_358
timestamp 1679585382
transform 1 0 34944 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_365
timestamp 1679585382
transform 1 0 35616 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_372
timestamp 1679585382
transform 1 0 36288 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_379
timestamp 1679585382
transform 1 0 36960 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_386
timestamp 1679585382
transform 1 0 37632 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_420
timestamp 1679585382
transform 1 0 40896 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_427
timestamp 1679585382
transform 1 0 41568 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_434
timestamp 1679585382
transform 1 0 42240 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_441
timestamp 1679585382
transform 1 0 42912 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_448
timestamp 1679581501
transform 1 0 43584 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_452
timestamp 1677583258
transform 1 0 43968 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_480
timestamp 1677583704
transform 1 0 46656 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_503
timestamp 1679585382
transform 1 0 48864 0 1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_12_510
timestamp 1677583258
transform 1 0 49536 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_519
timestamp 1679585382
transform 1 0 50400 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_526
timestamp 1679581501
transform 1 0 51072 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_570
timestamp 1677583704
transform 1 0 55296 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_576
timestamp 1679585382
transform 1 0 55872 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_592
timestamp 1679585382
transform 1 0 57408 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_599
timestamp 1679585382
transform 1 0 58080 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_606
timestamp 1679585382
transform 1 0 58752 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_613
timestamp 1679585382
transform 1 0 59424 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_620
timestamp 1679585382
transform 1 0 60096 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_627
timestamp 1679585382
transform 1 0 60768 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_634
timestamp 1679585382
transform 1 0 61440 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_641
timestamp 1679585382
transform 1 0 62112 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_648
timestamp 1679585382
transform 1 0 62784 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_655
timestamp 1679585382
transform 1 0 63456 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_662
timestamp 1679585382
transform 1 0 64128 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_669
timestamp 1679585382
transform 1 0 64800 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_676
timestamp 1679585382
transform 1 0 65472 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_683
timestamp 1679585382
transform 1 0 66144 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_690
timestamp 1679585382
transform 1 0 66816 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_697
timestamp 1679585382
transform 1 0 67488 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_704
timestamp 1679585382
transform 1 0 68160 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_711
timestamp 1679585382
transform 1 0 68832 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_718
timestamp 1679585382
transform 1 0 69504 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_725
timestamp 1679585382
transform 1 0 70176 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_732
timestamp 1679585382
transform 1 0 70848 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_739
timestamp 1679585382
transform 1 0 71520 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_746
timestamp 1679585382
transform 1 0 72192 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_753
timestamp 1679585382
transform 1 0 72864 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_760
timestamp 1679585382
transform 1 0 73536 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_767
timestamp 1679585382
transform 1 0 74208 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_774
timestamp 1679585382
transform 1 0 74880 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_781
timestamp 1679585382
transform 1 0 75552 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_788
timestamp 1679585382
transform 1 0 76224 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_795
timestamp 1679585382
transform 1 0 76896 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_802
timestamp 1679585382
transform 1 0 77568 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_809
timestamp 1679585382
transform 1 0 78240 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_816
timestamp 1679585382
transform 1 0 78912 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_823
timestamp 1679585382
transform 1 0 79584 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_830
timestamp 1679585382
transform 1 0 80256 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_837
timestamp 1679585382
transform 1 0 80928 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_844
timestamp 1679585382
transform 1 0 81600 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_851
timestamp 1679585382
transform 1 0 82272 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_858
timestamp 1679585382
transform 1 0 82944 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_865
timestamp 1679585382
transform 1 0 83616 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_872
timestamp 1679585382
transform 1 0 84288 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_879
timestamp 1679585382
transform 1 0 84960 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_886
timestamp 1679585382
transform 1 0 85632 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_893
timestamp 1679585382
transform 1 0 86304 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_900
timestamp 1679585382
transform 1 0 86976 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_907
timestamp 1679585382
transform 1 0 87648 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_914
timestamp 1679585382
transform 1 0 88320 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_921
timestamp 1679585382
transform 1 0 88992 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_928
timestamp 1679585382
transform 1 0 89664 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_935
timestamp 1679585382
transform 1 0 90336 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_942
timestamp 1679585382
transform 1 0 91008 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_949
timestamp 1679585382
transform 1 0 91680 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_956
timestamp 1679585382
transform 1 0 92352 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_963
timestamp 1679585382
transform 1 0 93024 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_970
timestamp 1679585382
transform 1 0 93696 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_977
timestamp 1679585382
transform 1 0 94368 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_984
timestamp 1679585382
transform 1 0 95040 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_991
timestamp 1679585382
transform 1 0 95712 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_998
timestamp 1679585382
transform 1 0 96384 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1005
timestamp 1679585382
transform 1 0 97056 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1012
timestamp 1679585382
transform 1 0 97728 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1019
timestamp 1679585382
transform 1 0 98400 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_1026
timestamp 1677583704
transform 1 0 99072 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_1028
timestamp 1677583258
transform 1 0 99264 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_4
timestamp 1679585382
transform 1 0 960 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_11
timestamp 1679585382
transform 1 0 1632 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_18
timestamp 1679585382
transform 1 0 2304 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_25
timestamp 1679585382
transform 1 0 2976 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_32
timestamp 1679585382
transform 1 0 3648 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_39
timestamp 1679585382
transform 1 0 4320 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_46
timestamp 1679585382
transform 1 0 4992 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_53
timestamp 1679585382
transform 1 0 5664 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_60
timestamp 1679585382
transform 1 0 6336 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_67
timestamp 1679585382
transform 1 0 7008 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_74
timestamp 1679585382
transform 1 0 7680 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_81
timestamp 1679585382
transform 1 0 8352 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_88
timestamp 1679585382
transform 1 0 9024 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_95
timestamp 1679585382
transform 1 0 9696 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_102
timestamp 1679585382
transform 1 0 10368 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_109
timestamp 1679585382
transform 1 0 11040 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_116
timestamp 1679585382
transform 1 0 11712 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_123
timestamp 1679585382
transform 1 0 12384 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_130
timestamp 1679585382
transform 1 0 13056 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_137
timestamp 1679585382
transform 1 0 13728 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_144
timestamp 1679585382
transform 1 0 14400 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_151
timestamp 1679585382
transform 1 0 15072 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_13_158
timestamp 1677583258
transform 1 0 15744 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_168
timestamp 1679585382
transform 1 0 16704 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_175
timestamp 1679585382
transform 1 0 17376 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_182
timestamp 1679585382
transform 1 0 18048 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_189
timestamp 1679585382
transform 1 0 18720 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_196
timestamp 1679585382
transform 1 0 19392 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_203
timestamp 1679585382
transform 1 0 20064 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_210
timestamp 1679585382
transform 1 0 20736 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_217
timestamp 1679585382
transform 1 0 21408 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_224
timestamp 1679585382
transform 1 0 22080 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_231
timestamp 1677583704
transform 1 0 22752 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_260
timestamp 1679585382
transform 1 0 25536 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_267
timestamp 1679585382
transform 1 0 26208 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_274
timestamp 1679585382
transform 1 0 26880 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_281
timestamp 1679585382
transform 1 0 27552 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_288
timestamp 1679585382
transform 1 0 28224 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_295
timestamp 1679585382
transform 1 0 28896 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_302
timestamp 1679585382
transform 1 0 29568 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_309
timestamp 1679585382
transform 1 0 30240 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_316
timestamp 1679585382
transform 1 0 30912 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_327
timestamp 1679585382
transform 1 0 31968 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_13_334
timestamp 1677583258
transform 1 0 32640 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_344
timestamp 1679585382
transform 1 0 33600 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_351
timestamp 1679585382
transform 1 0 34272 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_358
timestamp 1679585382
transform 1 0 34944 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_365
timestamp 1679581501
transform 1 0 35616 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_13_382
timestamp 1679585382
transform 1 0 37248 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_389
timestamp 1679585382
transform 1 0 37920 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_396
timestamp 1679585382
transform 1 0 38592 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_403
timestamp 1679581501
transform 1 0 39264 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_407
timestamp 1677583704
transform 1 0 39648 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_418
timestamp 1679585382
transform 1 0 40704 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_425
timestamp 1679585382
transform 1 0 41376 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_432
timestamp 1679585382
transform 1 0 42048 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_439
timestamp 1679585382
transform 1 0 42720 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_13_446
timestamp 1677583258
transform 1 0 43392 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_464
timestamp 1679585382
transform 1 0 45120 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_471
timestamp 1679585382
transform 1 0 45792 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_478
timestamp 1679585382
transform 1 0 46464 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_485
timestamp 1679585382
transform 1 0 47136 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_492
timestamp 1679585382
transform 1 0 47808 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_499
timestamp 1679585382
transform 1 0 48480 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_506
timestamp 1679585382
transform 1 0 49152 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_513
timestamp 1679585382
transform 1 0 49824 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_520
timestamp 1679585382
transform 1 0 50496 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_527
timestamp 1679585382
transform 1 0 51168 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_534
timestamp 1679585382
transform 1 0 51840 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_541
timestamp 1679585382
transform 1 0 52512 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_548
timestamp 1679581501
transform 1 0 53184 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_552
timestamp 1677583704
transform 1 0 53568 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_4  FILLER_13_558
timestamp 1679581501
transform 1 0 54144 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_562
timestamp 1677583258
transform 1 0 54528 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_572
timestamp 1677583704
transform 1 0 55488 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_578
timestamp 1679585382
transform 1 0 56064 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_585
timestamp 1679585382
transform 1 0 56736 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_592
timestamp 1679585382
transform 1 0 57408 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_599
timestamp 1679585382
transform 1 0 58080 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_606
timestamp 1679585382
transform 1 0 58752 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_613
timestamp 1679585382
transform 1 0 59424 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_620
timestamp 1679585382
transform 1 0 60096 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_627
timestamp 1679585382
transform 1 0 60768 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_634
timestamp 1679585382
transform 1 0 61440 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_641
timestamp 1679585382
transform 1 0 62112 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_648
timestamp 1679585382
transform 1 0 62784 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_655
timestamp 1679585382
transform 1 0 63456 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_662
timestamp 1679585382
transform 1 0 64128 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_669
timestamp 1679585382
transform 1 0 64800 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_676
timestamp 1679585382
transform 1 0 65472 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_683
timestamp 1679585382
transform 1 0 66144 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_690
timestamp 1679585382
transform 1 0 66816 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_697
timestamp 1679585382
transform 1 0 67488 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_704
timestamp 1679585382
transform 1 0 68160 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_711
timestamp 1679585382
transform 1 0 68832 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_718
timestamp 1679585382
transform 1 0 69504 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_725
timestamp 1679585382
transform 1 0 70176 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_732
timestamp 1679585382
transform 1 0 70848 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_739
timestamp 1679585382
transform 1 0 71520 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_746
timestamp 1679585382
transform 1 0 72192 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_753
timestamp 1679585382
transform 1 0 72864 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_760
timestamp 1679585382
transform 1 0 73536 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_767
timestamp 1679585382
transform 1 0 74208 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_774
timestamp 1679585382
transform 1 0 74880 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_781
timestamp 1679585382
transform 1 0 75552 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_788
timestamp 1679585382
transform 1 0 76224 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_795
timestamp 1679585382
transform 1 0 76896 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_802
timestamp 1679585382
transform 1 0 77568 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_809
timestamp 1679585382
transform 1 0 78240 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_816
timestamp 1679585382
transform 1 0 78912 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_823
timestamp 1679585382
transform 1 0 79584 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_830
timestamp 1679585382
transform 1 0 80256 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_837
timestamp 1679585382
transform 1 0 80928 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_844
timestamp 1679585382
transform 1 0 81600 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_851
timestamp 1679585382
transform 1 0 82272 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_858
timestamp 1679585382
transform 1 0 82944 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_865
timestamp 1679585382
transform 1 0 83616 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_872
timestamp 1679585382
transform 1 0 84288 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_879
timestamp 1679585382
transform 1 0 84960 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_886
timestamp 1679585382
transform 1 0 85632 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_893
timestamp 1679585382
transform 1 0 86304 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_900
timestamp 1679585382
transform 1 0 86976 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_907
timestamp 1679585382
transform 1 0 87648 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_914
timestamp 1679585382
transform 1 0 88320 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_921
timestamp 1679585382
transform 1 0 88992 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_928
timestamp 1679585382
transform 1 0 89664 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_935
timestamp 1679585382
transform 1 0 90336 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_942
timestamp 1679585382
transform 1 0 91008 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_949
timestamp 1679585382
transform 1 0 91680 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_956
timestamp 1679585382
transform 1 0 92352 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_963
timestamp 1679585382
transform 1 0 93024 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_970
timestamp 1679585382
transform 1 0 93696 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_977
timestamp 1679585382
transform 1 0 94368 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_984
timestamp 1679585382
transform 1 0 95040 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_991
timestamp 1679585382
transform 1 0 95712 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_998
timestamp 1679585382
transform 1 0 96384 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1005
timestamp 1679585382
transform 1 0 97056 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1012
timestamp 1679585382
transform 1 0 97728 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1019
timestamp 1679585382
transform 1 0 98400 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_1026
timestamp 1677583704
transform 1 0 99072 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_1028
timestamp 1677583258
transform 1 0 99264 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_4
timestamp 1679585382
transform 1 0 960 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_11
timestamp 1679585382
transform 1 0 1632 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_18
timestamp 1679585382
transform 1 0 2304 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_25
timestamp 1677583704
transform 1 0 2976 0 1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_14_31
timestamp 1677583704
transform 1 0 3552 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_33
timestamp 1677583258
transform 1 0 3744 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_55
timestamp 1679585382
transform 1 0 5856 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_62
timestamp 1679585382
transform 1 0 6528 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_69
timestamp 1679585382
transform 1 0 7200 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_76
timestamp 1679585382
transform 1 0 7872 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_83
timestamp 1679585382
transform 1 0 8544 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_90
timestamp 1679585382
transform 1 0 9216 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_97
timestamp 1679585382
transform 1 0 9888 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_104
timestamp 1679585382
transform 1 0 10560 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_111
timestamp 1679585382
transform 1 0 11232 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_118
timestamp 1679585382
transform 1 0 11904 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_125
timestamp 1679585382
transform 1 0 12576 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_132
timestamp 1679585382
transform 1 0 13248 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_139
timestamp 1679585382
transform 1 0 13920 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_146
timestamp 1679585382
transform 1 0 14592 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_153
timestamp 1679585382
transform 1 0 15264 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_169
timestamp 1677583704
transform 1 0 16800 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_171
timestamp 1677583258
transform 1 0 16992 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_176
timestamp 1679585382
transform 1 0 17472 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_183
timestamp 1679581501
transform 1 0 18144 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_187
timestamp 1677583704
transform 1 0 18528 0 1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_202
timestamp 1679585382
transform 1 0 19968 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_209
timestamp 1679585382
transform 1 0 20640 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_216
timestamp 1679585382
transform 1 0 21312 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_223
timestamp 1679585382
transform 1 0 21984 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_230
timestamp 1679585382
transform 1 0 22656 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_237
timestamp 1679585382
transform 1 0 23328 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_244
timestamp 1679585382
transform 1 0 24000 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_251
timestamp 1679585382
transform 1 0 24672 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_258
timestamp 1679585382
transform 1 0 25344 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_265
timestamp 1679585382
transform 1 0 26016 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_272
timestamp 1679585382
transform 1 0 26688 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_279
timestamp 1679585382
transform 1 0 27360 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_286
timestamp 1679585382
transform 1 0 28032 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_293
timestamp 1679585382
transform 1 0 28704 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_300
timestamp 1679585382
transform 1 0 29376 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_307
timestamp 1679585382
transform 1 0 30048 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_314
timestamp 1679581501
transform 1 0 30720 0 1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_14_349
timestamp 1679585382
transform 1 0 34080 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_356
timestamp 1679585382
transform 1 0 34752 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_363
timestamp 1679585382
transform 1 0 35424 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_370
timestamp 1679585382
transform 1 0 36096 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_377
timestamp 1679585382
transform 1 0 36768 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_384
timestamp 1679585382
transform 1 0 37440 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_391
timestamp 1679585382
transform 1 0 38112 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_398
timestamp 1679585382
transform 1 0 38784 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_405
timestamp 1679585382
transform 1 0 39456 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_412
timestamp 1679581501
transform 1 0 40128 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_416
timestamp 1677583258
transform 1 0 40512 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_426
timestamp 1679585382
transform 1 0 41472 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_433
timestamp 1679585382
transform 1 0 42144 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_440
timestamp 1679585382
transform 1 0 42816 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_447
timestamp 1679585382
transform 1 0 43488 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_454
timestamp 1679585382
transform 1 0 44160 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_461
timestamp 1679585382
transform 1 0 44832 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_468
timestamp 1679585382
transform 1 0 45504 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_475
timestamp 1679581501
transform 1 0 46176 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_479
timestamp 1677583704
transform 1 0 46560 0 1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_490
timestamp 1679585382
transform 1 0 47616 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_497
timestamp 1679585382
transform 1 0 48288 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_504
timestamp 1679585382
transform 1 0 48960 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_511
timestamp 1679585382
transform 1 0 49632 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_518
timestamp 1679585382
transform 1 0 50304 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_525
timestamp 1679585382
transform 1 0 50976 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_532
timestamp 1679585382
transform 1 0 51648 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_539
timestamp 1679585382
transform 1 0 52320 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_546
timestamp 1679585382
transform 1 0 52992 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_553
timestamp 1679585382
transform 1 0 53664 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_560
timestamp 1679585382
transform 1 0 54336 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_567
timestamp 1679585382
transform 1 0 55008 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_574
timestamp 1679585382
transform 1 0 55680 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_581
timestamp 1679585382
transform 1 0 56352 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_588
timestamp 1679585382
transform 1 0 57024 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_595
timestamp 1679585382
transform 1 0 57696 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_602
timestamp 1679585382
transform 1 0 58368 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_609
timestamp 1679585382
transform 1 0 59040 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_616
timestamp 1679585382
transform 1 0 59712 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_623
timestamp 1679585382
transform 1 0 60384 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_630
timestamp 1679585382
transform 1 0 61056 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_637
timestamp 1679585382
transform 1 0 61728 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_644
timestamp 1679585382
transform 1 0 62400 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_651
timestamp 1679585382
transform 1 0 63072 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_658
timestamp 1679585382
transform 1 0 63744 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_665
timestamp 1679585382
transform 1 0 64416 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_672
timestamp 1679585382
transform 1 0 65088 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_679
timestamp 1679585382
transform 1 0 65760 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_686
timestamp 1679585382
transform 1 0 66432 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_693
timestamp 1679585382
transform 1 0 67104 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_700
timestamp 1679585382
transform 1 0 67776 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_707
timestamp 1679585382
transform 1 0 68448 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_714
timestamp 1679585382
transform 1 0 69120 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_721
timestamp 1679585382
transform 1 0 69792 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_728
timestamp 1679585382
transform 1 0 70464 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_735
timestamp 1679585382
transform 1 0 71136 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_742
timestamp 1679585382
transform 1 0 71808 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_749
timestamp 1679585382
transform 1 0 72480 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_756
timestamp 1679585382
transform 1 0 73152 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_763
timestamp 1679585382
transform 1 0 73824 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_770
timestamp 1679585382
transform 1 0 74496 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_777
timestamp 1679585382
transform 1 0 75168 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_784
timestamp 1679585382
transform 1 0 75840 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_791
timestamp 1679585382
transform 1 0 76512 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_798
timestamp 1679585382
transform 1 0 77184 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_805
timestamp 1679585382
transform 1 0 77856 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_812
timestamp 1679585382
transform 1 0 78528 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_819
timestamp 1679585382
transform 1 0 79200 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_826
timestamp 1679585382
transform 1 0 79872 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_833
timestamp 1679585382
transform 1 0 80544 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_840
timestamp 1679585382
transform 1 0 81216 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_847
timestamp 1679585382
transform 1 0 81888 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_854
timestamp 1679585382
transform 1 0 82560 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_861
timestamp 1679585382
transform 1 0 83232 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_868
timestamp 1679585382
transform 1 0 83904 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_875
timestamp 1679585382
transform 1 0 84576 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_882
timestamp 1679585382
transform 1 0 85248 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_889
timestamp 1679585382
transform 1 0 85920 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_896
timestamp 1679585382
transform 1 0 86592 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_903
timestamp 1679585382
transform 1 0 87264 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_910
timestamp 1679585382
transform 1 0 87936 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_917
timestamp 1679585382
transform 1 0 88608 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_924
timestamp 1679585382
transform 1 0 89280 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_931
timestamp 1679585382
transform 1 0 89952 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_938
timestamp 1679585382
transform 1 0 90624 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_945
timestamp 1679585382
transform 1 0 91296 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_952
timestamp 1679585382
transform 1 0 91968 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_959
timestamp 1679585382
transform 1 0 92640 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_966
timestamp 1679585382
transform 1 0 93312 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_973
timestamp 1679585382
transform 1 0 93984 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_980
timestamp 1679585382
transform 1 0 94656 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_987
timestamp 1679585382
transform 1 0 95328 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_994
timestamp 1679585382
transform 1 0 96000 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1001
timestamp 1679585382
transform 1 0 96672 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1008
timestamp 1679585382
transform 1 0 97344 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1015
timestamp 1679585382
transform 1 0 98016 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1022
timestamp 1679585382
transform 1 0 98688 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_4
timestamp 1679585382
transform 1 0 960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_11
timestamp 1679581501
transform 1 0 1632 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_15
timestamp 1677583258
transform 1 0 2016 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_47
timestamp 1679585382
transform 1 0 5088 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_54
timestamp 1679581501
transform 1 0 5760 0 -1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_15_85
timestamp 1679585382
transform 1 0 8736 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_119
timestamp 1679585382
transform 1 0 12000 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_126
timestamp 1679585382
transform 1 0 12672 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_133
timestamp 1679585382
transform 1 0 13344 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_140
timestamp 1679585382
transform 1 0 14016 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_147
timestamp 1679585382
transform 1 0 14688 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_154
timestamp 1679585382
transform 1 0 15360 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_161
timestamp 1679585382
transform 1 0 16032 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_168
timestamp 1679585382
transform 1 0 16704 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_175
timestamp 1679585382
transform 1 0 17376 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_182
timestamp 1677583258
transform 1 0 18048 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_205
timestamp 1679585382
transform 1 0 20256 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_212
timestamp 1677583704
transform 1 0 20928 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_214
timestamp 1677583258
transform 1 0 21120 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_224
timestamp 1679585382
transform 1 0 22080 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_231
timestamp 1679585382
transform 1 0 22752 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_238
timestamp 1679585382
transform 1 0 23424 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_245
timestamp 1679585382
transform 1 0 24096 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_252
timestamp 1679585382
transform 1 0 24768 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_259
timestamp 1679585382
transform 1 0 25440 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_266
timestamp 1679585382
transform 1 0 26112 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_273
timestamp 1679585382
transform 1 0 26784 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_280
timestamp 1677583258
transform 1 0 27456 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_308
timestamp 1679585382
transform 1 0 30144 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_315
timestamp 1679585382
transform 1 0 30816 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_322
timestamp 1679581501
transform 1 0 31488 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_326
timestamp 1677583258
transform 1 0 31872 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_331
timestamp 1677583258
transform 1 0 32352 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_354
timestamp 1679585382
transform 1 0 34560 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_361
timestamp 1679585382
transform 1 0 35232 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_368
timestamp 1679585382
transform 1 0 35904 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_375
timestamp 1679585382
transform 1 0 36576 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_382
timestamp 1679585382
transform 1 0 37248 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_389
timestamp 1679585382
transform 1 0 37920 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_396
timestamp 1679585382
transform 1 0 38592 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_403
timestamp 1679585382
transform 1 0 39264 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_410
timestamp 1679585382
transform 1 0 39936 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_417
timestamp 1679585382
transform 1 0 40608 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_424
timestamp 1679585382
transform 1 0 41280 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_431
timestamp 1679585382
transform 1 0 41952 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_438
timestamp 1679585382
transform 1 0 42624 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_445
timestamp 1679585382
transform 1 0 43296 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_452
timestamp 1679585382
transform 1 0 43968 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_459
timestamp 1679585382
transform 1 0 44640 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_466
timestamp 1679585382
transform 1 0 45312 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_473
timestamp 1679585382
transform 1 0 45984 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_480
timestamp 1679585382
transform 1 0 46656 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_487
timestamp 1679585382
transform 1 0 47328 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_494
timestamp 1679585382
transform 1 0 48000 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_501
timestamp 1679585382
transform 1 0 48672 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_508
timestamp 1679585382
transform 1 0 49344 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_515
timestamp 1679585382
transform 1 0 50016 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_522
timestamp 1679585382
transform 1 0 50688 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_529
timestamp 1679585382
transform 1 0 51360 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_536
timestamp 1679585382
transform 1 0 52032 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_543
timestamp 1679585382
transform 1 0 52704 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_550
timestamp 1679585382
transform 1 0 53376 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_557
timestamp 1679585382
transform 1 0 54048 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_564
timestamp 1677583258
transform 1 0 54720 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_570
timestamp 1679585382
transform 1 0 55296 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_577
timestamp 1677583704
transform 1 0 55968 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_587
timestamp 1679585382
transform 1 0 56928 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_603
timestamp 1679585382
transform 1 0 58464 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_610
timestamp 1679585382
transform 1 0 59136 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_617
timestamp 1679585382
transform 1 0 59808 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_624
timestamp 1679585382
transform 1 0 60480 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_631
timestamp 1679585382
transform 1 0 61152 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_638
timestamp 1679585382
transform 1 0 61824 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_645
timestamp 1679585382
transform 1 0 62496 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_652
timestamp 1679585382
transform 1 0 63168 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_659
timestamp 1679585382
transform 1 0 63840 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_666
timestamp 1679585382
transform 1 0 64512 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_673
timestamp 1679585382
transform 1 0 65184 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_680
timestamp 1679585382
transform 1 0 65856 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_687
timestamp 1679585382
transform 1 0 66528 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_694
timestamp 1679585382
transform 1 0 67200 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_701
timestamp 1679585382
transform 1 0 67872 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_708
timestamp 1679585382
transform 1 0 68544 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_715
timestamp 1679585382
transform 1 0 69216 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_722
timestamp 1679585382
transform 1 0 69888 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_729
timestamp 1679585382
transform 1 0 70560 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_736
timestamp 1679585382
transform 1 0 71232 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_743
timestamp 1679585382
transform 1 0 71904 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_750
timestamp 1679585382
transform 1 0 72576 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_757
timestamp 1679585382
transform 1 0 73248 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_764
timestamp 1679585382
transform 1 0 73920 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_771
timestamp 1679585382
transform 1 0 74592 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_778
timestamp 1679585382
transform 1 0 75264 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_785
timestamp 1679585382
transform 1 0 75936 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_792
timestamp 1679585382
transform 1 0 76608 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_799
timestamp 1679585382
transform 1 0 77280 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_806
timestamp 1679585382
transform 1 0 77952 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_813
timestamp 1679585382
transform 1 0 78624 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_820
timestamp 1679585382
transform 1 0 79296 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_827
timestamp 1679585382
transform 1 0 79968 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_834
timestamp 1679585382
transform 1 0 80640 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_841
timestamp 1679585382
transform 1 0 81312 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_848
timestamp 1679585382
transform 1 0 81984 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_855
timestamp 1679585382
transform 1 0 82656 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_862
timestamp 1679585382
transform 1 0 83328 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_869
timestamp 1679585382
transform 1 0 84000 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_876
timestamp 1679585382
transform 1 0 84672 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_883
timestamp 1679585382
transform 1 0 85344 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_890
timestamp 1679585382
transform 1 0 86016 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_897
timestamp 1679585382
transform 1 0 86688 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_904
timestamp 1679585382
transform 1 0 87360 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_911
timestamp 1679585382
transform 1 0 88032 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_918
timestamp 1679585382
transform 1 0 88704 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_925
timestamp 1679585382
transform 1 0 89376 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_932
timestamp 1679585382
transform 1 0 90048 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_939
timestamp 1679585382
transform 1 0 90720 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_946
timestamp 1679585382
transform 1 0 91392 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_953
timestamp 1679585382
transform 1 0 92064 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_960
timestamp 1679585382
transform 1 0 92736 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_967
timestamp 1679585382
transform 1 0 93408 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_974
timestamp 1679585382
transform 1 0 94080 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_981
timestamp 1679585382
transform 1 0 94752 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_988
timestamp 1679585382
transform 1 0 95424 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_995
timestamp 1679585382
transform 1 0 96096 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1002
timestamp 1679585382
transform 1 0 96768 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1009
timestamp 1679585382
transform 1 0 97440 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1016
timestamp 1679585382
transform 1 0 98112 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_1023
timestamp 1679581501
transform 1 0 98784 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_1027
timestamp 1677583704
transform 1 0 99168 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_4
timestamp 1679585382
transform 1 0 960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_11
timestamp 1679581501
transform 1 0 1632 0 1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_16_42
timestamp 1679585382
transform 1 0 4608 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_49
timestamp 1679585382
transform 1 0 5280 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_56
timestamp 1679585382
transform 1 0 5952 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_63
timestamp 1679581501
transform 1 0 6624 0 1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_16_80
timestamp 1679585382
transform 1 0 8256 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_87
timestamp 1677583704
transform 1 0 8928 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_98
timestamp 1679585382
transform 1 0 9984 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_118
timestamp 1677583704
transform 1 0 11904 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_120
timestamp 1677583258
transform 1 0 12096 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_148
timestamp 1679585382
transform 1 0 14784 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_155
timestamp 1679585382
transform 1 0 15456 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_162
timestamp 1679585382
transform 1 0 16128 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_169
timestamp 1679585382
transform 1 0 16800 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_176
timestamp 1679585382
transform 1 0 17472 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_183
timestamp 1677583704
transform 1 0 18144 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_185
timestamp 1677583258
transform 1 0 18336 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_194
timestamp 1677583258
transform 1 0 19200 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_208
timestamp 1679585382
transform 1 0 20544 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_215
timestamp 1679585382
transform 1 0 21216 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_222
timestamp 1679585382
transform 1 0 21888 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_269
timestamp 1679585382
transform 1 0 26400 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_276
timestamp 1679585382
transform 1 0 27072 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_283
timestamp 1679581501
transform 1 0 27744 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_287
timestamp 1677583704
transform 1 0 28128 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_293
timestamp 1677583258
transform 1 0 28704 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_298
timestamp 1677583704
transform 1 0 29184 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_317
timestamp 1679585382
transform 1 0 31008 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_324
timestamp 1679581501
transform 1 0 31680 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_328
timestamp 1677583258
transform 1 0 32064 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_334
timestamp 1679585382
transform 1 0 32640 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_341
timestamp 1679585382
transform 1 0 33312 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_348
timestamp 1679585382
transform 1 0 33984 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_355
timestamp 1679585382
transform 1 0 34656 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_362
timestamp 1679585382
transform 1 0 35328 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_369
timestamp 1679585382
transform 1 0 36000 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_376
timestamp 1679581501
transform 1 0 36672 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_380
timestamp 1677583258
transform 1 0 37056 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_416
timestamp 1679585382
transform 1 0 40512 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_423
timestamp 1677583704
transform 1 0 41184 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_452
timestamp 1679585382
transform 1 0 43968 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_459
timestamp 1679585382
transform 1 0 44640 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_466
timestamp 1679581501
transform 1 0 45312 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_470
timestamp 1677583704
transform 1 0 45696 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_499
timestamp 1679585382
transform 1 0 48480 0 1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_16_506
timestamp 1677583258
transform 1 0 49152 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_520
timestamp 1679585382
transform 1 0 50496 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_527
timestamp 1679581501
transform 1 0 51168 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_531
timestamp 1677583704
transform 1 0 51552 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_560
timestamp 1677583258
transform 1 0 54336 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_574
timestamp 1679581501
transform 1 0 55680 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_578
timestamp 1677583258
transform 1 0 56064 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_606
timestamp 1679585382
transform 1 0 58752 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_613
timestamp 1679585382
transform 1 0 59424 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_620
timestamp 1679585382
transform 1 0 60096 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_627
timestamp 1679585382
transform 1 0 60768 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_634
timestamp 1679585382
transform 1 0 61440 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_641
timestamp 1679585382
transform 1 0 62112 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_648
timestamp 1679585382
transform 1 0 62784 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_655
timestamp 1679585382
transform 1 0 63456 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_662
timestamp 1679585382
transform 1 0 64128 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_669
timestamp 1679585382
transform 1 0 64800 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_676
timestamp 1679585382
transform 1 0 65472 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_683
timestamp 1679585382
transform 1 0 66144 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_690
timestamp 1679585382
transform 1 0 66816 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_697
timestamp 1679585382
transform 1 0 67488 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_704
timestamp 1679585382
transform 1 0 68160 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_711
timestamp 1679585382
transform 1 0 68832 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_718
timestamp 1679585382
transform 1 0 69504 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_725
timestamp 1679585382
transform 1 0 70176 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_732
timestamp 1679585382
transform 1 0 70848 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_739
timestamp 1679585382
transform 1 0 71520 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_746
timestamp 1679585382
transform 1 0 72192 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_753
timestamp 1679585382
transform 1 0 72864 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_760
timestamp 1679585382
transform 1 0 73536 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_767
timestamp 1679585382
transform 1 0 74208 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_774
timestamp 1679585382
transform 1 0 74880 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_781
timestamp 1679585382
transform 1 0 75552 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_788
timestamp 1679585382
transform 1 0 76224 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_795
timestamp 1679585382
transform 1 0 76896 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_802
timestamp 1679585382
transform 1 0 77568 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_809
timestamp 1679585382
transform 1 0 78240 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_816
timestamp 1679585382
transform 1 0 78912 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_823
timestamp 1679585382
transform 1 0 79584 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_830
timestamp 1679585382
transform 1 0 80256 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_837
timestamp 1679585382
transform 1 0 80928 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_844
timestamp 1679585382
transform 1 0 81600 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_851
timestamp 1679585382
transform 1 0 82272 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_858
timestamp 1679585382
transform 1 0 82944 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_865
timestamp 1679585382
transform 1 0 83616 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_872
timestamp 1679585382
transform 1 0 84288 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_879
timestamp 1679585382
transform 1 0 84960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_886
timestamp 1679585382
transform 1 0 85632 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_893
timestamp 1679585382
transform 1 0 86304 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_900
timestamp 1679585382
transform 1 0 86976 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_907
timestamp 1679585382
transform 1 0 87648 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_914
timestamp 1679585382
transform 1 0 88320 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_921
timestamp 1679585382
transform 1 0 88992 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_928
timestamp 1679585382
transform 1 0 89664 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_935
timestamp 1679585382
transform 1 0 90336 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_942
timestamp 1679585382
transform 1 0 91008 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_949
timestamp 1679585382
transform 1 0 91680 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_956
timestamp 1679585382
transform 1 0 92352 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_963
timestamp 1679585382
transform 1 0 93024 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_970
timestamp 1679585382
transform 1 0 93696 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_977
timestamp 1679585382
transform 1 0 94368 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_984
timestamp 1679585382
transform 1 0 95040 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_991
timestamp 1679585382
transform 1 0 95712 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_998
timestamp 1679585382
transform 1 0 96384 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1005
timestamp 1679585382
transform 1 0 97056 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1012
timestamp 1679585382
transform 1 0 97728 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1019
timestamp 1679585382
transform 1 0 98400 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_1026
timestamp 1677583704
transform 1 0 99072 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_1028
timestamp 1677583258
transform 1 0 99264 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_0
timestamp 1679585382
transform 1 0 576 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_7
timestamp 1679585382
transform 1 0 1248 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_14
timestamp 1679585382
transform 1 0 1920 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_21
timestamp 1679585382
transform 1 0 2592 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_28
timestamp 1677583704
transform 1 0 3264 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_39
timestamp 1679585382
transform 1 0 4320 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_46
timestamp 1679585382
transform 1 0 4992 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_53
timestamp 1679585382
transform 1 0 5664 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_60
timestamp 1679585382
transform 1 0 6336 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_67
timestamp 1679585382
transform 1 0 7008 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_74
timestamp 1679585382
transform 1 0 7680 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_81
timestamp 1679585382
transform 1 0 8352 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_88
timestamp 1679585382
transform 1 0 9024 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_95
timestamp 1679585382
transform 1 0 9696 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_102
timestamp 1679585382
transform 1 0 10368 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_109
timestamp 1679585382
transform 1 0 11040 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_116
timestamp 1679581501
transform 1 0 11712 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_17_129
timestamp 1677583258
transform 1 0 12960 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_143
timestamp 1679585382
transform 1 0 14304 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_150
timestamp 1677583258
transform 1 0 14976 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_200
timestamp 1679585382
transform 1 0 19776 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_207
timestamp 1679585382
transform 1 0 20448 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_214
timestamp 1679585382
transform 1 0 21120 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_221
timestamp 1679585382
transform 1 0 21792 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_228
timestamp 1679585382
transform 1 0 22464 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_235
timestamp 1679585382
transform 1 0 23136 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_242
timestamp 1679585382
transform 1 0 23808 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_249
timestamp 1679581501
transform 1 0 24480 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_253
timestamp 1677583704
transform 1 0 24864 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_17_259
timestamp 1679581501
transform 1 0 25440 0 -1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_17_272
timestamp 1679585382
transform 1 0 26688 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_279
timestamp 1679585382
transform 1 0 27360 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_286
timestamp 1679585382
transform 1 0 28032 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_293
timestamp 1679585382
transform 1 0 28704 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_300
timestamp 1679585382
transform 1 0 29376 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_307
timestamp 1679585382
transform 1 0 30048 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_314
timestamp 1679585382
transform 1 0 30720 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_321
timestamp 1679585382
transform 1 0 31392 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_328
timestamp 1679585382
transform 1 0 32064 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_335
timestamp 1679585382
transform 1 0 32736 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_342
timestamp 1677583704
transform 1 0 33408 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_371
timestamp 1679585382
transform 1 0 36192 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_387
timestamp 1679585382
transform 1 0 37728 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_394
timestamp 1679581501
transform 1 0 38400 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_411
timestamp 1677583704
transform 1 0 40032 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_17_422
timestamp 1677583704
transform 1 0 41088 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_424
timestamp 1677583258
transform 1 0 41280 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_434
timestamp 1679585382
transform 1 0 42240 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_441
timestamp 1679585382
transform 1 0 42912 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_448
timestamp 1679585382
transform 1 0 43584 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_455
timestamp 1679585382
transform 1 0 44256 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_462
timestamp 1679585382
transform 1 0 44928 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_469
timestamp 1679585382
transform 1 0 45600 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_476
timestamp 1679585382
transform 1 0 46272 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_483
timestamp 1679585382
transform 1 0 46944 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_490
timestamp 1677583704
transform 1 0 47616 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_492
timestamp 1677583258
transform 1 0 47808 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_17_529
timestamp 1679581501
transform 1 0 51360 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_533
timestamp 1677583704
transform 1 0 51744 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_552
timestamp 1679585382
transform 1 0 53568 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_559
timestamp 1677583704
transform 1 0 54240 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_564
timestamp 1679585382
transform 1 0 54720 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_579
timestamp 1677583258
transform 1 0 56160 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_607
timestamp 1679585382
transform 1 0 58848 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_614
timestamp 1679585382
transform 1 0 59520 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_621
timestamp 1679585382
transform 1 0 60192 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_628
timestamp 1679585382
transform 1 0 60864 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_635
timestamp 1679585382
transform 1 0 61536 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_642
timestamp 1679585382
transform 1 0 62208 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_649
timestamp 1679585382
transform 1 0 62880 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_656
timestamp 1679585382
transform 1 0 63552 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_663
timestamp 1679585382
transform 1 0 64224 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_670
timestamp 1679585382
transform 1 0 64896 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_677
timestamp 1679585382
transform 1 0 65568 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_684
timestamp 1679585382
transform 1 0 66240 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_691
timestamp 1679585382
transform 1 0 66912 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_698
timestamp 1679585382
transform 1 0 67584 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_705
timestamp 1679585382
transform 1 0 68256 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_712
timestamp 1679585382
transform 1 0 68928 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_719
timestamp 1679585382
transform 1 0 69600 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_726
timestamp 1679585382
transform 1 0 70272 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_733
timestamp 1679585382
transform 1 0 70944 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_740
timestamp 1679585382
transform 1 0 71616 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_747
timestamp 1679585382
transform 1 0 72288 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_754
timestamp 1679585382
transform 1 0 72960 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_761
timestamp 1679585382
transform 1 0 73632 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_768
timestamp 1679585382
transform 1 0 74304 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_775
timestamp 1679585382
transform 1 0 74976 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_782
timestamp 1679585382
transform 1 0 75648 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_789
timestamp 1679585382
transform 1 0 76320 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_796
timestamp 1679585382
transform 1 0 76992 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_803
timestamp 1679585382
transform 1 0 77664 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_810
timestamp 1679585382
transform 1 0 78336 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_817
timestamp 1679585382
transform 1 0 79008 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_824
timestamp 1679585382
transform 1 0 79680 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_831
timestamp 1679585382
transform 1 0 80352 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_838
timestamp 1679585382
transform 1 0 81024 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_845
timestamp 1679585382
transform 1 0 81696 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_852
timestamp 1679585382
transform 1 0 82368 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_859
timestamp 1679585382
transform 1 0 83040 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_866
timestamp 1679585382
transform 1 0 83712 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_873
timestamp 1679585382
transform 1 0 84384 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_880
timestamp 1679585382
transform 1 0 85056 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_887
timestamp 1679585382
transform 1 0 85728 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_894
timestamp 1679585382
transform 1 0 86400 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_901
timestamp 1679585382
transform 1 0 87072 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_908
timestamp 1679585382
transform 1 0 87744 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_915
timestamp 1679585382
transform 1 0 88416 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_922
timestamp 1679585382
transform 1 0 89088 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_929
timestamp 1679585382
transform 1 0 89760 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_936
timestamp 1679585382
transform 1 0 90432 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_943
timestamp 1679585382
transform 1 0 91104 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_950
timestamp 1679585382
transform 1 0 91776 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_957
timestamp 1679585382
transform 1 0 92448 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_964
timestamp 1679585382
transform 1 0 93120 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_971
timestamp 1679585382
transform 1 0 93792 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_978
timestamp 1679585382
transform 1 0 94464 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_985
timestamp 1679585382
transform 1 0 95136 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_992
timestamp 1679585382
transform 1 0 95808 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_999
timestamp 1679585382
transform 1 0 96480 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1006
timestamp 1679585382
transform 1 0 97152 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1013
timestamp 1679585382
transform 1 0 97824 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1020
timestamp 1679585382
transform 1 0 98496 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_1027
timestamp 1677583704
transform 1 0 99168 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_4
timestamp 1679585382
transform 1 0 960 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_11
timestamp 1679585382
transform 1 0 1632 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_18
timestamp 1679585382
transform 1 0 2304 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_25
timestamp 1679585382
transform 1 0 2976 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_32
timestamp 1679585382
transform 1 0 3648 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_39
timestamp 1679585382
transform 1 0 4320 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_46
timestamp 1679585382
transform 1 0 4992 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_53
timestamp 1679585382
transform 1 0 5664 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_60
timestamp 1679585382
transform 1 0 6336 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_67
timestamp 1679585382
transform 1 0 7008 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_74
timestamp 1679585382
transform 1 0 7680 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_81
timestamp 1679581501
transform 1 0 8352 0 1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_18_98
timestamp 1679585382
transform 1 0 9984 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_105
timestamp 1679585382
transform 1 0 10656 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_112
timestamp 1679585382
transform 1 0 11328 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_119
timestamp 1679585382
transform 1 0 12000 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_126
timestamp 1679585382
transform 1 0 12672 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_133
timestamp 1679585382
transform 1 0 13344 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_140
timestamp 1679585382
transform 1 0 14016 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_147
timestamp 1679585382
transform 1 0 14688 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_154
timestamp 1679585382
transform 1 0 15360 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_161
timestamp 1679581501
transform 1 0 16032 0 1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_18_174
timestamp 1679585382
transform 1 0 17280 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_181
timestamp 1679585382
transform 1 0 17952 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_188
timestamp 1679585382
transform 1 0 18624 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_195
timestamp 1679585382
transform 1 0 19296 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_202
timestamp 1679585382
transform 1 0 19968 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_209
timestamp 1679585382
transform 1 0 20640 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_216
timestamp 1677583258
transform 1 0 21312 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_243
timestamp 1679585382
transform 1 0 23904 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_250
timestamp 1679585382
transform 1 0 24576 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_257
timestamp 1679585382
transform 1 0 25248 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_264
timestamp 1679585382
transform 1 0 25920 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_271
timestamp 1679585382
transform 1 0 26592 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_278
timestamp 1679585382
transform 1 0 27264 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_285
timestamp 1679585382
transform 1 0 27936 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_292
timestamp 1679585382
transform 1 0 28608 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_299
timestamp 1679585382
transform 1 0 29280 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_306
timestamp 1679585382
transform 1 0 29952 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_313
timestamp 1679585382
transform 1 0 30624 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_320
timestamp 1679585382
transform 1 0 31296 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_327
timestamp 1679585382
transform 1 0 31968 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_334
timestamp 1679585382
transform 1 0 32640 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_341
timestamp 1679585382
transform 1 0 33312 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_348
timestamp 1679585382
transform 1 0 33984 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_355
timestamp 1679585382
transform 1 0 34656 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_362
timestamp 1679581501
transform 1 0 35328 0 1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_18_366
timestamp 1677583704
transform 1 0 35712 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_376
timestamp 1679585382
transform 1 0 36672 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_383
timestamp 1679585382
transform 1 0 37344 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_390
timestamp 1679585382
transform 1 0 38016 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_397
timestamp 1679585382
transform 1 0 38688 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_404
timestamp 1679585382
transform 1 0 39360 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_411
timestamp 1679585382
transform 1 0 40032 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_422
timestamp 1677583258
transform 1 0 41088 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_431
timestamp 1679585382
transform 1 0 41952 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_438
timestamp 1679585382
transform 1 0 42624 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_445
timestamp 1679585382
transform 1 0 43296 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_452
timestamp 1679585382
transform 1 0 43968 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_459
timestamp 1677583704
transform 1 0 44640 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_461
timestamp 1677583258
transform 1 0 44832 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_475
timestamp 1677583704
transform 1 0 46176 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_477
timestamp 1677583258
transform 1 0 46368 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_491
timestamp 1679585382
transform 1 0 47712 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_498
timestamp 1679585382
transform 1 0 48384 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_505
timestamp 1679585382
transform 1 0 49056 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_512
timestamp 1679585382
transform 1 0 49728 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_519
timestamp 1679585382
transform 1 0 50400 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_526
timestamp 1677583258
transform 1 0 51072 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_540
timestamp 1677583258
transform 1 0 52416 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_549
timestamp 1679585382
transform 1 0 53280 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_556
timestamp 1679585382
transform 1 0 53952 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_563
timestamp 1679585382
transform 1 0 54624 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_570
timestamp 1679585382
transform 1 0 55296 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_577
timestamp 1679585382
transform 1 0 55968 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_584
timestamp 1677583258
transform 1 0 56640 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_589
timestamp 1679585382
transform 1 0 57120 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_596
timestamp 1677583258
transform 1 0 57792 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_606
timestamp 1679585382
transform 1 0 58752 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_613
timestamp 1679585382
transform 1 0 59424 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_620
timestamp 1679585382
transform 1 0 60096 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_627
timestamp 1679585382
transform 1 0 60768 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_634
timestamp 1679585382
transform 1 0 61440 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_641
timestamp 1679585382
transform 1 0 62112 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_648
timestamp 1679585382
transform 1 0 62784 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_655
timestamp 1679585382
transform 1 0 63456 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_662
timestamp 1679585382
transform 1 0 64128 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_669
timestamp 1679585382
transform 1 0 64800 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_676
timestamp 1679585382
transform 1 0 65472 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_683
timestamp 1679585382
transform 1 0 66144 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_690
timestamp 1679585382
transform 1 0 66816 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_697
timestamp 1679585382
transform 1 0 67488 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_704
timestamp 1679585382
transform 1 0 68160 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_711
timestamp 1679585382
transform 1 0 68832 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_718
timestamp 1679585382
transform 1 0 69504 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_725
timestamp 1679585382
transform 1 0 70176 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_732
timestamp 1679585382
transform 1 0 70848 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_739
timestamp 1679585382
transform 1 0 71520 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_746
timestamp 1679585382
transform 1 0 72192 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_753
timestamp 1679585382
transform 1 0 72864 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_760
timestamp 1679585382
transform 1 0 73536 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_767
timestamp 1679585382
transform 1 0 74208 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_774
timestamp 1679585382
transform 1 0 74880 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_781
timestamp 1679585382
transform 1 0 75552 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_788
timestamp 1679585382
transform 1 0 76224 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_795
timestamp 1679585382
transform 1 0 76896 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_802
timestamp 1679585382
transform 1 0 77568 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_809
timestamp 1679585382
transform 1 0 78240 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_816
timestamp 1679585382
transform 1 0 78912 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_823
timestamp 1679585382
transform 1 0 79584 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_830
timestamp 1679585382
transform 1 0 80256 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_837
timestamp 1679585382
transform 1 0 80928 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_844
timestamp 1679585382
transform 1 0 81600 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_851
timestamp 1679585382
transform 1 0 82272 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_858
timestamp 1679585382
transform 1 0 82944 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_865
timestamp 1679585382
transform 1 0 83616 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_872
timestamp 1679585382
transform 1 0 84288 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_879
timestamp 1679585382
transform 1 0 84960 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_886
timestamp 1679585382
transform 1 0 85632 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_893
timestamp 1679585382
transform 1 0 86304 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_900
timestamp 1679585382
transform 1 0 86976 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_907
timestamp 1679585382
transform 1 0 87648 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_914
timestamp 1679585382
transform 1 0 88320 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_921
timestamp 1679585382
transform 1 0 88992 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_928
timestamp 1679585382
transform 1 0 89664 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_935
timestamp 1679585382
transform 1 0 90336 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_942
timestamp 1679585382
transform 1 0 91008 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_949
timestamp 1679585382
transform 1 0 91680 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_956
timestamp 1679585382
transform 1 0 92352 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_963
timestamp 1679585382
transform 1 0 93024 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_970
timestamp 1679585382
transform 1 0 93696 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_977
timestamp 1679585382
transform 1 0 94368 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_984
timestamp 1679585382
transform 1 0 95040 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_991
timestamp 1679585382
transform 1 0 95712 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_998
timestamp 1679585382
transform 1 0 96384 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1005
timestamp 1679585382
transform 1 0 97056 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1012
timestamp 1679585382
transform 1 0 97728 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1019
timestamp 1679585382
transform 1 0 98400 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_1026
timestamp 1677583704
transform 1 0 99072 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_1028
timestamp 1677583258
transform 1 0 99264 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_4
timestamp 1679585382
transform 1 0 960 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_11
timestamp 1679585382
transform 1 0 1632 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_18
timestamp 1679585382
transform 1 0 2304 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_25
timestamp 1679585382
transform 1 0 2976 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_32
timestamp 1679585382
transform 1 0 3648 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_39
timestamp 1679585382
transform 1 0 4320 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_46
timestamp 1679585382
transform 1 0 4992 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_53
timestamp 1679585382
transform 1 0 5664 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_60
timestamp 1679585382
transform 1 0 6336 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_67
timestamp 1679585382
transform 1 0 7008 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_74
timestamp 1679585382
transform 1 0 7680 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_81
timestamp 1679585382
transform 1 0 8352 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_88
timestamp 1679585382
transform 1 0 9024 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_95
timestamp 1679585382
transform 1 0 9696 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_102
timestamp 1679585382
transform 1 0 10368 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_109
timestamp 1679585382
transform 1 0 11040 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_116
timestamp 1679585382
transform 1 0 11712 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_123
timestamp 1679585382
transform 1 0 12384 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_130
timestamp 1679585382
transform 1 0 13056 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_137
timestamp 1679585382
transform 1 0 13728 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_144
timestamp 1679585382
transform 1 0 14400 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_151
timestamp 1679585382
transform 1 0 15072 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_158
timestamp 1679585382
transform 1 0 15744 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_165
timestamp 1679585382
transform 1 0 16416 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_172
timestamp 1679585382
transform 1 0 17088 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_179
timestamp 1679585382
transform 1 0 17760 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_186
timestamp 1679585382
transform 1 0 18432 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_193
timestamp 1679585382
transform 1 0 19104 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_200
timestamp 1679585382
transform 1 0 19776 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_207
timestamp 1679585382
transform 1 0 20448 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_214
timestamp 1679585382
transform 1 0 21120 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_221
timestamp 1679585382
transform 1 0 21792 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_228
timestamp 1679585382
transform 1 0 22464 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_235
timestamp 1679585382
transform 1 0 23136 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_242
timestamp 1679585382
transform 1 0 23808 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_249
timestamp 1679585382
transform 1 0 24480 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_256
timestamp 1679585382
transform 1 0 25152 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_263
timestamp 1679585382
transform 1 0 25824 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_270
timestamp 1679585382
transform 1 0 26496 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_277
timestamp 1679585382
transform 1 0 27168 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_284
timestamp 1679585382
transform 1 0 27840 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_291
timestamp 1679585382
transform 1 0 28512 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_298
timestamp 1679585382
transform 1 0 29184 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_305
timestamp 1679585382
transform 1 0 29856 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_339
timestamp 1679585382
transform 1 0 33120 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_346
timestamp 1679585382
transform 1 0 33792 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_353
timestamp 1679585382
transform 1 0 34464 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_360
timestamp 1679581501
transform 1 0 35136 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_364
timestamp 1677583258
transform 1 0 35520 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_378
timestamp 1679585382
transform 1 0 36864 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_385
timestamp 1679585382
transform 1 0 37536 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_392
timestamp 1679585382
transform 1 0 38208 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_399
timestamp 1679585382
transform 1 0 38880 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_406
timestamp 1679585382
transform 1 0 39552 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_413
timestamp 1679581501
transform 1 0 40224 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_417
timestamp 1677583704
transform 1 0 40608 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_441
timestamp 1679585382
transform 1 0 42912 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_448
timestamp 1679585382
transform 1 0 43584 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_455
timestamp 1679585382
transform 1 0 44256 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_462
timestamp 1679585382
transform 1 0 44928 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_469
timestamp 1679585382
transform 1 0 45600 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_476
timestamp 1679585382
transform 1 0 46272 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_483
timestamp 1679585382
transform 1 0 46944 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_490
timestamp 1679585382
transform 1 0 47616 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_497
timestamp 1679585382
transform 1 0 48288 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_504
timestamp 1677583704
transform 1 0 48960 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_533
timestamp 1677583704
transform 1 0 51744 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_535
timestamp 1677583258
transform 1 0 51936 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_545
timestamp 1679585382
transform 1 0 52896 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_552
timestamp 1679585382
transform 1 0 53568 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_559
timestamp 1679585382
transform 1 0 54240 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_566
timestamp 1679585382
transform 1 0 54912 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_573
timestamp 1679585382
transform 1 0 55584 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_580
timestamp 1679585382
transform 1 0 56256 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_587
timestamp 1679585382
transform 1 0 56928 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_594
timestamp 1679585382
transform 1 0 57600 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_601
timestamp 1679585382
transform 1 0 58272 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_608
timestamp 1679585382
transform 1 0 58944 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_615
timestamp 1679585382
transform 1 0 59616 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_622
timestamp 1679585382
transform 1 0 60288 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_629
timestamp 1679585382
transform 1 0 60960 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_636
timestamp 1679585382
transform 1 0 61632 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_643
timestamp 1679585382
transform 1 0 62304 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_650
timestamp 1679585382
transform 1 0 62976 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_657
timestamp 1679585382
transform 1 0 63648 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_664
timestamp 1679585382
transform 1 0 64320 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_671
timestamp 1679585382
transform 1 0 64992 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_678
timestamp 1679585382
transform 1 0 65664 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_685
timestamp 1679585382
transform 1 0 66336 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_692
timestamp 1679585382
transform 1 0 67008 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_699
timestamp 1679585382
transform 1 0 67680 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_706
timestamp 1679585382
transform 1 0 68352 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_713
timestamp 1679585382
transform 1 0 69024 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_720
timestamp 1679585382
transform 1 0 69696 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_727
timestamp 1679585382
transform 1 0 70368 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_734
timestamp 1679585382
transform 1 0 71040 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_741
timestamp 1679585382
transform 1 0 71712 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_748
timestamp 1679585382
transform 1 0 72384 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_755
timestamp 1679585382
transform 1 0 73056 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_762
timestamp 1679585382
transform 1 0 73728 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_769
timestamp 1679585382
transform 1 0 74400 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_776
timestamp 1679585382
transform 1 0 75072 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_783
timestamp 1679585382
transform 1 0 75744 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_790
timestamp 1679585382
transform 1 0 76416 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_797
timestamp 1679585382
transform 1 0 77088 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_804
timestamp 1679585382
transform 1 0 77760 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_811
timestamp 1679585382
transform 1 0 78432 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_818
timestamp 1679585382
transform 1 0 79104 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_825
timestamp 1679585382
transform 1 0 79776 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_832
timestamp 1679585382
transform 1 0 80448 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_839
timestamp 1679585382
transform 1 0 81120 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_846
timestamp 1679585382
transform 1 0 81792 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_853
timestamp 1679585382
transform 1 0 82464 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_860
timestamp 1679585382
transform 1 0 83136 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_867
timestamp 1679585382
transform 1 0 83808 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_874
timestamp 1679585382
transform 1 0 84480 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_881
timestamp 1679585382
transform 1 0 85152 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_888
timestamp 1679585382
transform 1 0 85824 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_895
timestamp 1679585382
transform 1 0 86496 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_902
timestamp 1679585382
transform 1 0 87168 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_909
timestamp 1679585382
transform 1 0 87840 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_916
timestamp 1679585382
transform 1 0 88512 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_923
timestamp 1679585382
transform 1 0 89184 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_930
timestamp 1679585382
transform 1 0 89856 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_937
timestamp 1679585382
transform 1 0 90528 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_944
timestamp 1679585382
transform 1 0 91200 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_951
timestamp 1679585382
transform 1 0 91872 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_958
timestamp 1679585382
transform 1 0 92544 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_965
timestamp 1679585382
transform 1 0 93216 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_972
timestamp 1679585382
transform 1 0 93888 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_979
timestamp 1679585382
transform 1 0 94560 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_986
timestamp 1679585382
transform 1 0 95232 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_993
timestamp 1679585382
transform 1 0 95904 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1000
timestamp 1679585382
transform 1 0 96576 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1007
timestamp 1679585382
transform 1 0 97248 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1014
timestamp 1679585382
transform 1 0 97920 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1021
timestamp 1679585382
transform 1 0 98592 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_1028
timestamp 1677583258
transform 1 0 99264 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_4
timestamp 1679585382
transform 1 0 960 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_11
timestamp 1679585382
transform 1 0 1632 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_18
timestamp 1679585382
transform 1 0 2304 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_25
timestamp 1679585382
transform 1 0 2976 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_32
timestamp 1679585382
transform 1 0 3648 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_39
timestamp 1679585382
transform 1 0 4320 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_46
timestamp 1679585382
transform 1 0 4992 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_53
timestamp 1679585382
transform 1 0 5664 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_60
timestamp 1679585382
transform 1 0 6336 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_67
timestamp 1679585382
transform 1 0 7008 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_74
timestamp 1679585382
transform 1 0 7680 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_81
timestamp 1679585382
transform 1 0 8352 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_88
timestamp 1679585382
transform 1 0 9024 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_95
timestamp 1679585382
transform 1 0 9696 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_102
timestamp 1679581501
transform 1 0 10368 0 1 15876
box -48 -56 432 834
use sg13g2_decap_4  FILLER_20_110
timestamp 1679581501
transform 1 0 11136 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_114
timestamp 1677583258
transform 1 0 11520 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_137
timestamp 1679585382
transform 1 0 13728 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_144
timestamp 1679585382
transform 1 0 14400 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_151
timestamp 1679585382
transform 1 0 15072 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_158
timestamp 1679585382
transform 1 0 15744 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_165
timestamp 1679585382
transform 1 0 16416 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_172
timestamp 1679585382
transform 1 0 17088 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_179
timestamp 1679585382
transform 1 0 17760 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_186
timestamp 1679585382
transform 1 0 18432 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_193
timestamp 1679585382
transform 1 0 19104 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_200
timestamp 1679585382
transform 1 0 19776 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_207
timestamp 1679585382
transform 1 0 20448 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_214
timestamp 1679585382
transform 1 0 21120 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_221
timestamp 1679585382
transform 1 0 21792 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_228
timestamp 1679585382
transform 1 0 22464 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_235
timestamp 1679585382
transform 1 0 23136 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_242
timestamp 1679585382
transform 1 0 23808 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_249
timestamp 1679585382
transform 1 0 24480 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_256
timestamp 1679585382
transform 1 0 25152 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_263
timestamp 1679585382
transform 1 0 25824 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_270
timestamp 1679585382
transform 1 0 26496 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_277
timestamp 1679585382
transform 1 0 27168 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_284
timestamp 1679585382
transform 1 0 27840 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_291
timestamp 1679585382
transform 1 0 28512 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_298
timestamp 1679585382
transform 1 0 29184 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_305
timestamp 1679585382
transform 1 0 29856 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_312
timestamp 1679585382
transform 1 0 30528 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_319
timestamp 1679585382
transform 1 0 31200 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_326
timestamp 1679585382
transform 1 0 31872 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_333
timestamp 1679585382
transform 1 0 32544 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_340
timestamp 1679585382
transform 1 0 33216 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_347
timestamp 1679585382
transform 1 0 33888 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_354
timestamp 1677583704
transform 1 0 34560 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_356
timestamp 1677583258
transform 1 0 34752 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_374
timestamp 1679585382
transform 1 0 36480 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_381
timestamp 1679585382
transform 1 0 37152 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_388
timestamp 1679585382
transform 1 0 37824 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_395
timestamp 1679585382
transform 1 0 38496 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_402
timestamp 1679585382
transform 1 0 39168 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_409
timestamp 1679585382
transform 1 0 39840 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_416
timestamp 1679585382
transform 1 0 40512 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_423
timestamp 1679585382
transform 1 0 41184 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_430
timestamp 1679585382
transform 1 0 41856 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_437
timestamp 1679585382
transform 1 0 42528 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_444
timestamp 1679585382
transform 1 0 43200 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_451
timestamp 1679585382
transform 1 0 43872 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_458
timestamp 1679585382
transform 1 0 44544 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_465
timestamp 1679585382
transform 1 0 45216 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_472
timestamp 1679585382
transform 1 0 45888 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_479
timestamp 1679585382
transform 1 0 46560 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_486
timestamp 1679585382
transform 1 0 47232 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_493
timestamp 1679585382
transform 1 0 47904 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_500
timestamp 1679585382
transform 1 0 48576 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_507
timestamp 1679585382
transform 1 0 49248 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_514
timestamp 1679585382
transform 1 0 49920 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_521
timestamp 1679585382
transform 1 0 50592 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_528
timestamp 1679585382
transform 1 0 51264 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_535
timestamp 1679585382
transform 1 0 51936 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_542
timestamp 1679585382
transform 1 0 52608 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_549
timestamp 1679585382
transform 1 0 53280 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_556
timestamp 1679585382
transform 1 0 53952 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_563
timestamp 1679585382
transform 1 0 54624 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_570
timestamp 1679585382
transform 1 0 55296 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_577
timestamp 1679585382
transform 1 0 55968 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_584
timestamp 1679585382
transform 1 0 56640 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_591
timestamp 1679585382
transform 1 0 57312 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_598
timestamp 1679585382
transform 1 0 57984 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_605
timestamp 1679585382
transform 1 0 58656 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_612
timestamp 1679585382
transform 1 0 59328 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_619
timestamp 1679585382
transform 1 0 60000 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_626
timestamp 1679585382
transform 1 0 60672 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_633
timestamp 1679585382
transform 1 0 61344 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_640
timestamp 1679585382
transform 1 0 62016 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_647
timestamp 1679585382
transform 1 0 62688 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_654
timestamp 1679585382
transform 1 0 63360 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_661
timestamp 1679585382
transform 1 0 64032 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_668
timestamp 1679585382
transform 1 0 64704 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_675
timestamp 1679585382
transform 1 0 65376 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_682
timestamp 1679585382
transform 1 0 66048 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_689
timestamp 1679585382
transform 1 0 66720 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_696
timestamp 1679585382
transform 1 0 67392 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_703
timestamp 1679585382
transform 1 0 68064 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_710
timestamp 1679585382
transform 1 0 68736 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_717
timestamp 1679585382
transform 1 0 69408 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_724
timestamp 1679585382
transform 1 0 70080 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_731
timestamp 1679585382
transform 1 0 70752 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_738
timestamp 1679585382
transform 1 0 71424 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_745
timestamp 1679585382
transform 1 0 72096 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_752
timestamp 1679585382
transform 1 0 72768 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_759
timestamp 1679585382
transform 1 0 73440 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_766
timestamp 1679585382
transform 1 0 74112 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_773
timestamp 1679585382
transform 1 0 74784 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_780
timestamp 1679585382
transform 1 0 75456 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_787
timestamp 1679585382
transform 1 0 76128 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_794
timestamp 1679585382
transform 1 0 76800 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_801
timestamp 1679585382
transform 1 0 77472 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_808
timestamp 1679585382
transform 1 0 78144 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_815
timestamp 1679585382
transform 1 0 78816 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_822
timestamp 1679585382
transform 1 0 79488 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_829
timestamp 1679585382
transform 1 0 80160 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_836
timestamp 1679585382
transform 1 0 80832 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_843
timestamp 1679585382
transform 1 0 81504 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_850
timestamp 1679585382
transform 1 0 82176 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_857
timestamp 1679585382
transform 1 0 82848 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_864
timestamp 1679585382
transform 1 0 83520 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_871
timestamp 1679585382
transform 1 0 84192 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_878
timestamp 1679585382
transform 1 0 84864 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_885
timestamp 1679585382
transform 1 0 85536 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_892
timestamp 1679585382
transform 1 0 86208 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_899
timestamp 1679585382
transform 1 0 86880 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_906
timestamp 1679585382
transform 1 0 87552 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_913
timestamp 1679585382
transform 1 0 88224 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_920
timestamp 1679585382
transform 1 0 88896 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_927
timestamp 1679585382
transform 1 0 89568 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_934
timestamp 1679585382
transform 1 0 90240 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_941
timestamp 1679585382
transform 1 0 90912 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_948
timestamp 1679585382
transform 1 0 91584 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_955
timestamp 1679585382
transform 1 0 92256 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_962
timestamp 1679585382
transform 1 0 92928 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_969
timestamp 1679585382
transform 1 0 93600 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_976
timestamp 1679585382
transform 1 0 94272 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_983
timestamp 1679585382
transform 1 0 94944 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_990
timestamp 1679585382
transform 1 0 95616 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_997
timestamp 1679585382
transform 1 0 96288 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1004
timestamp 1679585382
transform 1 0 96960 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1011
timestamp 1679585382
transform 1 0 97632 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1018
timestamp 1679585382
transform 1 0 98304 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_1025
timestamp 1679581501
transform 1 0 98976 0 1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_21_4
timestamp 1679585382
transform 1 0 960 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_11
timestamp 1679585382
transform 1 0 1632 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_18
timestamp 1679585382
transform 1 0 2304 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_25
timestamp 1679585382
transform 1 0 2976 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_32
timestamp 1679585382
transform 1 0 3648 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_39
timestamp 1679585382
transform 1 0 4320 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_46
timestamp 1677583704
transform 1 0 4992 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_83
timestamp 1679585382
transform 1 0 8544 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_90
timestamp 1679585382
transform 1 0 9216 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_97
timestamp 1679581501
transform 1 0 9888 0 -1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_21_132
timestamp 1679585382
transform 1 0 13248 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_139
timestamp 1679585382
transform 1 0 13920 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_146
timestamp 1679585382
transform 1 0 14592 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_153
timestamp 1679585382
transform 1 0 15264 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_160
timestamp 1679581501
transform 1 0 15936 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_164
timestamp 1677583258
transform 1 0 16320 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_205
timestamp 1679585382
transform 1 0 20256 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_212
timestamp 1679585382
transform 1 0 20928 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_21_219
timestamp 1677583258
transform 1 0 21600 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_21_224
timestamp 1679581501
transform 1 0 22080 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_21_228
timestamp 1677583704
transform 1 0 22464 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_257
timestamp 1679585382
transform 1 0 25248 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_264
timestamp 1679585382
transform 1 0 25920 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_271
timestamp 1679585382
transform 1 0 26592 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_278
timestamp 1679585382
transform 1 0 27264 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_285
timestamp 1679585382
transform 1 0 27936 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_292
timestamp 1679585382
transform 1 0 28608 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_299
timestamp 1679585382
transform 1 0 29280 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_306
timestamp 1679585382
transform 1 0 29952 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_313
timestamp 1677583704
transform 1 0 30624 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_315
timestamp 1677583258
transform 1 0 30816 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_351
timestamp 1679585382
transform 1 0 34272 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_358
timestamp 1679585382
transform 1 0 34944 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_365
timestamp 1679585382
transform 1 0 35616 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_408
timestamp 1677583704
transform 1 0 39744 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_437
timestamp 1679585382
transform 1 0 42528 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_444
timestamp 1679585382
transform 1 0 43200 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_451
timestamp 1679585382
transform 1 0 43872 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_458
timestamp 1679585382
transform 1 0 44544 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_465
timestamp 1679585382
transform 1 0 45216 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_472
timestamp 1679585382
transform 1 0 45888 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_479
timestamp 1679585382
transform 1 0 46560 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_486
timestamp 1679585382
transform 1 0 47232 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_493
timestamp 1679585382
transform 1 0 47904 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_500
timestamp 1679585382
transform 1 0 48576 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_507
timestamp 1679585382
transform 1 0 49248 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_514
timestamp 1679585382
transform 1 0 49920 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_521
timestamp 1679585382
transform 1 0 50592 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_528
timestamp 1679585382
transform 1 0 51264 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_535
timestamp 1679585382
transform 1 0 51936 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_542
timestamp 1679585382
transform 1 0 52608 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_549
timestamp 1679585382
transform 1 0 53280 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_556
timestamp 1679581501
transform 1 0 53952 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_560
timestamp 1677583258
transform 1 0 54336 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_596
timestamp 1679585382
transform 1 0 57792 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_603
timestamp 1679585382
transform 1 0 58464 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_610
timestamp 1679585382
transform 1 0 59136 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_617
timestamp 1679585382
transform 1 0 59808 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_624
timestamp 1679585382
transform 1 0 60480 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_631
timestamp 1679585382
transform 1 0 61152 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_638
timestamp 1679585382
transform 1 0 61824 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_645
timestamp 1679585382
transform 1 0 62496 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_652
timestamp 1679585382
transform 1 0 63168 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_659
timestamp 1679585382
transform 1 0 63840 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_666
timestamp 1679585382
transform 1 0 64512 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_673
timestamp 1679585382
transform 1 0 65184 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_680
timestamp 1679585382
transform 1 0 65856 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_687
timestamp 1679585382
transform 1 0 66528 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_694
timestamp 1679585382
transform 1 0 67200 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_701
timestamp 1679585382
transform 1 0 67872 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_708
timestamp 1679585382
transform 1 0 68544 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_715
timestamp 1679585382
transform 1 0 69216 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_722
timestamp 1679585382
transform 1 0 69888 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_729
timestamp 1679585382
transform 1 0 70560 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_736
timestamp 1679585382
transform 1 0 71232 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_743
timestamp 1679585382
transform 1 0 71904 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_750
timestamp 1679585382
transform 1 0 72576 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_757
timestamp 1679585382
transform 1 0 73248 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_764
timestamp 1679585382
transform 1 0 73920 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_771
timestamp 1679585382
transform 1 0 74592 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_778
timestamp 1679585382
transform 1 0 75264 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_785
timestamp 1679585382
transform 1 0 75936 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_792
timestamp 1679585382
transform 1 0 76608 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_799
timestamp 1679585382
transform 1 0 77280 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_806
timestamp 1679585382
transform 1 0 77952 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_813
timestamp 1679585382
transform 1 0 78624 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_820
timestamp 1679585382
transform 1 0 79296 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_827
timestamp 1679585382
transform 1 0 79968 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_834
timestamp 1679585382
transform 1 0 80640 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_841
timestamp 1679585382
transform 1 0 81312 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_848
timestamp 1679585382
transform 1 0 81984 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_855
timestamp 1679585382
transform 1 0 82656 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_862
timestamp 1679585382
transform 1 0 83328 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_869
timestamp 1679585382
transform 1 0 84000 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_876
timestamp 1679585382
transform 1 0 84672 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_883
timestamp 1679585382
transform 1 0 85344 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_890
timestamp 1679585382
transform 1 0 86016 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_897
timestamp 1679585382
transform 1 0 86688 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_904
timestamp 1679585382
transform 1 0 87360 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_911
timestamp 1679585382
transform 1 0 88032 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_918
timestamp 1679585382
transform 1 0 88704 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_925
timestamp 1679585382
transform 1 0 89376 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_932
timestamp 1679585382
transform 1 0 90048 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_939
timestamp 1679585382
transform 1 0 90720 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_946
timestamp 1679585382
transform 1 0 91392 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_953
timestamp 1679585382
transform 1 0 92064 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_960
timestamp 1679585382
transform 1 0 92736 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_967
timestamp 1679585382
transform 1 0 93408 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_974
timestamp 1679585382
transform 1 0 94080 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_981
timestamp 1679585382
transform 1 0 94752 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_988
timestamp 1679585382
transform 1 0 95424 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_995
timestamp 1679585382
transform 1 0 96096 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1002
timestamp 1679585382
transform 1 0 96768 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1009
timestamp 1679585382
transform 1 0 97440 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1016
timestamp 1679585382
transform 1 0 98112 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_1023
timestamp 1679581501
transform 1 0 98784 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_21_1027
timestamp 1677583704
transform 1 0 99168 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_4
timestamp 1679585382
transform 1 0 960 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_11
timestamp 1679585382
transform 1 0 1632 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_18
timestamp 1679585382
transform 1 0 2304 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_25
timestamp 1679585382
transform 1 0 2976 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_32
timestamp 1679581501
transform 1 0 3648 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_72
timestamp 1677583258
transform 1 0 7488 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_82
timestamp 1677583704
transform 1 0 8448 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_84
timestamp 1677583258
transform 1 0 8640 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_89
timestamp 1679585382
transform 1 0 9120 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_96
timestamp 1679585382
transform 1 0 9792 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_103
timestamp 1679581501
transform 1 0 10464 0 1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_22_134
timestamp 1679585382
transform 1 0 13440 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_141
timestamp 1679585382
transform 1 0 14112 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_148
timestamp 1679585382
transform 1 0 14784 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_155
timestamp 1679585382
transform 1 0 15456 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_162
timestamp 1679585382
transform 1 0 16128 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_169
timestamp 1679585382
transform 1 0 16800 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_176
timestamp 1679585382
transform 1 0 17472 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_183
timestamp 1679585382
transform 1 0 18144 0 1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_22_190
timestamp 1677583258
transform 1 0 18816 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_194
timestamp 1679585382
transform 1 0 19200 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_201
timestamp 1679585382
transform 1 0 19872 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_208
timestamp 1679581501
transform 1 0 20544 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_239
timestamp 1677583704
transform 1 0 23520 0 1 17388
box -48 -56 240 834
use sg13g2_decap_4  FILLER_22_245
timestamp 1679581501
transform 1 0 24096 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_249
timestamp 1677583258
transform 1 0 24480 0 1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_22_259
timestamp 1679581501
transform 1 0 25440 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_267
timestamp 1677583704
transform 1 0 26208 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_273
timestamp 1677583704
transform 1 0 26784 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_288
timestamp 1679585382
transform 1 0 28224 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_295
timestamp 1679585382
transform 1 0 28896 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_302
timestamp 1677583704
transform 1 0 29568 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_304
timestamp 1677583258
transform 1 0 29760 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_332
timestamp 1679585382
transform 1 0 32448 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_339
timestamp 1679585382
transform 1 0 33120 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_346
timestamp 1679585382
transform 1 0 33792 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_353
timestamp 1679585382
transform 1 0 34464 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_360
timestamp 1679585382
transform 1 0 35136 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_367
timestamp 1679585382
transform 1 0 35808 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_374
timestamp 1679585382
transform 1 0 36480 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_381
timestamp 1679585382
transform 1 0 37152 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_388
timestamp 1679585382
transform 1 0 37824 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_395
timestamp 1679585382
transform 1 0 38496 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_402
timestamp 1679585382
transform 1 0 39168 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_409
timestamp 1679585382
transform 1 0 39840 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_416
timestamp 1679585382
transform 1 0 40512 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_423
timestamp 1677583704
transform 1 0 41184 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_433
timestamp 1679585382
transform 1 0 42144 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_440
timestamp 1679585382
transform 1 0 42816 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_447
timestamp 1679585382
transform 1 0 43488 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_454
timestamp 1679585382
transform 1 0 44160 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_461
timestamp 1679585382
transform 1 0 44832 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_468
timestamp 1679585382
transform 1 0 45504 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_475
timestamp 1679585382
transform 1 0 46176 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_482
timestamp 1677583704
transform 1 0 46848 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_484
timestamp 1677583258
transform 1 0 47040 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_493
timestamp 1677583258
transform 1 0 47904 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_508
timestamp 1679585382
transform 1 0 49344 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_515
timestamp 1679585382
transform 1 0 50016 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_522
timestamp 1679585382
transform 1 0 50688 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_529
timestamp 1679585382
transform 1 0 51360 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_536
timestamp 1679585382
transform 1 0 52032 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_543
timestamp 1679585382
transform 1 0 52704 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_550
timestamp 1679585382
transform 1 0 53376 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_557
timestamp 1679585382
transform 1 0 54048 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_564
timestamp 1679585382
transform 1 0 54720 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_571
timestamp 1679585382
transform 1 0 55392 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_578
timestamp 1679585382
transform 1 0 56064 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_585
timestamp 1679585382
transform 1 0 56736 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_592
timestamp 1679585382
transform 1 0 57408 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_599
timestamp 1679585382
transform 1 0 58080 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_606
timestamp 1679585382
transform 1 0 58752 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_613
timestamp 1679585382
transform 1 0 59424 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_620
timestamp 1679585382
transform 1 0 60096 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_627
timestamp 1679585382
transform 1 0 60768 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_634
timestamp 1679585382
transform 1 0 61440 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_641
timestamp 1679585382
transform 1 0 62112 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_648
timestamp 1679585382
transform 1 0 62784 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_655
timestamp 1679585382
transform 1 0 63456 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_662
timestamp 1679585382
transform 1 0 64128 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_669
timestamp 1679585382
transform 1 0 64800 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_676
timestamp 1679585382
transform 1 0 65472 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_683
timestamp 1679585382
transform 1 0 66144 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_690
timestamp 1679585382
transform 1 0 66816 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_697
timestamp 1679585382
transform 1 0 67488 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_704
timestamp 1679585382
transform 1 0 68160 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_711
timestamp 1679585382
transform 1 0 68832 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_718
timestamp 1679585382
transform 1 0 69504 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_725
timestamp 1679585382
transform 1 0 70176 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_732
timestamp 1679585382
transform 1 0 70848 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_739
timestamp 1679585382
transform 1 0 71520 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_746
timestamp 1679585382
transform 1 0 72192 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_753
timestamp 1679585382
transform 1 0 72864 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_760
timestamp 1679585382
transform 1 0 73536 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_767
timestamp 1679585382
transform 1 0 74208 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_774
timestamp 1679585382
transform 1 0 74880 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_781
timestamp 1679585382
transform 1 0 75552 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_788
timestamp 1679585382
transform 1 0 76224 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_795
timestamp 1679585382
transform 1 0 76896 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_802
timestamp 1679585382
transform 1 0 77568 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_809
timestamp 1679585382
transform 1 0 78240 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_816
timestamp 1679585382
transform 1 0 78912 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_823
timestamp 1679585382
transform 1 0 79584 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_830
timestamp 1679585382
transform 1 0 80256 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_837
timestamp 1679585382
transform 1 0 80928 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_844
timestamp 1679585382
transform 1 0 81600 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_851
timestamp 1679585382
transform 1 0 82272 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_858
timestamp 1679585382
transform 1 0 82944 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_865
timestamp 1679585382
transform 1 0 83616 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_872
timestamp 1679585382
transform 1 0 84288 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_879
timestamp 1679585382
transform 1 0 84960 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_886
timestamp 1679585382
transform 1 0 85632 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_893
timestamp 1679585382
transform 1 0 86304 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_900
timestamp 1679585382
transform 1 0 86976 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_907
timestamp 1679585382
transform 1 0 87648 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_914
timestamp 1679585382
transform 1 0 88320 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_921
timestamp 1679585382
transform 1 0 88992 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_928
timestamp 1679585382
transform 1 0 89664 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_935
timestamp 1679585382
transform 1 0 90336 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_942
timestamp 1679585382
transform 1 0 91008 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_949
timestamp 1679585382
transform 1 0 91680 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_956
timestamp 1679585382
transform 1 0 92352 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_963
timestamp 1679585382
transform 1 0 93024 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_970
timestamp 1679585382
transform 1 0 93696 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_977
timestamp 1679585382
transform 1 0 94368 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_984
timestamp 1679585382
transform 1 0 95040 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_991
timestamp 1679585382
transform 1 0 95712 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_998
timestamp 1679585382
transform 1 0 96384 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1005
timestamp 1679585382
transform 1 0 97056 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1012
timestamp 1679585382
transform 1 0 97728 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1019
timestamp 1679585382
transform 1 0 98400 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_1026
timestamp 1677583704
transform 1 0 99072 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_1028
timestamp 1677583258
transform 1 0 99264 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_4
timestamp 1679585382
transform 1 0 960 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_38
timestamp 1679585382
transform 1 0 4224 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_45
timestamp 1679585382
transform 1 0 4896 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_52
timestamp 1679585382
transform 1 0 5568 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_59
timestamp 1677583704
transform 1 0 6240 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_61
timestamp 1677583258
transform 1 0 6432 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_87
timestamp 1679585382
transform 1 0 8928 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_94
timestamp 1679585382
transform 1 0 9600 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_101
timestamp 1679585382
transform 1 0 10272 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_108
timestamp 1679585382
transform 1 0 10944 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_23_115
timestamp 1677583258
transform 1 0 11616 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_130
timestamp 1679585382
transform 1 0 13056 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_137
timestamp 1679585382
transform 1 0 13728 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_144
timestamp 1679585382
transform 1 0 14400 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_151
timestamp 1679585382
transform 1 0 15072 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_158
timestamp 1679585382
transform 1 0 15744 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_165
timestamp 1679585382
transform 1 0 16416 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_172
timestamp 1677583704
transform 1 0 17088 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_201
timestamp 1679585382
transform 1 0 19872 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_208
timestamp 1679585382
transform 1 0 20544 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_215
timestamp 1679585382
transform 1 0 21216 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_222
timestamp 1679585382
transform 1 0 21888 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_229
timestamp 1677583704
transform 1 0 22560 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_240
timestamp 1679585382
transform 1 0 23616 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_247
timestamp 1679585382
transform 1 0 24288 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_23_254
timestamp 1677583258
transform 1 0 24960 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_282
timestamp 1679585382
transform 1 0 27648 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_289
timestamp 1679585382
transform 1 0 28320 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_296
timestamp 1679585382
transform 1 0 28992 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_303
timestamp 1679585382
transform 1 0 29664 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_310
timestamp 1679585382
transform 1 0 30336 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_317
timestamp 1679585382
transform 1 0 31008 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_324
timestamp 1679585382
transform 1 0 31680 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_331
timestamp 1679585382
transform 1 0 32352 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_338
timestamp 1679585382
transform 1 0 33024 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_345
timestamp 1679585382
transform 1 0 33696 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_352
timestamp 1679585382
transform 1 0 34368 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_359
timestamp 1679585382
transform 1 0 35040 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_366
timestamp 1679585382
transform 1 0 35712 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_373
timestamp 1679585382
transform 1 0 36384 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_380
timestamp 1679585382
transform 1 0 37056 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_387
timestamp 1679585382
transform 1 0 37728 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_394
timestamp 1679585382
transform 1 0 38400 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_401
timestamp 1679585382
transform 1 0 39072 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_408
timestamp 1677583704
transform 1 0 39744 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_419
timestamp 1677583704
transform 1 0 40800 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_448
timestamp 1679585382
transform 1 0 43584 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_455
timestamp 1679585382
transform 1 0 44256 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_462
timestamp 1679585382
transform 1 0 44928 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_469
timestamp 1679585382
transform 1 0 45600 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_476
timestamp 1679581501
transform 1 0 46272 0 -1 18900
box -48 -56 432 834
use sg13g2_decap_8  FILLER_23_507
timestamp 1679585382
transform 1 0 49248 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_514
timestamp 1679585382
transform 1 0 49920 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_521
timestamp 1679585382
transform 1 0 50592 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_528
timestamp 1679585382
transform 1 0 51264 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_562
timestamp 1679585382
transform 1 0 54528 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_569
timestamp 1679585382
transform 1 0 55200 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_576
timestamp 1679585382
transform 1 0 55872 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_583
timestamp 1679585382
transform 1 0 56544 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_590
timestamp 1679585382
transform 1 0 57216 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_597
timestamp 1679585382
transform 1 0 57888 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_604
timestamp 1679585382
transform 1 0 58560 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_611
timestamp 1679585382
transform 1 0 59232 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_618
timestamp 1679585382
transform 1 0 59904 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_625
timestamp 1679585382
transform 1 0 60576 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_632
timestamp 1679585382
transform 1 0 61248 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_639
timestamp 1679585382
transform 1 0 61920 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_646
timestamp 1679585382
transform 1 0 62592 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_653
timestamp 1679585382
transform 1 0 63264 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_660
timestamp 1679585382
transform 1 0 63936 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_667
timestamp 1679585382
transform 1 0 64608 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_674
timestamp 1679585382
transform 1 0 65280 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_681
timestamp 1679585382
transform 1 0 65952 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_688
timestamp 1679585382
transform 1 0 66624 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_695
timestamp 1679585382
transform 1 0 67296 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_702
timestamp 1679585382
transform 1 0 67968 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_709
timestamp 1679585382
transform 1 0 68640 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_716
timestamp 1679585382
transform 1 0 69312 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_723
timestamp 1679585382
transform 1 0 69984 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_730
timestamp 1679585382
transform 1 0 70656 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_737
timestamp 1679585382
transform 1 0 71328 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_744
timestamp 1679585382
transform 1 0 72000 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_751
timestamp 1679585382
transform 1 0 72672 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_758
timestamp 1679585382
transform 1 0 73344 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_765
timestamp 1679585382
transform 1 0 74016 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_772
timestamp 1679585382
transform 1 0 74688 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_779
timestamp 1679585382
transform 1 0 75360 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_786
timestamp 1679585382
transform 1 0 76032 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_793
timestamp 1679585382
transform 1 0 76704 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_800
timestamp 1679585382
transform 1 0 77376 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_807
timestamp 1679585382
transform 1 0 78048 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_814
timestamp 1679585382
transform 1 0 78720 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_821
timestamp 1679585382
transform 1 0 79392 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_828
timestamp 1679585382
transform 1 0 80064 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_835
timestamp 1679585382
transform 1 0 80736 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_842
timestamp 1679585382
transform 1 0 81408 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_849
timestamp 1679585382
transform 1 0 82080 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_856
timestamp 1679585382
transform 1 0 82752 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_863
timestamp 1679585382
transform 1 0 83424 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_870
timestamp 1679585382
transform 1 0 84096 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_877
timestamp 1679585382
transform 1 0 84768 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_884
timestamp 1679585382
transform 1 0 85440 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_891
timestamp 1679585382
transform 1 0 86112 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_898
timestamp 1679585382
transform 1 0 86784 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_905
timestamp 1679585382
transform 1 0 87456 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_912
timestamp 1679585382
transform 1 0 88128 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_919
timestamp 1679585382
transform 1 0 88800 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_926
timestamp 1679585382
transform 1 0 89472 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_933
timestamp 1679585382
transform 1 0 90144 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_940
timestamp 1679585382
transform 1 0 90816 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_947
timestamp 1679585382
transform 1 0 91488 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_954
timestamp 1679585382
transform 1 0 92160 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_961
timestamp 1679585382
transform 1 0 92832 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_968
timestamp 1679585382
transform 1 0 93504 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_975
timestamp 1679585382
transform 1 0 94176 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_982
timestamp 1679585382
transform 1 0 94848 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_989
timestamp 1679585382
transform 1 0 95520 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_996
timestamp 1679585382
transform 1 0 96192 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1003
timestamp 1679585382
transform 1 0 96864 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1010
timestamp 1679585382
transform 1 0 97536 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1017
timestamp 1679585382
transform 1 0 98208 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_1024
timestamp 1679581501
transform 1 0 98880 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_1028
timestamp 1677583258
transform 1 0 99264 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_4
timestamp 1679585382
transform 1 0 960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_11
timestamp 1679585382
transform 1 0 1632 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_18
timestamp 1677583704
transform 1 0 2304 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_20
timestamp 1677583258
transform 1 0 2496 0 1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_24_25
timestamp 1679581501
transform 1 0 2976 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_29
timestamp 1677583704
transform 1 0 3360 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_40
timestamp 1679585382
transform 1 0 4416 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_47
timestamp 1679585382
transform 1 0 5088 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_54
timestamp 1679585382
transform 1 0 5760 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_61
timestamp 1679585382
transform 1 0 6432 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_68
timestamp 1679585382
transform 1 0 7104 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_75
timestamp 1679585382
transform 1 0 7776 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_82
timestamp 1679585382
transform 1 0 8448 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_89
timestamp 1679585382
transform 1 0 9120 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_96
timestamp 1679585382
transform 1 0 9792 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_103
timestamp 1679585382
transform 1 0 10464 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_110
timestamp 1679585382
transform 1 0 11136 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_117
timestamp 1679585382
transform 1 0 11808 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_124
timestamp 1679585382
transform 1 0 12480 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_131
timestamp 1679585382
transform 1 0 13152 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_138
timestamp 1679585382
transform 1 0 13824 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_145
timestamp 1679585382
transform 1 0 14496 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_152
timestamp 1679585382
transform 1 0 15168 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_159
timestamp 1679585382
transform 1 0 15840 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_166
timestamp 1679585382
transform 1 0 16512 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_173
timestamp 1679585382
transform 1 0 17184 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_180
timestamp 1679585382
transform 1 0 17856 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_187
timestamp 1679585382
transform 1 0 18528 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_194
timestamp 1679585382
transform 1 0 19200 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_201
timestamp 1679585382
transform 1 0 19872 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_208
timestamp 1679585382
transform 1 0 20544 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_215
timestamp 1679585382
transform 1 0 21216 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_222
timestamp 1679585382
transform 1 0 21888 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_229
timestamp 1679585382
transform 1 0 22560 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_236
timestamp 1679585382
transform 1 0 23232 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_243
timestamp 1679585382
transform 1 0 23904 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_250
timestamp 1679585382
transform 1 0 24576 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_257
timestamp 1679585382
transform 1 0 25248 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_264
timestamp 1679581501
transform 1 0 25920 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_268
timestamp 1677583704
transform 1 0 26304 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_283
timestamp 1679585382
transform 1 0 27744 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_290
timestamp 1679585382
transform 1 0 28416 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_297
timestamp 1679585382
transform 1 0 29088 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_304
timestamp 1679585382
transform 1 0 29760 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_311
timestamp 1679585382
transform 1 0 30432 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_318
timestamp 1679585382
transform 1 0 31104 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_325
timestamp 1679585382
transform 1 0 31776 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_332
timestamp 1679585382
transform 1 0 32448 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_339
timestamp 1679585382
transform 1 0 33120 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_346
timestamp 1679585382
transform 1 0 33792 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_353
timestamp 1677583704
transform 1 0 34464 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_355
timestamp 1677583258
transform 1 0 34656 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_369
timestamp 1679585382
transform 1 0 36000 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_376
timestamp 1679585382
transform 1 0 36672 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_383
timestamp 1679585382
transform 1 0 37344 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_390
timestamp 1679585382
transform 1 0 38016 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_397
timestamp 1679581501
transform 1 0 38688 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_401
timestamp 1677583704
transform 1 0 39072 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_411
timestamp 1679585382
transform 1 0 40032 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_418
timestamp 1679585382
transform 1 0 40704 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_425
timestamp 1679585382
transform 1 0 41376 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_432
timestamp 1679585382
transform 1 0 42048 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_439
timestamp 1679585382
transform 1 0 42720 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_446
timestamp 1679585382
transform 1 0 43392 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_453
timestamp 1679585382
transform 1 0 44064 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_460
timestamp 1679585382
transform 1 0 44736 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_467
timestamp 1679585382
transform 1 0 45408 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_474
timestamp 1677583704
transform 1 0 46080 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_503
timestamp 1679585382
transform 1 0 48864 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_510
timestamp 1679581501
transform 1 0 49536 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_514
timestamp 1677583704
transform 1 0 49920 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_524
timestamp 1679585382
transform 1 0 50880 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_531
timestamp 1679585382
transform 1 0 51552 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_538
timestamp 1679585382
transform 1 0 52224 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_545
timestamp 1679585382
transform 1 0 52896 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_552
timestamp 1679585382
transform 1 0 53568 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_559
timestamp 1679585382
transform 1 0 54240 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_566
timestamp 1679585382
transform 1 0 54912 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_573
timestamp 1679585382
transform 1 0 55584 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_580
timestamp 1679585382
transform 1 0 56256 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_587
timestamp 1679585382
transform 1 0 56928 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_594
timestamp 1679585382
transform 1 0 57600 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_601
timestamp 1679585382
transform 1 0 58272 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_608
timestamp 1679585382
transform 1 0 58944 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_615
timestamp 1679585382
transform 1 0 59616 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_622
timestamp 1679585382
transform 1 0 60288 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_629
timestamp 1679585382
transform 1 0 60960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_636
timestamp 1679585382
transform 1 0 61632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_643
timestamp 1679585382
transform 1 0 62304 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_650
timestamp 1679585382
transform 1 0 62976 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_657
timestamp 1679585382
transform 1 0 63648 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_664
timestamp 1679585382
transform 1 0 64320 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_671
timestamp 1679585382
transform 1 0 64992 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_678
timestamp 1679585382
transform 1 0 65664 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_685
timestamp 1679585382
transform 1 0 66336 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_692
timestamp 1679585382
transform 1 0 67008 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_699
timestamp 1679585382
transform 1 0 67680 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_706
timestamp 1679585382
transform 1 0 68352 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_713
timestamp 1679585382
transform 1 0 69024 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_720
timestamp 1679585382
transform 1 0 69696 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_727
timestamp 1679585382
transform 1 0 70368 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_734
timestamp 1679585382
transform 1 0 71040 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_741
timestamp 1679585382
transform 1 0 71712 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_748
timestamp 1679585382
transform 1 0 72384 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_755
timestamp 1679585382
transform 1 0 73056 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_762
timestamp 1679585382
transform 1 0 73728 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_769
timestamp 1679585382
transform 1 0 74400 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_776
timestamp 1679585382
transform 1 0 75072 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_783
timestamp 1679585382
transform 1 0 75744 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_790
timestamp 1679585382
transform 1 0 76416 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_797
timestamp 1679585382
transform 1 0 77088 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_804
timestamp 1679585382
transform 1 0 77760 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_811
timestamp 1679585382
transform 1 0 78432 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_818
timestamp 1679585382
transform 1 0 79104 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_825
timestamp 1679585382
transform 1 0 79776 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_832
timestamp 1679585382
transform 1 0 80448 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_839
timestamp 1679585382
transform 1 0 81120 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_846
timestamp 1679585382
transform 1 0 81792 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_853
timestamp 1679585382
transform 1 0 82464 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_860
timestamp 1679585382
transform 1 0 83136 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_867
timestamp 1679585382
transform 1 0 83808 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_874
timestamp 1679585382
transform 1 0 84480 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_881
timestamp 1679585382
transform 1 0 85152 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_888
timestamp 1679585382
transform 1 0 85824 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_895
timestamp 1679585382
transform 1 0 86496 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_902
timestamp 1679585382
transform 1 0 87168 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_909
timestamp 1679585382
transform 1 0 87840 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_916
timestamp 1679585382
transform 1 0 88512 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_923
timestamp 1679585382
transform 1 0 89184 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_930
timestamp 1679585382
transform 1 0 89856 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_937
timestamp 1679585382
transform 1 0 90528 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_944
timestamp 1679585382
transform 1 0 91200 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_951
timestamp 1679585382
transform 1 0 91872 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_958
timestamp 1679585382
transform 1 0 92544 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_965
timestamp 1679585382
transform 1 0 93216 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_972
timestamp 1679585382
transform 1 0 93888 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_979
timestamp 1679585382
transform 1 0 94560 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_986
timestamp 1679585382
transform 1 0 95232 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_993
timestamp 1679585382
transform 1 0 95904 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1000
timestamp 1679585382
transform 1 0 96576 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1007
timestamp 1679585382
transform 1 0 97248 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1014
timestamp 1679585382
transform 1 0 97920 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1021
timestamp 1679585382
transform 1 0 98592 0 1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_24_1028
timestamp 1677583258
transform 1 0 99264 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_4
timestamp 1679585382
transform 1 0 960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_11
timestamp 1679585382
transform 1 0 1632 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_18
timestamp 1679585382
transform 1 0 2304 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_25
timestamp 1679585382
transform 1 0 2976 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_32
timestamp 1679585382
transform 1 0 3648 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_39
timestamp 1679585382
transform 1 0 4320 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_46
timestamp 1679585382
transform 1 0 4992 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_53
timestamp 1679585382
transform 1 0 5664 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_60
timestamp 1679585382
transform 1 0 6336 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_67
timestamp 1679585382
transform 1 0 7008 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_74
timestamp 1679585382
transform 1 0 7680 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_81
timestamp 1677583704
transform 1 0 8352 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_83
timestamp 1677583258
transform 1 0 8544 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_111
timestamp 1679585382
transform 1 0 11232 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_118
timestamp 1679585382
transform 1 0 11904 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_125
timestamp 1679581501
transform 1 0 12576 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_25_156
timestamp 1679585382
transform 1 0 15552 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_163
timestamp 1679585382
transform 1 0 16224 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_170
timestamp 1679585382
transform 1 0 16896 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_177
timestamp 1679585382
transform 1 0 17568 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_184
timestamp 1679585382
transform 1 0 18240 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_191
timestamp 1679585382
transform 1 0 18912 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_198
timestamp 1679585382
transform 1 0 19584 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_25_205
timestamp 1677583258
transform 1 0 20256 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_215
timestamp 1679585382
transform 1 0 21216 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_222
timestamp 1679585382
transform 1 0 21888 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_229
timestamp 1679585382
transform 1 0 22560 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_236
timestamp 1679585382
transform 1 0 23232 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_243
timestamp 1679585382
transform 1 0 23904 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_250
timestamp 1677583704
transform 1 0 24576 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_252
timestamp 1677583258
transform 1 0 24768 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_280
timestamp 1679585382
transform 1 0 27456 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_287
timestamp 1679585382
transform 1 0 28128 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_294
timestamp 1677583704
transform 1 0 28800 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_296
timestamp 1677583258
transform 1 0 28992 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_323
timestamp 1679585382
transform 1 0 31584 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_330
timestamp 1679585382
transform 1 0 32256 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_337
timestamp 1679585382
transform 1 0 32928 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_344
timestamp 1679585382
transform 1 0 33600 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_351
timestamp 1679585382
transform 1 0 34272 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_358
timestamp 1679585382
transform 1 0 34944 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_365
timestamp 1679581501
transform 1 0 35616 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_25_396
timestamp 1679585382
transform 1 0 38592 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_403
timestamp 1679581501
transform 1 0 39264 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_411
timestamp 1677583704
transform 1 0 40032 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_430
timestamp 1679585382
transform 1 0 41856 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_437
timestamp 1679585382
transform 1 0 42528 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_444
timestamp 1679585382
transform 1 0 43200 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_451
timestamp 1679585382
transform 1 0 43872 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_458
timestamp 1679585382
transform 1 0 44544 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_465
timestamp 1679585382
transform 1 0 45216 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_472
timestamp 1679585382
transform 1 0 45888 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_479
timestamp 1679585382
transform 1 0 46560 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_486
timestamp 1679585382
transform 1 0 47232 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_493
timestamp 1677583704
transform 1 0 47904 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_25_504
timestamp 1677583704
transform 1 0 48960 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_506
timestamp 1677583258
transform 1 0 49152 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_515
timestamp 1679585382
transform 1 0 50016 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_522
timestamp 1679585382
transform 1 0 50688 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_529
timestamp 1679585382
transform 1 0 51360 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_536
timestamp 1679585382
transform 1 0 52032 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_543
timestamp 1679585382
transform 1 0 52704 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_550
timestamp 1679585382
transform 1 0 53376 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_557
timestamp 1679585382
transform 1 0 54048 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_564
timestamp 1679585382
transform 1 0 54720 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_571
timestamp 1679585382
transform 1 0 55392 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_578
timestamp 1679585382
transform 1 0 56064 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_585
timestamp 1679585382
transform 1 0 56736 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_592
timestamp 1679585382
transform 1 0 57408 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_599
timestamp 1679585382
transform 1 0 58080 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_606
timestamp 1679585382
transform 1 0 58752 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_613
timestamp 1679585382
transform 1 0 59424 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_620
timestamp 1679585382
transform 1 0 60096 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_627
timestamp 1679585382
transform 1 0 60768 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_634
timestamp 1679585382
transform 1 0 61440 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_641
timestamp 1679585382
transform 1 0 62112 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_648
timestamp 1679585382
transform 1 0 62784 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_655
timestamp 1679585382
transform 1 0 63456 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_662
timestamp 1679585382
transform 1 0 64128 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_669
timestamp 1679585382
transform 1 0 64800 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_676
timestamp 1679585382
transform 1 0 65472 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_683
timestamp 1679585382
transform 1 0 66144 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_690
timestamp 1679585382
transform 1 0 66816 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_697
timestamp 1679585382
transform 1 0 67488 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_704
timestamp 1679585382
transform 1 0 68160 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_711
timestamp 1679585382
transform 1 0 68832 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_718
timestamp 1679585382
transform 1 0 69504 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_725
timestamp 1679585382
transform 1 0 70176 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_732
timestamp 1679585382
transform 1 0 70848 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_739
timestamp 1679585382
transform 1 0 71520 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_746
timestamp 1679585382
transform 1 0 72192 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_753
timestamp 1679585382
transform 1 0 72864 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_760
timestamp 1679585382
transform 1 0 73536 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_767
timestamp 1679585382
transform 1 0 74208 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_774
timestamp 1679585382
transform 1 0 74880 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_781
timestamp 1679585382
transform 1 0 75552 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_788
timestamp 1679585382
transform 1 0 76224 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_795
timestamp 1679585382
transform 1 0 76896 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_802
timestamp 1679585382
transform 1 0 77568 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_809
timestamp 1679585382
transform 1 0 78240 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_816
timestamp 1679585382
transform 1 0 78912 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_823
timestamp 1679585382
transform 1 0 79584 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_830
timestamp 1679585382
transform 1 0 80256 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_837
timestamp 1679585382
transform 1 0 80928 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_844
timestamp 1679585382
transform 1 0 81600 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_851
timestamp 1679585382
transform 1 0 82272 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_858
timestamp 1679585382
transform 1 0 82944 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_865
timestamp 1679585382
transform 1 0 83616 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_872
timestamp 1679585382
transform 1 0 84288 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_879
timestamp 1679585382
transform 1 0 84960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_886
timestamp 1679585382
transform 1 0 85632 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_893
timestamp 1679585382
transform 1 0 86304 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_900
timestamp 1679585382
transform 1 0 86976 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_907
timestamp 1679585382
transform 1 0 87648 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_914
timestamp 1679585382
transform 1 0 88320 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_921
timestamp 1679585382
transform 1 0 88992 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_928
timestamp 1679585382
transform 1 0 89664 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_935
timestamp 1679585382
transform 1 0 90336 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_942
timestamp 1679585382
transform 1 0 91008 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_949
timestamp 1679585382
transform 1 0 91680 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_956
timestamp 1679585382
transform 1 0 92352 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_963
timestamp 1679585382
transform 1 0 93024 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_970
timestamp 1679585382
transform 1 0 93696 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_977
timestamp 1679585382
transform 1 0 94368 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_984
timestamp 1679585382
transform 1 0 95040 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_991
timestamp 1679585382
transform 1 0 95712 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_998
timestamp 1679585382
transform 1 0 96384 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1005
timestamp 1679585382
transform 1 0 97056 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1012
timestamp 1679585382
transform 1 0 97728 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1019
timestamp 1679585382
transform 1 0 98400 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_1026
timestamp 1677583704
transform 1 0 99072 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_1028
timestamp 1677583258
transform 1 0 99264 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_4
timestamp 1679585382
transform 1 0 960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_11
timestamp 1679585382
transform 1 0 1632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_18
timestamp 1679585382
transform 1 0 2304 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_25
timestamp 1679585382
transform 1 0 2976 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_32
timestamp 1679585382
transform 1 0 3648 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_39
timestamp 1679585382
transform 1 0 4320 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_46
timestamp 1679585382
transform 1 0 4992 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_53
timestamp 1679585382
transform 1 0 5664 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_60
timestamp 1679585382
transform 1 0 6336 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_67
timestamp 1679585382
transform 1 0 7008 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_74
timestamp 1679585382
transform 1 0 7680 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_81
timestamp 1679585382
transform 1 0 8352 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_88
timestamp 1679585382
transform 1 0 9024 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_108
timestamp 1679585382
transform 1 0 10944 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_115
timestamp 1679585382
transform 1 0 11616 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_122
timestamp 1679585382
transform 1 0 12288 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_129
timestamp 1679585382
transform 1 0 12960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_149
timestamp 1679585382
transform 1 0 14880 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_156
timestamp 1679585382
transform 1 0 15552 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_163
timestamp 1679585382
transform 1 0 16224 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_170
timestamp 1679585382
transform 1 0 16896 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_177
timestamp 1679585382
transform 1 0 17568 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_184
timestamp 1679585382
transform 1 0 18240 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_191
timestamp 1679585382
transform 1 0 18912 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_198
timestamp 1679585382
transform 1 0 19584 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_205
timestamp 1679585382
transform 1 0 20256 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_212
timestamp 1679585382
transform 1 0 20928 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_219
timestamp 1679585382
transform 1 0 21600 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_226
timestamp 1679585382
transform 1 0 22272 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_233
timestamp 1679585382
transform 1 0 22944 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_240
timestamp 1679585382
transform 1 0 23616 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_247
timestamp 1679585382
transform 1 0 24288 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_254
timestamp 1679585382
transform 1 0 24960 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_261
timestamp 1677583704
transform 1 0 25632 0 1 20412
box -48 -56 240 834
use sg13g2_decap_4  FILLER_26_267
timestamp 1679581501
transform 1 0 26208 0 1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_26_271
timestamp 1677583704
transform 1 0 26592 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_282
timestamp 1679585382
transform 1 0 27648 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_289
timestamp 1679585382
transform 1 0 28320 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_296
timestamp 1679585382
transform 1 0 28992 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_303
timestamp 1679585382
transform 1 0 29664 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_310
timestamp 1679585382
transform 1 0 30336 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_317
timestamp 1679585382
transform 1 0 31008 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_324
timestamp 1679585382
transform 1 0 31680 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_331
timestamp 1679585382
transform 1 0 32352 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_338
timestamp 1679585382
transform 1 0 33024 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_345
timestamp 1679585382
transform 1 0 33696 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_352
timestamp 1679585382
transform 1 0 34368 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_359
timestamp 1679585382
transform 1 0 35040 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_366
timestamp 1679585382
transform 1 0 35712 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_373
timestamp 1679585382
transform 1 0 36384 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_380
timestamp 1679585382
transform 1 0 37056 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_387
timestamp 1679585382
transform 1 0 37728 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_394
timestamp 1679581501
transform 1 0 38400 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_398
timestamp 1677583258
transform 1 0 38784 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_417
timestamp 1679585382
transform 1 0 40608 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_424
timestamp 1679585382
transform 1 0 41280 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_431
timestamp 1679585382
transform 1 0 41952 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_438
timestamp 1679585382
transform 1 0 42624 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_445
timestamp 1679585382
transform 1 0 43296 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_452
timestamp 1679585382
transform 1 0 43968 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_459
timestamp 1679585382
transform 1 0 44640 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_466
timestamp 1679585382
transform 1 0 45312 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_473
timestamp 1679585382
transform 1 0 45984 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_480
timestamp 1679585382
transform 1 0 46656 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_487
timestamp 1679585382
transform 1 0 47328 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_494
timestamp 1679585382
transform 1 0 48000 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_501
timestamp 1679585382
transform 1 0 48672 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_508
timestamp 1679585382
transform 1 0 49344 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_515
timestamp 1679585382
transform 1 0 50016 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_522
timestamp 1679585382
transform 1 0 50688 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_529
timestamp 1679585382
transform 1 0 51360 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_536
timestamp 1679585382
transform 1 0 52032 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_543
timestamp 1679585382
transform 1 0 52704 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_550
timestamp 1679585382
transform 1 0 53376 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_557
timestamp 1679585382
transform 1 0 54048 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_564
timestamp 1679585382
transform 1 0 54720 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_571
timestamp 1679585382
transform 1 0 55392 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_578
timestamp 1679585382
transform 1 0 56064 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_585
timestamp 1679585382
transform 1 0 56736 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_592
timestamp 1679585382
transform 1 0 57408 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_599
timestamp 1679585382
transform 1 0 58080 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_606
timestamp 1679585382
transform 1 0 58752 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_613
timestamp 1679585382
transform 1 0 59424 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_620
timestamp 1679585382
transform 1 0 60096 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_627
timestamp 1679585382
transform 1 0 60768 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_634
timestamp 1679585382
transform 1 0 61440 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_641
timestamp 1679585382
transform 1 0 62112 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_648
timestamp 1679585382
transform 1 0 62784 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_655
timestamp 1679585382
transform 1 0 63456 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_662
timestamp 1679585382
transform 1 0 64128 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_669
timestamp 1679585382
transform 1 0 64800 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_676
timestamp 1679585382
transform 1 0 65472 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_683
timestamp 1679585382
transform 1 0 66144 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_690
timestamp 1679585382
transform 1 0 66816 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_697
timestamp 1679585382
transform 1 0 67488 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_704
timestamp 1679585382
transform 1 0 68160 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_711
timestamp 1679585382
transform 1 0 68832 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_718
timestamp 1679585382
transform 1 0 69504 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_725
timestamp 1679585382
transform 1 0 70176 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_732
timestamp 1679585382
transform 1 0 70848 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_739
timestamp 1679585382
transform 1 0 71520 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_746
timestamp 1679585382
transform 1 0 72192 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_753
timestamp 1679585382
transform 1 0 72864 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_760
timestamp 1679585382
transform 1 0 73536 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_767
timestamp 1679585382
transform 1 0 74208 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_774
timestamp 1679585382
transform 1 0 74880 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_781
timestamp 1679585382
transform 1 0 75552 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_788
timestamp 1679585382
transform 1 0 76224 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_795
timestamp 1679585382
transform 1 0 76896 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_802
timestamp 1679585382
transform 1 0 77568 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_809
timestamp 1679585382
transform 1 0 78240 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_816
timestamp 1679585382
transform 1 0 78912 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_823
timestamp 1679585382
transform 1 0 79584 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_830
timestamp 1679585382
transform 1 0 80256 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_837
timestamp 1679585382
transform 1 0 80928 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_844
timestamp 1679585382
transform 1 0 81600 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_851
timestamp 1679585382
transform 1 0 82272 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_858
timestamp 1679585382
transform 1 0 82944 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_865
timestamp 1679585382
transform 1 0 83616 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_872
timestamp 1679585382
transform 1 0 84288 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_879
timestamp 1679585382
transform 1 0 84960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_886
timestamp 1679585382
transform 1 0 85632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_893
timestamp 1679585382
transform 1 0 86304 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_900
timestamp 1679585382
transform 1 0 86976 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_907
timestamp 1679585382
transform 1 0 87648 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_914
timestamp 1679585382
transform 1 0 88320 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_921
timestamp 1679585382
transform 1 0 88992 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_928
timestamp 1679585382
transform 1 0 89664 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_935
timestamp 1679585382
transform 1 0 90336 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_942
timestamp 1679585382
transform 1 0 91008 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_949
timestamp 1679585382
transform 1 0 91680 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_956
timestamp 1679585382
transform 1 0 92352 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_963
timestamp 1679585382
transform 1 0 93024 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_970
timestamp 1679585382
transform 1 0 93696 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_977
timestamp 1679585382
transform 1 0 94368 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_984
timestamp 1679585382
transform 1 0 95040 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_991
timestamp 1679585382
transform 1 0 95712 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_998
timestamp 1679585382
transform 1 0 96384 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1005
timestamp 1679585382
transform 1 0 97056 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1012
timestamp 1679585382
transform 1 0 97728 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1019
timestamp 1679585382
transform 1 0 98400 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_1026
timestamp 1677583704
transform 1 0 99072 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_1028
timestamp 1677583258
transform 1 0 99264 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1679585382
transform 1 0 576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_7
timestamp 1679585382
transform 1 0 1248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_14
timestamp 1679585382
transform 1 0 1920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_48
timestamp 1679585382
transform 1 0 5184 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_55
timestamp 1679585382
transform 1 0 5856 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_62
timestamp 1679585382
transform 1 0 6528 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_69
timestamp 1679585382
transform 1 0 7200 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_76
timestamp 1679585382
transform 1 0 7872 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_83
timestamp 1679585382
transform 1 0 8544 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_90
timestamp 1679585382
transform 1 0 9216 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_97
timestamp 1679585382
transform 1 0 9888 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_104
timestamp 1679585382
transform 1 0 10560 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_111
timestamp 1679585382
transform 1 0 11232 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_118
timestamp 1679585382
transform 1 0 11904 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_125
timestamp 1679585382
transform 1 0 12576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_132
timestamp 1679585382
transform 1 0 13248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_139
timestamp 1679585382
transform 1 0 13920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_146
timestamp 1679581501
transform 1 0 14592 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_150
timestamp 1677583704
transform 1 0 14976 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_161
timestamp 1679585382
transform 1 0 16032 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_168
timestamp 1679585382
transform 1 0 16704 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_175
timestamp 1679585382
transform 1 0 17376 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_182
timestamp 1679585382
transform 1 0 18048 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_189
timestamp 1679585382
transform 1 0 18720 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_196
timestamp 1679585382
transform 1 0 19392 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_203
timestamp 1679585382
transform 1 0 20064 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_210
timestamp 1677583704
transform 1 0 20736 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_233
timestamp 1679585382
transform 1 0 22944 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_240
timestamp 1679585382
transform 1 0 23616 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_247
timestamp 1679585382
transform 1 0 24288 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_254
timestamp 1679585382
transform 1 0 24960 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_261
timestamp 1679585382
transform 1 0 25632 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_268
timestamp 1679585382
transform 1 0 26304 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_275
timestamp 1679585382
transform 1 0 26976 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_282
timestamp 1679585382
transform 1 0 27648 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_289
timestamp 1679585382
transform 1 0 28320 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_296
timestamp 1679585382
transform 1 0 28992 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_303
timestamp 1679581501
transform 1 0 29664 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_307
timestamp 1677583704
transform 1 0 30048 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_336
timestamp 1679585382
transform 1 0 32832 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_343
timestamp 1677583704
transform 1 0 33504 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_350
timestamp 1679585382
transform 1 0 34176 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_357
timestamp 1679585382
transform 1 0 34848 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_364
timestamp 1679585382
transform 1 0 35520 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_371
timestamp 1679585382
transform 1 0 36192 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_378
timestamp 1679581501
transform 1 0 36864 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_382
timestamp 1677583258
transform 1 0 37248 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_410
timestamp 1679585382
transform 1 0 39936 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_417
timestamp 1679585382
transform 1 0 40608 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_424
timestamp 1679585382
transform 1 0 41280 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_431
timestamp 1679585382
transform 1 0 41952 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_438
timestamp 1679585382
transform 1 0 42624 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_445
timestamp 1679585382
transform 1 0 43296 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_452
timestamp 1679585382
transform 1 0 43968 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_459
timestamp 1679585382
transform 1 0 44640 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_466
timestamp 1679585382
transform 1 0 45312 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_473
timestamp 1679585382
transform 1 0 45984 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_480
timestamp 1679585382
transform 1 0 46656 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_487
timestamp 1679585382
transform 1 0 47328 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_498
timestamp 1679581501
transform 1 0 48384 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_502
timestamp 1677583704
transform 1 0 48768 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_526
timestamp 1679585382
transform 1 0 51072 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_533
timestamp 1679585382
transform 1 0 51744 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_540
timestamp 1679585382
transform 1 0 52416 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_547
timestamp 1679585382
transform 1 0 53088 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_554
timestamp 1679585382
transform 1 0 53760 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_561
timestamp 1679585382
transform 1 0 54432 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_568
timestamp 1679585382
transform 1 0 55104 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_575
timestamp 1679585382
transform 1 0 55776 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_582
timestamp 1679585382
transform 1 0 56448 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_589
timestamp 1679585382
transform 1 0 57120 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_596
timestamp 1679585382
transform 1 0 57792 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_603
timestamp 1679585382
transform 1 0 58464 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_610
timestamp 1679585382
transform 1 0 59136 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_617
timestamp 1679585382
transform 1 0 59808 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_624
timestamp 1679585382
transform 1 0 60480 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_631
timestamp 1679585382
transform 1 0 61152 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_638
timestamp 1679585382
transform 1 0 61824 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_645
timestamp 1679585382
transform 1 0 62496 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_652
timestamp 1679585382
transform 1 0 63168 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_659
timestamp 1679585382
transform 1 0 63840 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_666
timestamp 1679585382
transform 1 0 64512 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_673
timestamp 1679585382
transform 1 0 65184 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_680
timestamp 1679585382
transform 1 0 65856 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_687
timestamp 1679585382
transform 1 0 66528 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_694
timestamp 1679585382
transform 1 0 67200 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_701
timestamp 1679585382
transform 1 0 67872 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_708
timestamp 1679585382
transform 1 0 68544 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_715
timestamp 1679585382
transform 1 0 69216 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_722
timestamp 1679585382
transform 1 0 69888 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_729
timestamp 1679585382
transform 1 0 70560 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_736
timestamp 1679585382
transform 1 0 71232 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_743
timestamp 1679585382
transform 1 0 71904 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_750
timestamp 1679585382
transform 1 0 72576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_757
timestamp 1679585382
transform 1 0 73248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_764
timestamp 1679585382
transform 1 0 73920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_771
timestamp 1679585382
transform 1 0 74592 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_778
timestamp 1679585382
transform 1 0 75264 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_785
timestamp 1679585382
transform 1 0 75936 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_792
timestamp 1679585382
transform 1 0 76608 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_799
timestamp 1679585382
transform 1 0 77280 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_806
timestamp 1679585382
transform 1 0 77952 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_813
timestamp 1679585382
transform 1 0 78624 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_820
timestamp 1679585382
transform 1 0 79296 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_827
timestamp 1679585382
transform 1 0 79968 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_834
timestamp 1679585382
transform 1 0 80640 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_841
timestamp 1679585382
transform 1 0 81312 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_848
timestamp 1679585382
transform 1 0 81984 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_855
timestamp 1679585382
transform 1 0 82656 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_862
timestamp 1679585382
transform 1 0 83328 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_869
timestamp 1679585382
transform 1 0 84000 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_876
timestamp 1679585382
transform 1 0 84672 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_883
timestamp 1679585382
transform 1 0 85344 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_890
timestamp 1679585382
transform 1 0 86016 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_897
timestamp 1679585382
transform 1 0 86688 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_904
timestamp 1679585382
transform 1 0 87360 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_911
timestamp 1679585382
transform 1 0 88032 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_918
timestamp 1679585382
transform 1 0 88704 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_925
timestamp 1679585382
transform 1 0 89376 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_932
timestamp 1679585382
transform 1 0 90048 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_939
timestamp 1679585382
transform 1 0 90720 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_946
timestamp 1679585382
transform 1 0 91392 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_953
timestamp 1679585382
transform 1 0 92064 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_960
timestamp 1679585382
transform 1 0 92736 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_967
timestamp 1679585382
transform 1 0 93408 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_974
timestamp 1679585382
transform 1 0 94080 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_981
timestamp 1679585382
transform 1 0 94752 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_988
timestamp 1679585382
transform 1 0 95424 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_995
timestamp 1679585382
transform 1 0 96096 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1002
timestamp 1679585382
transform 1 0 96768 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1009
timestamp 1679585382
transform 1 0 97440 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1016
timestamp 1679585382
transform 1 0 98112 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_1023
timestamp 1679581501
transform 1 0 98784 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_1027
timestamp 1677583704
transform 1 0 99168 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_4
timestamp 1679585382
transform 1 0 960 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_11
timestamp 1679585382
transform 1 0 1632 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_18
timestamp 1679585382
transform 1 0 2304 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_25
timestamp 1679581501
transform 1 0 2976 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_33
timestamp 1677583704
transform 1 0 3744 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_35
timestamp 1677583258
transform 1 0 3936 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_49
timestamp 1679585382
transform 1 0 5280 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_56
timestamp 1679585382
transform 1 0 5952 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_63
timestamp 1679585382
transform 1 0 6624 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_70
timestamp 1679585382
transform 1 0 7296 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_77
timestamp 1679585382
transform 1 0 7968 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_84
timestamp 1679585382
transform 1 0 8640 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_91
timestamp 1679585382
transform 1 0 9312 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_98
timestamp 1679585382
transform 1 0 9984 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_105
timestamp 1679581501
transform 1 0 10656 0 1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_28_117
timestamp 1679585382
transform 1 0 11808 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_124
timestamp 1679585382
transform 1 0 12480 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_131
timestamp 1679585382
transform 1 0 13152 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_142
timestamp 1677583704
transform 1 0 14208 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_188
timestamp 1679585382
transform 1 0 18624 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_195
timestamp 1679581501
transform 1 0 19296 0 1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_28_239
timestamp 1679585382
transform 1 0 23520 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_246
timestamp 1679585382
transform 1 0 24192 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_253
timestamp 1679585382
transform 1 0 24864 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_260
timestamp 1679585382
transform 1 0 25536 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_267
timestamp 1679585382
transform 1 0 26208 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_274
timestamp 1679585382
transform 1 0 26880 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_281
timestamp 1679581501
transform 1 0 27552 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_285
timestamp 1677583704
transform 1 0 27936 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_314
timestamp 1677583258
transform 1 0 30720 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_355
timestamp 1679585382
transform 1 0 34656 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_362
timestamp 1679585382
transform 1 0 35328 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_369
timestamp 1679585382
transform 1 0 36000 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_376
timestamp 1679585382
transform 1 0 36672 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_383
timestamp 1679585382
transform 1 0 37344 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_390
timestamp 1679585382
transform 1 0 38016 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_397
timestamp 1679585382
transform 1 0 38688 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_404
timestamp 1679585382
transform 1 0 39360 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_411
timestamp 1679585382
transform 1 0 40032 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_418
timestamp 1679585382
transform 1 0 40704 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_425
timestamp 1679585382
transform 1 0 41376 0 1 21924
box -48 -56 720 834
use sg13g2_fill_1  FILLER_28_432
timestamp 1677583258
transform 1 0 42048 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_464
timestamp 1679585382
transform 1 0 45120 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_471
timestamp 1679585382
transform 1 0 45792 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_478
timestamp 1679585382
transform 1 0 46464 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_525
timestamp 1679585382
transform 1 0 50976 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_532
timestamp 1679585382
transform 1 0 51648 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_539
timestamp 1679585382
transform 1 0 52320 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_546
timestamp 1679585382
transform 1 0 52992 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_553
timestamp 1679585382
transform 1 0 53664 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_560
timestamp 1679585382
transform 1 0 54336 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_567
timestamp 1679585382
transform 1 0 55008 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_574
timestamp 1679585382
transform 1 0 55680 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_581
timestamp 1679585382
transform 1 0 56352 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_588
timestamp 1679585382
transform 1 0 57024 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_595
timestamp 1679585382
transform 1 0 57696 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_602
timestamp 1679585382
transform 1 0 58368 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_609
timestamp 1679585382
transform 1 0 59040 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_616
timestamp 1679585382
transform 1 0 59712 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_623
timestamp 1679585382
transform 1 0 60384 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_630
timestamp 1679585382
transform 1 0 61056 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_637
timestamp 1679585382
transform 1 0 61728 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_644
timestamp 1679585382
transform 1 0 62400 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_651
timestamp 1679585382
transform 1 0 63072 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_658
timestamp 1679585382
transform 1 0 63744 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_665
timestamp 1679585382
transform 1 0 64416 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_672
timestamp 1679585382
transform 1 0 65088 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_679
timestamp 1679585382
transform 1 0 65760 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_686
timestamp 1679585382
transform 1 0 66432 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_693
timestamp 1679585382
transform 1 0 67104 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_700
timestamp 1679585382
transform 1 0 67776 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_707
timestamp 1679585382
transform 1 0 68448 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_714
timestamp 1679585382
transform 1 0 69120 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_721
timestamp 1679585382
transform 1 0 69792 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_728
timestamp 1679585382
transform 1 0 70464 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_735
timestamp 1679585382
transform 1 0 71136 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_742
timestamp 1679585382
transform 1 0 71808 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_749
timestamp 1679585382
transform 1 0 72480 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_756
timestamp 1679585382
transform 1 0 73152 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_763
timestamp 1679585382
transform 1 0 73824 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_770
timestamp 1679585382
transform 1 0 74496 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_777
timestamp 1679585382
transform 1 0 75168 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_784
timestamp 1679585382
transform 1 0 75840 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_791
timestamp 1679585382
transform 1 0 76512 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_798
timestamp 1679585382
transform 1 0 77184 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_805
timestamp 1679585382
transform 1 0 77856 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_812
timestamp 1679585382
transform 1 0 78528 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_819
timestamp 1679585382
transform 1 0 79200 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_826
timestamp 1679585382
transform 1 0 79872 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_833
timestamp 1679585382
transform 1 0 80544 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_840
timestamp 1679585382
transform 1 0 81216 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_847
timestamp 1679585382
transform 1 0 81888 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_854
timestamp 1679585382
transform 1 0 82560 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_861
timestamp 1679585382
transform 1 0 83232 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_868
timestamp 1679585382
transform 1 0 83904 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_875
timestamp 1679585382
transform 1 0 84576 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_882
timestamp 1679585382
transform 1 0 85248 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_889
timestamp 1679585382
transform 1 0 85920 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_896
timestamp 1679585382
transform 1 0 86592 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_903
timestamp 1679585382
transform 1 0 87264 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_910
timestamp 1679585382
transform 1 0 87936 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_917
timestamp 1679585382
transform 1 0 88608 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_924
timestamp 1679585382
transform 1 0 89280 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_931
timestamp 1679585382
transform 1 0 89952 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_938
timestamp 1679585382
transform 1 0 90624 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_945
timestamp 1679585382
transform 1 0 91296 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_952
timestamp 1679585382
transform 1 0 91968 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_959
timestamp 1679585382
transform 1 0 92640 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_966
timestamp 1679585382
transform 1 0 93312 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_973
timestamp 1679585382
transform 1 0 93984 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_980
timestamp 1679585382
transform 1 0 94656 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_987
timestamp 1679585382
transform 1 0 95328 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_994
timestamp 1679585382
transform 1 0 96000 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1001
timestamp 1679585382
transform 1 0 96672 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1008
timestamp 1679585382
transform 1 0 97344 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1015
timestamp 1679585382
transform 1 0 98016 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1022
timestamp 1679585382
transform 1 0 98688 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_0
timestamp 1679585382
transform 1 0 576 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_7
timestamp 1679585382
transform 1 0 1248 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_14
timestamp 1679585382
transform 1 0 1920 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_61
timestamp 1679585382
transform 1 0 6432 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_29_68
timestamp 1679581501
transform 1 0 7104 0 -1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_29_99
timestamp 1679585382
transform 1 0 10080 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_106
timestamp 1679585382
transform 1 0 10752 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_113
timestamp 1679585382
transform 1 0 11424 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_120
timestamp 1679585382
transform 1 0 12096 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_144
timestamp 1679585382
transform 1 0 14400 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_151
timestamp 1679585382
transform 1 0 15072 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_158
timestamp 1679585382
transform 1 0 15744 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_165
timestamp 1679585382
transform 1 0 16416 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_172
timestamp 1679585382
transform 1 0 17088 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_179
timestamp 1679585382
transform 1 0 17760 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_29_186
timestamp 1677583258
transform 1 0 18432 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_195
timestamp 1677583704
transform 1 0 19296 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_206
timestamp 1679585382
transform 1 0 20352 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_29_213
timestamp 1679581501
transform 1 0 21024 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_29_217
timestamp 1677583258
transform 1 0 21408 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_235
timestamp 1679585382
transform 1 0 23136 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_242
timestamp 1679585382
transform 1 0 23808 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_249
timestamp 1677583704
transform 1 0 24480 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_251
timestamp 1677583258
transform 1 0 24672 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_278
timestamp 1679585382
transform 1 0 27264 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_285
timestamp 1679585382
transform 1 0 27936 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_29_292
timestamp 1677583258
transform 1 0 28608 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_306
timestamp 1679585382
transform 1 0 29952 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_313
timestamp 1679585382
transform 1 0 30624 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_320
timestamp 1677583704
transform 1 0 31296 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_322
timestamp 1677583258
transform 1 0 31488 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_327
timestamp 1677583704
transform 1 0 31968 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_329
timestamp 1677583258
transform 1 0 32160 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_356
timestamp 1679585382
transform 1 0 34752 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_363
timestamp 1679585382
transform 1 0 35424 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_370
timestamp 1679585382
transform 1 0 36096 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_377
timestamp 1679585382
transform 1 0 36768 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_384
timestamp 1679585382
transform 1 0 37440 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_29_391
timestamp 1679581501
transform 1 0 38112 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_29_395
timestamp 1677583704
transform 1 0 38496 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_402
timestamp 1679585382
transform 1 0 39168 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_409
timestamp 1679585382
transform 1 0 39840 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_416
timestamp 1679585382
transform 1 0 40512 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_423
timestamp 1679585382
transform 1 0 41184 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_430
timestamp 1679585382
transform 1 0 41856 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_29_437
timestamp 1677583258
transform 1 0 42528 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_474
timestamp 1679585382
transform 1 0 46080 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_481
timestamp 1679585382
transform 1 0 46752 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_29_488
timestamp 1679581501
transform 1 0 47424 0 -1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_29_519
timestamp 1679585382
transform 1 0 50400 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_526
timestamp 1679585382
transform 1 0 51072 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_533
timestamp 1679585382
transform 1 0 51744 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_540
timestamp 1679585382
transform 1 0 52416 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_547
timestamp 1679585382
transform 1 0 53088 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_554
timestamp 1679585382
transform 1 0 53760 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_561
timestamp 1679585382
transform 1 0 54432 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_568
timestamp 1679585382
transform 1 0 55104 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_575
timestamp 1679585382
transform 1 0 55776 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_582
timestamp 1679585382
transform 1 0 56448 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_589
timestamp 1679585382
transform 1 0 57120 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_596
timestamp 1679585382
transform 1 0 57792 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_603
timestamp 1679585382
transform 1 0 58464 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_610
timestamp 1679585382
transform 1 0 59136 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_617
timestamp 1679585382
transform 1 0 59808 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_624
timestamp 1679585382
transform 1 0 60480 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_631
timestamp 1679585382
transform 1 0 61152 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_638
timestamp 1679585382
transform 1 0 61824 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_645
timestamp 1679585382
transform 1 0 62496 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_652
timestamp 1679585382
transform 1 0 63168 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_659
timestamp 1679585382
transform 1 0 63840 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_666
timestamp 1679585382
transform 1 0 64512 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_673
timestamp 1679585382
transform 1 0 65184 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_680
timestamp 1679585382
transform 1 0 65856 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_687
timestamp 1679585382
transform 1 0 66528 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_694
timestamp 1679585382
transform 1 0 67200 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_701
timestamp 1679585382
transform 1 0 67872 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_708
timestamp 1679585382
transform 1 0 68544 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_715
timestamp 1679585382
transform 1 0 69216 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_722
timestamp 1679585382
transform 1 0 69888 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_729
timestamp 1679585382
transform 1 0 70560 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_736
timestamp 1679585382
transform 1 0 71232 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_743
timestamp 1679585382
transform 1 0 71904 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_750
timestamp 1679585382
transform 1 0 72576 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_757
timestamp 1679585382
transform 1 0 73248 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_764
timestamp 1679585382
transform 1 0 73920 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_771
timestamp 1679585382
transform 1 0 74592 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_778
timestamp 1679585382
transform 1 0 75264 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_785
timestamp 1679585382
transform 1 0 75936 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_792
timestamp 1679585382
transform 1 0 76608 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_799
timestamp 1679585382
transform 1 0 77280 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_806
timestamp 1679585382
transform 1 0 77952 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_813
timestamp 1679585382
transform 1 0 78624 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_820
timestamp 1679585382
transform 1 0 79296 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_827
timestamp 1679585382
transform 1 0 79968 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_834
timestamp 1679585382
transform 1 0 80640 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_841
timestamp 1679585382
transform 1 0 81312 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_848
timestamp 1679585382
transform 1 0 81984 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_855
timestamp 1679585382
transform 1 0 82656 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_862
timestamp 1679585382
transform 1 0 83328 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_869
timestamp 1679585382
transform 1 0 84000 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_876
timestamp 1679585382
transform 1 0 84672 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_883
timestamp 1679585382
transform 1 0 85344 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_890
timestamp 1679585382
transform 1 0 86016 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_897
timestamp 1679585382
transform 1 0 86688 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_904
timestamp 1679585382
transform 1 0 87360 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_911
timestamp 1679585382
transform 1 0 88032 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_918
timestamp 1679585382
transform 1 0 88704 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_925
timestamp 1679585382
transform 1 0 89376 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_932
timestamp 1679585382
transform 1 0 90048 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_939
timestamp 1679585382
transform 1 0 90720 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_946
timestamp 1679585382
transform 1 0 91392 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_953
timestamp 1679585382
transform 1 0 92064 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_960
timestamp 1679585382
transform 1 0 92736 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_967
timestamp 1679585382
transform 1 0 93408 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_974
timestamp 1679585382
transform 1 0 94080 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_981
timestamp 1679585382
transform 1 0 94752 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_988
timestamp 1679585382
transform 1 0 95424 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_995
timestamp 1679585382
transform 1 0 96096 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1002
timestamp 1679585382
transform 1 0 96768 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1009
timestamp 1679585382
transform 1 0 97440 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1016
timestamp 1679585382
transform 1 0 98112 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_29_1023
timestamp 1679581501
transform 1 0 98784 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_29_1027
timestamp 1677583704
transform 1 0 99168 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_0
timestamp 1679585382
transform 1 0 576 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_7
timestamp 1679585382
transform 1 0 1248 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_14
timestamp 1679585382
transform 1 0 1920 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_21
timestamp 1679585382
transform 1 0 2592 0 1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_30_28
timestamp 1677583258
transform 1 0 3264 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_33
timestamp 1677583704
transform 1 0 3744 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_35
timestamp 1677583258
transform 1 0 3936 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_49
timestamp 1679585382
transform 1 0 5280 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_56
timestamp 1679585382
transform 1 0 5952 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_63
timestamp 1679585382
transform 1 0 6624 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_70
timestamp 1679585382
transform 1 0 7296 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_77
timestamp 1679585382
transform 1 0 7968 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_84
timestamp 1679581501
transform 1 0 8640 0 1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_30_115
timestamp 1679585382
transform 1 0 11616 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_122
timestamp 1679585382
transform 1 0 12288 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_129
timestamp 1679581501
transform 1 0 12960 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_133
timestamp 1677583258
transform 1 0 13344 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_170
timestamp 1679585382
transform 1 0 16896 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_177
timestamp 1679585382
transform 1 0 17568 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_184
timestamp 1679581501
transform 1 0 18240 0 1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_30_197
timestamp 1679585382
transform 1 0 19488 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_204
timestamp 1679585382
transform 1 0 20160 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_211
timestamp 1679585382
transform 1 0 20832 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_218
timestamp 1679585382
transform 1 0 21504 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_225
timestamp 1679585382
transform 1 0 22176 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_232
timestamp 1679585382
transform 1 0 22848 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_239
timestamp 1679585382
transform 1 0 23520 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_246
timestamp 1679585382
transform 1 0 24192 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_253
timestamp 1679585382
transform 1 0 24864 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_260
timestamp 1679585382
transform 1 0 25536 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_267
timestamp 1679585382
transform 1 0 26208 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_274
timestamp 1679585382
transform 1 0 26880 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_281
timestamp 1679585382
transform 1 0 27552 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_288
timestamp 1679585382
transform 1 0 28224 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_295
timestamp 1679585382
transform 1 0 28896 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_302
timestamp 1679585382
transform 1 0 29568 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_309
timestamp 1679585382
transform 1 0 30240 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_316
timestamp 1679585382
transform 1 0 30912 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_323
timestamp 1679585382
transform 1 0 31584 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_330
timestamp 1679585382
transform 1 0 32256 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_337
timestamp 1679585382
transform 1 0 32928 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_344
timestamp 1679585382
transform 1 0 33600 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_351
timestamp 1679585382
transform 1 0 34272 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_358
timestamp 1679585382
transform 1 0 34944 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_365
timestamp 1679585382
transform 1 0 35616 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_372
timestamp 1679581501
transform 1 0 36288 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_376
timestamp 1677583258
transform 1 0 36672 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_404
timestamp 1679585382
transform 1 0 39360 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_411
timestamp 1679585382
transform 1 0 40032 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_418
timestamp 1679585382
transform 1 0 40704 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_425
timestamp 1679585382
transform 1 0 41376 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_432
timestamp 1679585382
transform 1 0 42048 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_447
timestamp 1677583704
transform 1 0 43488 0 1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_458
timestamp 1679585382
transform 1 0 44544 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_465
timestamp 1679585382
transform 1 0 45216 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_472
timestamp 1679585382
transform 1 0 45888 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_479
timestamp 1679585382
transform 1 0 46560 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_486
timestamp 1679585382
transform 1 0 47232 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_493
timestamp 1679585382
transform 1 0 47904 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_500
timestamp 1679585382
transform 1 0 48576 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_507
timestamp 1679585382
transform 1 0 49248 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_514
timestamp 1679585382
transform 1 0 49920 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_521
timestamp 1679585382
transform 1 0 50592 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_528
timestamp 1679585382
transform 1 0 51264 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_535
timestamp 1679585382
transform 1 0 51936 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_542
timestamp 1679585382
transform 1 0 52608 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_549
timestamp 1679585382
transform 1 0 53280 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_556
timestamp 1679585382
transform 1 0 53952 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_563
timestamp 1679585382
transform 1 0 54624 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_570
timestamp 1679585382
transform 1 0 55296 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_577
timestamp 1679585382
transform 1 0 55968 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_584
timestamp 1679585382
transform 1 0 56640 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_591
timestamp 1679585382
transform 1 0 57312 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_598
timestamp 1679585382
transform 1 0 57984 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_605
timestamp 1679585382
transform 1 0 58656 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_612
timestamp 1679585382
transform 1 0 59328 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_619
timestamp 1679585382
transform 1 0 60000 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_626
timestamp 1679585382
transform 1 0 60672 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_633
timestamp 1679585382
transform 1 0 61344 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_640
timestamp 1679585382
transform 1 0 62016 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_647
timestamp 1679585382
transform 1 0 62688 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_654
timestamp 1679585382
transform 1 0 63360 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_661
timestamp 1679585382
transform 1 0 64032 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_668
timestamp 1679585382
transform 1 0 64704 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_675
timestamp 1679585382
transform 1 0 65376 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_682
timestamp 1679585382
transform 1 0 66048 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_689
timestamp 1679585382
transform 1 0 66720 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_696
timestamp 1679585382
transform 1 0 67392 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_703
timestamp 1679585382
transform 1 0 68064 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_710
timestamp 1679585382
transform 1 0 68736 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_717
timestamp 1679585382
transform 1 0 69408 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_724
timestamp 1679585382
transform 1 0 70080 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_731
timestamp 1679585382
transform 1 0 70752 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_738
timestamp 1679585382
transform 1 0 71424 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_745
timestamp 1679585382
transform 1 0 72096 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_752
timestamp 1679585382
transform 1 0 72768 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_759
timestamp 1679585382
transform 1 0 73440 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_766
timestamp 1679585382
transform 1 0 74112 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_773
timestamp 1679585382
transform 1 0 74784 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_780
timestamp 1679585382
transform 1 0 75456 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_787
timestamp 1679585382
transform 1 0 76128 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_794
timestamp 1679585382
transform 1 0 76800 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_801
timestamp 1679585382
transform 1 0 77472 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_808
timestamp 1679585382
transform 1 0 78144 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_815
timestamp 1679585382
transform 1 0 78816 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_822
timestamp 1679585382
transform 1 0 79488 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_829
timestamp 1679585382
transform 1 0 80160 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_836
timestamp 1679585382
transform 1 0 80832 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_843
timestamp 1679585382
transform 1 0 81504 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_850
timestamp 1679585382
transform 1 0 82176 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_857
timestamp 1679585382
transform 1 0 82848 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_864
timestamp 1679585382
transform 1 0 83520 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_871
timestamp 1679585382
transform 1 0 84192 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_878
timestamp 1679585382
transform 1 0 84864 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_885
timestamp 1679585382
transform 1 0 85536 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_892
timestamp 1679585382
transform 1 0 86208 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_899
timestamp 1679585382
transform 1 0 86880 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_906
timestamp 1679585382
transform 1 0 87552 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_913
timestamp 1679585382
transform 1 0 88224 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_920
timestamp 1679585382
transform 1 0 88896 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_927
timestamp 1679585382
transform 1 0 89568 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_934
timestamp 1679585382
transform 1 0 90240 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_941
timestamp 1679585382
transform 1 0 90912 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_948
timestamp 1679585382
transform 1 0 91584 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_955
timestamp 1679585382
transform 1 0 92256 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_962
timestamp 1679585382
transform 1 0 92928 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_969
timestamp 1679585382
transform 1 0 93600 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_976
timestamp 1679585382
transform 1 0 94272 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_983
timestamp 1679585382
transform 1 0 94944 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_990
timestamp 1679585382
transform 1 0 95616 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_997
timestamp 1679585382
transform 1 0 96288 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1004
timestamp 1679585382
transform 1 0 96960 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1011
timestamp 1679585382
transform 1 0 97632 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1018
timestamp 1679585382
transform 1 0 98304 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_1025
timestamp 1679581501
transform 1 0 98976 0 1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_31_0
timestamp 1679585382
transform 1 0 576 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_7
timestamp 1679585382
transform 1 0 1248 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_14
timestamp 1679585382
transform 1 0 1920 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_21
timestamp 1679585382
transform 1 0 2592 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_28
timestamp 1679585382
transform 1 0 3264 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_35
timestamp 1679585382
transform 1 0 3936 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_42
timestamp 1679585382
transform 1 0 4608 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_49
timestamp 1679585382
transform 1 0 5280 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_56
timestamp 1679585382
transform 1 0 5952 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_63
timestamp 1679585382
transform 1 0 6624 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_70
timestamp 1679585382
transform 1 0 7296 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_77
timestamp 1679585382
transform 1 0 7968 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_84
timestamp 1679585382
transform 1 0 8640 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_91
timestamp 1679585382
transform 1 0 9312 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_98
timestamp 1679585382
transform 1 0 9984 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_105
timestamp 1679585382
transform 1 0 10656 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_112
timestamp 1679585382
transform 1 0 11328 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_119
timestamp 1679585382
transform 1 0 12000 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_126
timestamp 1679585382
transform 1 0 12672 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_133
timestamp 1679585382
transform 1 0 13344 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_140
timestamp 1679585382
transform 1 0 14016 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_147
timestamp 1679585382
transform 1 0 14688 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_154
timestamp 1679585382
transform 1 0 15360 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_161
timestamp 1679585382
transform 1 0 16032 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_168
timestamp 1679585382
transform 1 0 16704 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_175
timestamp 1679585382
transform 1 0 17376 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_182
timestamp 1677583704
transform 1 0 18048 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_184
timestamp 1677583258
transform 1 0 18240 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_189
timestamp 1679585382
transform 1 0 18720 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_196
timestamp 1679585382
transform 1 0 19392 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_203
timestamp 1679585382
transform 1 0 20064 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_210
timestamp 1679585382
transform 1 0 20736 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_217
timestamp 1679585382
transform 1 0 21408 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_224
timestamp 1679585382
transform 1 0 22080 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_231
timestamp 1679585382
transform 1 0 22752 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_238
timestamp 1679585382
transform 1 0 23424 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_245
timestamp 1679585382
transform 1 0 24096 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_252
timestamp 1679585382
transform 1 0 24768 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_259
timestamp 1679585382
transform 1 0 25440 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_266
timestamp 1679585382
transform 1 0 26112 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_273
timestamp 1679585382
transform 1 0 26784 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_280
timestamp 1679585382
transform 1 0 27456 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_287
timestamp 1679585382
transform 1 0 28128 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_294
timestamp 1679585382
transform 1 0 28800 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_301
timestamp 1679585382
transform 1 0 29472 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_308
timestamp 1679585382
transform 1 0 30144 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_315
timestamp 1679585382
transform 1 0 30816 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_322
timestamp 1677583704
transform 1 0 31488 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_324
timestamp 1677583258
transform 1 0 31680 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_350
timestamp 1679585382
transform 1 0 34176 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_357
timestamp 1679585382
transform 1 0 34848 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_364
timestamp 1679585382
transform 1 0 35520 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_371
timestamp 1679585382
transform 1 0 36192 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_378
timestamp 1679585382
transform 1 0 36864 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_385
timestamp 1677583258
transform 1 0 37536 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_390
timestamp 1679581501
transform 1 0 38016 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_394
timestamp 1677583704
transform 1 0 38400 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_405
timestamp 1679585382
transform 1 0 39456 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_412
timestamp 1679585382
transform 1 0 40128 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_419
timestamp 1679585382
transform 1 0 40800 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_426
timestamp 1679585382
transform 1 0 41472 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_433
timestamp 1677583258
transform 1 0 42144 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_447
timestamp 1679585382
transform 1 0 43488 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_454
timestamp 1679585382
transform 1 0 44160 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_461
timestamp 1679585382
transform 1 0 44832 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_468
timestamp 1679585382
transform 1 0 45504 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_475
timestamp 1679585382
transform 1 0 46176 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_482
timestamp 1679585382
transform 1 0 46848 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_489
timestamp 1679585382
transform 1 0 47520 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_496
timestamp 1679585382
transform 1 0 48192 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_503
timestamp 1679585382
transform 1 0 48864 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_510
timestamp 1679585382
transform 1 0 49536 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_517
timestamp 1679585382
transform 1 0 50208 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_524
timestamp 1679585382
transform 1 0 50880 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_531
timestamp 1679585382
transform 1 0 51552 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_538
timestamp 1679585382
transform 1 0 52224 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_545
timestamp 1679585382
transform 1 0 52896 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_552
timestamp 1679585382
transform 1 0 53568 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_559
timestamp 1679585382
transform 1 0 54240 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_566
timestamp 1679585382
transform 1 0 54912 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_573
timestamp 1679585382
transform 1 0 55584 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_580
timestamp 1679585382
transform 1 0 56256 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_587
timestamp 1679585382
transform 1 0 56928 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_594
timestamp 1679585382
transform 1 0 57600 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_601
timestamp 1679585382
transform 1 0 58272 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_608
timestamp 1679585382
transform 1 0 58944 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_615
timestamp 1679585382
transform 1 0 59616 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_622
timestamp 1679585382
transform 1 0 60288 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_629
timestamp 1679585382
transform 1 0 60960 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_636
timestamp 1679585382
transform 1 0 61632 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_643
timestamp 1679585382
transform 1 0 62304 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_650
timestamp 1679585382
transform 1 0 62976 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_657
timestamp 1679585382
transform 1 0 63648 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_664
timestamp 1679585382
transform 1 0 64320 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_671
timestamp 1679585382
transform 1 0 64992 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_678
timestamp 1679585382
transform 1 0 65664 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_685
timestamp 1679585382
transform 1 0 66336 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_692
timestamp 1679585382
transform 1 0 67008 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_699
timestamp 1679585382
transform 1 0 67680 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_706
timestamp 1679585382
transform 1 0 68352 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_713
timestamp 1679585382
transform 1 0 69024 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_720
timestamp 1679585382
transform 1 0 69696 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_727
timestamp 1679585382
transform 1 0 70368 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_734
timestamp 1679585382
transform 1 0 71040 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_741
timestamp 1679585382
transform 1 0 71712 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_748
timestamp 1679585382
transform 1 0 72384 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_755
timestamp 1679585382
transform 1 0 73056 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_762
timestamp 1679585382
transform 1 0 73728 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_769
timestamp 1679585382
transform 1 0 74400 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_776
timestamp 1679585382
transform 1 0 75072 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_783
timestamp 1679585382
transform 1 0 75744 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_790
timestamp 1679585382
transform 1 0 76416 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_797
timestamp 1679585382
transform 1 0 77088 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_804
timestamp 1679585382
transform 1 0 77760 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_811
timestamp 1679585382
transform 1 0 78432 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_818
timestamp 1679585382
transform 1 0 79104 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_825
timestamp 1679585382
transform 1 0 79776 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_832
timestamp 1679585382
transform 1 0 80448 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_839
timestamp 1679585382
transform 1 0 81120 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_846
timestamp 1679585382
transform 1 0 81792 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_853
timestamp 1679585382
transform 1 0 82464 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_860
timestamp 1679585382
transform 1 0 83136 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_867
timestamp 1679585382
transform 1 0 83808 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_874
timestamp 1679585382
transform 1 0 84480 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_881
timestamp 1679585382
transform 1 0 85152 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_888
timestamp 1679585382
transform 1 0 85824 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_895
timestamp 1679585382
transform 1 0 86496 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_902
timestamp 1679585382
transform 1 0 87168 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_909
timestamp 1679585382
transform 1 0 87840 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_916
timestamp 1679585382
transform 1 0 88512 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_923
timestamp 1679585382
transform 1 0 89184 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_930
timestamp 1679585382
transform 1 0 89856 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_937
timestamp 1679585382
transform 1 0 90528 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_944
timestamp 1679585382
transform 1 0 91200 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_951
timestamp 1679585382
transform 1 0 91872 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_958
timestamp 1679585382
transform 1 0 92544 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_965
timestamp 1679585382
transform 1 0 93216 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_972
timestamp 1679585382
transform 1 0 93888 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_979
timestamp 1679585382
transform 1 0 94560 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_986
timestamp 1679585382
transform 1 0 95232 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_993
timestamp 1679585382
transform 1 0 95904 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1000
timestamp 1679585382
transform 1 0 96576 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1007
timestamp 1679585382
transform 1 0 97248 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1014
timestamp 1679585382
transform 1 0 97920 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1021
timestamp 1679585382
transform 1 0 98592 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_1028
timestamp 1677583258
transform 1 0 99264 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_0
timestamp 1679585382
transform 1 0 576 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_7
timestamp 1679585382
transform 1 0 1248 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_14
timestamp 1679581501
transform 1 0 1920 0 1 24948
box -48 -56 432 834
use sg13g2_decap_8  FILLER_32_45
timestamp 1679585382
transform 1 0 4896 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_52
timestamp 1679585382
transform 1 0 5568 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_59
timestamp 1679585382
transform 1 0 6240 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_66
timestamp 1679585382
transform 1 0 6912 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_73
timestamp 1679585382
transform 1 0 7584 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_80
timestamp 1679585382
transform 1 0 8256 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_87
timestamp 1679585382
transform 1 0 8928 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_94
timestamp 1679585382
transform 1 0 9600 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_101
timestamp 1679585382
transform 1 0 10272 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_108
timestamp 1679585382
transform 1 0 10944 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_115
timestamp 1679585382
transform 1 0 11616 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_122
timestamp 1679585382
transform 1 0 12288 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_129
timestamp 1679585382
transform 1 0 12960 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_136
timestamp 1679585382
transform 1 0 13632 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_143
timestamp 1679585382
transform 1 0 14304 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_150
timestamp 1679585382
transform 1 0 14976 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_157
timestamp 1679585382
transform 1 0 15648 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_164
timestamp 1679581501
transform 1 0 16320 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_176
timestamp 1677583258
transform 1 0 17472 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_194
timestamp 1677583704
transform 1 0 19200 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_200
timestamp 1679585382
transform 1 0 19776 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_207
timestamp 1679585382
transform 1 0 20448 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_214
timestamp 1679585382
transform 1 0 21120 0 1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_32_230
timestamp 1677583258
transform 1 0 22656 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_267
timestamp 1679585382
transform 1 0 26208 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_274
timestamp 1679585382
transform 1 0 26880 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_281
timestamp 1679585382
transform 1 0 27552 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_288
timestamp 1679585382
transform 1 0 28224 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_295
timestamp 1679585382
transform 1 0 28896 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_302
timestamp 1679585382
transform 1 0 29568 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_309
timestamp 1679585382
transform 1 0 30240 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_316
timestamp 1679585382
transform 1 0 30912 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_323
timestamp 1677583704
transform 1 0 31584 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_329
timestamp 1679585382
transform 1 0 32160 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_336
timestamp 1679585382
transform 1 0 32832 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_343
timestamp 1679581501
transform 1 0 33504 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_347
timestamp 1677583258
transform 1 0 33888 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_361
timestamp 1679585382
transform 1 0 35232 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_368
timestamp 1679585382
transform 1 0 35904 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_375
timestamp 1679585382
transform 1 0 36576 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_382
timestamp 1679585382
transform 1 0 37248 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_389
timestamp 1679585382
transform 1 0 37920 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_396
timestamp 1679585382
transform 1 0 38592 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_403
timestamp 1677583704
transform 1 0 39264 0 1 24948
box -48 -56 240 834
use sg13g2_decap_4  FILLER_32_409
timestamp 1679581501
transform 1 0 39840 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_421
timestamp 1677583704
transform 1 0 40992 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_431
timestamp 1679585382
transform 1 0 41952 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_438
timestamp 1679585382
transform 1 0 42624 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_445
timestamp 1679585382
transform 1 0 43296 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_452
timestamp 1679585382
transform 1 0 43968 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_459
timestamp 1679585382
transform 1 0 44640 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_466
timestamp 1679585382
transform 1 0 45312 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_473
timestamp 1679585382
transform 1 0 45984 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_480
timestamp 1679585382
transform 1 0 46656 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_487
timestamp 1679585382
transform 1 0 47328 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_494
timestamp 1679585382
transform 1 0 48000 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_501
timestamp 1679585382
transform 1 0 48672 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_508
timestamp 1679585382
transform 1 0 49344 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_515
timestamp 1679585382
transform 1 0 50016 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_522
timestamp 1679585382
transform 1 0 50688 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_529
timestamp 1679585382
transform 1 0 51360 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_536
timestamp 1679585382
transform 1 0 52032 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_543
timestamp 1679585382
transform 1 0 52704 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_550
timestamp 1679585382
transform 1 0 53376 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_557
timestamp 1679585382
transform 1 0 54048 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_564
timestamp 1679585382
transform 1 0 54720 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_571
timestamp 1679585382
transform 1 0 55392 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_578
timestamp 1679585382
transform 1 0 56064 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_585
timestamp 1679585382
transform 1 0 56736 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_592
timestamp 1679585382
transform 1 0 57408 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_599
timestamp 1679585382
transform 1 0 58080 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_606
timestamp 1679585382
transform 1 0 58752 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_613
timestamp 1679585382
transform 1 0 59424 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_620
timestamp 1679585382
transform 1 0 60096 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_627
timestamp 1679585382
transform 1 0 60768 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_634
timestamp 1679585382
transform 1 0 61440 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_641
timestamp 1679585382
transform 1 0 62112 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_648
timestamp 1679585382
transform 1 0 62784 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_655
timestamp 1679585382
transform 1 0 63456 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_662
timestamp 1679585382
transform 1 0 64128 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_669
timestamp 1679585382
transform 1 0 64800 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_676
timestamp 1679585382
transform 1 0 65472 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_683
timestamp 1679585382
transform 1 0 66144 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_690
timestamp 1679585382
transform 1 0 66816 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_697
timestamp 1679585382
transform 1 0 67488 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_704
timestamp 1679585382
transform 1 0 68160 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_711
timestamp 1679585382
transform 1 0 68832 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_718
timestamp 1679585382
transform 1 0 69504 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_725
timestamp 1679585382
transform 1 0 70176 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_732
timestamp 1679585382
transform 1 0 70848 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_739
timestamp 1679585382
transform 1 0 71520 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_746
timestamp 1679585382
transform 1 0 72192 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_753
timestamp 1679585382
transform 1 0 72864 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_760
timestamp 1679585382
transform 1 0 73536 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_767
timestamp 1679585382
transform 1 0 74208 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_774
timestamp 1679585382
transform 1 0 74880 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_781
timestamp 1679585382
transform 1 0 75552 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_788
timestamp 1679585382
transform 1 0 76224 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_795
timestamp 1679585382
transform 1 0 76896 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_802
timestamp 1679585382
transform 1 0 77568 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_809
timestamp 1679585382
transform 1 0 78240 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_816
timestamp 1679585382
transform 1 0 78912 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_823
timestamp 1679585382
transform 1 0 79584 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_830
timestamp 1679585382
transform 1 0 80256 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_837
timestamp 1679585382
transform 1 0 80928 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_844
timestamp 1679585382
transform 1 0 81600 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_851
timestamp 1679585382
transform 1 0 82272 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_858
timestamp 1679585382
transform 1 0 82944 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_865
timestamp 1679585382
transform 1 0 83616 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_872
timestamp 1679585382
transform 1 0 84288 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_879
timestamp 1679585382
transform 1 0 84960 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_886
timestamp 1679585382
transform 1 0 85632 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_893
timestamp 1679585382
transform 1 0 86304 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_900
timestamp 1679585382
transform 1 0 86976 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_907
timestamp 1679585382
transform 1 0 87648 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_914
timestamp 1679585382
transform 1 0 88320 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_921
timestamp 1679585382
transform 1 0 88992 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_928
timestamp 1679585382
transform 1 0 89664 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_935
timestamp 1679585382
transform 1 0 90336 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_942
timestamp 1679585382
transform 1 0 91008 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_949
timestamp 1679585382
transform 1 0 91680 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_956
timestamp 1679585382
transform 1 0 92352 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_963
timestamp 1679585382
transform 1 0 93024 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_970
timestamp 1679585382
transform 1 0 93696 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_977
timestamp 1679585382
transform 1 0 94368 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_984
timestamp 1679585382
transform 1 0 95040 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_991
timestamp 1679585382
transform 1 0 95712 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_998
timestamp 1679585382
transform 1 0 96384 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1005
timestamp 1679585382
transform 1 0 97056 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1012
timestamp 1679585382
transform 1 0 97728 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1019
timestamp 1679585382
transform 1 0 98400 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_1026
timestamp 1677583704
transform 1 0 99072 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_1028
timestamp 1677583258
transform 1 0 99264 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_0
timestamp 1679585382
transform 1 0 576 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_7
timestamp 1679585382
transform 1 0 1248 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_14
timestamp 1679585382
transform 1 0 1920 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_21
timestamp 1679581501
transform 1 0 2592 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_25
timestamp 1677583704
transform 1 0 2976 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_33_31
timestamp 1679581501
transform 1 0 3552 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_35
timestamp 1677583704
transform 1 0 3936 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_46
timestamp 1679585382
transform 1 0 4992 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_53
timestamp 1679585382
transform 1 0 5664 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_60
timestamp 1679585382
transform 1 0 6336 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_67
timestamp 1679585382
transform 1 0 7008 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_74
timestamp 1679585382
transform 1 0 7680 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_81
timestamp 1679585382
transform 1 0 8352 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_88
timestamp 1679585382
transform 1 0 9024 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_95
timestamp 1679585382
transform 1 0 9696 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_102
timestamp 1679585382
transform 1 0 10368 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_33_109
timestamp 1677583258
transform 1 0 11040 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_123
timestamp 1679585382
transform 1 0 12384 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_130
timestamp 1679585382
transform 1 0 13056 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_137
timestamp 1679585382
transform 1 0 13728 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_144
timestamp 1679585382
transform 1 0 14400 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_151
timestamp 1679585382
transform 1 0 15072 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_158
timestamp 1679585382
transform 1 0 15744 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_165
timestamp 1679585382
transform 1 0 16416 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_172
timestamp 1679585382
transform 1 0 17088 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_179
timestamp 1679585382
transform 1 0 17760 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_186
timestamp 1679581501
transform 1 0 18432 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_33_190
timestamp 1677583258
transform 1 0 18816 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_227
timestamp 1679585382
transform 1 0 22368 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_234
timestamp 1679581501
transform 1 0 23040 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_33_238
timestamp 1677583258
transform 1 0 23424 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_243
timestamp 1679585382
transform 1 0 23904 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_250
timestamp 1679585382
transform 1 0 24576 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_257
timestamp 1679585382
transform 1 0 25248 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_264
timestamp 1679585382
transform 1 0 25920 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_271
timestamp 1679585382
transform 1 0 26592 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_278
timestamp 1679585382
transform 1 0 27264 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_285
timestamp 1679585382
transform 1 0 27936 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_292
timestamp 1679585382
transform 1 0 28608 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_299
timestamp 1677583704
transform 1 0 29280 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_301
timestamp 1677583258
transform 1 0 29472 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_342
timestamp 1679585382
transform 1 0 33408 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_349
timestamp 1679581501
transform 1 0 34080 0 -1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_33_380
timestamp 1679585382
transform 1 0 37056 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_387
timestamp 1679581501
transform 1 0 37728 0 -1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_33_395
timestamp 1679585382
transform 1 0 38496 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_402
timestamp 1679585382
transform 1 0 39168 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_409
timestamp 1679585382
transform 1 0 39840 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_416
timestamp 1679585382
transform 1 0 40512 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_33_423
timestamp 1677583258
transform 1 0 41184 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_451
timestamp 1679585382
transform 1 0 43872 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_458
timestamp 1679585382
transform 1 0 44544 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_465
timestamp 1679581501
transform 1 0 45216 0 -1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_33_482
timestamp 1679585382
transform 1 0 46848 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_489
timestamp 1679585382
transform 1 0 47520 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_496
timestamp 1679585382
transform 1 0 48192 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_503
timestamp 1679585382
transform 1 0 48864 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_510
timestamp 1679585382
transform 1 0 49536 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_517
timestamp 1679585382
transform 1 0 50208 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_524
timestamp 1679585382
transform 1 0 50880 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_531
timestamp 1679585382
transform 1 0 51552 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_538
timestamp 1679585382
transform 1 0 52224 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_545
timestamp 1679585382
transform 1 0 52896 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_552
timestamp 1679585382
transform 1 0 53568 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_559
timestamp 1679585382
transform 1 0 54240 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_566
timestamp 1679585382
transform 1 0 54912 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_573
timestamp 1679585382
transform 1 0 55584 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_580
timestamp 1679585382
transform 1 0 56256 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_587
timestamp 1679585382
transform 1 0 56928 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_594
timestamp 1679585382
transform 1 0 57600 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_601
timestamp 1679585382
transform 1 0 58272 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_608
timestamp 1679585382
transform 1 0 58944 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_615
timestamp 1679585382
transform 1 0 59616 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_622
timestamp 1679585382
transform 1 0 60288 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_629
timestamp 1679585382
transform 1 0 60960 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_636
timestamp 1679585382
transform 1 0 61632 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_643
timestamp 1679585382
transform 1 0 62304 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_650
timestamp 1679585382
transform 1 0 62976 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_657
timestamp 1679585382
transform 1 0 63648 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_664
timestamp 1679585382
transform 1 0 64320 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_671
timestamp 1679585382
transform 1 0 64992 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_678
timestamp 1679585382
transform 1 0 65664 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_685
timestamp 1679585382
transform 1 0 66336 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_692
timestamp 1679585382
transform 1 0 67008 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_699
timestamp 1679585382
transform 1 0 67680 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_706
timestamp 1679585382
transform 1 0 68352 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_713
timestamp 1679585382
transform 1 0 69024 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_720
timestamp 1679585382
transform 1 0 69696 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_727
timestamp 1679585382
transform 1 0 70368 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_734
timestamp 1679585382
transform 1 0 71040 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_741
timestamp 1679585382
transform 1 0 71712 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_748
timestamp 1679585382
transform 1 0 72384 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_755
timestamp 1679585382
transform 1 0 73056 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_762
timestamp 1679585382
transform 1 0 73728 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_769
timestamp 1679585382
transform 1 0 74400 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_776
timestamp 1679585382
transform 1 0 75072 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_783
timestamp 1679585382
transform 1 0 75744 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_790
timestamp 1679585382
transform 1 0 76416 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_797
timestamp 1679585382
transform 1 0 77088 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_804
timestamp 1679585382
transform 1 0 77760 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_811
timestamp 1679585382
transform 1 0 78432 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_818
timestamp 1679585382
transform 1 0 79104 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_825
timestamp 1679585382
transform 1 0 79776 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_832
timestamp 1679585382
transform 1 0 80448 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_839
timestamp 1679585382
transform 1 0 81120 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_846
timestamp 1679585382
transform 1 0 81792 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_853
timestamp 1679585382
transform 1 0 82464 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_860
timestamp 1679585382
transform 1 0 83136 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_867
timestamp 1679585382
transform 1 0 83808 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_874
timestamp 1679585382
transform 1 0 84480 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_881
timestamp 1679585382
transform 1 0 85152 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_888
timestamp 1679585382
transform 1 0 85824 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_895
timestamp 1679585382
transform 1 0 86496 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_902
timestamp 1679585382
transform 1 0 87168 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_909
timestamp 1679585382
transform 1 0 87840 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_916
timestamp 1679585382
transform 1 0 88512 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_923
timestamp 1679585382
transform 1 0 89184 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_930
timestamp 1679585382
transform 1 0 89856 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_937
timestamp 1679585382
transform 1 0 90528 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_944
timestamp 1679585382
transform 1 0 91200 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_951
timestamp 1679585382
transform 1 0 91872 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_958
timestamp 1679585382
transform 1 0 92544 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_965
timestamp 1679585382
transform 1 0 93216 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_972
timestamp 1679585382
transform 1 0 93888 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_979
timestamp 1679585382
transform 1 0 94560 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_986
timestamp 1679585382
transform 1 0 95232 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_993
timestamp 1679585382
transform 1 0 95904 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1000
timestamp 1679585382
transform 1 0 96576 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1007
timestamp 1679585382
transform 1 0 97248 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1014
timestamp 1679585382
transform 1 0 97920 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1021
timestamp 1679585382
transform 1 0 98592 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_33_1028
timestamp 1677583258
transform 1 0 99264 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_0
timestamp 1679585382
transform 1 0 576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_7
timestamp 1679585382
transform 1 0 1248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_14
timestamp 1679585382
transform 1 0 1920 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_21
timestamp 1679585382
transform 1 0 2592 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_28
timestamp 1679585382
transform 1 0 3264 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_35
timestamp 1679581501
transform 1 0 3936 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_39
timestamp 1677583258
transform 1 0 4320 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_44
timestamp 1679585382
transform 1 0 4800 0 1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_34_51
timestamp 1677583258
transform 1 0 5472 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_61
timestamp 1679585382
transform 1 0 6432 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_68
timestamp 1679585382
transform 1 0 7104 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_75
timestamp 1679585382
transform 1 0 7776 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_82
timestamp 1679585382
transform 1 0 8448 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_102
timestamp 1679585382
transform 1 0 10368 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_109
timestamp 1679585382
transform 1 0 11040 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_116
timestamp 1679585382
transform 1 0 11712 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_123
timestamp 1677583704
transform 1 0 12384 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_125
timestamp 1677583258
transform 1 0 12576 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_180
timestamp 1679585382
transform 1 0 17856 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_187
timestamp 1679585382
transform 1 0 18528 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_194
timestamp 1677583704
transform 1 0 19200 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_196
timestamp 1677583258
transform 1 0 19392 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_210
timestamp 1679585382
transform 1 0 20736 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_217
timestamp 1679585382
transform 1 0 21408 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_224
timestamp 1679585382
transform 1 0 22080 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_231
timestamp 1679585382
transform 1 0 22752 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_238
timestamp 1679585382
transform 1 0 23424 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_245
timestamp 1679585382
transform 1 0 24096 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_252
timestamp 1679585382
transform 1 0 24768 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_259
timestamp 1679585382
transform 1 0 25440 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_266
timestamp 1679585382
transform 1 0 26112 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_273
timestamp 1679585382
transform 1 0 26784 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_280
timestamp 1677583704
transform 1 0 27456 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_282
timestamp 1677583258
transform 1 0 27648 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_310
timestamp 1679585382
transform 1 0 30336 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_317
timestamp 1679581501
transform 1 0 31008 0 1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_34_330
timestamp 1679585382
transform 1 0 32256 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_337
timestamp 1679585382
transform 1 0 32928 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_344
timestamp 1679585382
transform 1 0 33600 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_351
timestamp 1679585382
transform 1 0 34272 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_358
timestamp 1679585382
transform 1 0 34944 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_365
timestamp 1679585382
transform 1 0 35616 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_372
timestamp 1679585382
transform 1 0 36288 0 1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_34_379
timestamp 1677583258
transform 1 0 36960 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_416
timestamp 1679585382
transform 1 0 40512 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_423
timestamp 1679585382
transform 1 0 41184 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_430
timestamp 1679585382
transform 1 0 41856 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_437
timestamp 1679585382
transform 1 0 42528 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_444
timestamp 1677583704
transform 1 0 43200 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_446
timestamp 1677583258
transform 1 0 43392 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_460
timestamp 1679585382
transform 1 0 44736 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_467
timestamp 1679585382
transform 1 0 45408 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_474
timestamp 1679585382
transform 1 0 46080 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_481
timestamp 1677583704
transform 1 0 46752 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_510
timestamp 1679585382
transform 1 0 49536 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_517
timestamp 1679585382
transform 1 0 50208 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_524
timestamp 1679585382
transform 1 0 50880 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_531
timestamp 1679585382
transform 1 0 51552 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_538
timestamp 1679585382
transform 1 0 52224 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_545
timestamp 1679585382
transform 1 0 52896 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_552
timestamp 1679585382
transform 1 0 53568 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_559
timestamp 1679585382
transform 1 0 54240 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_566
timestamp 1679585382
transform 1 0 54912 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_573
timestamp 1679585382
transform 1 0 55584 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_580
timestamp 1679585382
transform 1 0 56256 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_587
timestamp 1679585382
transform 1 0 56928 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_594
timestamp 1679585382
transform 1 0 57600 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_601
timestamp 1679585382
transform 1 0 58272 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_608
timestamp 1679585382
transform 1 0 58944 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_615
timestamp 1679585382
transform 1 0 59616 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_622
timestamp 1679585382
transform 1 0 60288 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_629
timestamp 1679585382
transform 1 0 60960 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_636
timestamp 1679585382
transform 1 0 61632 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_643
timestamp 1679585382
transform 1 0 62304 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_650
timestamp 1679585382
transform 1 0 62976 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_657
timestamp 1679585382
transform 1 0 63648 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_664
timestamp 1679585382
transform 1 0 64320 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_671
timestamp 1679585382
transform 1 0 64992 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_678
timestamp 1679585382
transform 1 0 65664 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_685
timestamp 1679585382
transform 1 0 66336 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_692
timestamp 1679585382
transform 1 0 67008 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_699
timestamp 1679585382
transform 1 0 67680 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_706
timestamp 1679585382
transform 1 0 68352 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_713
timestamp 1679585382
transform 1 0 69024 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_720
timestamp 1679585382
transform 1 0 69696 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_727
timestamp 1679585382
transform 1 0 70368 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_734
timestamp 1679585382
transform 1 0 71040 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_741
timestamp 1679585382
transform 1 0 71712 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_748
timestamp 1679585382
transform 1 0 72384 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_755
timestamp 1679585382
transform 1 0 73056 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_762
timestamp 1679585382
transform 1 0 73728 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_769
timestamp 1679585382
transform 1 0 74400 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_776
timestamp 1679585382
transform 1 0 75072 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_783
timestamp 1679585382
transform 1 0 75744 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_790
timestamp 1679585382
transform 1 0 76416 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_797
timestamp 1679585382
transform 1 0 77088 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_804
timestamp 1679585382
transform 1 0 77760 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_811
timestamp 1679585382
transform 1 0 78432 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_818
timestamp 1679585382
transform 1 0 79104 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_825
timestamp 1679585382
transform 1 0 79776 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_832
timestamp 1679585382
transform 1 0 80448 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_839
timestamp 1679585382
transform 1 0 81120 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_846
timestamp 1679585382
transform 1 0 81792 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_853
timestamp 1679585382
transform 1 0 82464 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_860
timestamp 1679585382
transform 1 0 83136 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_867
timestamp 1679585382
transform 1 0 83808 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_874
timestamp 1679585382
transform 1 0 84480 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_881
timestamp 1679585382
transform 1 0 85152 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_888
timestamp 1679585382
transform 1 0 85824 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_895
timestamp 1679585382
transform 1 0 86496 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_902
timestamp 1679585382
transform 1 0 87168 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_909
timestamp 1679585382
transform 1 0 87840 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_916
timestamp 1679585382
transform 1 0 88512 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_923
timestamp 1679585382
transform 1 0 89184 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_930
timestamp 1679585382
transform 1 0 89856 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_937
timestamp 1679585382
transform 1 0 90528 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_944
timestamp 1679585382
transform 1 0 91200 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_951
timestamp 1679585382
transform 1 0 91872 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_958
timestamp 1679585382
transform 1 0 92544 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_965
timestamp 1679585382
transform 1 0 93216 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_972
timestamp 1679585382
transform 1 0 93888 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_979
timestamp 1679585382
transform 1 0 94560 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_986
timestamp 1679585382
transform 1 0 95232 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_993
timestamp 1679585382
transform 1 0 95904 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1000
timestamp 1679585382
transform 1 0 96576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1007
timestamp 1679585382
transform 1 0 97248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1014
timestamp 1679585382
transform 1 0 97920 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1021
timestamp 1679585382
transform 1 0 98592 0 1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_34_1028
timestamp 1677583258
transform 1 0 99264 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_0
timestamp 1679585382
transform 1 0 576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_7
timestamp 1679585382
transform 1 0 1248 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_14
timestamp 1679585382
transform 1 0 1920 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_21
timestamp 1679581501
transform 1 0 2592 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_25
timestamp 1677583704
transform 1 0 2976 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_35_31
timestamp 1677583704
transform 1 0 3552 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_33
timestamp 1677583258
transform 1 0 3744 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_61
timestamp 1679585382
transform 1 0 6432 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_68
timestamp 1679585382
transform 1 0 7104 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_75
timestamp 1679585382
transform 1 0 7776 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_35_82
timestamp 1677583258
transform 1 0 8448 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_110
timestamp 1679585382
transform 1 0 11136 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_117
timestamp 1679585382
transform 1 0 11808 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_124
timestamp 1677583704
transform 1 0 12480 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_126
timestamp 1677583258
transform 1 0 12672 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_35_144
timestamp 1677583258
transform 1 0 14400 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_154
timestamp 1679585382
transform 1 0 15360 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_161
timestamp 1679585382
transform 1 0 16032 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_168
timestamp 1679585382
transform 1 0 16704 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_175
timestamp 1679585382
transform 1 0 17376 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_182
timestamp 1679585382
transform 1 0 18048 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_189
timestamp 1679585382
transform 1 0 18720 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_196
timestamp 1679585382
transform 1 0 19392 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_203
timestamp 1679585382
transform 1 0 20064 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_35_210
timestamp 1677583258
transform 1 0 20736 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_238
timestamp 1679585382
transform 1 0 23424 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_245
timestamp 1679585382
transform 1 0 24096 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_252
timestamp 1679585382
transform 1 0 24768 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_259
timestamp 1679585382
transform 1 0 25440 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_266
timestamp 1679585382
transform 1 0 26112 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_273
timestamp 1679585382
transform 1 0 26784 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_280
timestamp 1679585382
transform 1 0 27456 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_287
timestamp 1679585382
transform 1 0 28128 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_294
timestamp 1679585382
transform 1 0 28800 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_301
timestamp 1677583704
transform 1 0 29472 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_312
timestamp 1679585382
transform 1 0 30528 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_319
timestamp 1679585382
transform 1 0 31200 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_326
timestamp 1679585382
transform 1 0 31872 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_333
timestamp 1679585382
transform 1 0 32544 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_340
timestamp 1679585382
transform 1 0 33216 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_347
timestamp 1679585382
transform 1 0 33888 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_354
timestamp 1679585382
transform 1 0 34560 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_361
timestamp 1679585382
transform 1 0 35232 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_368
timestamp 1679585382
transform 1 0 35904 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_375
timestamp 1679585382
transform 1 0 36576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_382
timestamp 1679585382
transform 1 0 37248 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_389
timestamp 1679585382
transform 1 0 37920 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_396
timestamp 1679585382
transform 1 0 38592 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_403
timestamp 1679585382
transform 1 0 39264 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_410
timestamp 1679585382
transform 1 0 39936 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_417
timestamp 1679585382
transform 1 0 40608 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_424
timestamp 1679585382
transform 1 0 41280 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_431
timestamp 1679581501
transform 1 0 41952 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_435
timestamp 1677583258
transform 1 0 42336 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_35_476
timestamp 1679581501
transform 1 0 46272 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_35_480
timestamp 1677583258
transform 1 0 46656 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_494
timestamp 1679585382
transform 1 0 48000 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_501
timestamp 1679585382
transform 1 0 48672 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_508
timestamp 1679585382
transform 1 0 49344 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_515
timestamp 1679585382
transform 1 0 50016 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_522
timestamp 1679585382
transform 1 0 50688 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_529
timestamp 1679585382
transform 1 0 51360 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_536
timestamp 1679585382
transform 1 0 52032 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_543
timestamp 1679585382
transform 1 0 52704 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_550
timestamp 1679585382
transform 1 0 53376 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_557
timestamp 1679585382
transform 1 0 54048 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_564
timestamp 1679585382
transform 1 0 54720 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_571
timestamp 1679585382
transform 1 0 55392 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_578
timestamp 1679585382
transform 1 0 56064 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_585
timestamp 1679585382
transform 1 0 56736 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_592
timestamp 1679585382
transform 1 0 57408 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_599
timestamp 1679585382
transform 1 0 58080 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_606
timestamp 1679585382
transform 1 0 58752 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_613
timestamp 1679585382
transform 1 0 59424 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_620
timestamp 1679585382
transform 1 0 60096 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_627
timestamp 1679585382
transform 1 0 60768 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_634
timestamp 1679585382
transform 1 0 61440 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_641
timestamp 1679585382
transform 1 0 62112 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_648
timestamp 1679585382
transform 1 0 62784 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_655
timestamp 1679585382
transform 1 0 63456 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_662
timestamp 1679585382
transform 1 0 64128 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_669
timestamp 1679585382
transform 1 0 64800 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_676
timestamp 1679585382
transform 1 0 65472 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_683
timestamp 1679585382
transform 1 0 66144 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_690
timestamp 1679585382
transform 1 0 66816 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_697
timestamp 1679585382
transform 1 0 67488 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_704
timestamp 1679585382
transform 1 0 68160 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_711
timestamp 1679585382
transform 1 0 68832 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_718
timestamp 1679585382
transform 1 0 69504 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_725
timestamp 1679585382
transform 1 0 70176 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_732
timestamp 1679585382
transform 1 0 70848 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_739
timestamp 1679585382
transform 1 0 71520 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_746
timestamp 1679585382
transform 1 0 72192 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_753
timestamp 1679585382
transform 1 0 72864 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_760
timestamp 1679585382
transform 1 0 73536 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_767
timestamp 1679585382
transform 1 0 74208 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_774
timestamp 1679585382
transform 1 0 74880 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_781
timestamp 1679585382
transform 1 0 75552 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_788
timestamp 1679585382
transform 1 0 76224 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_795
timestamp 1679585382
transform 1 0 76896 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_802
timestamp 1679585382
transform 1 0 77568 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_809
timestamp 1679585382
transform 1 0 78240 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_816
timestamp 1679585382
transform 1 0 78912 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_823
timestamp 1679585382
transform 1 0 79584 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_830
timestamp 1679585382
transform 1 0 80256 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_837
timestamp 1679585382
transform 1 0 80928 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_844
timestamp 1679585382
transform 1 0 81600 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_851
timestamp 1679585382
transform 1 0 82272 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_858
timestamp 1679585382
transform 1 0 82944 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_865
timestamp 1679585382
transform 1 0 83616 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_872
timestamp 1679585382
transform 1 0 84288 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_879
timestamp 1679585382
transform 1 0 84960 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_886
timestamp 1679585382
transform 1 0 85632 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_893
timestamp 1679585382
transform 1 0 86304 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_900
timestamp 1679585382
transform 1 0 86976 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_907
timestamp 1679585382
transform 1 0 87648 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_914
timestamp 1679585382
transform 1 0 88320 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_921
timestamp 1679585382
transform 1 0 88992 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_928
timestamp 1679585382
transform 1 0 89664 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_935
timestamp 1679585382
transform 1 0 90336 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_942
timestamp 1679585382
transform 1 0 91008 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_949
timestamp 1679585382
transform 1 0 91680 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_956
timestamp 1679585382
transform 1 0 92352 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_963
timestamp 1679585382
transform 1 0 93024 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_970
timestamp 1679585382
transform 1 0 93696 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_977
timestamp 1679585382
transform 1 0 94368 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_984
timestamp 1679585382
transform 1 0 95040 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_991
timestamp 1679585382
transform 1 0 95712 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_998
timestamp 1679585382
transform 1 0 96384 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1005
timestamp 1679585382
transform 1 0 97056 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1012
timestamp 1679585382
transform 1 0 97728 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1019
timestamp 1679585382
transform 1 0 98400 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_1026
timestamp 1677583704
transform 1 0 99072 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_1028
timestamp 1677583258
transform 1 0 99264 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_0
timestamp 1679585382
transform 1 0 576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_7
timestamp 1679585382
transform 1 0 1248 0 1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_36_14
timestamp 1677583704
transform 1 0 1920 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_16
timestamp 1677583258
transform 1 0 2112 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_44
timestamp 1677583704
transform 1 0 4800 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_46
timestamp 1677583258
transform 1 0 4992 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_65
timestamp 1679585382
transform 1 0 6816 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_72
timestamp 1679585382
transform 1 0 7488 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_79
timestamp 1679585382
transform 1 0 8160 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_86
timestamp 1679585382
transform 1 0 8832 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_93
timestamp 1679585382
transform 1 0 9504 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_100
timestamp 1679585382
transform 1 0 10176 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_107
timestamp 1679585382
transform 1 0 10848 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_114
timestamp 1679581501
transform 1 0 11520 0 1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_36_118
timestamp 1677583258
transform 1 0 11904 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_132
timestamp 1679585382
transform 1 0 13248 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_139
timestamp 1679585382
transform 1 0 13920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_146
timestamp 1679585382
transform 1 0 14592 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_153
timestamp 1679585382
transform 1 0 15264 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_160
timestamp 1679585382
transform 1 0 15936 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_167
timestamp 1679585382
transform 1 0 16608 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_174
timestamp 1679585382
transform 1 0 17280 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_181
timestamp 1679585382
transform 1 0 17952 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_188
timestamp 1679585382
transform 1 0 18624 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_195
timestamp 1679585382
transform 1 0 19296 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_202
timestamp 1679585382
transform 1 0 19968 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_209
timestamp 1679585382
transform 1 0 20640 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_216
timestamp 1679585382
transform 1 0 21312 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_223
timestamp 1679585382
transform 1 0 21984 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_230
timestamp 1679585382
transform 1 0 22656 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_237
timestamp 1679585382
transform 1 0 23328 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_244
timestamp 1679585382
transform 1 0 24000 0 1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_36_251
timestamp 1677583704
transform 1 0 24672 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_253
timestamp 1677583258
transform 1 0 24864 0 1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_36_276
timestamp 1679581501
transform 1 0 27072 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_280
timestamp 1677583704
transform 1 0 27456 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_298
timestamp 1679585382
transform 1 0 29184 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_305
timestamp 1679585382
transform 1 0 29856 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_312
timestamp 1679585382
transform 1 0 30528 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_319
timestamp 1679585382
transform 1 0 31200 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_326
timestamp 1679585382
transform 1 0 31872 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_333
timestamp 1679585382
transform 1 0 32544 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_340
timestamp 1679585382
transform 1 0 33216 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_347
timestamp 1679585382
transform 1 0 33888 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_354
timestamp 1679585382
transform 1 0 34560 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_361
timestamp 1679585382
transform 1 0 35232 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_368
timestamp 1679585382
transform 1 0 35904 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_375
timestamp 1679585382
transform 1 0 36576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_382
timestamp 1679585382
transform 1 0 37248 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_389
timestamp 1679585382
transform 1 0 37920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_396
timestamp 1679585382
transform 1 0 38592 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_403
timestamp 1679585382
transform 1 0 39264 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_410
timestamp 1679585382
transform 1 0 39936 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_417
timestamp 1679585382
transform 1 0 40608 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_424
timestamp 1679581501
transform 1 0 41280 0 1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_36_441
timestamp 1679585382
transform 1 0 42912 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_448
timestamp 1679585382
transform 1 0 43584 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_455
timestamp 1679581501
transform 1 0 44256 0 1 27972
box -48 -56 432 834
use sg13g2_decap_4  FILLER_36_463
timestamp 1679581501
transform 1 0 45024 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_467
timestamp 1677583704
transform 1 0 45408 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_478
timestamp 1679585382
transform 1 0 46464 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_485
timestamp 1679585382
transform 1 0 47136 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_492
timestamp 1679585382
transform 1 0 47808 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_499
timestamp 1679585382
transform 1 0 48480 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_506
timestamp 1679585382
transform 1 0 49152 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_513
timestamp 1679585382
transform 1 0 49824 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_520
timestamp 1679585382
transform 1 0 50496 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_527
timestamp 1679585382
transform 1 0 51168 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_534
timestamp 1679585382
transform 1 0 51840 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_541
timestamp 1679585382
transform 1 0 52512 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_548
timestamp 1679585382
transform 1 0 53184 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_555
timestamp 1679585382
transform 1 0 53856 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_562
timestamp 1679585382
transform 1 0 54528 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_569
timestamp 1679585382
transform 1 0 55200 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_576
timestamp 1679585382
transform 1 0 55872 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_583
timestamp 1679585382
transform 1 0 56544 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_590
timestamp 1679585382
transform 1 0 57216 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_597
timestamp 1679585382
transform 1 0 57888 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_604
timestamp 1679585382
transform 1 0 58560 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_611
timestamp 1679585382
transform 1 0 59232 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_618
timestamp 1679585382
transform 1 0 59904 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_625
timestamp 1679585382
transform 1 0 60576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_632
timestamp 1679585382
transform 1 0 61248 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_639
timestamp 1679585382
transform 1 0 61920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_646
timestamp 1679585382
transform 1 0 62592 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_653
timestamp 1679585382
transform 1 0 63264 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_660
timestamp 1679585382
transform 1 0 63936 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_667
timestamp 1679585382
transform 1 0 64608 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_674
timestamp 1679585382
transform 1 0 65280 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_681
timestamp 1679585382
transform 1 0 65952 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_688
timestamp 1679585382
transform 1 0 66624 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_695
timestamp 1679585382
transform 1 0 67296 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_702
timestamp 1679585382
transform 1 0 67968 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_709
timestamp 1679585382
transform 1 0 68640 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_716
timestamp 1679585382
transform 1 0 69312 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_723
timestamp 1679585382
transform 1 0 69984 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_730
timestamp 1679585382
transform 1 0 70656 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_737
timestamp 1679585382
transform 1 0 71328 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_744
timestamp 1679585382
transform 1 0 72000 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_751
timestamp 1679585382
transform 1 0 72672 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_758
timestamp 1679585382
transform 1 0 73344 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_765
timestamp 1679585382
transform 1 0 74016 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_772
timestamp 1679585382
transform 1 0 74688 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_779
timestamp 1679585382
transform 1 0 75360 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_786
timestamp 1679585382
transform 1 0 76032 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_793
timestamp 1679585382
transform 1 0 76704 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_800
timestamp 1679585382
transform 1 0 77376 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_807
timestamp 1679585382
transform 1 0 78048 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_814
timestamp 1679585382
transform 1 0 78720 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_821
timestamp 1679585382
transform 1 0 79392 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_828
timestamp 1679585382
transform 1 0 80064 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_835
timestamp 1679585382
transform 1 0 80736 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_842
timestamp 1679585382
transform 1 0 81408 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_849
timestamp 1679585382
transform 1 0 82080 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_856
timestamp 1679585382
transform 1 0 82752 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_863
timestamp 1679585382
transform 1 0 83424 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_870
timestamp 1679585382
transform 1 0 84096 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_877
timestamp 1679585382
transform 1 0 84768 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_884
timestamp 1679585382
transform 1 0 85440 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_891
timestamp 1679585382
transform 1 0 86112 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_898
timestamp 1679585382
transform 1 0 86784 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_905
timestamp 1679585382
transform 1 0 87456 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_912
timestamp 1679585382
transform 1 0 88128 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_919
timestamp 1679585382
transform 1 0 88800 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_926
timestamp 1679585382
transform 1 0 89472 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_933
timestamp 1679585382
transform 1 0 90144 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_940
timestamp 1679585382
transform 1 0 90816 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_947
timestamp 1679585382
transform 1 0 91488 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_954
timestamp 1679585382
transform 1 0 92160 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_961
timestamp 1679585382
transform 1 0 92832 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_968
timestamp 1679585382
transform 1 0 93504 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_975
timestamp 1679585382
transform 1 0 94176 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_982
timestamp 1679585382
transform 1 0 94848 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_989
timestamp 1679585382
transform 1 0 95520 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_996
timestamp 1679585382
transform 1 0 96192 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1003
timestamp 1679585382
transform 1 0 96864 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1010
timestamp 1679585382
transform 1 0 97536 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1017
timestamp 1679585382
transform 1 0 98208 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_1024
timestamp 1679581501
transform 1 0 98880 0 1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_36_1028
timestamp 1677583258
transform 1 0 99264 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_0
timestamp 1679585382
transform 1 0 576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_7
timestamp 1679585382
transform 1 0 1248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_14
timestamp 1679585382
transform 1 0 1920 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_21
timestamp 1679585382
transform 1 0 2592 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_28
timestamp 1679585382
transform 1 0 3264 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_35
timestamp 1677583704
transform 1 0 3936 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_37_50
timestamp 1679585382
transform 1 0 5376 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_57
timestamp 1679585382
transform 1 0 6048 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_64
timestamp 1679585382
transform 1 0 6720 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_71
timestamp 1679585382
transform 1 0 7392 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_78
timestamp 1679585382
transform 1 0 8064 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_98
timestamp 1679585382
transform 1 0 9984 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_105
timestamp 1679585382
transform 1 0 10656 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_112
timestamp 1679585382
transform 1 0 11328 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_119
timestamp 1677583258
transform 1 0 12000 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_128
timestamp 1679585382
transform 1 0 12864 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_135
timestamp 1679585382
transform 1 0 13536 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_142
timestamp 1679585382
transform 1 0 14208 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_149
timestamp 1679585382
transform 1 0 14880 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_156
timestamp 1679585382
transform 1 0 15552 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_163
timestamp 1679585382
transform 1 0 16224 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_170
timestamp 1679585382
transform 1 0 16896 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_177
timestamp 1679585382
transform 1 0 17568 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_184
timestamp 1679585382
transform 1 0 18240 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_191
timestamp 1679585382
transform 1 0 18912 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_198
timestamp 1679585382
transform 1 0 19584 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_205
timestamp 1679585382
transform 1 0 20256 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_212
timestamp 1679585382
transform 1 0 20928 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_219
timestamp 1679581501
transform 1 0 21600 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_37_223
timestamp 1677583258
transform 1 0 21984 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_237
timestamp 1679585382
transform 1 0 23328 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_244
timestamp 1679585382
transform 1 0 24000 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_251
timestamp 1679585382
transform 1 0 24672 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_258
timestamp 1679585382
transform 1 0 25344 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_265
timestamp 1679585382
transform 1 0 26016 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_272
timestamp 1679585382
transform 1 0 26688 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_279
timestamp 1679585382
transform 1 0 27360 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_286
timestamp 1679581501
transform 1 0 28032 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_37_294
timestamp 1677583704
transform 1 0 28800 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_296
timestamp 1677583258
transform 1 0 28992 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_319
timestamp 1679585382
transform 1 0 31200 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_326
timestamp 1677583704
transform 1 0 31872 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_37_355
timestamp 1679585382
transform 1 0 34656 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_362
timestamp 1679585382
transform 1 0 35328 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_369
timestamp 1679585382
transform 1 0 36000 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_376
timestamp 1679585382
transform 1 0 36672 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_383
timestamp 1679585382
transform 1 0 37344 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_390
timestamp 1679585382
transform 1 0 38016 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_397
timestamp 1679585382
transform 1 0 38688 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_404
timestamp 1679585382
transform 1 0 39360 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_411
timestamp 1679585382
transform 1 0 40032 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_418
timestamp 1679585382
transform 1 0 40704 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_425
timestamp 1679585382
transform 1 0 41376 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_432
timestamp 1679585382
transform 1 0 42048 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_439
timestamp 1679585382
transform 1 0 42720 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_446
timestamp 1679585382
transform 1 0 43392 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_453
timestamp 1679585382
transform 1 0 44064 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_460
timestamp 1679585382
transform 1 0 44736 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_467
timestamp 1679585382
transform 1 0 45408 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_474
timestamp 1679585382
transform 1 0 46080 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_485
timestamp 1679585382
transform 1 0 47136 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_492
timestamp 1679585382
transform 1 0 47808 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_499
timestamp 1679585382
transform 1 0 48480 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_506
timestamp 1679585382
transform 1 0 49152 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_513
timestamp 1679585382
transform 1 0 49824 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_520
timestamp 1679585382
transform 1 0 50496 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_527
timestamp 1679585382
transform 1 0 51168 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_534
timestamp 1679585382
transform 1 0 51840 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_541
timestamp 1679585382
transform 1 0 52512 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_548
timestamp 1679585382
transform 1 0 53184 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_555
timestamp 1679585382
transform 1 0 53856 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_562
timestamp 1679585382
transform 1 0 54528 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_569
timestamp 1679585382
transform 1 0 55200 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_576
timestamp 1679585382
transform 1 0 55872 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_583
timestamp 1679585382
transform 1 0 56544 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_590
timestamp 1679585382
transform 1 0 57216 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_597
timestamp 1679585382
transform 1 0 57888 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_604
timestamp 1679585382
transform 1 0 58560 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_611
timestamp 1679585382
transform 1 0 59232 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_618
timestamp 1679585382
transform 1 0 59904 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_625
timestamp 1679585382
transform 1 0 60576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_632
timestamp 1679585382
transform 1 0 61248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_639
timestamp 1679585382
transform 1 0 61920 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_646
timestamp 1679585382
transform 1 0 62592 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_653
timestamp 1679585382
transform 1 0 63264 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_660
timestamp 1679585382
transform 1 0 63936 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_667
timestamp 1679585382
transform 1 0 64608 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_674
timestamp 1679585382
transform 1 0 65280 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_681
timestamp 1679585382
transform 1 0 65952 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_688
timestamp 1679585382
transform 1 0 66624 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_695
timestamp 1679585382
transform 1 0 67296 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_702
timestamp 1679585382
transform 1 0 67968 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_709
timestamp 1679585382
transform 1 0 68640 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_716
timestamp 1679585382
transform 1 0 69312 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_723
timestamp 1679585382
transform 1 0 69984 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_730
timestamp 1679585382
transform 1 0 70656 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_737
timestamp 1679585382
transform 1 0 71328 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_744
timestamp 1679585382
transform 1 0 72000 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_751
timestamp 1679585382
transform 1 0 72672 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_758
timestamp 1679585382
transform 1 0 73344 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_765
timestamp 1679585382
transform 1 0 74016 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_772
timestamp 1679585382
transform 1 0 74688 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_779
timestamp 1679585382
transform 1 0 75360 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_786
timestamp 1679585382
transform 1 0 76032 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_793
timestamp 1679585382
transform 1 0 76704 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_800
timestamp 1679585382
transform 1 0 77376 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_807
timestamp 1679585382
transform 1 0 78048 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_814
timestamp 1679585382
transform 1 0 78720 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_821
timestamp 1679585382
transform 1 0 79392 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_828
timestamp 1679585382
transform 1 0 80064 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_835
timestamp 1679585382
transform 1 0 80736 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_842
timestamp 1679585382
transform 1 0 81408 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_849
timestamp 1679585382
transform 1 0 82080 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_856
timestamp 1679585382
transform 1 0 82752 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_863
timestamp 1679585382
transform 1 0 83424 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_870
timestamp 1679585382
transform 1 0 84096 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_877
timestamp 1679585382
transform 1 0 84768 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_884
timestamp 1679585382
transform 1 0 85440 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_891
timestamp 1679585382
transform 1 0 86112 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_898
timestamp 1679585382
transform 1 0 86784 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_905
timestamp 1679585382
transform 1 0 87456 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_912
timestamp 1679585382
transform 1 0 88128 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_919
timestamp 1679585382
transform 1 0 88800 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_926
timestamp 1679585382
transform 1 0 89472 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_933
timestamp 1679585382
transform 1 0 90144 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_940
timestamp 1679585382
transform 1 0 90816 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_947
timestamp 1679585382
transform 1 0 91488 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_954
timestamp 1679585382
transform 1 0 92160 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_961
timestamp 1679585382
transform 1 0 92832 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_968
timestamp 1679585382
transform 1 0 93504 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_975
timestamp 1679585382
transform 1 0 94176 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_982
timestamp 1679585382
transform 1 0 94848 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_989
timestamp 1679585382
transform 1 0 95520 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_996
timestamp 1679585382
transform 1 0 96192 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1003
timestamp 1679585382
transform 1 0 96864 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1010
timestamp 1679585382
transform 1 0 97536 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1017
timestamp 1679585382
transform 1 0 98208 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_1024
timestamp 1679581501
transform 1 0 98880 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_37_1028
timestamp 1677583258
transform 1 0 99264 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_0
timestamp 1679585382
transform 1 0 576 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_7
timestamp 1679585382
transform 1 0 1248 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_14
timestamp 1679585382
transform 1 0 1920 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_21
timestamp 1679585382
transform 1 0 2592 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_28
timestamp 1679585382
transform 1 0 3264 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_35
timestamp 1679585382
transform 1 0 3936 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_42
timestamp 1679581501
transform 1 0 4608 0 1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_38_46
timestamp 1677583258
transform 1 0 4992 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_55
timestamp 1679585382
transform 1 0 5856 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_62
timestamp 1679585382
transform 1 0 6528 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_69
timestamp 1679585382
transform 1 0 7200 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_76
timestamp 1679585382
transform 1 0 7872 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_83
timestamp 1679585382
transform 1 0 8544 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_90
timestamp 1679585382
transform 1 0 9216 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_97
timestamp 1679585382
transform 1 0 9888 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_104
timestamp 1679581501
transform 1 0 10560 0 1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_38_108
timestamp 1677583258
transform 1 0 10944 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_117
timestamp 1679585382
transform 1 0 11808 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_124
timestamp 1679585382
transform 1 0 12480 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_131
timestamp 1679585382
transform 1 0 13152 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_138
timestamp 1679585382
transform 1 0 13824 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_145
timestamp 1679585382
transform 1 0 14496 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_152
timestamp 1679581501
transform 1 0 15168 0 1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_38_156
timestamp 1677583258
transform 1 0 15552 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_170
timestamp 1679585382
transform 1 0 16896 0 1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_38_177
timestamp 1677583704
transform 1 0 17568 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_179
timestamp 1677583258
transform 1 0 17760 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_184
timestamp 1679585382
transform 1 0 18240 0 1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_38_191
timestamp 1677583704
transform 1 0 18912 0 1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_38_202
timestamp 1679585382
transform 1 0 19968 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_209
timestamp 1679585382
transform 1 0 20640 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_216
timestamp 1679585382
transform 1 0 21312 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_223
timestamp 1679585382
transform 1 0 21984 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_230
timestamp 1679585382
transform 1 0 22656 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_237
timestamp 1679585382
transform 1 0 23328 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_244
timestamp 1679585382
transform 1 0 24000 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_251
timestamp 1679585382
transform 1 0 24672 0 1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_38_258
timestamp 1677583704
transform 1 0 25344 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_260
timestamp 1677583258
transform 1 0 25536 0 1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_38_288
timestamp 1677583258
transform 1 0 28224 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_298
timestamp 1679585382
transform 1 0 29184 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_305
timestamp 1679585382
transform 1 0 29856 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_312
timestamp 1679585382
transform 1 0 30528 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_319
timestamp 1679585382
transform 1 0 31200 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_326
timestamp 1679585382
transform 1 0 31872 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_333
timestamp 1679585382
transform 1 0 32544 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_340
timestamp 1679585382
transform 1 0 33216 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_347
timestamp 1679585382
transform 1 0 33888 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_354
timestamp 1679585382
transform 1 0 34560 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_361
timestamp 1679585382
transform 1 0 35232 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_368
timestamp 1679585382
transform 1 0 35904 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_375
timestamp 1679581501
transform 1 0 36576 0 1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_38_379
timestamp 1677583258
transform 1 0 36960 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_392
timestamp 1679585382
transform 1 0 38208 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_399
timestamp 1679585382
transform 1 0 38880 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_406
timestamp 1679585382
transform 1 0 39552 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_413
timestamp 1679585382
transform 1 0 40224 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_420
timestamp 1679585382
transform 1 0 40896 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_427
timestamp 1679585382
transform 1 0 41568 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_434
timestamp 1679581501
transform 1 0 42240 0 1 29484
box -48 -56 432 834
use sg13g2_decap_8  FILLER_38_451
timestamp 1679585382
transform 1 0 43872 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_458
timestamp 1679585382
transform 1 0 44544 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_465
timestamp 1679581501
transform 1 0 45216 0 1 29484
box -48 -56 432 834
use sg13g2_decap_8  FILLER_38_495
timestamp 1679585382
transform 1 0 48096 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_502
timestamp 1679585382
transform 1 0 48768 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_509
timestamp 1679585382
transform 1 0 49440 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_516
timestamp 1679585382
transform 1 0 50112 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_523
timestamp 1679585382
transform 1 0 50784 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_530
timestamp 1679585382
transform 1 0 51456 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_537
timestamp 1679585382
transform 1 0 52128 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_544
timestamp 1679585382
transform 1 0 52800 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_551
timestamp 1679585382
transform 1 0 53472 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_558
timestamp 1679585382
transform 1 0 54144 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_565
timestamp 1679585382
transform 1 0 54816 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_572
timestamp 1679585382
transform 1 0 55488 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_579
timestamp 1679585382
transform 1 0 56160 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_586
timestamp 1679585382
transform 1 0 56832 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_593
timestamp 1679585382
transform 1 0 57504 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_600
timestamp 1679585382
transform 1 0 58176 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_607
timestamp 1679585382
transform 1 0 58848 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_614
timestamp 1679585382
transform 1 0 59520 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_621
timestamp 1679585382
transform 1 0 60192 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_628
timestamp 1679585382
transform 1 0 60864 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_635
timestamp 1679585382
transform 1 0 61536 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_642
timestamp 1679585382
transform 1 0 62208 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_649
timestamp 1679585382
transform 1 0 62880 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_656
timestamp 1679585382
transform 1 0 63552 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_663
timestamp 1679585382
transform 1 0 64224 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_670
timestamp 1679585382
transform 1 0 64896 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_677
timestamp 1679585382
transform 1 0 65568 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_684
timestamp 1679585382
transform 1 0 66240 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_691
timestamp 1679585382
transform 1 0 66912 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_698
timestamp 1679585382
transform 1 0 67584 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_705
timestamp 1679585382
transform 1 0 68256 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_712
timestamp 1679585382
transform 1 0 68928 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_719
timestamp 1679585382
transform 1 0 69600 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_726
timestamp 1679585382
transform 1 0 70272 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_733
timestamp 1679585382
transform 1 0 70944 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_740
timestamp 1679585382
transform 1 0 71616 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_747
timestamp 1679585382
transform 1 0 72288 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_754
timestamp 1679585382
transform 1 0 72960 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_761
timestamp 1679585382
transform 1 0 73632 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_768
timestamp 1679585382
transform 1 0 74304 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_775
timestamp 1679585382
transform 1 0 74976 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_782
timestamp 1679585382
transform 1 0 75648 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_789
timestamp 1679585382
transform 1 0 76320 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_796
timestamp 1679585382
transform 1 0 76992 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_803
timestamp 1679585382
transform 1 0 77664 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_810
timestamp 1679585382
transform 1 0 78336 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_817
timestamp 1679585382
transform 1 0 79008 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_824
timestamp 1679585382
transform 1 0 79680 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_831
timestamp 1679585382
transform 1 0 80352 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_838
timestamp 1679585382
transform 1 0 81024 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_845
timestamp 1679585382
transform 1 0 81696 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_852
timestamp 1679585382
transform 1 0 82368 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_859
timestamp 1679585382
transform 1 0 83040 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_866
timestamp 1679585382
transform 1 0 83712 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_873
timestamp 1679585382
transform 1 0 84384 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_880
timestamp 1679585382
transform 1 0 85056 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_887
timestamp 1679585382
transform 1 0 85728 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_894
timestamp 1679585382
transform 1 0 86400 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_901
timestamp 1679585382
transform 1 0 87072 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_908
timestamp 1679585382
transform 1 0 87744 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_915
timestamp 1679585382
transform 1 0 88416 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_922
timestamp 1679585382
transform 1 0 89088 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_929
timestamp 1679585382
transform 1 0 89760 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_936
timestamp 1679585382
transform 1 0 90432 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_943
timestamp 1679585382
transform 1 0 91104 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_950
timestamp 1679585382
transform 1 0 91776 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_957
timestamp 1679585382
transform 1 0 92448 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_964
timestamp 1679585382
transform 1 0 93120 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_971
timestamp 1679585382
transform 1 0 93792 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_978
timestamp 1679585382
transform 1 0 94464 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_985
timestamp 1679585382
transform 1 0 95136 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_992
timestamp 1679585382
transform 1 0 95808 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_999
timestamp 1679585382
transform 1 0 96480 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1006
timestamp 1679585382
transform 1 0 97152 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1013
timestamp 1679585382
transform 1 0 97824 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1020
timestamp 1679585382
transform 1 0 98496 0 1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_38_1027
timestamp 1677583704
transform 1 0 99168 0 1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_0
timestamp 1679585382
transform 1 0 576 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_7
timestamp 1679585382
transform 1 0 1248 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_14
timestamp 1679585382
transform 1 0 1920 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_21
timestamp 1679585382
transform 1 0 2592 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_32
timestamp 1677583704
transform 1 0 3648 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_34
timestamp 1677583258
transform 1 0 3840 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_48
timestamp 1679585382
transform 1 0 5184 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_55
timestamp 1679585382
transform 1 0 5856 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_62
timestamp 1679585382
transform 1 0 6528 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_96
timestamp 1679585382
transform 1 0 9792 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_103
timestamp 1679585382
transform 1 0 10464 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_110
timestamp 1679585382
transform 1 0 11136 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_117
timestamp 1679585382
transform 1 0 11808 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_124
timestamp 1679585382
transform 1 0 12480 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_131
timestamp 1677583704
transform 1 0 13152 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_133
timestamp 1677583258
transform 1 0 13344 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_143
timestamp 1679585382
transform 1 0 14304 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_150
timestamp 1679585382
transform 1 0 14976 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_157
timestamp 1679585382
transform 1 0 15648 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_164
timestamp 1679585382
transform 1 0 16320 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_171
timestamp 1679581501
transform 1 0 16992 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_39_175
timestamp 1677583258
transform 1 0 17376 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_203
timestamp 1679585382
transform 1 0 20064 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_210
timestamp 1679585382
transform 1 0 20736 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_217
timestamp 1679581501
transform 1 0 21408 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_39_221
timestamp 1677583258
transform 1 0 21792 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_4  FILLER_39_249
timestamp 1679581501
transform 1 0 24480 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_39_253
timestamp 1677583704
transform 1 0 24864 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_281
timestamp 1679585382
transform 1 0 27552 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_288
timestamp 1679585382
transform 1 0 28224 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_295
timestamp 1679585382
transform 1 0 28896 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_302
timestamp 1679585382
transform 1 0 29568 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_309
timestamp 1677583704
transform 1 0 30240 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_311
timestamp 1677583258
transform 1 0 30432 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_320
timestamp 1679585382
transform 1 0 31296 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_327
timestamp 1679585382
transform 1 0 31968 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_334
timestamp 1679585382
transform 1 0 32640 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_341
timestamp 1679585382
transform 1 0 33312 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_39_348
timestamp 1677583258
transform 1 0 33984 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_365
timestamp 1677583704
transform 1 0 35616 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_367
timestamp 1677583258
transform 1 0 35808 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_377
timestamp 1677583704
transform 1 0 36768 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_406
timestamp 1679585382
transform 1 0 39552 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_413
timestamp 1679585382
transform 1 0 40224 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_39_420
timestamp 1677583258
transform 1 0 40896 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_461
timestamp 1679585382
transform 1 0 44832 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_468
timestamp 1679581501
transform 1 0 45504 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_39_472
timestamp 1677583704
transform 1 0 45888 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_477
timestamp 1679585382
transform 1 0 46368 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_484
timestamp 1679585382
transform 1 0 47040 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_491
timestamp 1679581501
transform 1 0 47712 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_39_495
timestamp 1677583704
transform 1 0 48096 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_532
timestamp 1679585382
transform 1 0 51648 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_539
timestamp 1679585382
transform 1 0 52320 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_546
timestamp 1679585382
transform 1 0 52992 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_553
timestamp 1679585382
transform 1 0 53664 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_560
timestamp 1679585382
transform 1 0 54336 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_567
timestamp 1679585382
transform 1 0 55008 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_574
timestamp 1679585382
transform 1 0 55680 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_581
timestamp 1679585382
transform 1 0 56352 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_588
timestamp 1679585382
transform 1 0 57024 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_595
timestamp 1679585382
transform 1 0 57696 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_602
timestamp 1679585382
transform 1 0 58368 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_609
timestamp 1679585382
transform 1 0 59040 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_616
timestamp 1679585382
transform 1 0 59712 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_623
timestamp 1679585382
transform 1 0 60384 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_630
timestamp 1679585382
transform 1 0 61056 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_637
timestamp 1679585382
transform 1 0 61728 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_644
timestamp 1679585382
transform 1 0 62400 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_651
timestamp 1679585382
transform 1 0 63072 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_658
timestamp 1679585382
transform 1 0 63744 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_665
timestamp 1679585382
transform 1 0 64416 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_672
timestamp 1679585382
transform 1 0 65088 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_679
timestamp 1679585382
transform 1 0 65760 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_686
timestamp 1679585382
transform 1 0 66432 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_693
timestamp 1679585382
transform 1 0 67104 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_700
timestamp 1679585382
transform 1 0 67776 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_707
timestamp 1679585382
transform 1 0 68448 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_714
timestamp 1679585382
transform 1 0 69120 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_721
timestamp 1679585382
transform 1 0 69792 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_728
timestamp 1679585382
transform 1 0 70464 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_735
timestamp 1679585382
transform 1 0 71136 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_742
timestamp 1679585382
transform 1 0 71808 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_749
timestamp 1679585382
transform 1 0 72480 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_756
timestamp 1679585382
transform 1 0 73152 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_763
timestamp 1679585382
transform 1 0 73824 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_770
timestamp 1679585382
transform 1 0 74496 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_777
timestamp 1679585382
transform 1 0 75168 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_784
timestamp 1679585382
transform 1 0 75840 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_791
timestamp 1679585382
transform 1 0 76512 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_798
timestamp 1679585382
transform 1 0 77184 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_805
timestamp 1679585382
transform 1 0 77856 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_812
timestamp 1679585382
transform 1 0 78528 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_819
timestamp 1679585382
transform 1 0 79200 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_826
timestamp 1679585382
transform 1 0 79872 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_833
timestamp 1679585382
transform 1 0 80544 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_840
timestamp 1679585382
transform 1 0 81216 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_847
timestamp 1679585382
transform 1 0 81888 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_854
timestamp 1679585382
transform 1 0 82560 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_861
timestamp 1679585382
transform 1 0 83232 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_868
timestamp 1679585382
transform 1 0 83904 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_875
timestamp 1679585382
transform 1 0 84576 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_882
timestamp 1679585382
transform 1 0 85248 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_889
timestamp 1679585382
transform 1 0 85920 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_896
timestamp 1679585382
transform 1 0 86592 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_903
timestamp 1679585382
transform 1 0 87264 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_910
timestamp 1679585382
transform 1 0 87936 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_917
timestamp 1679585382
transform 1 0 88608 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_924
timestamp 1679585382
transform 1 0 89280 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_931
timestamp 1679585382
transform 1 0 89952 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_938
timestamp 1679585382
transform 1 0 90624 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_945
timestamp 1679585382
transform 1 0 91296 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_952
timestamp 1679585382
transform 1 0 91968 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_959
timestamp 1679585382
transform 1 0 92640 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_966
timestamp 1679585382
transform 1 0 93312 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_973
timestamp 1679585382
transform 1 0 93984 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_980
timestamp 1679585382
transform 1 0 94656 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_987
timestamp 1679585382
transform 1 0 95328 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_994
timestamp 1679585382
transform 1 0 96000 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1001
timestamp 1679585382
transform 1 0 96672 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1008
timestamp 1679585382
transform 1 0 97344 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1015
timestamp 1679585382
transform 1 0 98016 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1022
timestamp 1679585382
transform 1 0 98688 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_0
timestamp 1679585382
transform 1 0 576 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_7
timestamp 1679585382
transform 1 0 1248 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_14
timestamp 1677583704
transform 1 0 1920 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_47
timestamp 1679585382
transform 1 0 5088 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_54
timestamp 1679585382
transform 1 0 5760 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_61
timestamp 1679585382
transform 1 0 6432 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_68
timestamp 1679585382
transform 1 0 7104 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_75
timestamp 1679585382
transform 1 0 7776 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_82
timestamp 1679585382
transform 1 0 8448 0 1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_40_89
timestamp 1677583258
transform 1 0 9120 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_117
timestamp 1679585382
transform 1 0 11808 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_124
timestamp 1679585382
transform 1 0 12480 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_131
timestamp 1679585382
transform 1 0 13152 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_138
timestamp 1679585382
transform 1 0 13824 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_145
timestamp 1679585382
transform 1 0 14496 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_152
timestamp 1679585382
transform 1 0 15168 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_159
timestamp 1679585382
transform 1 0 15840 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_166
timestamp 1679585382
transform 1 0 16512 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_173
timestamp 1677583704
transform 1 0 17184 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_207
timestamp 1679585382
transform 1 0 20448 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_214
timestamp 1679585382
transform 1 0 21120 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_221
timestamp 1679581501
transform 1 0 21792 0 1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_40_225
timestamp 1677583704
transform 1 0 22176 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_240
timestamp 1679585382
transform 1 0 23616 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_247
timestamp 1679585382
transform 1 0 24288 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_254
timestamp 1677583704
transform 1 0 24960 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_256
timestamp 1677583258
transform 1 0 25152 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_270
timestamp 1679585382
transform 1 0 26496 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_277
timestamp 1679585382
transform 1 0 27168 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_284
timestamp 1679585382
transform 1 0 27840 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_291
timestamp 1679585382
transform 1 0 28512 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_298
timestamp 1679585382
transform 1 0 29184 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_305
timestamp 1679585382
transform 1 0 29856 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_312
timestamp 1679585382
transform 1 0 30528 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_319
timestamp 1679585382
transform 1 0 31200 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_326
timestamp 1679581501
transform 1 0 31872 0 1 30996
box -48 -56 432 834
use sg13g2_decap_8  FILLER_40_357
timestamp 1679585382
transform 1 0 34848 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_364
timestamp 1679585382
transform 1 0 35520 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_398
timestamp 1679585382
transform 1 0 38784 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_405
timestamp 1679585382
transform 1 0 39456 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_412
timestamp 1679585382
transform 1 0 40128 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_419
timestamp 1679581501
transform 1 0 40800 0 1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_40_423
timestamp 1677583704
transform 1 0 41184 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_438
timestamp 1679585382
transform 1 0 42624 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_445
timestamp 1679585382
transform 1 0 43296 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_452
timestamp 1679585382
transform 1 0 43968 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_459
timestamp 1679585382
transform 1 0 44640 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_466
timestamp 1679585382
transform 1 0 45312 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_473
timestamp 1679585382
transform 1 0 45984 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_511
timestamp 1679581501
transform 1 0 49632 0 1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_40_515
timestamp 1677583704
transform 1 0 50016 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_526
timestamp 1679585382
transform 1 0 51072 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_533
timestamp 1679585382
transform 1 0 51744 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_540
timestamp 1679585382
transform 1 0 52416 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_547
timestamp 1679585382
transform 1 0 53088 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_554
timestamp 1679585382
transform 1 0 53760 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_561
timestamp 1679585382
transform 1 0 54432 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_568
timestamp 1679585382
transform 1 0 55104 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_575
timestamp 1679585382
transform 1 0 55776 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_582
timestamp 1679585382
transform 1 0 56448 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_589
timestamp 1679585382
transform 1 0 57120 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_596
timestamp 1679585382
transform 1 0 57792 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_603
timestamp 1679585382
transform 1 0 58464 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_610
timestamp 1679585382
transform 1 0 59136 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_617
timestamp 1679585382
transform 1 0 59808 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_624
timestamp 1679585382
transform 1 0 60480 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_631
timestamp 1679585382
transform 1 0 61152 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_638
timestamp 1679585382
transform 1 0 61824 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_645
timestamp 1679585382
transform 1 0 62496 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_652
timestamp 1679585382
transform 1 0 63168 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_659
timestamp 1679585382
transform 1 0 63840 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_666
timestamp 1679585382
transform 1 0 64512 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_673
timestamp 1679585382
transform 1 0 65184 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_680
timestamp 1679585382
transform 1 0 65856 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_687
timestamp 1679585382
transform 1 0 66528 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_694
timestamp 1679585382
transform 1 0 67200 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_701
timestamp 1679585382
transform 1 0 67872 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_708
timestamp 1679585382
transform 1 0 68544 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_715
timestamp 1679585382
transform 1 0 69216 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_722
timestamp 1679585382
transform 1 0 69888 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_729
timestamp 1679585382
transform 1 0 70560 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_736
timestamp 1679585382
transform 1 0 71232 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_743
timestamp 1679585382
transform 1 0 71904 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_750
timestamp 1679585382
transform 1 0 72576 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_757
timestamp 1679585382
transform 1 0 73248 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_764
timestamp 1679585382
transform 1 0 73920 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_771
timestamp 1679585382
transform 1 0 74592 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_778
timestamp 1679585382
transform 1 0 75264 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_785
timestamp 1679585382
transform 1 0 75936 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_792
timestamp 1679585382
transform 1 0 76608 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_799
timestamp 1679585382
transform 1 0 77280 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_806
timestamp 1679585382
transform 1 0 77952 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_813
timestamp 1679585382
transform 1 0 78624 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_820
timestamp 1679585382
transform 1 0 79296 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_827
timestamp 1679585382
transform 1 0 79968 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_834
timestamp 1679585382
transform 1 0 80640 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_841
timestamp 1679585382
transform 1 0 81312 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_848
timestamp 1679585382
transform 1 0 81984 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_855
timestamp 1679585382
transform 1 0 82656 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_862
timestamp 1679585382
transform 1 0 83328 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_869
timestamp 1679585382
transform 1 0 84000 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_876
timestamp 1679585382
transform 1 0 84672 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_883
timestamp 1679585382
transform 1 0 85344 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_890
timestamp 1679585382
transform 1 0 86016 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_897
timestamp 1679585382
transform 1 0 86688 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_904
timestamp 1679585382
transform 1 0 87360 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_911
timestamp 1679585382
transform 1 0 88032 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_918
timestamp 1679585382
transform 1 0 88704 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_925
timestamp 1679585382
transform 1 0 89376 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_932
timestamp 1679585382
transform 1 0 90048 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_939
timestamp 1679585382
transform 1 0 90720 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_946
timestamp 1679585382
transform 1 0 91392 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_953
timestamp 1679585382
transform 1 0 92064 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_960
timestamp 1679585382
transform 1 0 92736 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_967
timestamp 1679585382
transform 1 0 93408 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_974
timestamp 1679585382
transform 1 0 94080 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_981
timestamp 1679585382
transform 1 0 94752 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_988
timestamp 1679585382
transform 1 0 95424 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_995
timestamp 1679585382
transform 1 0 96096 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1002
timestamp 1679585382
transform 1 0 96768 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1009
timestamp 1679585382
transform 1 0 97440 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1016
timestamp 1679585382
transform 1 0 98112 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_1023
timestamp 1679581501
transform 1 0 98784 0 1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_40_1027
timestamp 1677583704
transform 1 0 99168 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_41_0
timestamp 1679585382
transform 1 0 576 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_7
timestamp 1679581501
transform 1 0 1248 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_41_11
timestamp 1677583704
transform 1 0 1632 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_41_40
timestamp 1679585382
transform 1 0 4416 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_47
timestamp 1679585382
transform 1 0 5088 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_54
timestamp 1679585382
transform 1 0 5760 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_61
timestamp 1679585382
transform 1 0 6432 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_68
timestamp 1679585382
transform 1 0 7104 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_75
timestamp 1679585382
transform 1 0 7776 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_82
timestamp 1679585382
transform 1 0 8448 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_89
timestamp 1679581501
transform 1 0 9120 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_41_106
timestamp 1677583704
transform 1 0 10752 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_41_135
timestamp 1679585382
transform 1 0 13536 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_142
timestamp 1679585382
transform 1 0 14208 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_149
timestamp 1679585382
transform 1 0 14880 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_156
timestamp 1679585382
transform 1 0 15552 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_163
timestamp 1679585382
transform 1 0 16224 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_170
timestamp 1679585382
transform 1 0 16896 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_177
timestamp 1679581501
transform 1 0 17568 0 -1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_41_185
timestamp 1679585382
transform 1 0 18336 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_41_192
timestamp 1677583258
transform 1 0 19008 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_202
timestamp 1679585382
transform 1 0 19968 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_209
timestamp 1679585382
transform 1 0 20640 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_216
timestamp 1679585382
transform 1 0 21312 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_223
timestamp 1679585382
transform 1 0 21984 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_230
timestamp 1679585382
transform 1 0 22656 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_237
timestamp 1679585382
transform 1 0 23328 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_244
timestamp 1679585382
transform 1 0 24000 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_251
timestamp 1679585382
transform 1 0 24672 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_258
timestamp 1679581501
transform 1 0 25344 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_41_262
timestamp 1677583704
transform 1 0 25728 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_41_272
timestamp 1679585382
transform 1 0 26688 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_279
timestamp 1679585382
transform 1 0 27360 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_313
timestamp 1679585382
transform 1 0 30624 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_320
timestamp 1679585382
transform 1 0 31296 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_327
timestamp 1679585382
transform 1 0 31968 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_334
timestamp 1679585382
transform 1 0 32640 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_341
timestamp 1679585382
transform 1 0 33312 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_348
timestamp 1679585382
transform 1 0 33984 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_355
timestamp 1679585382
transform 1 0 34656 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_41_362
timestamp 1677583258
transform 1 0 35328 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_398
timestamp 1679585382
transform 1 0 38784 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_405
timestamp 1679585382
transform 1 0 39456 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_412
timestamp 1679585382
transform 1 0 40128 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_419
timestamp 1679585382
transform 1 0 40800 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_426
timestamp 1679585382
transform 1 0 41472 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_433
timestamp 1679581501
transform 1 0 42144 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_41_437
timestamp 1677583704
transform 1 0 42528 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_41_447
timestamp 1679585382
transform 1 0 43488 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_454
timestamp 1679585382
transform 1 0 44160 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_461
timestamp 1679585382
transform 1 0 44832 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_468
timestamp 1679585382
transform 1 0 45504 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_475
timestamp 1679585382
transform 1 0 46176 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_482
timestamp 1679585382
transform 1 0 46848 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_489
timestamp 1679585382
transform 1 0 47520 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_505
timestamp 1679585382
transform 1 0 49056 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_512
timestamp 1679585382
transform 1 0 49728 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_519
timestamp 1679585382
transform 1 0 50400 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_526
timestamp 1679585382
transform 1 0 51072 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_533
timestamp 1679585382
transform 1 0 51744 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_540
timestamp 1679585382
transform 1 0 52416 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_547
timestamp 1679585382
transform 1 0 53088 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_554
timestamp 1679585382
transform 1 0 53760 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_561
timestamp 1679585382
transform 1 0 54432 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_568
timestamp 1679585382
transform 1 0 55104 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_575
timestamp 1679585382
transform 1 0 55776 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_582
timestamp 1679585382
transform 1 0 56448 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_589
timestamp 1679585382
transform 1 0 57120 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_596
timestamp 1679585382
transform 1 0 57792 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_603
timestamp 1679585382
transform 1 0 58464 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_610
timestamp 1679585382
transform 1 0 59136 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_617
timestamp 1679585382
transform 1 0 59808 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_624
timestamp 1679585382
transform 1 0 60480 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_631
timestamp 1679585382
transform 1 0 61152 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_638
timestamp 1679585382
transform 1 0 61824 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_645
timestamp 1679585382
transform 1 0 62496 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_652
timestamp 1679585382
transform 1 0 63168 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_659
timestamp 1679585382
transform 1 0 63840 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_666
timestamp 1679585382
transform 1 0 64512 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_673
timestamp 1679585382
transform 1 0 65184 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_680
timestamp 1679585382
transform 1 0 65856 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_687
timestamp 1679585382
transform 1 0 66528 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_694
timestamp 1679585382
transform 1 0 67200 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_701
timestamp 1679585382
transform 1 0 67872 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_708
timestamp 1679585382
transform 1 0 68544 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_715
timestamp 1679585382
transform 1 0 69216 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_722
timestamp 1679585382
transform 1 0 69888 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_729
timestamp 1679585382
transform 1 0 70560 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_736
timestamp 1679585382
transform 1 0 71232 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_743
timestamp 1679585382
transform 1 0 71904 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_750
timestamp 1679585382
transform 1 0 72576 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_757
timestamp 1679585382
transform 1 0 73248 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_764
timestamp 1679585382
transform 1 0 73920 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_771
timestamp 1679585382
transform 1 0 74592 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_778
timestamp 1679585382
transform 1 0 75264 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_785
timestamp 1679585382
transform 1 0 75936 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_792
timestamp 1679585382
transform 1 0 76608 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_799
timestamp 1679585382
transform 1 0 77280 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_806
timestamp 1679585382
transform 1 0 77952 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_813
timestamp 1679585382
transform 1 0 78624 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_820
timestamp 1679585382
transform 1 0 79296 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_827
timestamp 1679585382
transform 1 0 79968 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_834
timestamp 1679585382
transform 1 0 80640 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_841
timestamp 1679585382
transform 1 0 81312 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_848
timestamp 1679585382
transform 1 0 81984 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_855
timestamp 1679585382
transform 1 0 82656 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_862
timestamp 1679585382
transform 1 0 83328 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_869
timestamp 1679585382
transform 1 0 84000 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_876
timestamp 1679585382
transform 1 0 84672 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_883
timestamp 1679585382
transform 1 0 85344 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_890
timestamp 1679585382
transform 1 0 86016 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_897
timestamp 1679585382
transform 1 0 86688 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_904
timestamp 1679585382
transform 1 0 87360 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_911
timestamp 1679585382
transform 1 0 88032 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_918
timestamp 1679585382
transform 1 0 88704 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_925
timestamp 1679585382
transform 1 0 89376 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_932
timestamp 1679585382
transform 1 0 90048 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_939
timestamp 1679585382
transform 1 0 90720 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_946
timestamp 1679585382
transform 1 0 91392 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_953
timestamp 1679585382
transform 1 0 92064 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_960
timestamp 1679585382
transform 1 0 92736 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_967
timestamp 1679585382
transform 1 0 93408 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_974
timestamp 1679585382
transform 1 0 94080 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_981
timestamp 1679585382
transform 1 0 94752 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_988
timestamp 1679585382
transform 1 0 95424 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_995
timestamp 1679585382
transform 1 0 96096 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1002
timestamp 1679585382
transform 1 0 96768 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1009
timestamp 1679585382
transform 1 0 97440 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1016
timestamp 1679585382
transform 1 0 98112 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_1023
timestamp 1679581501
transform 1 0 98784 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_41_1027
timestamp 1677583704
transform 1 0 99168 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_0
timestamp 1679585382
transform 1 0 576 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_7
timestamp 1679585382
transform 1 0 1248 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_14
timestamp 1679585382
transform 1 0 1920 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_21
timestamp 1679585382
transform 1 0 2592 0 1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_42_28
timestamp 1677583258
transform 1 0 3264 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_38
timestamp 1679585382
transform 1 0 4224 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_45
timestamp 1679585382
transform 1 0 4896 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_52
timestamp 1679585382
transform 1 0 5568 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_59
timestamp 1679585382
transform 1 0 6240 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_66
timestamp 1679585382
transform 1 0 6912 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_73
timestamp 1679585382
transform 1 0 7584 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_80
timestamp 1679585382
transform 1 0 8256 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_87
timestamp 1679585382
transform 1 0 8928 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_94
timestamp 1679585382
transform 1 0 9600 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_101
timestamp 1679585382
transform 1 0 10272 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_108
timestamp 1679585382
transform 1 0 10944 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_115
timestamp 1679585382
transform 1 0 11616 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_122
timestamp 1679585382
transform 1 0 12288 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_129
timestamp 1679585382
transform 1 0 12960 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_136
timestamp 1679585382
transform 1 0 13632 0 1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_42_143
timestamp 1677583258
transform 1 0 14304 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_171
timestamp 1679585382
transform 1 0 16992 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_178
timestamp 1677583704
transform 1 0 17664 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_180
timestamp 1677583258
transform 1 0 17856 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_185
timestamp 1679585382
transform 1 0 18336 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_192
timestamp 1679585382
transform 1 0 19008 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_199
timestamp 1679585382
transform 1 0 19680 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_206
timestamp 1679585382
transform 1 0 20352 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_213
timestamp 1679585382
transform 1 0 21024 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_220
timestamp 1679585382
transform 1 0 21696 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_227
timestamp 1679585382
transform 1 0 22368 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_234
timestamp 1679585382
transform 1 0 23040 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_241
timestamp 1679585382
transform 1 0 23712 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_248
timestamp 1679585382
transform 1 0 24384 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_255
timestamp 1679585382
transform 1 0 25056 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_262
timestamp 1679585382
transform 1 0 25728 0 1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_42_269
timestamp 1677583258
transform 1 0 26400 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_288
timestamp 1679585382
transform 1 0 28224 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_295
timestamp 1679585382
transform 1 0 28896 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_302
timestamp 1679585382
transform 1 0 29568 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_309
timestamp 1679585382
transform 1 0 30240 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_316
timestamp 1679585382
transform 1 0 30912 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_323
timestamp 1679585382
transform 1 0 31584 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_330
timestamp 1679585382
transform 1 0 32256 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_337
timestamp 1679585382
transform 1 0 32928 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_344
timestamp 1679585382
transform 1 0 33600 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_351
timestamp 1679585382
transform 1 0 34272 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_358
timestamp 1679585382
transform 1 0 34944 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_365
timestamp 1679585382
transform 1 0 35616 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_372
timestamp 1679585382
transform 1 0 36288 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_379
timestamp 1679585382
transform 1 0 36960 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_386
timestamp 1679585382
transform 1 0 37632 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_393
timestamp 1679585382
transform 1 0 38304 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_400
timestamp 1679585382
transform 1 0 38976 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_407
timestamp 1679585382
transform 1 0 39648 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_414
timestamp 1679585382
transform 1 0 40320 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_421
timestamp 1679585382
transform 1 0 40992 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_428
timestamp 1679585382
transform 1 0 41664 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_435
timestamp 1679585382
transform 1 0 42336 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_442
timestamp 1679585382
transform 1 0 43008 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_449
timestamp 1679585382
transform 1 0 43680 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_456
timestamp 1679585382
transform 1 0 44352 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_463
timestamp 1679585382
transform 1 0 45024 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_470
timestamp 1679585382
transform 1 0 45696 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_477
timestamp 1679585382
transform 1 0 46368 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_484
timestamp 1679585382
transform 1 0 47040 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_491
timestamp 1679585382
transform 1 0 47712 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_498
timestamp 1679585382
transform 1 0 48384 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_505
timestamp 1679585382
transform 1 0 49056 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_512
timestamp 1679585382
transform 1 0 49728 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_519
timestamp 1679585382
transform 1 0 50400 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_526
timestamp 1679585382
transform 1 0 51072 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_533
timestamp 1679585382
transform 1 0 51744 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_540
timestamp 1679585382
transform 1 0 52416 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_547
timestamp 1679585382
transform 1 0 53088 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_554
timestamp 1679585382
transform 1 0 53760 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_561
timestamp 1679585382
transform 1 0 54432 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_568
timestamp 1679585382
transform 1 0 55104 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_575
timestamp 1679585382
transform 1 0 55776 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_582
timestamp 1679585382
transform 1 0 56448 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_589
timestamp 1679585382
transform 1 0 57120 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_596
timestamp 1679585382
transform 1 0 57792 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_603
timestamp 1679585382
transform 1 0 58464 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_610
timestamp 1679585382
transform 1 0 59136 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_617
timestamp 1679585382
transform 1 0 59808 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_624
timestamp 1679585382
transform 1 0 60480 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_631
timestamp 1679585382
transform 1 0 61152 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_638
timestamp 1679585382
transform 1 0 61824 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_645
timestamp 1679585382
transform 1 0 62496 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_652
timestamp 1679585382
transform 1 0 63168 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_659
timestamp 1679585382
transform 1 0 63840 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_666
timestamp 1679585382
transform 1 0 64512 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_673
timestamp 1679585382
transform 1 0 65184 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_680
timestamp 1679585382
transform 1 0 65856 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_687
timestamp 1679585382
transform 1 0 66528 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_694
timestamp 1679585382
transform 1 0 67200 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_701
timestamp 1679585382
transform 1 0 67872 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_708
timestamp 1679585382
transform 1 0 68544 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_715
timestamp 1679585382
transform 1 0 69216 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_722
timestamp 1679585382
transform 1 0 69888 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_729
timestamp 1679585382
transform 1 0 70560 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_736
timestamp 1679585382
transform 1 0 71232 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_743
timestamp 1679585382
transform 1 0 71904 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_750
timestamp 1679585382
transform 1 0 72576 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_757
timestamp 1679585382
transform 1 0 73248 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_764
timestamp 1679585382
transform 1 0 73920 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_771
timestamp 1679585382
transform 1 0 74592 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_778
timestamp 1679585382
transform 1 0 75264 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_785
timestamp 1679585382
transform 1 0 75936 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_792
timestamp 1679585382
transform 1 0 76608 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_799
timestamp 1679585382
transform 1 0 77280 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_806
timestamp 1679585382
transform 1 0 77952 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_813
timestamp 1679585382
transform 1 0 78624 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_820
timestamp 1679585382
transform 1 0 79296 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_827
timestamp 1679585382
transform 1 0 79968 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_834
timestamp 1679585382
transform 1 0 80640 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_841
timestamp 1679585382
transform 1 0 81312 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_848
timestamp 1679585382
transform 1 0 81984 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_855
timestamp 1679585382
transform 1 0 82656 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_862
timestamp 1679585382
transform 1 0 83328 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_869
timestamp 1679585382
transform 1 0 84000 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_876
timestamp 1679585382
transform 1 0 84672 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_883
timestamp 1679585382
transform 1 0 85344 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_890
timestamp 1679585382
transform 1 0 86016 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_897
timestamp 1679585382
transform 1 0 86688 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_904
timestamp 1679585382
transform 1 0 87360 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_911
timestamp 1679585382
transform 1 0 88032 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_918
timestamp 1679585382
transform 1 0 88704 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_925
timestamp 1679585382
transform 1 0 89376 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_932
timestamp 1679585382
transform 1 0 90048 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_939
timestamp 1679585382
transform 1 0 90720 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_946
timestamp 1679585382
transform 1 0 91392 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_953
timestamp 1679585382
transform 1 0 92064 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_960
timestamp 1679585382
transform 1 0 92736 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_967
timestamp 1679585382
transform 1 0 93408 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_974
timestamp 1679585382
transform 1 0 94080 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_981
timestamp 1679585382
transform 1 0 94752 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_988
timestamp 1679585382
transform 1 0 95424 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_995
timestamp 1679585382
transform 1 0 96096 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1002
timestamp 1679585382
transform 1 0 96768 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1009
timestamp 1679585382
transform 1 0 97440 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1016
timestamp 1679585382
transform 1 0 98112 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_1023
timestamp 1679581501
transform 1 0 98784 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_1027
timestamp 1677583704
transform 1 0 99168 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_43_0
timestamp 1679585382
transform 1 0 576 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_7
timestamp 1679585382
transform 1 0 1248 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_14
timestamp 1679585382
transform 1 0 1920 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_21
timestamp 1679585382
transform 1 0 2592 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_28
timestamp 1679585382
transform 1 0 3264 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_35
timestamp 1679585382
transform 1 0 3936 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_42
timestamp 1679585382
transform 1 0 4608 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_49
timestamp 1679585382
transform 1 0 5280 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_43_56
timestamp 1677583704
transform 1 0 5952 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_43_71
timestamp 1679585382
transform 1 0 7392 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_78
timestamp 1679585382
transform 1 0 8064 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_85
timestamp 1679585382
transform 1 0 8736 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_92
timestamp 1679585382
transform 1 0 9408 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_99
timestamp 1679585382
transform 1 0 10080 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_106
timestamp 1679585382
transform 1 0 10752 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_113
timestamp 1679585382
transform 1 0 11424 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_120
timestamp 1679585382
transform 1 0 12096 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_127
timestamp 1679585382
transform 1 0 12768 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_134
timestamp 1679585382
transform 1 0 13440 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_141
timestamp 1679585382
transform 1 0 14112 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_148
timestamp 1679585382
transform 1 0 14784 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_159
timestamp 1679581501
transform 1 0 15840 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_43_163
timestamp 1677583258
transform 1 0 16224 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_173
timestamp 1679585382
transform 1 0 17184 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_180
timestamp 1679581501
transform 1 0 17856 0 -1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_43_196
timestamp 1679585382
transform 1 0 19392 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_203
timestamp 1679585382
transform 1 0 20064 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_210
timestamp 1679585382
transform 1 0 20736 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_217
timestamp 1679585382
transform 1 0 21408 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_224
timestamp 1679585382
transform 1 0 22080 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_231
timestamp 1679585382
transform 1 0 22752 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_238
timestamp 1679585382
transform 1 0 23424 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_245
timestamp 1679585382
transform 1 0 24096 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_252
timestamp 1679581501
transform 1 0 24768 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_43_259
timestamp 1677583704
transform 1 0 25440 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_43_288
timestamp 1679585382
transform 1 0 28224 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_295
timestamp 1679585382
transform 1 0 28896 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_302
timestamp 1679585382
transform 1 0 29568 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_309
timestamp 1679585382
transform 1 0 30240 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_316
timestamp 1679585382
transform 1 0 30912 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_323
timestamp 1679585382
transform 1 0 31584 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_330
timestamp 1679585382
transform 1 0 32256 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_337
timestamp 1679585382
transform 1 0 32928 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_344
timestamp 1679585382
transform 1 0 33600 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_351
timestamp 1679585382
transform 1 0 34272 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_358
timestamp 1679585382
transform 1 0 34944 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_365
timestamp 1679585382
transform 1 0 35616 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_372
timestamp 1679585382
transform 1 0 36288 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_379
timestamp 1679585382
transform 1 0 36960 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_386
timestamp 1679585382
transform 1 0 37632 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_393
timestamp 1679585382
transform 1 0 38304 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_400
timestamp 1679585382
transform 1 0 38976 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_407
timestamp 1679581501
transform 1 0 39648 0 -1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_43_411
timestamp 1677583704
transform 1 0 40032 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_43_440
timestamp 1679585382
transform 1 0 42816 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_447
timestamp 1679585382
transform 1 0 43488 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_454
timestamp 1679585382
transform 1 0 44160 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_461
timestamp 1679585382
transform 1 0 44832 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_468
timestamp 1679585382
transform 1 0 45504 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_475
timestamp 1679585382
transform 1 0 46176 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_482
timestamp 1679585382
transform 1 0 46848 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_489
timestamp 1679585382
transform 1 0 47520 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_496
timestamp 1679585382
transform 1 0 48192 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_503
timestamp 1679585382
transform 1 0 48864 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_510
timestamp 1679585382
transform 1 0 49536 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_517
timestamp 1679585382
transform 1 0 50208 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_524
timestamp 1679585382
transform 1 0 50880 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_531
timestamp 1679585382
transform 1 0 51552 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_538
timestamp 1679585382
transform 1 0 52224 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_545
timestamp 1679585382
transform 1 0 52896 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_552
timestamp 1679585382
transform 1 0 53568 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_559
timestamp 1679585382
transform 1 0 54240 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_566
timestamp 1679585382
transform 1 0 54912 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_573
timestamp 1679585382
transform 1 0 55584 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_580
timestamp 1679585382
transform 1 0 56256 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_587
timestamp 1679585382
transform 1 0 56928 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_594
timestamp 1679585382
transform 1 0 57600 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_601
timestamp 1679585382
transform 1 0 58272 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_608
timestamp 1679585382
transform 1 0 58944 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_615
timestamp 1679585382
transform 1 0 59616 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_622
timestamp 1679585382
transform 1 0 60288 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_629
timestamp 1679585382
transform 1 0 60960 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_636
timestamp 1679585382
transform 1 0 61632 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_643
timestamp 1679585382
transform 1 0 62304 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_650
timestamp 1679585382
transform 1 0 62976 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_657
timestamp 1679585382
transform 1 0 63648 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_664
timestamp 1679585382
transform 1 0 64320 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_671
timestamp 1679585382
transform 1 0 64992 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_678
timestamp 1679585382
transform 1 0 65664 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_685
timestamp 1679585382
transform 1 0 66336 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_692
timestamp 1679585382
transform 1 0 67008 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_699
timestamp 1679585382
transform 1 0 67680 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_706
timestamp 1679585382
transform 1 0 68352 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_713
timestamp 1679585382
transform 1 0 69024 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_720
timestamp 1679585382
transform 1 0 69696 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_727
timestamp 1679585382
transform 1 0 70368 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_734
timestamp 1679585382
transform 1 0 71040 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_741
timestamp 1679585382
transform 1 0 71712 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_748
timestamp 1679585382
transform 1 0 72384 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_755
timestamp 1679585382
transform 1 0 73056 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_762
timestamp 1679585382
transform 1 0 73728 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_769
timestamp 1679585382
transform 1 0 74400 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_776
timestamp 1679585382
transform 1 0 75072 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_783
timestamp 1679585382
transform 1 0 75744 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_790
timestamp 1679585382
transform 1 0 76416 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_797
timestamp 1679585382
transform 1 0 77088 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_804
timestamp 1679585382
transform 1 0 77760 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_811
timestamp 1679585382
transform 1 0 78432 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_818
timestamp 1679585382
transform 1 0 79104 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_825
timestamp 1679585382
transform 1 0 79776 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_832
timestamp 1679585382
transform 1 0 80448 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_839
timestamp 1679585382
transform 1 0 81120 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_846
timestamp 1679585382
transform 1 0 81792 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_853
timestamp 1679585382
transform 1 0 82464 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_860
timestamp 1679585382
transform 1 0 83136 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_867
timestamp 1679585382
transform 1 0 83808 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_874
timestamp 1679585382
transform 1 0 84480 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_881
timestamp 1679585382
transform 1 0 85152 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_888
timestamp 1679585382
transform 1 0 85824 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_895
timestamp 1679585382
transform 1 0 86496 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_902
timestamp 1679585382
transform 1 0 87168 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_909
timestamp 1679585382
transform 1 0 87840 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_916
timestamp 1679585382
transform 1 0 88512 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_923
timestamp 1679585382
transform 1 0 89184 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_930
timestamp 1679585382
transform 1 0 89856 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_937
timestamp 1679585382
transform 1 0 90528 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_944
timestamp 1679585382
transform 1 0 91200 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_951
timestamp 1679585382
transform 1 0 91872 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_958
timestamp 1679585382
transform 1 0 92544 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_965
timestamp 1679585382
transform 1 0 93216 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_972
timestamp 1679585382
transform 1 0 93888 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_979
timestamp 1679585382
transform 1 0 94560 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_986
timestamp 1679585382
transform 1 0 95232 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_993
timestamp 1679585382
transform 1 0 95904 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1000
timestamp 1679585382
transform 1 0 96576 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1007
timestamp 1679585382
transform 1 0 97248 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1014
timestamp 1679585382
transform 1 0 97920 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1021
timestamp 1679585382
transform 1 0 98592 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_43_1028
timestamp 1677583258
transform 1 0 99264 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_0
timestamp 1679585382
transform 1 0 576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_7
timestamp 1679585382
transform 1 0 1248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_14
timestamp 1679585382
transform 1 0 1920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_21
timestamp 1679585382
transform 1 0 2592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_28
timestamp 1679585382
transform 1 0 3264 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_35
timestamp 1679585382
transform 1 0 3936 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_42
timestamp 1679585382
transform 1 0 4608 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_49
timestamp 1679585382
transform 1 0 5280 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_56
timestamp 1679585382
transform 1 0 5952 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_63
timestamp 1679581501
transform 1 0 6624 0 1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_44_67
timestamp 1677583258
transform 1 0 7008 0 1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_44_72
timestamp 1679581501
transform 1 0 7488 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_44_76
timestamp 1677583704
transform 1 0 7872 0 1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_44_87
timestamp 1677583704
transform 1 0 8928 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_89
timestamp 1677583258
transform 1 0 9120 0 1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_44_98
timestamp 1679581501
transform 1 0 9984 0 1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_44_107
timestamp 1679585382
transform 1 0 10848 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_114
timestamp 1677583704
transform 1 0 11520 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_132
timestamp 1679585382
transform 1 0 13248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_139
timestamp 1679585382
transform 1 0 13920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_146
timestamp 1679585382
transform 1 0 14592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_153
timestamp 1679585382
transform 1 0 15264 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_160
timestamp 1679585382
transform 1 0 15936 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_167
timestamp 1679585382
transform 1 0 16608 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_174
timestamp 1679585382
transform 1 0 17280 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_181
timestamp 1679585382
transform 1 0 17952 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_188
timestamp 1679585382
transform 1 0 18624 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_195
timestamp 1679585382
transform 1 0 19296 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_202
timestamp 1679585382
transform 1 0 19968 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_209
timestamp 1677583704
transform 1 0 20640 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_238
timestamp 1679585382
transform 1 0 23424 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_253
timestamp 1677583704
transform 1 0 24864 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_255
timestamp 1677583258
transform 1 0 25056 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_269
timestamp 1679585382
transform 1 0 26400 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_276
timestamp 1679585382
transform 1 0 27072 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_283
timestamp 1679585382
transform 1 0 27744 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_290
timestamp 1679585382
transform 1 0 28416 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_297
timestamp 1679585382
transform 1 0 29088 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_304
timestamp 1679585382
transform 1 0 29760 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_311
timestamp 1679585382
transform 1 0 30432 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_318
timestamp 1679585382
transform 1 0 31104 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_325
timestamp 1679585382
transform 1 0 31776 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_332
timestamp 1679585382
transform 1 0 32448 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_339
timestamp 1679585382
transform 1 0 33120 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_346
timestamp 1677583704
transform 1 0 33792 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_348
timestamp 1677583258
transform 1 0 33984 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_353
timestamp 1679585382
transform 1 0 34464 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_360
timestamp 1679585382
transform 1 0 35136 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_367
timestamp 1679585382
transform 1 0 35808 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_374
timestamp 1679585382
transform 1 0 36480 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_381
timestamp 1679585382
transform 1 0 37152 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_388
timestamp 1679585382
transform 1 0 37824 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_395
timestamp 1679585382
transform 1 0 38496 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_402
timestamp 1679585382
transform 1 0 39168 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_409
timestamp 1679585382
transform 1 0 39840 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_416
timestamp 1679585382
transform 1 0 40512 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_423
timestamp 1679585382
transform 1 0 41184 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_430
timestamp 1679585382
transform 1 0 41856 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_437
timestamp 1679585382
transform 1 0 42528 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_444
timestamp 1679585382
transform 1 0 43200 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_451
timestamp 1679585382
transform 1 0 43872 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_458
timestamp 1679585382
transform 1 0 44544 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_465
timestamp 1679585382
transform 1 0 45216 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_472
timestamp 1679585382
transform 1 0 45888 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_479
timestamp 1679585382
transform 1 0 46560 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_486
timestamp 1679585382
transform 1 0 47232 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_493
timestamp 1679585382
transform 1 0 47904 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_500
timestamp 1679585382
transform 1 0 48576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_507
timestamp 1679585382
transform 1 0 49248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_514
timestamp 1679585382
transform 1 0 49920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_521
timestamp 1679585382
transform 1 0 50592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_528
timestamp 1679585382
transform 1 0 51264 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_535
timestamp 1679585382
transform 1 0 51936 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_542
timestamp 1679585382
transform 1 0 52608 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_549
timestamp 1679585382
transform 1 0 53280 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_556
timestamp 1679585382
transform 1 0 53952 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_563
timestamp 1679585382
transform 1 0 54624 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_570
timestamp 1679585382
transform 1 0 55296 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_577
timestamp 1679585382
transform 1 0 55968 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_584
timestamp 1679585382
transform 1 0 56640 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_591
timestamp 1679585382
transform 1 0 57312 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_598
timestamp 1679585382
transform 1 0 57984 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_605
timestamp 1679585382
transform 1 0 58656 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_612
timestamp 1679585382
transform 1 0 59328 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_619
timestamp 1679585382
transform 1 0 60000 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_626
timestamp 1679585382
transform 1 0 60672 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_633
timestamp 1679585382
transform 1 0 61344 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_640
timestamp 1679585382
transform 1 0 62016 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_647
timestamp 1679585382
transform 1 0 62688 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_654
timestamp 1679585382
transform 1 0 63360 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_661
timestamp 1679585382
transform 1 0 64032 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_668
timestamp 1679585382
transform 1 0 64704 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_675
timestamp 1679585382
transform 1 0 65376 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_682
timestamp 1679585382
transform 1 0 66048 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_689
timestamp 1679585382
transform 1 0 66720 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_696
timestamp 1679585382
transform 1 0 67392 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_703
timestamp 1679585382
transform 1 0 68064 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_710
timestamp 1679585382
transform 1 0 68736 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_717
timestamp 1679585382
transform 1 0 69408 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_724
timestamp 1679585382
transform 1 0 70080 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_731
timestamp 1679585382
transform 1 0 70752 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_738
timestamp 1679585382
transform 1 0 71424 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_745
timestamp 1679585382
transform 1 0 72096 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_752
timestamp 1679585382
transform 1 0 72768 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_759
timestamp 1679585382
transform 1 0 73440 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_766
timestamp 1679585382
transform 1 0 74112 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_773
timestamp 1679585382
transform 1 0 74784 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_780
timestamp 1679585382
transform 1 0 75456 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_787
timestamp 1679585382
transform 1 0 76128 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_794
timestamp 1679585382
transform 1 0 76800 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_801
timestamp 1679585382
transform 1 0 77472 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_808
timestamp 1679585382
transform 1 0 78144 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_815
timestamp 1679585382
transform 1 0 78816 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_822
timestamp 1679585382
transform 1 0 79488 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_829
timestamp 1679585382
transform 1 0 80160 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_836
timestamp 1679585382
transform 1 0 80832 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_843
timestamp 1679585382
transform 1 0 81504 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_850
timestamp 1679585382
transform 1 0 82176 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_857
timestamp 1679585382
transform 1 0 82848 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_864
timestamp 1679585382
transform 1 0 83520 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_871
timestamp 1679585382
transform 1 0 84192 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_878
timestamp 1679585382
transform 1 0 84864 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_885
timestamp 1679585382
transform 1 0 85536 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_892
timestamp 1679585382
transform 1 0 86208 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_899
timestamp 1679585382
transform 1 0 86880 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_906
timestamp 1679585382
transform 1 0 87552 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_913
timestamp 1679585382
transform 1 0 88224 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_920
timestamp 1679585382
transform 1 0 88896 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_927
timestamp 1679585382
transform 1 0 89568 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_934
timestamp 1679585382
transform 1 0 90240 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_941
timestamp 1679585382
transform 1 0 90912 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_948
timestamp 1679585382
transform 1 0 91584 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_955
timestamp 1679585382
transform 1 0 92256 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_962
timestamp 1679585382
transform 1 0 92928 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_969
timestamp 1679585382
transform 1 0 93600 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_976
timestamp 1679585382
transform 1 0 94272 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_983
timestamp 1679585382
transform 1 0 94944 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_990
timestamp 1679585382
transform 1 0 95616 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_997
timestamp 1679585382
transform 1 0 96288 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1004
timestamp 1679585382
transform 1 0 96960 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1011
timestamp 1679585382
transform 1 0 97632 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1018
timestamp 1679585382
transform 1 0 98304 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_1025
timestamp 1679581501
transform 1 0 98976 0 1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_45_0
timestamp 1679585382
transform 1 0 576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_7
timestamp 1679585382
transform 1 0 1248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_14
timestamp 1679585382
transform 1 0 1920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_21
timestamp 1679585382
transform 1 0 2592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_28
timestamp 1679585382
transform 1 0 3264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_35
timestamp 1679585382
transform 1 0 3936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_42
timestamp 1679585382
transform 1 0 4608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_49
timestamp 1679581501
transform 1 0 5280 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_45_53
timestamp 1677583704
transform 1 0 5664 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_90
timestamp 1679585382
transform 1 0 9216 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_97
timestamp 1679585382
transform 1 0 9888 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_104
timestamp 1679585382
transform 1 0 10560 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_111
timestamp 1679585382
transform 1 0 11232 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_118
timestamp 1679585382
transform 1 0 11904 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_125
timestamp 1679585382
transform 1 0 12576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_132
timestamp 1679585382
transform 1 0 13248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_139
timestamp 1679585382
transform 1 0 13920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_146
timestamp 1679585382
transform 1 0 14592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_153
timestamp 1679585382
transform 1 0 15264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_160
timestamp 1679585382
transform 1 0 15936 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_167
timestamp 1677583704
transform 1 0 16608 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_173
timestamp 1679585382
transform 1 0 17184 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_180
timestamp 1679585382
transform 1 0 17856 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_187
timestamp 1679585382
transform 1 0 18528 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_194
timestamp 1679585382
transform 1 0 19200 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_201
timestamp 1679581501
transform 1 0 19872 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_45_205
timestamp 1677583704
transform 1 0 20256 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_220
timestamp 1679585382
transform 1 0 21696 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_227
timestamp 1679585382
transform 1 0 22368 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_234
timestamp 1679585382
transform 1 0 23040 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_241
timestamp 1679585382
transform 1 0 23712 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_248
timestamp 1679585382
transform 1 0 24384 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_255
timestamp 1679581501
transform 1 0 25056 0 -1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_45_264
timestamp 1679585382
transform 1 0 25920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_271
timestamp 1679585382
transform 1 0 26592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_278
timestamp 1679585382
transform 1 0 27264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_285
timestamp 1679585382
transform 1 0 27936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_292
timestamp 1679585382
transform 1 0 28608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_299
timestamp 1679585382
transform 1 0 29280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_306
timestamp 1679585382
transform 1 0 29952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_313
timestamp 1679585382
transform 1 0 30624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_320
timestamp 1679585382
transform 1 0 31296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_327
timestamp 1679585382
transform 1 0 31968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_334
timestamp 1679581501
transform 1 0 32640 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_45_338
timestamp 1677583258
transform 1 0 33024 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_384
timestamp 1679585382
transform 1 0 37440 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_391
timestamp 1679585382
transform 1 0 38112 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_398
timestamp 1677583704
transform 1 0 38784 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_408
timestamp 1679585382
transform 1 0 39744 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_415
timestamp 1679585382
transform 1 0 40416 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_422
timestamp 1679585382
transform 1 0 41088 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_429
timestamp 1679585382
transform 1 0 41760 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_436
timestamp 1679585382
transform 1 0 42432 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_443
timestamp 1679585382
transform 1 0 43104 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_450
timestamp 1679585382
transform 1 0 43776 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_457
timestamp 1679585382
transform 1 0 44448 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_464
timestamp 1679585382
transform 1 0 45120 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_471
timestamp 1679585382
transform 1 0 45792 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_478
timestamp 1679585382
transform 1 0 46464 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_485
timestamp 1679585382
transform 1 0 47136 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_492
timestamp 1679585382
transform 1 0 47808 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_499
timestamp 1679585382
transform 1 0 48480 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_506
timestamp 1679585382
transform 1 0 49152 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_513
timestamp 1679585382
transform 1 0 49824 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_520
timestamp 1679585382
transform 1 0 50496 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_527
timestamp 1679585382
transform 1 0 51168 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_534
timestamp 1679585382
transform 1 0 51840 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_541
timestamp 1679585382
transform 1 0 52512 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_548
timestamp 1679585382
transform 1 0 53184 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_555
timestamp 1679585382
transform 1 0 53856 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_562
timestamp 1679585382
transform 1 0 54528 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_569
timestamp 1679585382
transform 1 0 55200 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_576
timestamp 1679585382
transform 1 0 55872 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_583
timestamp 1679585382
transform 1 0 56544 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_590
timestamp 1679585382
transform 1 0 57216 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_597
timestamp 1679585382
transform 1 0 57888 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_604
timestamp 1679585382
transform 1 0 58560 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_611
timestamp 1679585382
transform 1 0 59232 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_618
timestamp 1679585382
transform 1 0 59904 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_625
timestamp 1679585382
transform 1 0 60576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_632
timestamp 1679585382
transform 1 0 61248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_639
timestamp 1679585382
transform 1 0 61920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_646
timestamp 1679585382
transform 1 0 62592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_653
timestamp 1679585382
transform 1 0 63264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_660
timestamp 1679585382
transform 1 0 63936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_667
timestamp 1679585382
transform 1 0 64608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_674
timestamp 1679585382
transform 1 0 65280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_681
timestamp 1679585382
transform 1 0 65952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_688
timestamp 1679585382
transform 1 0 66624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_695
timestamp 1679585382
transform 1 0 67296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_702
timestamp 1679585382
transform 1 0 67968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_709
timestamp 1679585382
transform 1 0 68640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_716
timestamp 1679585382
transform 1 0 69312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_723
timestamp 1679585382
transform 1 0 69984 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_730
timestamp 1679585382
transform 1 0 70656 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_737
timestamp 1679585382
transform 1 0 71328 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_744
timestamp 1679585382
transform 1 0 72000 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_751
timestamp 1679585382
transform 1 0 72672 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_758
timestamp 1679585382
transform 1 0 73344 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_765
timestamp 1679585382
transform 1 0 74016 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_772
timestamp 1679585382
transform 1 0 74688 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_779
timestamp 1679585382
transform 1 0 75360 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_786
timestamp 1679585382
transform 1 0 76032 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_793
timestamp 1679585382
transform 1 0 76704 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_800
timestamp 1679585382
transform 1 0 77376 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_807
timestamp 1679585382
transform 1 0 78048 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_814
timestamp 1679585382
transform 1 0 78720 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_821
timestamp 1679585382
transform 1 0 79392 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_828
timestamp 1679585382
transform 1 0 80064 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_835
timestamp 1679585382
transform 1 0 80736 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_842
timestamp 1679585382
transform 1 0 81408 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_849
timestamp 1679585382
transform 1 0 82080 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_856
timestamp 1679585382
transform 1 0 82752 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_863
timestamp 1679585382
transform 1 0 83424 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_870
timestamp 1679585382
transform 1 0 84096 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_877
timestamp 1679585382
transform 1 0 84768 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_884
timestamp 1679585382
transform 1 0 85440 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_891
timestamp 1679585382
transform 1 0 86112 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_898
timestamp 1679585382
transform 1 0 86784 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_905
timestamp 1679585382
transform 1 0 87456 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_912
timestamp 1679585382
transform 1 0 88128 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_919
timestamp 1679585382
transform 1 0 88800 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_926
timestamp 1679585382
transform 1 0 89472 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_933
timestamp 1679585382
transform 1 0 90144 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_940
timestamp 1679585382
transform 1 0 90816 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_947
timestamp 1679585382
transform 1 0 91488 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_954
timestamp 1679585382
transform 1 0 92160 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_961
timestamp 1679585382
transform 1 0 92832 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_968
timestamp 1679585382
transform 1 0 93504 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_975
timestamp 1679585382
transform 1 0 94176 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_982
timestamp 1679585382
transform 1 0 94848 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_989
timestamp 1679585382
transform 1 0 95520 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_996
timestamp 1679585382
transform 1 0 96192 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1003
timestamp 1679585382
transform 1 0 96864 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1010
timestamp 1679585382
transform 1 0 97536 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1017
timestamp 1679585382
transform 1 0 98208 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_1024
timestamp 1679581501
transform 1 0 98880 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_45_1028
timestamp 1677583258
transform 1 0 99264 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_0
timestamp 1679585382
transform 1 0 576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_7
timestamp 1679585382
transform 1 0 1248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_14
timestamp 1679585382
transform 1 0 1920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_21
timestamp 1679585382
transform 1 0 2592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_28
timestamp 1679585382
transform 1 0 3264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_35
timestamp 1679585382
transform 1 0 3936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_42
timestamp 1679585382
transform 1 0 4608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_49
timestamp 1679581501
transform 1 0 5280 0 1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_46_80
timestamp 1679585382
transform 1 0 8256 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_87
timestamp 1679585382
transform 1 0 8928 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_94
timestamp 1679585382
transform 1 0 9600 0 1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_101
timestamp 1677583258
transform 1 0 10272 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_119
timestamp 1679585382
transform 1 0 12000 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_126
timestamp 1679585382
transform 1 0 12672 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_133
timestamp 1679585382
transform 1 0 13344 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_140
timestamp 1679585382
transform 1 0 14016 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_147
timestamp 1679585382
transform 1 0 14688 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_154
timestamp 1679581501
transform 1 0 15360 0 1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_46_194
timestamp 1679585382
transform 1 0 19200 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_201
timestamp 1679585382
transform 1 0 19872 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_208
timestamp 1679585382
transform 1 0 20544 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_215
timestamp 1679581501
transform 1 0 21216 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_219
timestamp 1677583258
transform 1 0 21600 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_224
timestamp 1679585382
transform 1 0 22080 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_231
timestamp 1679585382
transform 1 0 22752 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_238
timestamp 1679585382
transform 1 0 23424 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_245
timestamp 1679585382
transform 1 0 24096 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_252
timestamp 1679585382
transform 1 0 24768 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_259
timestamp 1679585382
transform 1 0 25440 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_270
timestamp 1679585382
transform 1 0 26496 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_277
timestamp 1677583704
transform 1 0 27168 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_310
timestamp 1679585382
transform 1 0 30336 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_317
timestamp 1679585382
transform 1 0 31008 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_324
timestamp 1679585382
transform 1 0 31680 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_331
timestamp 1679585382
transform 1 0 32352 0 1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_338
timestamp 1677583258
transform 1 0 33024 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_366
timestamp 1679585382
transform 1 0 35712 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_373
timestamp 1679585382
transform 1 0 36384 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_380
timestamp 1677583704
transform 1 0 37056 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_382
timestamp 1677583258
transform 1 0 37248 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_387
timestamp 1679585382
transform 1 0 37728 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_394
timestamp 1679585382
transform 1 0 38400 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_401
timestamp 1679581501
transform 1 0 39072 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_405
timestamp 1677583258
transform 1 0 39456 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_410
timestamp 1679585382
transform 1 0 39936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_417
timestamp 1679585382
transform 1 0 40608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_424
timestamp 1679585382
transform 1 0 41280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_431
timestamp 1679585382
transform 1 0 41952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_438
timestamp 1679585382
transform 1 0 42624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_445
timestamp 1679585382
transform 1 0 43296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_452
timestamp 1679585382
transform 1 0 43968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_459
timestamp 1679585382
transform 1 0 44640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_466
timestamp 1679585382
transform 1 0 45312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_473
timestamp 1679585382
transform 1 0 45984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_480
timestamp 1679585382
transform 1 0 46656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_487
timestamp 1679585382
transform 1 0 47328 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_494
timestamp 1679585382
transform 1 0 48000 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_501
timestamp 1679585382
transform 1 0 48672 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_508
timestamp 1679585382
transform 1 0 49344 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_515
timestamp 1679585382
transform 1 0 50016 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_522
timestamp 1679585382
transform 1 0 50688 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_529
timestamp 1679585382
transform 1 0 51360 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_536
timestamp 1679585382
transform 1 0 52032 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_543
timestamp 1679585382
transform 1 0 52704 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_550
timestamp 1679585382
transform 1 0 53376 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_557
timestamp 1679585382
transform 1 0 54048 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_564
timestamp 1679585382
transform 1 0 54720 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_571
timestamp 1679585382
transform 1 0 55392 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_578
timestamp 1679585382
transform 1 0 56064 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_585
timestamp 1679585382
transform 1 0 56736 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_592
timestamp 1679585382
transform 1 0 57408 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_599
timestamp 1679585382
transform 1 0 58080 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_606
timestamp 1679585382
transform 1 0 58752 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_613
timestamp 1679585382
transform 1 0 59424 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_620
timestamp 1679585382
transform 1 0 60096 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_627
timestamp 1679585382
transform 1 0 60768 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_634
timestamp 1679585382
transform 1 0 61440 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_641
timestamp 1679585382
transform 1 0 62112 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_648
timestamp 1679585382
transform 1 0 62784 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_655
timestamp 1679585382
transform 1 0 63456 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_662
timestamp 1679585382
transform 1 0 64128 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_669
timestamp 1679585382
transform 1 0 64800 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_676
timestamp 1679585382
transform 1 0 65472 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_683
timestamp 1679585382
transform 1 0 66144 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_690
timestamp 1679585382
transform 1 0 66816 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_697
timestamp 1679585382
transform 1 0 67488 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_704
timestamp 1679585382
transform 1 0 68160 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_711
timestamp 1679585382
transform 1 0 68832 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_718
timestamp 1679585382
transform 1 0 69504 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_725
timestamp 1679585382
transform 1 0 70176 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_732
timestamp 1679585382
transform 1 0 70848 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_739
timestamp 1679585382
transform 1 0 71520 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_746
timestamp 1679585382
transform 1 0 72192 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_753
timestamp 1679585382
transform 1 0 72864 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_760
timestamp 1679585382
transform 1 0 73536 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_767
timestamp 1679585382
transform 1 0 74208 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_774
timestamp 1679585382
transform 1 0 74880 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_781
timestamp 1679585382
transform 1 0 75552 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_788
timestamp 1679585382
transform 1 0 76224 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_795
timestamp 1679585382
transform 1 0 76896 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_802
timestamp 1679585382
transform 1 0 77568 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_809
timestamp 1679585382
transform 1 0 78240 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_816
timestamp 1679585382
transform 1 0 78912 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_823
timestamp 1679585382
transform 1 0 79584 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_830
timestamp 1679585382
transform 1 0 80256 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_837
timestamp 1679585382
transform 1 0 80928 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_844
timestamp 1679585382
transform 1 0 81600 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_851
timestamp 1679585382
transform 1 0 82272 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_858
timestamp 1679585382
transform 1 0 82944 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_865
timestamp 1679585382
transform 1 0 83616 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_872
timestamp 1679585382
transform 1 0 84288 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_879
timestamp 1679585382
transform 1 0 84960 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_886
timestamp 1679585382
transform 1 0 85632 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_893
timestamp 1679585382
transform 1 0 86304 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_900
timestamp 1679585382
transform 1 0 86976 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_907
timestamp 1679585382
transform 1 0 87648 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_914
timestamp 1679585382
transform 1 0 88320 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_921
timestamp 1679585382
transform 1 0 88992 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_928
timestamp 1679585382
transform 1 0 89664 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_935
timestamp 1679585382
transform 1 0 90336 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_942
timestamp 1679585382
transform 1 0 91008 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_949
timestamp 1679585382
transform 1 0 91680 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_956
timestamp 1679585382
transform 1 0 92352 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_963
timestamp 1679585382
transform 1 0 93024 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_970
timestamp 1679585382
transform 1 0 93696 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_977
timestamp 1679585382
transform 1 0 94368 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_984
timestamp 1679585382
transform 1 0 95040 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_991
timestamp 1679585382
transform 1 0 95712 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_998
timestamp 1679585382
transform 1 0 96384 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1005
timestamp 1679585382
transform 1 0 97056 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1012
timestamp 1679585382
transform 1 0 97728 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1019
timestamp 1679585382
transform 1 0 98400 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_1026
timestamp 1677583704
transform 1 0 99072 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_1028
timestamp 1677583258
transform 1 0 99264 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_0
timestamp 1679585382
transform 1 0 576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_7
timestamp 1679585382
transform 1 0 1248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_14
timestamp 1679585382
transform 1 0 1920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_21
timestamp 1679585382
transform 1 0 2592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_28
timestamp 1679585382
transform 1 0 3264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_35
timestamp 1679585382
transform 1 0 3936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_42
timestamp 1679585382
transform 1 0 4608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_49
timestamp 1679585382
transform 1 0 5280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_56
timestamp 1679585382
transform 1 0 5952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_63
timestamp 1679581501
transform 1 0 6624 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_47_67
timestamp 1677583704
transform 1 0 7008 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_78
timestamp 1679585382
transform 1 0 8064 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_85
timestamp 1679585382
transform 1 0 8736 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_92
timestamp 1679585382
transform 1 0 9408 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_99
timestamp 1679581501
transform 1 0 10080 0 -1 37044
box -48 -56 432 834
use sg13g2_decap_8  FILLER_47_134
timestamp 1679585382
transform 1 0 13440 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_141
timestamp 1679585382
transform 1 0 14112 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_148
timestamp 1679585382
transform 1 0 14784 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_155
timestamp 1679585382
transform 1 0 15456 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_162
timestamp 1679581501
transform 1 0 16128 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_47_166
timestamp 1677583704
transform 1 0 16512 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_195
timestamp 1679585382
transform 1 0 19296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_202
timestamp 1679585382
transform 1 0 19968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_209
timestamp 1679585382
transform 1 0 20640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_216
timestamp 1679581501
transform 1 0 21312 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_47_220
timestamp 1677583258
transform 1 0 21696 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_248
timestamp 1679585382
transform 1 0 24384 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_282
timestamp 1679585382
transform 1 0 27648 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_289
timestamp 1679581501
transform 1 0 28320 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_47_293
timestamp 1677583704
transform 1 0 28704 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_304
timestamp 1679585382
transform 1 0 29760 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_311
timestamp 1679585382
transform 1 0 30432 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_318
timestamp 1679585382
transform 1 0 31104 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_325
timestamp 1679585382
transform 1 0 31776 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_332
timestamp 1679585382
transform 1 0 32448 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_339
timestamp 1679585382
transform 1 0 33120 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_47_346
timestamp 1677583704
transform 1 0 33792 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_348
timestamp 1677583258
transform 1 0 33984 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_4  FILLER_47_353
timestamp 1679581501
transform 1 0 34464 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_47_357
timestamp 1677583704
transform 1 0 34848 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_368
timestamp 1679585382
transform 1 0 35904 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_375
timestamp 1679581501
transform 1 0 36576 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_47_379
timestamp 1677583258
transform 1 0 36960 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_434
timestamp 1679585382
transform 1 0 42240 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_441
timestamp 1679585382
transform 1 0 42912 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_448
timestamp 1679585382
transform 1 0 43584 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_455
timestamp 1679585382
transform 1 0 44256 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_462
timestamp 1679585382
transform 1 0 44928 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_469
timestamp 1679585382
transform 1 0 45600 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_476
timestamp 1679585382
transform 1 0 46272 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_483
timestamp 1679585382
transform 1 0 46944 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_490
timestamp 1679585382
transform 1 0 47616 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_497
timestamp 1679585382
transform 1 0 48288 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_504
timestamp 1679585382
transform 1 0 48960 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_511
timestamp 1679585382
transform 1 0 49632 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_518
timestamp 1679585382
transform 1 0 50304 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_525
timestamp 1679585382
transform 1 0 50976 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_532
timestamp 1679585382
transform 1 0 51648 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_539
timestamp 1679585382
transform 1 0 52320 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_546
timestamp 1679585382
transform 1 0 52992 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_553
timestamp 1679585382
transform 1 0 53664 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_560
timestamp 1679585382
transform 1 0 54336 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_567
timestamp 1679585382
transform 1 0 55008 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_574
timestamp 1679585382
transform 1 0 55680 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_581
timestamp 1679585382
transform 1 0 56352 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_588
timestamp 1679585382
transform 1 0 57024 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_595
timestamp 1679585382
transform 1 0 57696 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_602
timestamp 1679585382
transform 1 0 58368 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_609
timestamp 1679585382
transform 1 0 59040 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_616
timestamp 1679585382
transform 1 0 59712 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_623
timestamp 1679585382
transform 1 0 60384 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_630
timestamp 1679585382
transform 1 0 61056 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_637
timestamp 1679585382
transform 1 0 61728 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_644
timestamp 1679585382
transform 1 0 62400 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_651
timestamp 1679585382
transform 1 0 63072 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_658
timestamp 1679585382
transform 1 0 63744 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_665
timestamp 1679585382
transform 1 0 64416 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_672
timestamp 1679585382
transform 1 0 65088 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_679
timestamp 1679585382
transform 1 0 65760 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_686
timestamp 1679585382
transform 1 0 66432 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_693
timestamp 1679585382
transform 1 0 67104 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_700
timestamp 1679585382
transform 1 0 67776 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_707
timestamp 1679585382
transform 1 0 68448 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_714
timestamp 1679585382
transform 1 0 69120 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_721
timestamp 1679585382
transform 1 0 69792 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_728
timestamp 1679585382
transform 1 0 70464 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_735
timestamp 1679585382
transform 1 0 71136 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_742
timestamp 1679585382
transform 1 0 71808 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_749
timestamp 1679585382
transform 1 0 72480 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_756
timestamp 1679585382
transform 1 0 73152 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_763
timestamp 1679585382
transform 1 0 73824 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_770
timestamp 1679585382
transform 1 0 74496 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_777
timestamp 1679585382
transform 1 0 75168 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_784
timestamp 1679585382
transform 1 0 75840 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_791
timestamp 1679585382
transform 1 0 76512 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_798
timestamp 1679585382
transform 1 0 77184 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_805
timestamp 1679585382
transform 1 0 77856 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_812
timestamp 1679585382
transform 1 0 78528 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_819
timestamp 1679585382
transform 1 0 79200 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_826
timestamp 1679585382
transform 1 0 79872 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_833
timestamp 1679585382
transform 1 0 80544 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_840
timestamp 1679585382
transform 1 0 81216 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_847
timestamp 1679585382
transform 1 0 81888 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_854
timestamp 1679585382
transform 1 0 82560 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_861
timestamp 1679585382
transform 1 0 83232 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_868
timestamp 1679585382
transform 1 0 83904 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_875
timestamp 1679585382
transform 1 0 84576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_882
timestamp 1679585382
transform 1 0 85248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_889
timestamp 1679585382
transform 1 0 85920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_896
timestamp 1679585382
transform 1 0 86592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_903
timestamp 1679585382
transform 1 0 87264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_910
timestamp 1679585382
transform 1 0 87936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_917
timestamp 1679585382
transform 1 0 88608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_924
timestamp 1679585382
transform 1 0 89280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_931
timestamp 1679585382
transform 1 0 89952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_938
timestamp 1679585382
transform 1 0 90624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_945
timestamp 1679585382
transform 1 0 91296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_952
timestamp 1679585382
transform 1 0 91968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_959
timestamp 1679585382
transform 1 0 92640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_966
timestamp 1679585382
transform 1 0 93312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_973
timestamp 1679585382
transform 1 0 93984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_980
timestamp 1679585382
transform 1 0 94656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_987
timestamp 1679585382
transform 1 0 95328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_994
timestamp 1679585382
transform 1 0 96000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1001
timestamp 1679585382
transform 1 0 96672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1008
timestamp 1679585382
transform 1 0 97344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1015
timestamp 1679585382
transform 1 0 98016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1022
timestamp 1679585382
transform 1 0 98688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_0
timestamp 1679585382
transform 1 0 576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_7
timestamp 1679585382
transform 1 0 1248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_14
timestamp 1679585382
transform 1 0 1920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_21
timestamp 1679585382
transform 1 0 2592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_28
timestamp 1679585382
transform 1 0 3264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_35
timestamp 1679585382
transform 1 0 3936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_42
timestamp 1679585382
transform 1 0 4608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_49
timestamp 1679585382
transform 1 0 5280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_56
timestamp 1679585382
transform 1 0 5952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_63
timestamp 1679585382
transform 1 0 6624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_70
timestamp 1679585382
transform 1 0 7296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_77
timestamp 1679585382
transform 1 0 7968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_84
timestamp 1679585382
transform 1 0 8640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_91
timestamp 1679585382
transform 1 0 9312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_98
timestamp 1679585382
transform 1 0 9984 0 1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_48_105
timestamp 1677583704
transform 1 0 10656 0 1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_48_134
timestamp 1679585382
transform 1 0 13440 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_141
timestamp 1679585382
transform 1 0 14112 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_148
timestamp 1679585382
transform 1 0 14784 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_155
timestamp 1679585382
transform 1 0 15456 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_162
timestamp 1679585382
transform 1 0 16128 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_169
timestamp 1679585382
transform 1 0 16800 0 1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_48_176
timestamp 1679581501
transform 1 0 17472 0 1 37044
box -48 -56 432 834
use sg13g2_decap_4  FILLER_48_184
timestamp 1679581501
transform 1 0 18240 0 1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_48_188
timestamp 1677583258
transform 1 0 18624 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_198
timestamp 1679585382
transform 1 0 19584 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_205
timestamp 1679585382
transform 1 0 20256 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_212
timestamp 1679585382
transform 1 0 20928 0 1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_48_219
timestamp 1679581501
transform 1 0 21600 0 1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_48_223
timestamp 1677583258
transform 1 0 21984 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_232
timestamp 1679585382
transform 1 0 22848 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_239
timestamp 1679585382
transform 1 0 23520 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_246
timestamp 1679585382
transform 1 0 24192 0 1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_48_253
timestamp 1679581501
transform 1 0 24864 0 1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_48_257
timestamp 1677583704
transform 1 0 25248 0 1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_48_263
timestamp 1679585382
transform 1 0 25824 0 1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_48_270
timestamp 1677583704
transform 1 0 26496 0 1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_48_281
timestamp 1679585382
transform 1 0 27552 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_288
timestamp 1679585382
transform 1 0 28224 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_295
timestamp 1679585382
transform 1 0 28896 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_302
timestamp 1679585382
transform 1 0 29568 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_309
timestamp 1679585382
transform 1 0 30240 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_316
timestamp 1679585382
transform 1 0 30912 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_323
timestamp 1679585382
transform 1 0 31584 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_330
timestamp 1679585382
transform 1 0 32256 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_337
timestamp 1679585382
transform 1 0 32928 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_344
timestamp 1679585382
transform 1 0 33600 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_351
timestamp 1679585382
transform 1 0 34272 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_358
timestamp 1679585382
transform 1 0 34944 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_365
timestamp 1679585382
transform 1 0 35616 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_372
timestamp 1679585382
transform 1 0 36288 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_379
timestamp 1679585382
transform 1 0 36960 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_386
timestamp 1679585382
transform 1 0 37632 0 1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_48_393
timestamp 1677583704
transform 1 0 38304 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_395
timestamp 1677583258
transform 1 0 38496 0 1 37044
box -48 -56 144 834
use sg13g2_fill_1  FILLER_48_405
timestamp 1677583258
transform 1 0 39456 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_419
timestamp 1679585382
transform 1 0 40800 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_426
timestamp 1679585382
transform 1 0 41472 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_433
timestamp 1679585382
transform 1 0 42144 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_440
timestamp 1679585382
transform 1 0 42816 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_447
timestamp 1679585382
transform 1 0 43488 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_454
timestamp 1679585382
transform 1 0 44160 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_461
timestamp 1679585382
transform 1 0 44832 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_468
timestamp 1679585382
transform 1 0 45504 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_475
timestamp 1679585382
transform 1 0 46176 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_482
timestamp 1679585382
transform 1 0 46848 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_489
timestamp 1679585382
transform 1 0 47520 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_496
timestamp 1679585382
transform 1 0 48192 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_503
timestamp 1679585382
transform 1 0 48864 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_510
timestamp 1679585382
transform 1 0 49536 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_517
timestamp 1679585382
transform 1 0 50208 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_524
timestamp 1679585382
transform 1 0 50880 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_531
timestamp 1679585382
transform 1 0 51552 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_538
timestamp 1679585382
transform 1 0 52224 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_545
timestamp 1679585382
transform 1 0 52896 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_552
timestamp 1679585382
transform 1 0 53568 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_559
timestamp 1679585382
transform 1 0 54240 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_566
timestamp 1679585382
transform 1 0 54912 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_573
timestamp 1679585382
transform 1 0 55584 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_580
timestamp 1679585382
transform 1 0 56256 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_587
timestamp 1679585382
transform 1 0 56928 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_594
timestamp 1679585382
transform 1 0 57600 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_601
timestamp 1679585382
transform 1 0 58272 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_608
timestamp 1679585382
transform 1 0 58944 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_615
timestamp 1679585382
transform 1 0 59616 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_622
timestamp 1679585382
transform 1 0 60288 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_629
timestamp 1679585382
transform 1 0 60960 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_636
timestamp 1679585382
transform 1 0 61632 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_643
timestamp 1679585382
transform 1 0 62304 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_650
timestamp 1679585382
transform 1 0 62976 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_657
timestamp 1679585382
transform 1 0 63648 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_664
timestamp 1679585382
transform 1 0 64320 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_671
timestamp 1679585382
transform 1 0 64992 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_678
timestamp 1679585382
transform 1 0 65664 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_685
timestamp 1679585382
transform 1 0 66336 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_692
timestamp 1679585382
transform 1 0 67008 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_699
timestamp 1679585382
transform 1 0 67680 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_706
timestamp 1679585382
transform 1 0 68352 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_713
timestamp 1679585382
transform 1 0 69024 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_720
timestamp 1679585382
transform 1 0 69696 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_727
timestamp 1679585382
transform 1 0 70368 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_734
timestamp 1679585382
transform 1 0 71040 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_741
timestamp 1679585382
transform 1 0 71712 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_748
timestamp 1679585382
transform 1 0 72384 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_755
timestamp 1679585382
transform 1 0 73056 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_762
timestamp 1679585382
transform 1 0 73728 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_769
timestamp 1679585382
transform 1 0 74400 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_776
timestamp 1679585382
transform 1 0 75072 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_783
timestamp 1679585382
transform 1 0 75744 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_790
timestamp 1679585382
transform 1 0 76416 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_797
timestamp 1679585382
transform 1 0 77088 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_804
timestamp 1679585382
transform 1 0 77760 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_811
timestamp 1679585382
transform 1 0 78432 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_818
timestamp 1679585382
transform 1 0 79104 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_825
timestamp 1679585382
transform 1 0 79776 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_832
timestamp 1679585382
transform 1 0 80448 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_839
timestamp 1679585382
transform 1 0 81120 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_846
timestamp 1679585382
transform 1 0 81792 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_853
timestamp 1679585382
transform 1 0 82464 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_860
timestamp 1679585382
transform 1 0 83136 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_867
timestamp 1679585382
transform 1 0 83808 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_874
timestamp 1679585382
transform 1 0 84480 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_881
timestamp 1679585382
transform 1 0 85152 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_888
timestamp 1679585382
transform 1 0 85824 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_895
timestamp 1679585382
transform 1 0 86496 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_902
timestamp 1679585382
transform 1 0 87168 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_909
timestamp 1679585382
transform 1 0 87840 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_916
timestamp 1679585382
transform 1 0 88512 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_923
timestamp 1679585382
transform 1 0 89184 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_930
timestamp 1679585382
transform 1 0 89856 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_937
timestamp 1679585382
transform 1 0 90528 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_944
timestamp 1679585382
transform 1 0 91200 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_951
timestamp 1679585382
transform 1 0 91872 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_958
timestamp 1679585382
transform 1 0 92544 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_965
timestamp 1679585382
transform 1 0 93216 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_972
timestamp 1679585382
transform 1 0 93888 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_979
timestamp 1679585382
transform 1 0 94560 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_986
timestamp 1679585382
transform 1 0 95232 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_993
timestamp 1679585382
transform 1 0 95904 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1000
timestamp 1679585382
transform 1 0 96576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1007
timestamp 1679585382
transform 1 0 97248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1014
timestamp 1679585382
transform 1 0 97920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1021
timestamp 1679585382
transform 1 0 98592 0 1 37044
box -48 -56 720 834
use sg13g2_fill_1  FILLER_48_1028
timestamp 1677583258
transform 1 0 99264 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_0
timestamp 1679585382
transform 1 0 576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_7
timestamp 1679585382
transform 1 0 1248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_14
timestamp 1679585382
transform 1 0 1920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_21
timestamp 1679585382
transform 1 0 2592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_28
timestamp 1679585382
transform 1 0 3264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_35
timestamp 1679585382
transform 1 0 3936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_42
timestamp 1679585382
transform 1 0 4608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_49
timestamp 1679585382
transform 1 0 5280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_56
timestamp 1679585382
transform 1 0 5952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_63
timestamp 1679585382
transform 1 0 6624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_70
timestamp 1679585382
transform 1 0 7296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_77
timestamp 1679585382
transform 1 0 7968 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_84
timestamp 1679585382
transform 1 0 8640 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_91
timestamp 1679585382
transform 1 0 9312 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_98
timestamp 1679585382
transform 1 0 9984 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_105
timestamp 1679585382
transform 1 0 10656 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_112
timestamp 1679585382
transform 1 0 11328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_128
timestamp 1679585382
transform 1 0 12864 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_135
timestamp 1679585382
transform 1 0 13536 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_142
timestamp 1679585382
transform 1 0 14208 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_149
timestamp 1679585382
transform 1 0 14880 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_156
timestamp 1679585382
transform 1 0 15552 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_163
timestamp 1679585382
transform 1 0 16224 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_170
timestamp 1679585382
transform 1 0 16896 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_177
timestamp 1679585382
transform 1 0 17568 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_184
timestamp 1679585382
transform 1 0 18240 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_191
timestamp 1679585382
transform 1 0 18912 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_198
timestamp 1679585382
transform 1 0 19584 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_205
timestamp 1679585382
transform 1 0 20256 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_212
timestamp 1679585382
transform 1 0 20928 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_219
timestamp 1679585382
transform 1 0 21600 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_226
timestamp 1679585382
transform 1 0 22272 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_233
timestamp 1679585382
transform 1 0 22944 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_240
timestamp 1679585382
transform 1 0 23616 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_247
timestamp 1679585382
transform 1 0 24288 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_254
timestamp 1679585382
transform 1 0 24960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_261
timestamp 1679585382
transform 1 0 25632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_268
timestamp 1679585382
transform 1 0 26304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_275
timestamp 1679585382
transform 1 0 26976 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_282
timestamp 1679585382
transform 1 0 27648 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_289
timestamp 1679585382
transform 1 0 28320 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_296
timestamp 1679585382
transform 1 0 28992 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_303
timestamp 1679585382
transform 1 0 29664 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_310
timestamp 1679585382
transform 1 0 30336 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_317
timestamp 1679585382
transform 1 0 31008 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_324
timestamp 1679585382
transform 1 0 31680 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_331
timestamp 1679585382
transform 1 0 32352 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_338
timestamp 1679585382
transform 1 0 33024 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_345
timestamp 1679585382
transform 1 0 33696 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_352
timestamp 1679585382
transform 1 0 34368 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_359
timestamp 1679585382
transform 1 0 35040 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_366
timestamp 1679585382
transform 1 0 35712 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_373
timestamp 1679585382
transform 1 0 36384 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_380
timestamp 1679585382
transform 1 0 37056 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_387
timestamp 1679585382
transform 1 0 37728 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_394
timestamp 1679585382
transform 1 0 38400 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_401
timestamp 1679585382
transform 1 0 39072 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_408
timestamp 1679585382
transform 1 0 39744 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_415
timestamp 1679585382
transform 1 0 40416 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_422
timestamp 1679585382
transform 1 0 41088 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_429
timestamp 1679585382
transform 1 0 41760 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_436
timestamp 1679585382
transform 1 0 42432 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_443
timestamp 1679585382
transform 1 0 43104 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_450
timestamp 1679585382
transform 1 0 43776 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_457
timestamp 1679585382
transform 1 0 44448 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_464
timestamp 1679585382
transform 1 0 45120 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_471
timestamp 1679585382
transform 1 0 45792 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_478
timestamp 1679585382
transform 1 0 46464 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_485
timestamp 1679585382
transform 1 0 47136 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_492
timestamp 1679585382
transform 1 0 47808 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_499
timestamp 1679585382
transform 1 0 48480 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_506
timestamp 1679585382
transform 1 0 49152 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_513
timestamp 1679585382
transform 1 0 49824 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_520
timestamp 1679585382
transform 1 0 50496 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_527
timestamp 1679585382
transform 1 0 51168 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_534
timestamp 1679585382
transform 1 0 51840 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_541
timestamp 1679585382
transform 1 0 52512 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_548
timestamp 1679585382
transform 1 0 53184 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_555
timestamp 1679585382
transform 1 0 53856 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_562
timestamp 1679585382
transform 1 0 54528 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_569
timestamp 1679585382
transform 1 0 55200 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_576
timestamp 1679585382
transform 1 0 55872 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_583
timestamp 1679585382
transform 1 0 56544 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_590
timestamp 1679585382
transform 1 0 57216 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_597
timestamp 1679585382
transform 1 0 57888 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_604
timestamp 1679585382
transform 1 0 58560 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_611
timestamp 1679585382
transform 1 0 59232 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_618
timestamp 1679585382
transform 1 0 59904 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_625
timestamp 1679585382
transform 1 0 60576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_632
timestamp 1679585382
transform 1 0 61248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_639
timestamp 1679585382
transform 1 0 61920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_646
timestamp 1679585382
transform 1 0 62592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_653
timestamp 1679585382
transform 1 0 63264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_660
timestamp 1679585382
transform 1 0 63936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_667
timestamp 1679585382
transform 1 0 64608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_674
timestamp 1679585382
transform 1 0 65280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_681
timestamp 1679585382
transform 1 0 65952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_688
timestamp 1679585382
transform 1 0 66624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_695
timestamp 1679585382
transform 1 0 67296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_702
timestamp 1679585382
transform 1 0 67968 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_709
timestamp 1679585382
transform 1 0 68640 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_716
timestamp 1679585382
transform 1 0 69312 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_723
timestamp 1679585382
transform 1 0 69984 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_730
timestamp 1679585382
transform 1 0 70656 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_737
timestamp 1679585382
transform 1 0 71328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_744
timestamp 1679585382
transform 1 0 72000 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_751
timestamp 1679585382
transform 1 0 72672 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_758
timestamp 1679585382
transform 1 0 73344 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_765
timestamp 1679585382
transform 1 0 74016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_772
timestamp 1679585382
transform 1 0 74688 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_779
timestamp 1679585382
transform 1 0 75360 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_786
timestamp 1679585382
transform 1 0 76032 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_793
timestamp 1679585382
transform 1 0 76704 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_800
timestamp 1679585382
transform 1 0 77376 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_807
timestamp 1679585382
transform 1 0 78048 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_814
timestamp 1679585382
transform 1 0 78720 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_821
timestamp 1679585382
transform 1 0 79392 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_828
timestamp 1679585382
transform 1 0 80064 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_835
timestamp 1679585382
transform 1 0 80736 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_842
timestamp 1679585382
transform 1 0 81408 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_849
timestamp 1679585382
transform 1 0 82080 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_856
timestamp 1679585382
transform 1 0 82752 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_863
timestamp 1679585382
transform 1 0 83424 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_870
timestamp 1679585382
transform 1 0 84096 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_877
timestamp 1679585382
transform 1 0 84768 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_884
timestamp 1679585382
transform 1 0 85440 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_891
timestamp 1679585382
transform 1 0 86112 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_898
timestamp 1679585382
transform 1 0 86784 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_905
timestamp 1679585382
transform 1 0 87456 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_912
timestamp 1679585382
transform 1 0 88128 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_919
timestamp 1679585382
transform 1 0 88800 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_926
timestamp 1679585382
transform 1 0 89472 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_933
timestamp 1679585382
transform 1 0 90144 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_940
timestamp 1679585382
transform 1 0 90816 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_947
timestamp 1679585382
transform 1 0 91488 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_954
timestamp 1679585382
transform 1 0 92160 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_961
timestamp 1679585382
transform 1 0 92832 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_968
timestamp 1679585382
transform 1 0 93504 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_975
timestamp 1679585382
transform 1 0 94176 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_982
timestamp 1679585382
transform 1 0 94848 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_989
timestamp 1679585382
transform 1 0 95520 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_996
timestamp 1679585382
transform 1 0 96192 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1003
timestamp 1679585382
transform 1 0 96864 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1010
timestamp 1679585382
transform 1 0 97536 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1017
timestamp 1679585382
transform 1 0 98208 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_1024
timestamp 1679581501
transform 1 0 98880 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_49_1028
timestamp 1677583258
transform 1 0 99264 0 -1 38556
box -48 -56 144 834
use sg13g2_tielo  heichips25_template_5
timestamp 1680004237
transform -1 0 960 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_6
timestamp 1680004237
transform -1 0 960 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_7
timestamp 1680004237
transform -1 0 960 0 -1 11340
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_8
timestamp 1680004237
transform -1 0 960 0 1 11340
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_9
timestamp 1680004237
transform -1 0 960 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_10
timestamp 1680004237
transform -1 0 960 0 1 12852
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_11
timestamp 1680004237
transform -1 0 960 0 1 14364
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_12
timestamp 1680004237
transform -1 0 960 0 -1 15876
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_13
timestamp 1680004237
transform -1 0 960 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_14
timestamp 1680004237
transform -1 0 960 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_15
timestamp 1680004237
transform -1 0 960 0 -1 8316
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_16
timestamp 1680004237
transform -1 0 960 0 1 8316
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_17
timestamp 1680004251
transform -1 0 960 0 1 15876
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_18
timestamp 1680004251
transform -1 0 960 0 -1 17388
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_19
timestamp 1680004251
transform -1 0 960 0 1 17388
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_20
timestamp 1680004251
transform -1 0 960 0 -1 18900
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_21
timestamp 1680004251
transform -1 0 960 0 1 18900
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_22
timestamp 1680004251
transform -1 0 960 0 -1 20412
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_23
timestamp 1680004251
transform -1 0 960 0 1 20412
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_24
timestamp 1680004251
transform -1 0 960 0 1 21924
box -48 -56 432 834
use sg13g2_dlygate4sd3_1  hold1
timestamp 1677675658
transform -1 0 8160 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold2
timestamp 1677675658
transform -1 0 10752 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold3
timestamp 1677675658
transform 1 0 16992 0 -1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold4
timestamp 1677675658
transform 1 0 12096 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold5
timestamp 1677675658
transform 1 0 9120 0 1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold6
timestamp 1677675658
transform 1 0 26976 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold7
timestamp 1677675658
transform 1 0 24288 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold8
timestamp 1677675658
transform -1 0 13056 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold9
timestamp 1677675658
transform 1 0 20448 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold10
timestamp 1677675658
transform 1 0 15072 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold11
timestamp 1677675658
transform 1 0 21024 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold12
timestamp 1677675658
transform 1 0 25536 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold13
timestamp 1677675658
transform -1 0 51072 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold14
timestamp 1677675658
transform -1 0 43488 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold15
timestamp 1677675658
transform -1 0 29760 0 -1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold16
timestamp 1677675658
transform -1 0 56736 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold17
timestamp 1677675658
transform -1 0 4320 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold18
timestamp 1677675658
transform -1 0 8448 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold19
timestamp 1677675658
transform -1 0 4320 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold20
timestamp 1677675658
transform -1 0 57408 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold21
timestamp 1677675658
transform -1 0 8064 0 -1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold22
timestamp 1677675658
transform -1 0 40512 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold23
timestamp 1677675658
transform -1 0 27648 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold24
timestamp 1677675658
transform -1 0 32256 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold25
timestamp 1677675658
transform -1 0 4992 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold26
timestamp 1677675658
transform -1 0 4224 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold27
timestamp 1677675658
transform -1 0 40800 0 1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold28
timestamp 1677675658
transform -1 0 17184 0 -1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold29
timestamp 1677675658
transform -1 0 25440 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold30
timestamp 1677675658
transform 1 0 38784 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold31
timestamp 1677675658
transform -1 0 33600 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold32
timestamp 1677675658
transform -1 0 12864 0 -1 38556
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold33
timestamp 1677675658
transform 1 0 6624 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold34
timestamp 1677675658
transform -1 0 19200 0 1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold35
timestamp 1677675658
transform -1 0 51072 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold36
timestamp 1677675658
transform -1 0 35904 0 -1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold37
timestamp 1677675658
transform -1 0 58752 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold38
timestamp 1677675658
transform -1 0 4992 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold39
timestamp 1677675658
transform -1 0 48000 0 -1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold40
timestamp 1677675658
transform -1 0 40320 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold41
timestamp 1677675658
transform 1 0 9792 0 1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold42
timestamp 1677675658
transform -1 0 56640 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold43
timestamp 1677675658
transform -1 0 40608 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold44
timestamp 1677675658
transform -1 0 40800 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold45
timestamp 1677675658
transform -1 0 16032 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold46
timestamp 1677675658
transform 1 0 15168 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold47
timestamp 1677675658
transform 1 0 28704 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold48
timestamp 1677675658
transform -1 0 26688 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold49
timestamp 1677675658
transform 1 0 45504 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold50
timestamp 1677675658
transform -1 0 46368 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold51
timestamp 1677675658
transform -1 0 4416 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold52
timestamp 1677675658
transform -1 0 19584 0 1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold53
timestamp 1677675658
transform -1 0 27360 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold54
timestamp 1677675658
transform -1 0 25920 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold55
timestamp 1677675658
transform -1 0 50208 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold56
timestamp 1677675658
transform -1 0 9696 0 -1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold57
timestamp 1677675658
transform 1 0 18336 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold58
timestamp 1677675658
transform 1 0 19488 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold59
timestamp 1677675658
transform 1 0 13440 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold60
timestamp 1677675658
transform 1 0 14496 0 -1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold61
timestamp 1677675658
transform 1 0 34848 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold62
timestamp 1677675658
transform 1 0 36864 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold63
timestamp 1677675658
transform 1 0 51936 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold64
timestamp 1677675658
transform -1 0 51360 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold65
timestamp 1677675658
transform 1 0 16416 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold66
timestamp 1677675658
transform -1 0 16800 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold67
timestamp 1677675658
transform -1 0 27744 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold68
timestamp 1677675658
transform -1 0 13152 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold69
timestamp 1677675658
transform -1 0 5280 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold70
timestamp 1677675658
transform -1 0 41760 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold71
timestamp 1677675658
transform 1 0 35712 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold72
timestamp 1677675658
transform -1 0 58464 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold73
timestamp 1677675658
transform 1 0 37056 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold74
timestamp 1677675658
transform -1 0 36768 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold75
timestamp 1677675658
transform -1 0 27552 0 1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold76
timestamp 1677675658
transform -1 0 53856 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold77
timestamp 1677675658
transform -1 0 5184 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold78
timestamp 1677675658
transform -1 0 32064 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold79
timestamp 1677675658
transform -1 0 34560 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold80
timestamp 1677675658
transform -1 0 12000 0 1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold81
timestamp 1677675658
transform -1 0 19968 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold82
timestamp 1677675658
transform -1 0 5280 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold83
timestamp 1677675658
transform -1 0 13824 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold84
timestamp 1677675658
transform -1 0 30240 0 1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold85
timestamp 1677675658
transform -1 0 53088 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold86
timestamp 1677675658
transform -1 0 31200 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold87
timestamp 1677675658
transform -1 0 27072 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold88
timestamp 1677675658
transform -1 0 49344 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold89
timestamp 1677675658
transform -1 0 55488 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold90
timestamp 1677675658
transform -1 0 5088 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold91
timestamp 1677675658
transform -1 0 39456 0 1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold92
timestamp 1677675658
transform -1 0 39456 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold93
timestamp 1677675658
transform -1 0 46464 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold94
timestamp 1677675658
transform -1 0 49056 0 -1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold95
timestamp 1677675658
transform -1 0 41664 0 -1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold96
timestamp 1677675658
transform 1 0 40608 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold97
timestamp 1677675658
transform -1 0 34752 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold98
timestamp 1677675658
transform -1 0 8928 0 1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold99
timestamp 1677675658
transform -1 0 6432 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold100
timestamp 1677675658
transform -1 0 48960 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold101
timestamp 1677675658
transform 1 0 38208 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold102
timestamp 1677675658
transform -1 0 12480 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold103
timestamp 1677675658
transform 1 0 39456 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold104
timestamp 1677675658
transform -1 0 38784 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold105
timestamp 1677675658
transform -1 0 5184 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold106
timestamp 1677675658
transform -1 0 19968 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold107
timestamp 1677675658
transform -1 0 13056 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold108
timestamp 1677675658
transform -1 0 26784 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold109
timestamp 1677675658
transform -1 0 44544 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold110
timestamp 1677675658
transform -1 0 23616 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold111
timestamp 1677675658
transform 1 0 46752 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold112
timestamp 1677675658
transform -1 0 45120 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold113
timestamp 1677675658
transform 1 0 22272 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold114
timestamp 1677675658
transform -1 0 21216 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold115
timestamp 1677675658
transform 1 0 28704 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold116
timestamp 1677675658
transform -1 0 23712 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold117
timestamp 1677675658
transform -1 0 33024 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold118
timestamp 1677675658
transform -1 0 31104 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold119
timestamp 1677675658
transform -1 0 29472 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold120
timestamp 1677675658
transform 1 0 18912 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold121
timestamp 1677675658
transform 1 0 19296 0 1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold122
timestamp 1677675658
transform 1 0 21216 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold123
timestamp 1677675658
transform -1 0 48672 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold124
timestamp 1677675658
transform -1 0 48096 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold125
timestamp 1677675658
transform 1 0 40224 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold126
timestamp 1677675658
transform -1 0 42240 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold127
timestamp 1677675658
transform 1 0 38880 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold128
timestamp 1677675658
transform -1 0 41856 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold129
timestamp 1677675658
transform 1 0 12000 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold130
timestamp 1677675658
transform -1 0 13632 0 -1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold131
timestamp 1677675658
transform 1 0 25248 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold132
timestamp 1677675658
transform 1 0 27360 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold133
timestamp 1677675658
transform -1 0 36864 0 -1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold134
timestamp 1677675658
transform 1 0 36288 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold135
timestamp 1677675658
transform -1 0 19488 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold136
timestamp 1677675658
transform 1 0 18912 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold137
timestamp 1677675658
transform -1 0 52896 0 -1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold138
timestamp 1677675658
transform -1 0 52416 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold139
timestamp 1677675658
transform 1 0 28320 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold140
timestamp 1677675658
transform 1 0 29664 0 -1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold141
timestamp 1677675658
transform 1 0 12768 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold142
timestamp 1677675658
transform 1 0 13440 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold143
timestamp 1677675658
transform 1 0 45216 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold144
timestamp 1677675658
transform 1 0 47904 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold145
timestamp 1677675658
transform 1 0 37920 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold146
timestamp 1677675658
transform -1 0 37056 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold147
timestamp 1677675658
transform 1 0 39840 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold148
timestamp 1677675658
transform -1 0 39168 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold149
timestamp 1677675658
transform 1 0 21792 0 1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold150
timestamp 1677675658
transform -1 0 21792 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold151
timestamp 1677675658
transform 1 0 15840 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold152
timestamp 1677675658
transform -1 0 19776 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold153
timestamp 1677675658
transform -1 0 32448 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold154
timestamp 1677675658
transform -1 0 26784 0 1 6804
box -48 -56 912 834
use sg13g2_buf_1  output1
timestamp 1676385511
transform -1 0 960 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  output2
timestamp 1676385511
transform -1 0 960 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  output3
timestamp 1676385511
transform -1 0 960 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  output4
timestamp 1676385511
transform -1 0 960 0 -1 5292
box -48 -56 432 834
<< labels >>
flabel metal6 s 4316 630 4756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 19436 630 19876 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 34556 630 34996 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 49676 630 50116 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 64796 630 65236 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 79916 630 80356 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 95036 630 95476 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 3076 712 3516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 18196 712 18636 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 33316 712 33756 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 48436 712 48876 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 63556 712 63996 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 78676 712 79116 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 93796 712 94236 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 36668 80 36748 0 FreeSans 320 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 0 35828 80 35908 0 FreeSans 320 0 0 0 ena
port 3 nsew signal input
flabel metal3 s 0 37508 80 37588 0 FreeSans 320 0 0 0 rst_n
port 4 nsew signal input
flabel metal3 s 0 22388 80 22468 0 FreeSans 320 0 0 0 ui_in[0]
port 5 nsew signal input
flabel metal3 s 0 23228 80 23308 0 FreeSans 320 0 0 0 ui_in[1]
port 6 nsew signal input
flabel metal3 s 0 24068 80 24148 0 FreeSans 320 0 0 0 ui_in[2]
port 7 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 ui_in[3]
port 8 nsew signal input
flabel metal3 s 0 25748 80 25828 0 FreeSans 320 0 0 0 ui_in[4]
port 9 nsew signal input
flabel metal3 s 0 26588 80 26668 0 FreeSans 320 0 0 0 ui_in[5]
port 10 nsew signal input
flabel metal3 s 0 27428 80 27508 0 FreeSans 320 0 0 0 ui_in[6]
port 11 nsew signal input
flabel metal3 s 0 28268 80 28348 0 FreeSans 320 0 0 0 ui_in[7]
port 12 nsew signal input
flabel metal3 s 0 29108 80 29188 0 FreeSans 320 0 0 0 uio_in[0]
port 13 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 uio_in[1]
port 14 nsew signal input
flabel metal3 s 0 30788 80 30868 0 FreeSans 320 0 0 0 uio_in[2]
port 15 nsew signal input
flabel metal3 s 0 31628 80 31708 0 FreeSans 320 0 0 0 uio_in[3]
port 16 nsew signal input
flabel metal3 s 0 32468 80 32548 0 FreeSans 320 0 0 0 uio_in[4]
port 17 nsew signal input
flabel metal3 s 0 33308 80 33388 0 FreeSans 320 0 0 0 uio_in[5]
port 18 nsew signal input
flabel metal3 s 0 34148 80 34228 0 FreeSans 320 0 0 0 uio_in[6]
port 19 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 uio_in[7]
port 20 nsew signal input
flabel metal3 s 0 15668 80 15748 0 FreeSans 320 0 0 0 uio_oe[0]
port 21 nsew signal output
flabel metal3 s 0 16508 80 16588 0 FreeSans 320 0 0 0 uio_oe[1]
port 22 nsew signal output
flabel metal3 s 0 17348 80 17428 0 FreeSans 320 0 0 0 uio_oe[2]
port 23 nsew signal output
flabel metal3 s 0 18188 80 18268 0 FreeSans 320 0 0 0 uio_oe[3]
port 24 nsew signal output
flabel metal3 s 0 19028 80 19108 0 FreeSans 320 0 0 0 uio_oe[4]
port 25 nsew signal output
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 uio_oe[5]
port 26 nsew signal output
flabel metal3 s 0 20708 80 20788 0 FreeSans 320 0 0 0 uio_oe[6]
port 27 nsew signal output
flabel metal3 s 0 21548 80 21628 0 FreeSans 320 0 0 0 uio_oe[7]
port 28 nsew signal output
flabel metal3 s 0 8948 80 9028 0 FreeSans 320 0 0 0 uio_out[0]
port 29 nsew signal output
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 uio_out[1]
port 30 nsew signal output
flabel metal3 s 0 10628 80 10708 0 FreeSans 320 0 0 0 uio_out[2]
port 31 nsew signal output
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 uio_out[3]
port 32 nsew signal output
flabel metal3 s 0 12308 80 12388 0 FreeSans 320 0 0 0 uio_out[4]
port 33 nsew signal output
flabel metal3 s 0 13148 80 13228 0 FreeSans 320 0 0 0 uio_out[5]
port 34 nsew signal output
flabel metal3 s 0 13988 80 14068 0 FreeSans 320 0 0 0 uio_out[6]
port 35 nsew signal output
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 uio_out[7]
port 36 nsew signal output
flabel metal3 s 0 2228 80 2308 0 FreeSans 320 0 0 0 uo_out[0]
port 37 nsew signal output
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 uo_out[1]
port 38 nsew signal output
flabel metal3 s 0 3908 80 3988 0 FreeSans 320 0 0 0 uo_out[2]
port 39 nsew signal output
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 uo_out[3]
port 40 nsew signal output
flabel metal3 s 0 5588 80 5668 0 FreeSans 320 0 0 0 uo_out[4]
port 41 nsew signal output
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 uo_out[5]
port 42 nsew signal output
flabel metal3 s 0 7268 80 7348 0 FreeSans 320 0 0 0 uo_out[6]
port 43 nsew signal output
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 uo_out[7]
port 44 nsew signal output
rlabel via1 49968 38556 49968 38556 0 VGND
rlabel metal1 49968 37800 49968 37800 0 VPWR
rlabel metal2 44832 22512 44832 22512 0 DP_1.matrix\[0\]
rlabel metal2 28224 22806 28224 22806 0 DP_1.matrix\[10\]
rlabel metal2 30096 12684 30096 12684 0 DP_1.matrix\[18\]
rlabel metal2 33648 10416 33648 10416 0 DP_1.matrix\[19\]
rlabel metal2 40416 26838 40416 26838 0 DP_1.matrix\[1\]
rlabel metal2 27600 18732 27600 18732 0 DP_1.matrix\[27\]
rlabel metal2 27360 20496 27360 20496 0 DP_1.matrix\[28\]
rlabel metal2 55200 10710 55200 10710 0 DP_1.matrix\[36\]
rlabel metal2 58704 14196 58704 14196 0 DP_1.matrix\[37\]
rlabel metal2 49248 18018 49248 18018 0 DP_1.matrix\[45\]
rlabel metal2 50160 21588 50160 21588 0 DP_1.matrix\[46\]
rlabel metal3 37056 3612 37056 3612 0 DP_1.matrix\[54\]
rlabel metal2 39024 2856 39024 2856 0 DP_1.matrix\[55\]
rlabel metal3 54384 6636 54384 6636 0 DP_1.matrix\[63\]
rlabel metal2 56832 3864 56832 3864 0 DP_1.matrix\[64\]
rlabel metal2 13728 4074 13728 4074 0 DP_1.matrix\[72\]
rlabel metal2 9888 2646 9888 2646 0 DP_1.matrix\[73\]
rlabel metal2 34608 22512 34608 22512 0 DP_1.matrix\[9\]
rlabel metal2 39312 24024 39312 24024 0 DP_2.matrix\[0\]
rlabel metal2 33312 26544 33312 26544 0 DP_2.matrix\[10\]
rlabel metal3 34224 11928 34224 11928 0 DP_2.matrix\[18\]
rlabel metal2 26304 13734 26304 13734 0 DP_2.matrix\[19\]
rlabel metal2 43392 23058 43392 23058 0 DP_2.matrix\[1\]
rlabel metal2 23472 17976 23472 17976 0 DP_2.matrix\[27\]
rlabel metal2 25152 17472 25152 17472 0 DP_2.matrix\[28\]
rlabel metal2 58368 12768 58368 12768 0 DP_2.matrix\[36\]
rlabel metal2 57312 9912 57312 9912 0 DP_2.matrix\[37\]
rlabel metal2 48864 19488 48864 19488 0 DP_2.matrix\[45\]
rlabel metal2 50928 21588 50928 21588 0 DP_2.matrix\[46\]
rlabel metal2 41712 2856 41712 2856 0 DP_2.matrix\[54\]
rlabel metal2 40176 5880 40176 5880 0 DP_2.matrix\[55\]
rlabel metal2 52944 2856 52944 2856 0 DP_2.matrix\[63\]
rlabel metal2 57216 5250 57216 5250 0 DP_2.matrix\[64\]
rlabel metal2 13632 4998 13632 4998 0 DP_2.matrix\[72\]
rlabel metal2 9600 2562 9600 2562 0 DP_2.matrix\[73\]
rlabel metal2 32400 21756 32400 21756 0 DP_2.matrix\[9\]
rlabel metal2 5136 21756 5136 21756 0 DP_3.matrix\[0\]
rlabel metal2 6720 17766 6720 17766 0 DP_3.matrix\[10\]
rlabel metal2 8784 34356 8784 34356 0 DP_3.matrix\[18\]
rlabel metal2 13344 37926 13344 37926 0 DP_3.matrix\[19\]
rlabel metal2 4848 25536 4848 25536 0 DP_3.matrix\[1\]
rlabel metal2 6336 27090 6336 27090 0 DP_3.matrix\[27\]
rlabel metal2 4224 32340 4224 32340 0 DP_3.matrix\[28\]
rlabel metal2 19920 29820 19920 29820 0 DP_3.matrix\[36\]
rlabel metal2 19104 35910 19104 35910 0 DP_3.matrix\[37\]
rlabel metal2 27504 36876 27504 36876 0 DP_3.matrix\[45\]
rlabel metal2 19200 37128 19200 37128 0 DP_3.matrix\[46\]
rlabel metal3 49248 31500 49248 31500 0 DP_3.matrix\[54\]
rlabel metal3 48672 27048 48672 27048 0 DP_3.matrix\[55\]
rlabel metal2 39552 37128 39552 37128 0 DP_3.matrix\[63\]
rlabel metal2 35616 36414 35616 36414 0 DP_3.matrix\[64\]
rlabel metal2 5088 8820 5088 8820 0 DP_3.matrix\[72\]
rlabel metal2 4512 13734 4512 13734 0 DP_3.matrix\[73\]
rlabel metal2 13344 18270 13344 18270 0 DP_3.matrix\[9\]
rlabel metal2 5136 23268 5136 23268 0 DP_4.matrix\[0\]
rlabel metal2 8064 17472 8064 17472 0 DP_4.matrix\[10\]
rlabel metal2 11904 36204 11904 36204 0 DP_4.matrix\[18\]
rlabel metal2 8064 36120 8064 36120 0 DP_4.matrix\[19\]
rlabel metal2 4128 18984 4128 18984 0 DP_4.matrix\[1\]
rlabel metal2 5088 30912 5088 30912 0 DP_4.matrix\[27\]
rlabel metal2 4704 28854 4704 28854 0 DP_4.matrix\[28\]
rlabel metal2 19872 31878 19872 31878 0 DP_4.matrix\[36\]
rlabel metal2 16896 33390 16896 33390 0 DP_4.matrix\[37\]
rlabel metal3 26352 25536 26352 25536 0 DP_4.matrix\[45\]
rlabel metal2 30240 36414 30240 36414 0 DP_4.matrix\[46\]
rlabel metal2 46176 28056 46176 28056 0 DP_4.matrix\[54\]
rlabel metal2 51552 31080 51552 31080 0 DP_4.matrix\[55\]
rlabel metal2 35808 35154 35808 35154 0 DP_4.matrix\[63\]
rlabel metal2 40704 37128 40704 37128 0 DP_4.matrix\[64\]
rlabel metal2 4992 11970 4992 11970 0 DP_4.matrix\[72\]
rlabel metal2 4368 8904 4368 8904 0 DP_4.matrix\[73\]
rlabel metal2 12384 16506 12384 16506 0 DP_4.matrix\[9\]
rlabel metal2 21120 20454 21120 20454 0 _000_
rlabel metal2 21696 22218 21696 22218 0 _001_
rlabel metal2 40704 18816 40704 18816 0 _002_
rlabel metal3 41238 19992 41238 19992 0 _003_
rlabel metal2 36960 14280 36960 14280 0 _004_
rlabel metal2 36384 16674 36384 16674 0 _005_
rlabel metal2 51264 14070 51264 14070 0 _006_
rlabel metal2 52320 14742 52320 14742 0 _007_
rlabel metal2 45360 6636 45360 6636 0 _008_
rlabel metal3 47712 6468 47712 6468 0 _009_
rlabel metal2 40704 12348 40704 12348 0 _010_
rlabel metal2 41280 14280 41280 14280 0 _011_
rlabel metal3 46128 9660 46128 9660 0 _012_
rlabel metal2 48000 10206 48000 10206 0 _013_
rlabel metal2 38688 7602 38688 7602 0 _014_
rlabel metal2 39072 8694 39072 8694 0 _015_
rlabel metal2 29472 8148 29472 8148 0 _016_
rlabel metal3 26016 6972 26016 6972 0 _017_
rlabel metal3 26688 7182 26688 7182 0 _018_
rlabel metal3 20736 12516 20736 12516 0 _019_
rlabel metal2 16512 10878 16512 10878 0 _020_
rlabel metal2 19680 12474 19680 12474 0 _021_
rlabel metal2 14976 22218 14976 22218 0 _022_
rlabel metal2 13728 23520 13728 23520 0 _023_
rlabel metal2 14592 27678 14592 27678 0 _024_
rlabel metal2 13104 27636 13104 27636 0 _025_
rlabel metal2 25824 30702 25824 30702 0 _026_
rlabel metal2 27456 32802 27456 32802 0 _027_
rlabel metal2 37248 30198 37248 30198 0 _028_
rlabel metal2 36960 31626 36960 31626 0 _029_
rlabel metal2 19584 23142 19584 23142 0 _030_
rlabel metal3 18576 25536 18576 25536 0 _031_
rlabel metal2 27744 28224 27744 28224 0 _032_
rlabel metal2 29760 27888 29760 27888 0 _033_
rlabel metal3 36096 33180 36096 33180 0 _034_
rlabel metal2 40320 34524 40320 34524 0 _035_
rlabel metal3 21168 30744 21168 30744 0 _036_
rlabel metal2 19200 34062 19200 34062 0 _037_
rlabel metal2 4800 8946 4800 8946 0 _038_
rlabel metal2 5664 12054 5664 12054 0 _039_
rlabel metal2 12096 18858 12096 18858 0 _040_
rlabel metal2 8736 19404 8736 19404 0 _041_
rlabel metal2 37440 22260 37440 22260 0 _042_
rlabel metal2 41376 25662 41376 25662 0 _043_
rlabel metal3 35088 20076 35088 20076 0 _044_
rlabel metal2 32832 25074 32832 25074 0 _045_
rlabel metal2 32544 13734 32544 13734 0 _046_
rlabel metal2 30624 15330 30624 15330 0 _047_
rlabel metal3 29184 17136 29184 17136 0 _048_
rlabel metal3 28992 17640 28992 17640 0 _049_
rlabel metal2 54720 12684 54720 12684 0 _050_
rlabel metal3 56832 15792 56832 15792 0 _051_
rlabel metal3 48816 15624 48816 15624 0 _052_
rlabel metal2 52032 18858 52032 18858 0 _053_
rlabel metal2 40704 4662 40704 4662 0 _054_
rlabel metal2 44064 3276 44064 3276 0 _055_
rlabel metal3 49824 5040 49824 5040 0 _056_
rlabel metal2 53472 3150 53472 3150 0 _057_
rlabel metal3 7680 27720 7680 27720 0 _058_
rlabel metal2 5664 30198 5664 30198 0 _059_
rlabel metal2 25728 34356 25728 34356 0 _060_
rlabel metal3 22272 36792 22272 36792 0 _061_
rlabel metal3 40518 30660 40518 30660 0 _062_
rlabel metal3 46320 29736 46320 29736 0 _063_
rlabel metal2 6336 23478 6336 23478 0 _064_
rlabel metal3 6672 23184 6672 23184 0 _065_
rlabel metal2 10752 33474 10752 33474 0 _066_
rlabel metal2 9792 33474 9792 33474 0 _067_
rlabel metal3 13488 2604 13488 2604 0 _068_
rlabel metal3 17664 2604 17664 2604 0 _069_
rlabel metal2 42624 22134 42624 22134 0 _070_
rlabel metal2 38208 26502 38208 26502 0 _071_
rlabel metal2 32160 22554 32160 22554 0 _072_
rlabel metal2 30624 22554 30624 22554 0 _073_
rlabel metal2 27648 12810 27648 12810 0 _074_
rlabel metal3 31392 10164 31392 10164 0 _075_
rlabel metal3 25536 17976 25536 17976 0 _076_
rlabel metal3 25440 20160 25440 20160 0 _077_
rlabel metal2 52800 10458 52800 10458 0 _078_
rlabel metal3 56592 14112 56592 14112 0 _079_
rlabel metal3 47184 17976 47184 17976 0 _080_
rlabel metal3 48000 21756 48000 21756 0 _081_
rlabel metal2 33408 3738 33408 3738 0 _082_
rlabel metal3 37488 2604 37488 2604 0 _083_
rlabel metal2 52608 5502 52608 5502 0 _084_
rlabel metal2 54480 2856 54480 2856 0 _085_
rlabel metal2 11808 4284 11808 4284 0 _086_
rlabel metal3 7776 2100 7776 2100 0 _087_
rlabel metal3 37296 24360 37296 24360 0 _088_
rlabel metal2 45984 23394 45984 23394 0 _089_
rlabel metal2 30336 21756 30336 21756 0 _090_
rlabel metal3 31392 25536 31392 25536 0 _091_
rlabel metal2 31584 11970 31584 11970 0 _092_
rlabel metal2 23904 13524 23904 13524 0 _093_
rlabel metal2 21792 17430 21792 17430 0 _094_
rlabel metal3 23280 17136 23280 17136 0 _095_
rlabel metal2 56256 12894 56256 12894 0 _096_
rlabel metal2 54912 9954 54912 9954 0 _097_
rlabel metal2 47232 18564 47232 18564 0 _098_
rlabel metal2 48912 21756 48912 21756 0 _099_
rlabel metal2 39504 2604 39504 2604 0 _100_
rlabel metal2 37728 5922 37728 5922 0 _101_
rlabel metal2 50496 2898 50496 2898 0 _102_
rlabel metal2 54816 4872 54816 4872 0 _103_
rlabel metal2 11136 4032 11136 4032 0 _104_
rlabel metal2 7872 2268 7872 2268 0 _105_
rlabel metal3 3072 21672 3072 21672 0 _106_
rlabel metal2 2400 25578 2400 25578 0 _107_
rlabel metal2 10896 16380 10896 16380 0 _108_
rlabel metal2 5280 17430 5280 17430 0 _109_
rlabel metal3 6768 34608 6768 34608 0 _110_
rlabel metal2 10848 36876 10848 36876 0 _111_
rlabel metal2 4320 27048 4320 27048 0 _112_
rlabel metal2 2208 31878 2208 31878 0 _113_
rlabel metal2 17952 30156 17952 30156 0 _114_
rlabel metal2 16896 35406 16896 35406 0 _115_
rlabel metal2 25152 37002 25152 37002 0 _116_
rlabel metal3 17376 36792 17376 36792 0 _117_
rlabel metal2 47040 31248 47040 31248 0 _118_
rlabel metal2 47040 27090 47040 27090 0 _119_
rlabel metal2 37296 36120 37296 36120 0 _120_
rlabel metal2 33216 36204 33216 36204 0 _121_
rlabel metal2 2736 8064 2736 8064 0 _122_
rlabel metal2 2160 12684 2160 12684 0 _123_
rlabel metal2 2688 23394 2688 23394 0 _124_
rlabel metal2 1728 18858 1728 18858 0 _125_
rlabel metal2 10752 17178 10752 17178 0 _126_
rlabel metal2 5664 17724 5664 17724 0 _127_
rlabel metal2 10896 36120 10896 36120 0 _128_
rlabel metal2 5952 35574 5952 35574 0 _129_
rlabel metal2 3120 30828 3120 30828 0 _130_
rlabel metal3 2784 27468 2784 27468 0 _131_
rlabel metal2 17472 31626 17472 31626 0 _132_
rlabel metal2 15552 33138 15552 33138 0 _133_
rlabel metal2 23616 25578 23616 25578 0 _134_
rlabel metal2 27840 35742 27840 35742 0 _135_
rlabel metal3 44256 27720 44256 27720 0 _136_
rlabel metal2 49152 30786 49152 30786 0 _137_
rlabel metal3 33696 34608 33696 34608 0 _138_
rlabel metal2 39696 36792 39696 36792 0 _139_
rlabel metal2 3072 11928 3072 11928 0 _140_
rlabel metal2 2304 8358 2304 8358 0 _141_
rlabel metal2 29376 7224 29376 7224 0 _142_
rlabel metal2 30864 7392 30864 7392 0 _143_
rlabel metal2 29760 8400 29760 8400 0 _144_
rlabel metal3 29712 6972 29712 6972 0 _145_
rlabel metal2 40896 8946 40896 8946 0 _146_
rlabel metal2 40800 8988 40800 8988 0 _147_
rlabel metal2 18240 24444 18240 24444 0 _148_
rlabel metal2 17280 25242 17280 25242 0 _149_
rlabel metal2 22752 22386 22752 22386 0 _150_
rlabel metal3 22656 25116 22656 25116 0 _151_
rlabel metal2 21600 8610 21600 8610 0 _152_
rlabel metal3 22656 7980 22656 7980 0 _153_
rlabel metal2 23040 8232 23040 8232 0 _154_
rlabel metal2 21888 8400 21888 8400 0 _155_
rlabel metal2 25728 9156 25728 9156 0 _156_
rlabel metal2 25824 9387 25824 9387 0 _157_
rlabel metal2 26016 9450 26016 9450 0 _158_
rlabel metal2 25824 8694 25824 8694 0 _159_
rlabel metal2 40608 20118 40608 20118 0 _160_
rlabel metal2 40704 22008 40704 22008 0 _161_
rlabel metal2 35808 15918 35808 15918 0 _162_
rlabel metal2 36192 16674 36192 16674 0 _163_
rlabel metal2 52896 14658 52896 14658 0 _164_
rlabel metal2 54912 17220 54912 17220 0 _165_
rlabel metal3 46896 5628 46896 5628 0 _166_
rlabel metal2 47616 4620 47616 4620 0 _167_
rlabel metal3 41232 14700 41232 14700 0 _168_
rlabel metal2 41520 16968 41520 16968 0 _169_
rlabel metal2 48480 10206 48480 10206 0 _170_
rlabel metal2 49824 10122 49824 10122 0 _171_
rlabel metal3 17904 12516 17904 12516 0 _172_
rlabel metal3 19872 13188 19872 13188 0 _173_
rlabel metal2 19968 12558 19968 12558 0 _174_
rlabel metal2 18624 12768 18624 12768 0 _175_
rlabel metal2 13056 28770 13056 28770 0 _176_
rlabel metal2 11616 29400 11616 29400 0 _177_
rlabel metal2 26304 31878 26304 31878 0 _178_
rlabel metal3 25440 32172 25440 32172 0 _179_
rlabel metal2 38016 30450 38016 30450 0 _180_
rlabel metal3 42816 32214 42816 32214 0 _181_
rlabel metal2 28800 28602 28800 28602 0 _182_
rlabel metal3 30000 30744 30000 30744 0 _183_
rlabel metal2 14016 22806 14016 22806 0 _184_
rlabel metal2 11616 22302 11616 22302 0 _185_
rlabel metal2 9312 34860 9312 34860 0 _186_
rlabel metal2 9696 35070 9696 35070 0 _187_
rlabel metal3 11376 2604 11376 2604 0 _188_
rlabel metal2 12000 2730 12000 2730 0 _189_
rlabel metal3 38160 35196 38160 35196 0 _190_
rlabel metal2 39456 35322 39456 35322 0 _191_
rlabel metal2 18720 33768 18720 33768 0 _192_
rlabel metal3 18576 32928 18576 32928 0 _193_
rlabel metal3 4608 11676 4608 11676 0 _194_
rlabel metal3 4368 9576 4368 9576 0 _195_
rlabel metal2 8352 17346 8352 17346 0 _196_
rlabel metal2 8928 18102 8928 18102 0 _197_
rlabel metal2 41280 25326 41280 25326 0 _198_
rlabel metal3 42288 23856 42288 23856 0 _199_
rlabel metal3 32016 24612 32016 24612 0 _200_
rlabel metal2 31968 24738 31968 24738 0 _201_
rlabel metal2 31296 12558 31296 12558 0 _202_
rlabel metal3 29760 13188 29760 13188 0 _203_
rlabel metal2 27552 17850 27552 17850 0 _204_
rlabel metal3 27216 17724 27216 17724 0 _205_
rlabel metal3 56112 12600 56112 12600 0 _206_
rlabel metal2 55872 12558 55872 12558 0 _207_
rlabel metal3 49824 19236 49824 19236 0 _208_
rlabel metal2 50496 19698 50496 19698 0 _209_
rlabel metal3 40704 3528 40704 3528 0 _210_
rlabel metal3 40752 4116 40752 4116 0 _211_
rlabel metal2 53184 3486 53184 3486 0 _212_
rlabel metal2 53568 3360 53568 3360 0 _213_
rlabel metal2 5184 30114 5184 30114 0 _214_
rlabel metal2 5184 29274 5184 29274 0 _215_
rlabel metal2 21936 36120 21936 36120 0 _216_
rlabel metal2 22560 37002 22560 37002 0 _217_
rlabel metal2 46944 29526 46944 29526 0 _218_
rlabel metal2 47808 30114 47808 30114 0 _219_
rlabel metal3 4752 23100 4752 23100 0 _220_
rlabel metal2 4224 22596 4224 22596 0 _221_
rlabel via2 78 36708 78 36708 0 clk
rlabel metal2 33744 23100 33744 23100 0 clknet_0_clk
rlabel metal2 4224 10710 4224 10710 0 clknet_4_0_0_clk
rlabel metal3 52608 6468 52608 6468 0 clknet_4_10_0_clk
rlabel metal2 52320 11802 52320 11802 0 clknet_4_11_0_clk
rlabel metal2 34944 19698 34944 19698 0 clknet_4_12_0_clk
rlabel metal2 34368 28098 34368 28098 0 clknet_4_13_0_clk
rlabel metal2 46368 25536 46368 25536 0 clknet_4_14_0_clk
rlabel metal2 42480 27636 42480 27636 0 clknet_4_15_0_clk
rlabel metal3 8736 18564 8736 18564 0 clknet_4_1_0_clk
rlabel metal2 18144 5922 18144 5922 0 clknet_4_2_0_clk
rlabel metal2 19344 8652 19344 8652 0 clknet_4_3_0_clk
rlabel metal3 10464 28980 10464 28980 0 clknet_4_4_0_clk
rlabel metal3 11136 33600 11136 33600 0 clknet_4_5_0_clk
rlabel metal2 22176 27972 22176 27972 0 clknet_4_6_0_clk
rlabel metal2 21504 34776 21504 34776 0 clknet_4_7_0_clk
rlabel metal3 35232 5628 35232 5628 0 clknet_4_8_0_clk
rlabel metal2 36192 11214 36192 11214 0 clknet_4_9_0_clk
rlabel metal3 3600 12516 3600 12516 0 clknet_5_0__leaf_clk
rlabel metal2 3840 31752 3840 31752 0 clknet_5_10__leaf_clk
rlabel metal2 15648 33432 15648 33432 0 clknet_5_11__leaf_clk
rlabel metal3 19200 22260 19200 22260 0 clknet_5_12__leaf_clk
rlabel metal2 22080 27678 22080 27678 0 clknet_5_13__leaf_clk
rlabel metal2 22176 34440 22176 34440 0 clknet_5_14__leaf_clk
rlabel metal3 28176 33684 28176 33684 0 clknet_5_15__leaf_clk
rlabel metal2 33408 5250 33408 5250 0 clknet_5_16__leaf_clk
rlabel metal2 40608 3192 40608 3192 0 clknet_5_17__leaf_clk
rlabel metal2 35040 13314 35040 13314 0 clknet_5_18__leaf_clk
rlabel metal2 39936 13944 39936 13944 0 clknet_5_19__leaf_clk
rlabel metal2 8544 3024 8544 3024 0 clknet_5_1__leaf_clk
rlabel metal2 48288 3192 48288 3192 0 clknet_5_20__leaf_clk
rlabel metal3 53712 3444 53712 3444 0 clknet_5_21__leaf_clk
rlabel metal2 52992 13314 52992 13314 0 clknet_5_22__leaf_clk
rlabel metal3 55632 13020 55632 13020 0 clknet_5_23__leaf_clk
rlabel metal2 26400 18102 26400 18102 0 clknet_5_24__leaf_clk
rlabel metal2 37344 19572 37344 19572 0 clknet_5_25__leaf_clk
rlabel metal2 33216 27636 33216 27636 0 clknet_5_26__leaf_clk
rlabel metal2 34464 35532 34464 35532 0 clknet_5_27__leaf_clk
rlabel metal3 46944 23100 46944 23100 0 clknet_5_28__leaf_clk
rlabel metal3 47808 19236 47808 19236 0 clknet_5_29__leaf_clk
rlabel metal3 3456 18564 3456 18564 0 clknet_5_2__leaf_clk
rlabel metal3 39696 36708 39696 36708 0 clknet_5_30__leaf_clk
rlabel metal3 43104 30660 43104 30660 0 clknet_5_31__leaf_clk
rlabel metal2 12192 17682 12192 17682 0 clknet_5_3__leaf_clk
rlabel metal3 18096 3444 18096 3444 0 clknet_5_4__leaf_clk
rlabel metal2 26064 3444 26064 3444 0 clknet_5_5__leaf_clk
rlabel metal2 17184 9156 17184 9156 0 clknet_5_6__leaf_clk
rlabel metal3 17472 17052 17472 17052 0 clknet_5_7__leaf_clk
rlabel metal2 3936 23520 3936 23520 0 clknet_5_8__leaf_clk
rlabel metal2 15648 24486 15648 24486 0 clknet_5_9__leaf_clk
rlabel metal2 40512 21084 40512 21084 0 mac1.products_ff\[0\]
rlabel metal3 44496 5628 44496 5628 0 mac1.products_ff\[102\]
rlabel metal3 47280 2856 47280 2856 0 mac1.products_ff\[103\]
rlabel metal2 45312 4956 45312 4956 0 mac1.products_ff\[119\]
rlabel metal2 47136 3150 47136 3150 0 mac1.products_ff\[120\]
rlabel metal2 17088 2184 17088 2184 0 mac1.products_ff\[136\]
rlabel metal2 20064 3864 20064 3864 0 mac1.products_ff\[137\]
rlabel metal3 38928 19824 38928 19824 0 mac1.products_ff\[17\]
rlabel metal2 40320 25578 40320 25578 0 mac1.products_ff\[18\]
rlabel metal2 40704 25578 40704 25578 0 mac1.products_ff\[1\]
rlabel metal3 36384 15288 36384 15288 0 mac1.products_ff\[34\]
rlabel metal2 33024 16380 33024 16380 0 mac1.products_ff\[35\]
rlabel metal2 34944 16506 34944 16506 0 mac1.products_ff\[51\]
rlabel metal2 33888 17388 33888 17388 0 mac1.products_ff\[52\]
rlabel metal2 51840 13734 51840 13734 0 mac1.products_ff\[68\]
rlabel metal2 54912 17010 54912 17010 0 mac1.products_ff\[69\]
rlabel metal2 52800 15498 52800 15498 0 mac1.products_ff\[85\]
rlabel metal2 54480 17052 54480 17052 0 mac1.products_ff\[86\]
rlabel metal2 41568 16170 41568 16170 0 mac1.sum_lvl1_ff\[0\]
rlabel metal2 46848 12348 46848 12348 0 mac1.sum_lvl1_ff\[16\]
rlabel metal2 49920 10668 49920 10668 0 mac1.sum_lvl1_ff\[17\]
rlabel metal3 42672 17724 42672 17724 0 mac1.sum_lvl1_ff\[1\]
rlabel metal3 48144 9492 48144 9492 0 mac1.sum_lvl1_ff\[24\]
rlabel metal2 50784 8778 50784 8778 0 mac1.sum_lvl1_ff\[25\]
rlabel metal2 21120 3150 21120 3150 0 mac1.sum_lvl1_ff\[32\]
rlabel metal2 24384 4158 24384 4158 0 mac1.sum_lvl1_ff\[33\]
rlabel metal2 39648 13734 39648 13734 0 mac1.sum_lvl1_ff\[8\]
rlabel metal2 39648 17472 39648 17472 0 mac1.sum_lvl1_ff\[9\]
rlabel metal3 40128 11004 40128 11004 0 mac1.sum_lvl2_ff\[0\]
rlabel metal2 44112 11004 44112 11004 0 mac1.sum_lvl2_ff\[1\]
rlabel metal2 39552 8946 39552 8946 0 mac1.sum_lvl2_ff\[4\]
rlabel metal2 44064 10416 44064 10416 0 mac1.sum_lvl2_ff\[5\]
rlabel metal2 24576 4284 24576 4284 0 mac1.sum_lvl2_ff\[8\]
rlabel metal2 27120 3612 27120 3612 0 mac1.sum_lvl2_ff\[9\]
rlabel metal3 33132 6972 33132 6972 0 mac1.sum_lvl3_ff\[0\]
rlabel metal2 33216 7980 33216 7980 0 mac1.sum_lvl3_ff\[1\]
rlabel metal2 28896 5670 28896 5670 0 mac1.sum_lvl3_ff\[2\]
rlabel metal2 30288 4368 30288 4368 0 mac1.sum_lvl3_ff\[3\]
rlabel metal2 19200 7938 19200 7938 0 mac1.total_sum\[0\]
rlabel metal3 20640 8652 20640 8652 0 mac1.total_sum\[1\]
rlabel metal2 26496 9240 26496 9240 0 mac1.total_sum\[2\]
rlabel metal2 12864 23352 12864 23352 0 mac2.products_ff\[0\]
rlabel metal2 37104 30828 37104 30828 0 mac2.products_ff\[102\]
rlabel metal2 42336 31164 42336 31164 0 mac2.products_ff\[103\]
rlabel metal2 37872 31332 37872 31332 0 mac2.products_ff\[119\]
rlabel metal3 43056 33432 43056 33432 0 mac2.products_ff\[120\]
rlabel metal3 7632 8820 7632 8820 0 mac2.products_ff\[136\]
rlabel metal2 8640 12516 8640 12516 0 mac2.products_ff\[137\]
rlabel metal2 15456 20790 15456 20790 0 mac2.products_ff\[17\]
rlabel metal2 11136 20076 11136 20076 0 mac2.products_ff\[18\]
rlabel metal2 11136 22554 11136 22554 0 mac2.products_ff\[1\]
rlabel metal2 13488 30660 13488 30660 0 mac2.products_ff\[34\]
rlabel metal2 11520 30492 11520 30492 0 mac2.products_ff\[35\]
rlabel metal2 12096 27930 12096 27930 0 mac2.products_ff\[51\]
rlabel metal2 11136 30114 11136 30114 0 mac2.products_ff\[52\]
rlabel metal2 25344 30996 25344 30996 0 mac2.products_ff\[68\]
rlabel metal2 24144 34440 24144 34440 0 mac2.products_ff\[69\]
rlabel metal3 27696 32844 27696 32844 0 mac2.products_ff\[85\]
rlabel metal2 24480 35406 24480 35406 0 mac2.products_ff\[86\]
rlabel metal2 18624 23436 18624 23436 0 mac2.sum_lvl1_ff\[0\]
rlabel metal2 28128 28980 28128 28980 0 mac2.sum_lvl1_ff\[16\]
rlabel metal2 30576 30660 30576 30660 0 mac2.sum_lvl1_ff\[17\]
rlabel metal2 16800 24612 16800 24612 0 mac2.sum_lvl1_ff\[1\]
rlabel metal2 31104 29106 31104 29106 0 mac2.sum_lvl1_ff\[24\]
rlabel metal3 31680 30660 31680 30660 0 mac2.sum_lvl1_ff\[25\]
rlabel metal3 10224 8820 10224 8820 0 mac2.sum_lvl1_ff\[32\]
rlabel metal2 11904 13230 11904 13230 0 mac2.sum_lvl1_ff\[33\]
rlabel metal2 18240 25284 18240 25284 0 mac2.sum_lvl1_ff\[8\]
rlabel metal2 17088 25956 17088 25956 0 mac2.sum_lvl1_ff\[9\]
rlabel metal2 22272 22512 22272 22512 0 mac2.sum_lvl2_ff\[0\]
rlabel metal3 22560 25284 22560 25284 0 mac2.sum_lvl2_ff\[1\]
rlabel metal2 21888 26334 21888 26334 0 mac2.sum_lvl2_ff\[4\]
rlabel metal2 27840 25956 27840 25956 0 mac2.sum_lvl2_ff\[5\]
rlabel metal3 12672 8820 12672 8820 0 mac2.sum_lvl2_ff\[8\]
rlabel metal2 14688 13734 14688 13734 0 mac2.sum_lvl2_ff\[9\]
rlabel metal2 16512 15750 16512 15750 0 mac2.sum_lvl3_ff\[0\]
rlabel metal2 18768 14028 18768 14028 0 mac2.sum_lvl3_ff\[1\]
rlabel metal2 15936 10584 15936 10584 0 mac2.sum_lvl3_ff\[2\]
rlabel metal2 19008 13986 19008 13986 0 mac2.sum_lvl3_ff\[3\]
rlabel metal2 18816 8610 18816 8610 0 mac2.total_sum\[0\]
rlabel metal2 21120 9324 21120 9324 0 mac2.total_sum\[1\]
rlabel metal3 25968 9492 25968 9492 0 mac2.total_sum\[2\]
rlabel metal3 16512 2730 16512 2730 0 net1
rlabel metal3 366 13188 366 13188 0 net10
rlabel metal2 45552 8148 45552 8148 0 net100
rlabel metal2 3648 19824 3648 19824 0 net101
rlabel metal3 20304 37212 20304 37212 0 net102
rlabel metal3 26736 31332 26736 31332 0 net103
rlabel metal2 25728 30114 25728 30114 0 net104
rlabel metal2 49488 21420 49488 21420 0 net105
rlabel metal3 10128 2100 10128 2100 0 net106
rlabel metal2 19008 23520 19008 23520 0 net107
rlabel metal2 19776 22554 19776 22554 0 net108
rlabel metal2 14112 29022 14112 29022 0 net109
rlabel metal3 366 14028 366 14028 0 net11
rlabel metal2 15312 26796 15312 26796 0 net110
rlabel metal2 35712 15792 35712 15792 0 net111
rlabel metal2 37248 13482 37248 13482 0 net112
rlabel metal2 52704 14238 52704 14238 0 net113
rlabel metal2 48384 13482 48384 13482 0 net114
rlabel metal2 17184 13104 17184 13104 0 net115
rlabel metal2 15888 9576 15888 9576 0 net116
rlabel metal2 27171 17766 27171 17766 0 net117
rlabel metal2 12480 3612 12480 3612 0 net118
rlabel metal3 5328 23604 5328 23604 0 net119
rlabel metal3 366 14868 366 14868 0 net12
rlabel metal3 40704 3444 40704 3444 0 net120
rlabel metal2 36480 34692 36480 34692 0 net121
rlabel metal2 56448 12558 56448 12558 0 net122
rlabel metal2 37872 29820 37872 29820 0 net123
rlabel metal2 34512 29232 34512 29232 0 net124
rlabel metal3 26256 37464 26256 37464 0 net125
rlabel via2 53088 4956 53088 4956 0 net126
rlabel metal3 4848 9660 4848 9660 0 net127
rlabel metal2 31296 21924 31296 21924 0 net128
rlabel metal3 31728 12432 31728 12432 0 net129
rlabel metal3 366 5628 366 5628 0 net13
rlabel metal2 10464 35112 10464 35112 0 net130
rlabel metal2 18624 33432 18624 33432 0 net131
rlabel metal3 5280 22512 5280 22512 0 net132
rlabel metal2 12672 3486 12672 3486 0 net133
rlabel metal3 30912 13020 30912 13020 0 net134
rlabel metal2 52272 3612 52272 3612 0 net135
rlabel metal2 28512 29190 28512 29190 0 net136
rlabel metal2 23328 27552 23328 27552 0 net137
rlabel metal3 49104 17976 49104 17976 0 net138
rlabel metal3 54912 11172 54912 11172 0 net139
rlabel metal3 366 6468 366 6468 0 net14
rlabel metal3 4848 11508 4848 11508 0 net140
rlabel metal2 37632 35658 37632 35658 0 net141
rlabel metal3 39120 24780 39120 24780 0 net142
rlabel metal3 45312 28392 45312 28392 0 net143
rlabel metal2 46704 31416 46704 31416 0 net144
rlabel metal2 40896 15204 40896 15204 0 net145
rlabel metal2 40800 10836 40800 10836 0 net146
rlabel metal2 33888 22176 33888 22176 0 net147
rlabel metal3 9312 34188 9312 34188 0 net148
rlabel metal3 5472 27048 5472 27048 0 net149
rlabel metal3 366 7308 366 7308 0 net15
rlabel metal3 48768 20076 48768 20076 0 net150
rlabel metal3 36720 4200 36720 4200 0 net151
rlabel metal2 11712 16422 11712 16422 0 net152
rlabel metal2 40224 9156 40224 9156 0 net153
rlabel metal3 36960 7056 36960 7056 0 net154
rlabel metal2 4464 30492 4464 30492 0 net155
rlabel metal2 18144 31080 18144 31080 0 net156
rlabel metal3 12048 18732 12048 18732 0 net157
rlabel metal2 25728 35532 25728 35532 0 net158
rlabel metal3 40326 23268 40326 23268 0 net159
rlabel metal3 318 8148 318 8148 0 net16
rlabel metal3 22416 18312 22416 18312 0 net160
rlabel metal2 46944 10836 46944 10836 0 net161
rlabel metal2 41184 10164 41184 10164 0 net162
rlabel metal2 22848 22218 22848 22218 0 net163
rlabel metal2 18912 17388 18912 17388 0 net164
rlabel metal2 29664 6552 29664 6552 0 net165
rlabel metal3 19584 7140 19584 7140 0 net166
rlabel metal2 30960 7140 30960 7140 0 net167
rlabel metal3 30000 7980 30000 7980 0 net168
rlabel metal3 28032 8064 28032 8064 0 net169
rlabel metal3 318 15708 318 15708 0 net17
rlabel metal3 19152 14028 19152 14028 0 net170
rlabel metal2 20064 12768 20064 12768 0 net171
rlabel metal3 22512 12264 22512 12264 0 net172
rlabel metal2 47904 9912 47904 9912 0 net173
rlabel metal3 46944 10080 46944 10080 0 net174
rlabel metal2 40992 14448 40992 14448 0 net175
rlabel metal2 41472 13482 41472 13482 0 net176
rlabel metal2 39936 20412 39936 20412 0 net177
rlabel metal2 41088 19236 41088 19236 0 net178
rlabel metal2 12864 28308 12864 28308 0 net179
rlabel metal3 366 16548 366 16548 0 net18
rlabel metal2 12816 26796 12816 26796 0 net180
rlabel metal3 26112 31332 26112 31332 0 net181
rlabel metal2 28128 32466 28128 32466 0 net182
rlabel metal2 36000 15540 36000 15540 0 net183
rlabel metal2 37152 17052 37152 17052 0 net184
rlabel metal2 18720 24402 18720 24402 0 net185
rlabel metal2 19776 26124 19776 26124 0 net186
rlabel metal3 51792 15288 51792 15288 0 net187
rlabel metal3 51024 14532 51024 14532 0 net188
rlabel metal3 28896 29148 28896 29148 0 net189
rlabel metal3 366 17388 366 17388 0 net19
rlabel metal2 30240 27090 30240 27090 0 net190
rlabel metal2 13920 22554 13920 22554 0 net191
rlabel metal2 14304 23688 14304 23688 0 net192
rlabel metal2 46656 5586 46656 5586 0 net193
rlabel metal2 48672 6846 48672 6846 0 net194
rlabel metal3 38400 29820 38400 29820 0 net195
rlabel metal3 35520 31248 35520 31248 0 net196
rlabel metal2 41376 9576 41376 9576 0 net197
rlabel metal2 36000 8232 36000 8232 0 net198
rlabel metal2 22656 22764 22656 22764 0 net199
rlabel metal2 864 3444 864 3444 0 net2
rlabel metal3 366 18228 366 18228 0 net20
rlabel metal2 19776 18690 19776 18690 0 net200
rlabel metal2 16608 11214 16608 11214 0 net201
rlabel metal2 19008 11214 19008 11214 0 net202
rlabel metal3 30768 6468 30768 6468 0 net203
rlabel metal3 24384 7056 24384 7056 0 net204
rlabel metal3 366 19068 366 19068 0 net21
rlabel metal3 366 19908 366 19908 0 net22
rlabel metal3 366 20748 366 20748 0 net23
rlabel metal3 366 21588 366 21588 0 net24
rlabel metal2 7392 8946 7392 8946 0 net25
rlabel metal2 9984 8946 9984 8946 0 net26
rlabel metal2 17760 2310 17760 2310 0 net27
rlabel metal2 12288 13524 12288 13524 0 net28
rlabel metal2 9504 12810 9504 12810 0 net29
rlabel metal2 912 4200 912 4200 0 net3
rlabel metal2 27936 3990 27936 3990 0 net30
rlabel metal2 24768 3738 24768 3738 0 net31
rlabel metal2 11904 9786 11904 9786 0 net32
rlabel metal2 21312 4032 21312 4032 0 net33
rlabel metal2 15936 14028 15936 14028 0 net34
rlabel metal2 21984 3444 21984 3444 0 net35
rlabel metal2 26400 4956 26400 4956 0 net36
rlabel metal3 49536 30576 49536 30576 0 net37
rlabel metal2 43008 23520 43008 23520 0 net38
rlabel metal3 28224 35952 28224 35952 0 net39
rlabel metal2 864 7014 864 7014 0 net4
rlabel metal2 54432 5166 54432 5166 0 net40
rlabel metal2 3936 11718 3936 11718 0 net41
rlabel metal2 7680 18228 7680 18228 0 net42
rlabel metal3 2832 9492 2832 9492 0 net43
rlabel metal3 56208 10248 56208 10248 0 net44
rlabel metal2 7296 35826 7296 35826 0 net45
rlabel metal2 39744 25956 39744 25956 0 net46
rlabel metal3 26496 20832 26496 20832 0 net47
rlabel metal2 32064 25998 32064 25998 0 net48
rlabel metal3 3888 28980 3888 28980 0 net49
rlabel metal3 366 8988 366 8988 0 net5
rlabel metal3 3216 31416 3216 31416 0 net50
rlabel metal2 39840 36666 39840 36666 0 net51
rlabel metal2 16416 33138 16416 33138 0 net52
rlabel metal3 25584 17892 25584 17892 0 net53
rlabel metal3 38976 3360 38976 3360 0 net54
rlabel metal2 32832 11256 32832 11256 0 net55
rlabel metal3 11328 36624 11328 36624 0 net56
rlabel metal2 7392 17304 7392 17304 0 net57
rlabel metal3 17760 35112 17760 35112 0 net58
rlabel metal3 49776 21504 49776 21504 0 net59
rlabel metal3 366 9828 366 9828 0 net6
rlabel metal2 15648 5208 15648 5208 0 net60
rlabel metal2 15168 4200 15168 4200 0 net61
rlabel metal2 2976 12432 2976 12432 0 net62
rlabel metal3 12912 13188 12912 13188 0 net63
rlabel metal2 23328 13230 23328 13230 0 net64
rlabel metal2 18528 17262 18528 17262 0 net65
rlabel metal3 22272 17052 22272 17052 0 net66
rlabel metal2 3072 23058 3072 23058 0 net67
rlabel metal2 2304 31752 2304 31752 0 net68
rlabel metal2 13440 20118 13440 20118 0 net69
rlabel metal3 366 10668 366 10668 0 net7
rlabel metal2 17184 36624 17184 36624 0 net70
rlabel metal2 16512 23016 16512 23016 0 net71
rlabel metal2 22944 21504 22944 21504 0 net72
rlabel metal2 37152 2646 37152 2646 0 net73
rlabel metal2 37632 17976 37632 17976 0 net74
rlabel metal2 51840 8190 51840 8190 0 net75
rlabel metal2 55200 4788 55200 4788 0 net76
rlabel metal2 52368 18480 52368 18480 0 net77
rlabel metal2 53856 13230 53856 13230 0 net78
rlabel via2 37536 23772 37536 23772 0 net79
rlabel metal3 366 11508 366 11508 0 net8
rlabel metal3 21840 34020 21840 34020 0 net80
rlabel metal2 34944 26166 34944 26166 0 net81
rlabel metal3 33936 35196 33936 35196 0 net82
rlabel metal2 48288 23058 48288 23058 0 net83
rlabel metal2 42816 29400 42816 29400 0 net84
rlabel metal2 34080 14742 34080 14742 0 net85
rlabel metal2 35136 36246 35136 36246 0 net86
rlabel metal2 57024 13650 57024 13650 0 net87
rlabel metal2 4176 25872 4176 25872 0 net88
rlabel metal2 47040 28350 47040 28350 0 net89
rlabel metal3 366 12348 366 12348 0 net9
rlabel metal3 39792 6972 39792 6972 0 net90
rlabel metal3 9504 2520 9504 2520 0 net91
rlabel metal3 55296 2688 55296 2688 0 net92
rlabel metal2 39744 20202 39744 20202 0 net93
rlabel metal2 40032 17724 40032 17724 0 net94
rlabel metal2 14880 22008 14880 22008 0 net95
rlabel metal2 16032 22176 16032 22176 0 net96
rlabel metal2 29664 23058 29664 23058 0 net97
rlabel metal3 27408 13860 27408 13860 0 net98
rlabel metal3 45744 6468 45744 6468 0 net99
rlabel metal3 174 37548 174 37548 0 rst_n
rlabel metal3 366 2268 366 2268 0 uo_out[0]
rlabel metal3 366 3108 366 3108 0 uo_out[1]
rlabel metal3 366 3948 366 3948 0 uo_out[2]
rlabel metal3 366 4788 366 4788 0 uo_out[3]
<< properties >>
string FIXED_BBOX 0 0 100000 40000
<< end >>
