module heichips25_template (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \DP_1.I_range.data_plus_4[6] ;
 wire \DP_1.I_range.out_data[2] ;
 wire \DP_1.I_range.out_data[3] ;
 wire \DP_1.I_range.out_data[4] ;
 wire \DP_1.I_range.out_data[5] ;
 wire \DP_1.Q_range.data_plus_4[6] ;
 wire \DP_1.Q_range.out_data[2] ;
 wire \DP_1.Q_range.out_data[3] ;
 wire \DP_1.Q_range.out_data[4] ;
 wire \DP_1.Q_range.out_data[5] ;
 wire \DP_1.matrix[0] ;
 wire \DP_1.matrix[1] ;
 wire \DP_1.matrix[2] ;
 wire \DP_1.matrix[36] ;
 wire \DP_1.matrix[37] ;
 wire \DP_1.matrix[38] ;
 wire \DP_1.matrix[39] ;
 wire \DP_1.matrix[3] ;
 wire \DP_1.matrix[40] ;
 wire \DP_1.matrix[41] ;
 wire \DP_1.matrix[42] ;
 wire \DP_1.matrix[43] ;
 wire \DP_1.matrix[44] ;
 wire \DP_1.matrix[4] ;
 wire \DP_1.matrix[5] ;
 wire \DP_1.matrix[6] ;
 wire \DP_1.matrix[72] ;
 wire \DP_1.matrix[73] ;
 wire \DP_1.matrix[74] ;
 wire \DP_1.matrix[75] ;
 wire \DP_1.matrix[76] ;
 wire \DP_1.matrix[77] ;
 wire \DP_1.matrix[78] ;
 wire \DP_1.matrix[79] ;
 wire \DP_1.matrix[7] ;
 wire \DP_1.matrix[80] ;
 wire \DP_1.matrix[8] ;
 wire \DP_2.matrix[0] ;
 wire \DP_2.matrix[1] ;
 wire \DP_2.matrix[2] ;
 wire \DP_2.matrix[36] ;
 wire \DP_2.matrix[37] ;
 wire \DP_2.matrix[38] ;
 wire \DP_2.matrix[39] ;
 wire \DP_2.matrix[3] ;
 wire \DP_2.matrix[40] ;
 wire \DP_2.matrix[41] ;
 wire \DP_2.matrix[42] ;
 wire \DP_2.matrix[43] ;
 wire \DP_2.matrix[44] ;
 wire \DP_2.matrix[4] ;
 wire \DP_2.matrix[5] ;
 wire \DP_2.matrix[6] ;
 wire \DP_2.matrix[72] ;
 wire \DP_2.matrix[73] ;
 wire \DP_2.matrix[74] ;
 wire \DP_2.matrix[75] ;
 wire \DP_2.matrix[76] ;
 wire \DP_2.matrix[77] ;
 wire \DP_2.matrix[78] ;
 wire \DP_2.matrix[79] ;
 wire \DP_2.matrix[7] ;
 wire \DP_2.matrix[80] ;
 wire \DP_2.matrix[8] ;
 wire \DP_3.I_range.data_plus_4[6] ;
 wire \DP_3.I_range.out_data[2] ;
 wire \DP_3.I_range.out_data[3] ;
 wire \DP_3.I_range.out_data[4] ;
 wire \DP_3.I_range.out_data[5] ;
 wire \DP_3.Q_range.data_plus_4[6] ;
 wire \DP_3.Q_range.out_data[2] ;
 wire \DP_3.Q_range.out_data[3] ;
 wire \DP_3.Q_range.out_data[4] ;
 wire \DP_3.Q_range.out_data[5] ;
 wire \DP_3.matrix[0] ;
 wire \DP_3.matrix[1] ;
 wire \DP_3.matrix[2] ;
 wire \DP_3.matrix[36] ;
 wire \DP_3.matrix[37] ;
 wire \DP_3.matrix[38] ;
 wire \DP_3.matrix[39] ;
 wire \DP_3.matrix[3] ;
 wire \DP_3.matrix[40] ;
 wire \DP_3.matrix[41] ;
 wire \DP_3.matrix[42] ;
 wire \DP_3.matrix[43] ;
 wire \DP_3.matrix[44] ;
 wire \DP_3.matrix[4] ;
 wire \DP_3.matrix[5] ;
 wire \DP_3.matrix[6] ;
 wire \DP_3.matrix[72] ;
 wire \DP_3.matrix[73] ;
 wire \DP_3.matrix[74] ;
 wire \DP_3.matrix[75] ;
 wire \DP_3.matrix[76] ;
 wire \DP_3.matrix[77] ;
 wire \DP_3.matrix[78] ;
 wire \DP_3.matrix[79] ;
 wire \DP_3.matrix[7] ;
 wire \DP_3.matrix[80] ;
 wire \DP_3.matrix[8] ;
 wire \DP_4.matrix[0] ;
 wire \DP_4.matrix[1] ;
 wire \DP_4.matrix[2] ;
 wire \DP_4.matrix[36] ;
 wire \DP_4.matrix[37] ;
 wire \DP_4.matrix[38] ;
 wire \DP_4.matrix[39] ;
 wire \DP_4.matrix[3] ;
 wire \DP_4.matrix[40] ;
 wire \DP_4.matrix[41] ;
 wire \DP_4.matrix[42] ;
 wire \DP_4.matrix[43] ;
 wire \DP_4.matrix[44] ;
 wire \DP_4.matrix[4] ;
 wire \DP_4.matrix[5] ;
 wire \DP_4.matrix[6] ;
 wire \DP_4.matrix[72] ;
 wire \DP_4.matrix[73] ;
 wire \DP_4.matrix[74] ;
 wire \DP_4.matrix[75] ;
 wire \DP_4.matrix[76] ;
 wire \DP_4.matrix[77] ;
 wire \DP_4.matrix[78] ;
 wire \DP_4.matrix[79] ;
 wire \DP_4.matrix[7] ;
 wire \DP_4.matrix[80] ;
 wire \DP_4.matrix[8] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire \mac1.products_ff[0] ;
 wire \mac1.products_ff[10] ;
 wire \mac1.products_ff[11] ;
 wire \mac1.products_ff[12] ;
 wire \mac1.products_ff[136] ;
 wire \mac1.products_ff[137] ;
 wire \mac1.products_ff[138] ;
 wire \mac1.products_ff[139] ;
 wire \mac1.products_ff[13] ;
 wire \mac1.products_ff[140] ;
 wire \mac1.products_ff[141] ;
 wire \mac1.products_ff[142] ;
 wire \mac1.products_ff[143] ;
 wire \mac1.products_ff[144] ;
 wire \mac1.products_ff[145] ;
 wire \mac1.products_ff[146] ;
 wire \mac1.products_ff[147] ;
 wire \mac1.products_ff[148] ;
 wire \mac1.products_ff[149] ;
 wire \mac1.products_ff[14] ;
 wire \mac1.products_ff[150] ;
 wire \mac1.products_ff[151] ;
 wire \mac1.products_ff[15] ;
 wire \mac1.products_ff[1] ;
 wire \mac1.products_ff[2] ;
 wire \mac1.products_ff[3] ;
 wire \mac1.products_ff[4] ;
 wire \mac1.products_ff[5] ;
 wire \mac1.products_ff[68] ;
 wire \mac1.products_ff[69] ;
 wire \mac1.products_ff[6] ;
 wire \mac1.products_ff[70] ;
 wire \mac1.products_ff[71] ;
 wire \mac1.products_ff[72] ;
 wire \mac1.products_ff[73] ;
 wire \mac1.products_ff[74] ;
 wire \mac1.products_ff[75] ;
 wire \mac1.products_ff[76] ;
 wire \mac1.products_ff[77] ;
 wire \mac1.products_ff[78] ;
 wire \mac1.products_ff[79] ;
 wire \mac1.products_ff[7] ;
 wire \mac1.products_ff[80] ;
 wire \mac1.products_ff[81] ;
 wire \mac1.products_ff[82] ;
 wire \mac1.products_ff[83] ;
 wire \mac1.products_ff[8] ;
 wire \mac1.products_ff[9] ;
 wire \mac1.sum_lvl1_ff[0] ;
 wire \mac1.sum_lvl1_ff[10] ;
 wire \mac1.sum_lvl1_ff[11] ;
 wire \mac1.sum_lvl1_ff[12] ;
 wire \mac1.sum_lvl1_ff[13] ;
 wire \mac1.sum_lvl1_ff[14] ;
 wire \mac1.sum_lvl1_ff[15] ;
 wire \mac1.sum_lvl1_ff[1] ;
 wire \mac1.sum_lvl1_ff[2] ;
 wire \mac1.sum_lvl1_ff[36] ;
 wire \mac1.sum_lvl1_ff[37] ;
 wire \mac1.sum_lvl1_ff[38] ;
 wire \mac1.sum_lvl1_ff[39] ;
 wire \mac1.sum_lvl1_ff[3] ;
 wire \mac1.sum_lvl1_ff[40] ;
 wire \mac1.sum_lvl1_ff[41] ;
 wire \mac1.sum_lvl1_ff[42] ;
 wire \mac1.sum_lvl1_ff[43] ;
 wire \mac1.sum_lvl1_ff[44] ;
 wire \mac1.sum_lvl1_ff[45] ;
 wire \mac1.sum_lvl1_ff[46] ;
 wire \mac1.sum_lvl1_ff[47] ;
 wire \mac1.sum_lvl1_ff[48] ;
 wire \mac1.sum_lvl1_ff[49] ;
 wire \mac1.sum_lvl1_ff[4] ;
 wire \mac1.sum_lvl1_ff[50] ;
 wire \mac1.sum_lvl1_ff[51] ;
 wire \mac1.sum_lvl1_ff[5] ;
 wire \mac1.sum_lvl1_ff[6] ;
 wire \mac1.sum_lvl1_ff[72] ;
 wire \mac1.sum_lvl1_ff[73] ;
 wire \mac1.sum_lvl1_ff[74] ;
 wire \mac1.sum_lvl1_ff[75] ;
 wire \mac1.sum_lvl1_ff[76] ;
 wire \mac1.sum_lvl1_ff[77] ;
 wire \mac1.sum_lvl1_ff[78] ;
 wire \mac1.sum_lvl1_ff[79] ;
 wire \mac1.sum_lvl1_ff[7] ;
 wire \mac1.sum_lvl1_ff[80] ;
 wire \mac1.sum_lvl1_ff[81] ;
 wire \mac1.sum_lvl1_ff[82] ;
 wire \mac1.sum_lvl1_ff[83] ;
 wire \mac1.sum_lvl1_ff[84] ;
 wire \mac1.sum_lvl1_ff[85] ;
 wire \mac1.sum_lvl1_ff[86] ;
 wire \mac1.sum_lvl1_ff[87] ;
 wire \mac1.sum_lvl1_ff[8] ;
 wire \mac1.sum_lvl1_ff[9] ;
 wire \mac1.sum_lvl2_ff[0] ;
 wire \mac1.sum_lvl2_ff[10] ;
 wire \mac1.sum_lvl2_ff[11] ;
 wire \mac1.sum_lvl2_ff[12] ;
 wire \mac1.sum_lvl2_ff[13] ;
 wire \mac1.sum_lvl2_ff[14] ;
 wire \mac1.sum_lvl2_ff[15] ;
 wire \mac1.sum_lvl2_ff[19] ;
 wire \mac1.sum_lvl2_ff[1] ;
 wire \mac1.sum_lvl2_ff[20] ;
 wire \mac1.sum_lvl2_ff[21] ;
 wire \mac1.sum_lvl2_ff[22] ;
 wire \mac1.sum_lvl2_ff[23] ;
 wire \mac1.sum_lvl2_ff[24] ;
 wire \mac1.sum_lvl2_ff[25] ;
 wire \mac1.sum_lvl2_ff[26] ;
 wire \mac1.sum_lvl2_ff[27] ;
 wire \mac1.sum_lvl2_ff[28] ;
 wire \mac1.sum_lvl2_ff[29] ;
 wire \mac1.sum_lvl2_ff[2] ;
 wire \mac1.sum_lvl2_ff[30] ;
 wire \mac1.sum_lvl2_ff[31] ;
 wire \mac1.sum_lvl2_ff[32] ;
 wire \mac1.sum_lvl2_ff[33] ;
 wire \mac1.sum_lvl2_ff[34] ;
 wire \mac1.sum_lvl2_ff[38] ;
 wire \mac1.sum_lvl2_ff[39] ;
 wire \mac1.sum_lvl2_ff[3] ;
 wire \mac1.sum_lvl2_ff[40] ;
 wire \mac1.sum_lvl2_ff[41] ;
 wire \mac1.sum_lvl2_ff[42] ;
 wire \mac1.sum_lvl2_ff[43] ;
 wire \mac1.sum_lvl2_ff[44] ;
 wire \mac1.sum_lvl2_ff[45] ;
 wire \mac1.sum_lvl2_ff[46] ;
 wire \mac1.sum_lvl2_ff[47] ;
 wire \mac1.sum_lvl2_ff[48] ;
 wire \mac1.sum_lvl2_ff[49] ;
 wire \mac1.sum_lvl2_ff[4] ;
 wire \mac1.sum_lvl2_ff[50] ;
 wire \mac1.sum_lvl2_ff[51] ;
 wire \mac1.sum_lvl2_ff[52] ;
 wire \mac1.sum_lvl2_ff[53] ;
 wire \mac1.sum_lvl2_ff[5] ;
 wire \mac1.sum_lvl2_ff[6] ;
 wire \mac1.sum_lvl2_ff[7] ;
 wire \mac1.sum_lvl2_ff[8] ;
 wire \mac1.sum_lvl2_ff[9] ;
 wire \mac1.sum_lvl3_ff[0] ;
 wire \mac1.sum_lvl3_ff[10] ;
 wire \mac1.sum_lvl3_ff[11] ;
 wire \mac1.sum_lvl3_ff[12] ;
 wire \mac1.sum_lvl3_ff[13] ;
 wire \mac1.sum_lvl3_ff[14] ;
 wire \mac1.sum_lvl3_ff[15] ;
 wire \mac1.sum_lvl3_ff[1] ;
 wire \mac1.sum_lvl3_ff[20] ;
 wire \mac1.sum_lvl3_ff[21] ;
 wire \mac1.sum_lvl3_ff[22] ;
 wire \mac1.sum_lvl3_ff[23] ;
 wire \mac1.sum_lvl3_ff[24] ;
 wire \mac1.sum_lvl3_ff[25] ;
 wire \mac1.sum_lvl3_ff[26] ;
 wire \mac1.sum_lvl3_ff[27] ;
 wire \mac1.sum_lvl3_ff[28] ;
 wire \mac1.sum_lvl3_ff[29] ;
 wire \mac1.sum_lvl3_ff[2] ;
 wire \mac1.sum_lvl3_ff[30] ;
 wire \mac1.sum_lvl3_ff[31] ;
 wire \mac1.sum_lvl3_ff[32] ;
 wire \mac1.sum_lvl3_ff[33] ;
 wire \mac1.sum_lvl3_ff[34] ;
 wire \mac1.sum_lvl3_ff[35] ;
 wire \mac1.sum_lvl3_ff[3] ;
 wire \mac1.sum_lvl3_ff[4] ;
 wire \mac1.sum_lvl3_ff[5] ;
 wire \mac1.sum_lvl3_ff[6] ;
 wire \mac1.sum_lvl3_ff[7] ;
 wire \mac1.sum_lvl3_ff[8] ;
 wire \mac1.sum_lvl3_ff[9] ;
 wire \mac1.total_sum[0] ;
 wire \mac1.total_sum[10] ;
 wire \mac1.total_sum[11] ;
 wire \mac1.total_sum[12] ;
 wire \mac1.total_sum[13] ;
 wire \mac1.total_sum[14] ;
 wire \mac1.total_sum[15] ;
 wire \mac1.total_sum[1] ;
 wire \mac1.total_sum[2] ;
 wire \mac1.total_sum[3] ;
 wire \mac1.total_sum[4] ;
 wire \mac1.total_sum[5] ;
 wire \mac1.total_sum[6] ;
 wire \mac1.total_sum[7] ;
 wire \mac1.total_sum[8] ;
 wire \mac1.total_sum[9] ;
 wire \mac2.products_ff[0] ;
 wire \mac2.products_ff[10] ;
 wire \mac2.products_ff[11] ;
 wire \mac2.products_ff[12] ;
 wire \mac2.products_ff[136] ;
 wire \mac2.products_ff[137] ;
 wire \mac2.products_ff[138] ;
 wire \mac2.products_ff[139] ;
 wire \mac2.products_ff[13] ;
 wire \mac2.products_ff[140] ;
 wire \mac2.products_ff[141] ;
 wire \mac2.products_ff[142] ;
 wire \mac2.products_ff[143] ;
 wire \mac2.products_ff[144] ;
 wire \mac2.products_ff[145] ;
 wire \mac2.products_ff[146] ;
 wire \mac2.products_ff[147] ;
 wire \mac2.products_ff[148] ;
 wire \mac2.products_ff[149] ;
 wire \mac2.products_ff[14] ;
 wire \mac2.products_ff[150] ;
 wire \mac2.products_ff[151] ;
 wire \mac2.products_ff[15] ;
 wire \mac2.products_ff[1] ;
 wire \mac2.products_ff[2] ;
 wire \mac2.products_ff[3] ;
 wire \mac2.products_ff[4] ;
 wire \mac2.products_ff[5] ;
 wire \mac2.products_ff[68] ;
 wire \mac2.products_ff[69] ;
 wire \mac2.products_ff[6] ;
 wire \mac2.products_ff[70] ;
 wire \mac2.products_ff[71] ;
 wire \mac2.products_ff[72] ;
 wire \mac2.products_ff[73] ;
 wire \mac2.products_ff[74] ;
 wire \mac2.products_ff[75] ;
 wire \mac2.products_ff[76] ;
 wire \mac2.products_ff[77] ;
 wire \mac2.products_ff[78] ;
 wire \mac2.products_ff[79] ;
 wire \mac2.products_ff[7] ;
 wire \mac2.products_ff[80] ;
 wire \mac2.products_ff[81] ;
 wire \mac2.products_ff[82] ;
 wire \mac2.products_ff[83] ;
 wire \mac2.products_ff[8] ;
 wire \mac2.products_ff[9] ;
 wire \mac2.sum_lvl1_ff[0] ;
 wire \mac2.sum_lvl1_ff[10] ;
 wire \mac2.sum_lvl1_ff[11] ;
 wire \mac2.sum_lvl1_ff[12] ;
 wire \mac2.sum_lvl1_ff[13] ;
 wire \mac2.sum_lvl1_ff[14] ;
 wire \mac2.sum_lvl1_ff[15] ;
 wire \mac2.sum_lvl1_ff[1] ;
 wire \mac2.sum_lvl1_ff[2] ;
 wire \mac2.sum_lvl1_ff[36] ;
 wire \mac2.sum_lvl1_ff[37] ;
 wire \mac2.sum_lvl1_ff[38] ;
 wire \mac2.sum_lvl1_ff[39] ;
 wire \mac2.sum_lvl1_ff[3] ;
 wire \mac2.sum_lvl1_ff[40] ;
 wire \mac2.sum_lvl1_ff[41] ;
 wire \mac2.sum_lvl1_ff[42] ;
 wire \mac2.sum_lvl1_ff[43] ;
 wire \mac2.sum_lvl1_ff[44] ;
 wire \mac2.sum_lvl1_ff[45] ;
 wire \mac2.sum_lvl1_ff[46] ;
 wire \mac2.sum_lvl1_ff[47] ;
 wire \mac2.sum_lvl1_ff[48] ;
 wire \mac2.sum_lvl1_ff[49] ;
 wire \mac2.sum_lvl1_ff[4] ;
 wire \mac2.sum_lvl1_ff[50] ;
 wire \mac2.sum_lvl1_ff[51] ;
 wire \mac2.sum_lvl1_ff[5] ;
 wire \mac2.sum_lvl1_ff[6] ;
 wire \mac2.sum_lvl1_ff[72] ;
 wire \mac2.sum_lvl1_ff[73] ;
 wire \mac2.sum_lvl1_ff[74] ;
 wire \mac2.sum_lvl1_ff[75] ;
 wire \mac2.sum_lvl1_ff[76] ;
 wire \mac2.sum_lvl1_ff[77] ;
 wire \mac2.sum_lvl1_ff[78] ;
 wire \mac2.sum_lvl1_ff[79] ;
 wire \mac2.sum_lvl1_ff[7] ;
 wire \mac2.sum_lvl1_ff[80] ;
 wire \mac2.sum_lvl1_ff[81] ;
 wire \mac2.sum_lvl1_ff[82] ;
 wire \mac2.sum_lvl1_ff[83] ;
 wire \mac2.sum_lvl1_ff[84] ;
 wire \mac2.sum_lvl1_ff[85] ;
 wire \mac2.sum_lvl1_ff[86] ;
 wire \mac2.sum_lvl1_ff[87] ;
 wire \mac2.sum_lvl1_ff[8] ;
 wire \mac2.sum_lvl1_ff[9] ;
 wire \mac2.sum_lvl2_ff[0] ;
 wire \mac2.sum_lvl2_ff[10] ;
 wire \mac2.sum_lvl2_ff[11] ;
 wire \mac2.sum_lvl2_ff[12] ;
 wire \mac2.sum_lvl2_ff[13] ;
 wire \mac2.sum_lvl2_ff[14] ;
 wire \mac2.sum_lvl2_ff[15] ;
 wire \mac2.sum_lvl2_ff[19] ;
 wire \mac2.sum_lvl2_ff[1] ;
 wire \mac2.sum_lvl2_ff[20] ;
 wire \mac2.sum_lvl2_ff[21] ;
 wire \mac2.sum_lvl2_ff[22] ;
 wire \mac2.sum_lvl2_ff[23] ;
 wire \mac2.sum_lvl2_ff[24] ;
 wire \mac2.sum_lvl2_ff[25] ;
 wire \mac2.sum_lvl2_ff[26] ;
 wire \mac2.sum_lvl2_ff[27] ;
 wire \mac2.sum_lvl2_ff[28] ;
 wire \mac2.sum_lvl2_ff[29] ;
 wire \mac2.sum_lvl2_ff[2] ;
 wire \mac2.sum_lvl2_ff[30] ;
 wire \mac2.sum_lvl2_ff[31] ;
 wire \mac2.sum_lvl2_ff[32] ;
 wire \mac2.sum_lvl2_ff[33] ;
 wire \mac2.sum_lvl2_ff[34] ;
 wire \mac2.sum_lvl2_ff[38] ;
 wire \mac2.sum_lvl2_ff[39] ;
 wire \mac2.sum_lvl2_ff[3] ;
 wire \mac2.sum_lvl2_ff[40] ;
 wire \mac2.sum_lvl2_ff[41] ;
 wire \mac2.sum_lvl2_ff[42] ;
 wire \mac2.sum_lvl2_ff[43] ;
 wire \mac2.sum_lvl2_ff[44] ;
 wire \mac2.sum_lvl2_ff[45] ;
 wire \mac2.sum_lvl2_ff[46] ;
 wire \mac2.sum_lvl2_ff[47] ;
 wire \mac2.sum_lvl2_ff[48] ;
 wire \mac2.sum_lvl2_ff[49] ;
 wire \mac2.sum_lvl2_ff[4] ;
 wire \mac2.sum_lvl2_ff[50] ;
 wire \mac2.sum_lvl2_ff[51] ;
 wire \mac2.sum_lvl2_ff[52] ;
 wire \mac2.sum_lvl2_ff[53] ;
 wire \mac2.sum_lvl2_ff[5] ;
 wire \mac2.sum_lvl2_ff[6] ;
 wire \mac2.sum_lvl2_ff[7] ;
 wire \mac2.sum_lvl2_ff[8] ;
 wire \mac2.sum_lvl2_ff[9] ;
 wire \mac2.sum_lvl3_ff[0] ;
 wire \mac2.sum_lvl3_ff[10] ;
 wire \mac2.sum_lvl3_ff[11] ;
 wire \mac2.sum_lvl3_ff[12] ;
 wire \mac2.sum_lvl3_ff[13] ;
 wire \mac2.sum_lvl3_ff[14] ;
 wire \mac2.sum_lvl3_ff[15] ;
 wire \mac2.sum_lvl3_ff[1] ;
 wire \mac2.sum_lvl3_ff[20] ;
 wire \mac2.sum_lvl3_ff[21] ;
 wire \mac2.sum_lvl3_ff[22] ;
 wire \mac2.sum_lvl3_ff[23] ;
 wire \mac2.sum_lvl3_ff[24] ;
 wire \mac2.sum_lvl3_ff[25] ;
 wire \mac2.sum_lvl3_ff[26] ;
 wire \mac2.sum_lvl3_ff[27] ;
 wire \mac2.sum_lvl3_ff[28] ;
 wire \mac2.sum_lvl3_ff[29] ;
 wire \mac2.sum_lvl3_ff[2] ;
 wire \mac2.sum_lvl3_ff[30] ;
 wire \mac2.sum_lvl3_ff[31] ;
 wire \mac2.sum_lvl3_ff[32] ;
 wire \mac2.sum_lvl3_ff[33] ;
 wire \mac2.sum_lvl3_ff[34] ;
 wire \mac2.sum_lvl3_ff[35] ;
 wire \mac2.sum_lvl3_ff[3] ;
 wire \mac2.sum_lvl3_ff[4] ;
 wire \mac2.sum_lvl3_ff[5] ;
 wire \mac2.sum_lvl3_ff[6] ;
 wire \mac2.sum_lvl3_ff[7] ;
 wire \mac2.sum_lvl3_ff[8] ;
 wire \mac2.sum_lvl3_ff[9] ;
 wire \mac2.total_sum[0] ;
 wire \mac2.total_sum[10] ;
 wire \mac2.total_sum[11] ;
 wire \mac2.total_sum[12] ;
 wire \mac2.total_sum[13] ;
 wire \mac2.total_sum[14] ;
 wire \mac2.total_sum[15] ;
 wire \mac2.total_sum[1] ;
 wire \mac2.total_sum[2] ;
 wire \mac2.total_sum[3] ;
 wire \mac2.total_sum[4] ;
 wire \mac2.total_sum[5] ;
 wire \mac2.total_sum[6] ;
 wire \mac2.total_sum[7] ;
 wire \mac2.total_sum[8] ;
 wire \mac2.total_sum[9] ;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire clknet_leaf_0_clk;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net33;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;

 sg13g2_inv_1 _3032_ (.Y(\DP_1.I_range.data_plus_4[6] ),
    .A(net4));
 sg13g2_inv_1 _3033_ (.Y(\DP_3.I_range.data_plus_4[6] ),
    .A(net16));
 sg13g2_inv_1 _3034_ (.Y(\DP_3.Q_range.data_plus_4[6] ),
    .A(net12));
 sg13g2_inv_1 _3035_ (.Y(\DP_1.Q_range.data_plus_4[6] ),
    .A(net8));
 sg13g2_inv_1 _3036_ (.Y(_2633_),
    .A(\DP_3.I_range.out_data[5] ));
 sg13g2_inv_1 _3037_ (.Y(_2634_),
    .A(net906));
 sg13g2_inv_1 _3038_ (.Y(_2635_),
    .A(net850));
 sg13g2_and2_1 _3039_ (.A(net1003),
    .B(net946),
    .X(_0064_));
 sg13g2_and3_2 _3040_ (.X(_2636_),
    .A(net1002),
    .B(net942),
    .C(_0064_));
 sg13g2_a22oi_1 _3041_ (.Y(_2637_),
    .B1(net942),
    .B2(net1003),
    .A2(net1002),
    .A1(net946));
 sg13g2_nor2_2 _3042_ (.A(_2636_),
    .B(net516),
    .Y(_0065_));
 sg13g2_nand2_1 _3043_ (.Y(_2638_),
    .A(net1003),
    .B(net937));
 sg13g2_and4_1 _3044_ (.A(net946),
    .B(net1002),
    .C(net942),
    .D(net999),
    .X(_2639_));
 sg13g2_a22oi_1 _3045_ (.Y(_2640_),
    .B1(net999),
    .B2(net946),
    .A2(net942),
    .A1(net1002));
 sg13g2_nor3_1 _3046_ (.A(_2638_),
    .B(_2639_),
    .C(_2640_),
    .Y(_2641_));
 sg13g2_o21ai_1 _3047_ (.B1(_2638_),
    .Y(_2642_),
    .A1(_2639_),
    .A2(_2640_));
 sg13g2_nor2b_1 _3048_ (.A(_2641_),
    .B_N(_2642_),
    .Y(_2643_));
 sg13g2_nand2_1 _3049_ (.Y(_2644_),
    .A(_2636_),
    .B(_2643_));
 sg13g2_xor2_1 _3050_ (.B(_2643_),
    .A(_2636_),
    .X(_0066_));
 sg13g2_nand2_1 _3051_ (.Y(_2645_),
    .A(net1003),
    .B(\DP_2.matrix[75] ));
 sg13g2_or2_1 _3052_ (.X(_2646_),
    .B(_2641_),
    .A(_2639_));
 sg13g2_nand2_1 _3053_ (.Y(_2647_),
    .A(net1001),
    .B(net937));
 sg13g2_and4_1 _3054_ (.A(net946),
    .B(net942),
    .C(net999),
    .D(net997),
    .X(_2648_));
 sg13g2_nand4_1 _3055_ (.B(net942),
    .C(net999),
    .A(net946),
    .Y(_2649_),
    .D(net996));
 sg13g2_a22oi_1 _3056_ (.Y(_2650_),
    .B1(net997),
    .B2(net946),
    .A2(net999),
    .A1(net942));
 sg13g2_nor3_1 _3057_ (.A(_2647_),
    .B(_2648_),
    .C(_2650_),
    .Y(_2651_));
 sg13g2_o21ai_1 _3058_ (.B1(_2647_),
    .Y(_2652_),
    .A1(_2648_),
    .A2(_2650_));
 sg13g2_nor2b_2 _3059_ (.A(_2651_),
    .B_N(_2652_),
    .Y(_2653_));
 sg13g2_nand2_1 _3060_ (.Y(_2654_),
    .A(_2646_),
    .B(_2653_));
 sg13g2_xnor2_1 _3061_ (.Y(_2655_),
    .A(_2646_),
    .B(_2653_));
 sg13g2_xor2_1 _3062_ (.B(_2655_),
    .A(_2645_),
    .X(_2656_));
 sg13g2_nand2b_2 _3063_ (.Y(_2657_),
    .B(_2656_),
    .A_N(_2644_));
 sg13g2_xnor2_1 _3064_ (.Y(_0067_),
    .A(_2644_),
    .B(_2656_));
 sg13g2_a22oi_1 _3065_ (.Y(_2658_),
    .B1(net932),
    .B2(net1004),
    .A2(net934),
    .A1(net1000));
 sg13g2_nand2_1 _3066_ (.Y(_2659_),
    .A(net1000),
    .B(net932));
 sg13g2_and4_1 _3067_ (.A(net1004),
    .B(net1000),
    .C(net934),
    .D(net932),
    .X(_2660_));
 sg13g2_nor2_1 _3068_ (.A(_2658_),
    .B(_2660_),
    .Y(_2661_));
 sg13g2_inv_1 _3069_ (.Y(_2662_),
    .A(_2661_));
 sg13g2_o21ai_1 _3070_ (.B1(_2649_),
    .Y(_2663_),
    .A1(_2647_),
    .A2(_2650_));
 sg13g2_nand2_1 _3071_ (.Y(_2664_),
    .A(net998),
    .B(net936));
 sg13g2_and4_1 _3072_ (.A(net945),
    .B(net941),
    .C(net996),
    .D(net995),
    .X(_2665_));
 sg13g2_nand4_1 _3073_ (.B(net941),
    .C(net996),
    .A(net945),
    .Y(_2666_),
    .D(net995));
 sg13g2_a22oi_1 _3074_ (.Y(_2667_),
    .B1(net995),
    .B2(net945),
    .A2(net996),
    .A1(net941));
 sg13g2_or3_1 _3075_ (.A(_2664_),
    .B(_2665_),
    .C(_2667_),
    .X(_2668_));
 sg13g2_o21ai_1 _3076_ (.B1(_2664_),
    .Y(_2669_),
    .A1(_2665_),
    .A2(_2667_));
 sg13g2_nand3_1 _3077_ (.B(_2668_),
    .C(_2669_),
    .A(_2663_),
    .Y(_2670_));
 sg13g2_a21oi_1 _3078_ (.A1(_2668_),
    .A2(_2669_),
    .Y(_2671_),
    .B1(_2663_));
 sg13g2_a21o_1 _3079_ (.A2(_2669_),
    .A1(_2668_),
    .B1(_2663_),
    .X(_2672_));
 sg13g2_nand2_1 _3080_ (.Y(_2673_),
    .A(_2670_),
    .B(_2672_));
 sg13g2_xnor2_1 _3081_ (.Y(_2674_),
    .A(_2662_),
    .B(_2673_));
 sg13g2_o21ai_1 _3082_ (.B1(_2654_),
    .Y(_2675_),
    .A1(_2645_),
    .A2(_2655_));
 sg13g2_nor2b_2 _3083_ (.A(_2674_),
    .B_N(_2675_),
    .Y(_2676_));
 sg13g2_xor2_1 _3084_ (.B(_2675_),
    .A(_2674_),
    .X(_2677_));
 sg13g2_or2_1 _3085_ (.X(_2678_),
    .B(_2677_),
    .A(_2657_));
 sg13g2_xor2_1 _3086_ (.B(_2677_),
    .A(_2657_),
    .X(_0068_));
 sg13g2_o21ai_1 _3087_ (.B1(_2670_),
    .Y(_2679_),
    .A1(_2662_),
    .A2(_2671_));
 sg13g2_nand2_1 _3088_ (.Y(_2680_),
    .A(net1003),
    .B(net930));
 sg13g2_nand2_1 _3089_ (.Y(_2681_),
    .A(net998),
    .B(net933));
 sg13g2_nand2_1 _3090_ (.Y(_2682_),
    .A(net999),
    .B(net934));
 sg13g2_xor2_1 _3091_ (.B(_2682_),
    .A(_2659_),
    .X(_2683_));
 sg13g2_nand2b_1 _3092_ (.Y(_2684_),
    .B(_2683_),
    .A_N(_2680_));
 sg13g2_xor2_1 _3093_ (.B(_2683_),
    .A(_2680_),
    .X(_2685_));
 sg13g2_o21ai_1 _3094_ (.B1(_2666_),
    .Y(_2686_),
    .A1(_2664_),
    .A2(_2667_));
 sg13g2_nand2_1 _3095_ (.Y(_2687_),
    .A(net936),
    .B(net997));
 sg13g2_and4_1 _3096_ (.A(net945),
    .B(net940),
    .C(net994),
    .D(net993),
    .X(_2688_));
 sg13g2_nand4_1 _3097_ (.B(net940),
    .C(net994),
    .A(net944),
    .Y(_2689_),
    .D(net991));
 sg13g2_a22oi_1 _3098_ (.Y(_2690_),
    .B1(net991),
    .B2(net944),
    .A2(net994),
    .A1(net940));
 sg13g2_or3_1 _3099_ (.A(_2687_),
    .B(_2688_),
    .C(_2690_),
    .X(_2691_));
 sg13g2_o21ai_1 _3100_ (.B1(_2687_),
    .Y(_2692_),
    .A1(_2688_),
    .A2(_2690_));
 sg13g2_and3_1 _3101_ (.X(_2693_),
    .A(_2686_),
    .B(_2691_),
    .C(_2692_));
 sg13g2_nand3_1 _3102_ (.B(_2691_),
    .C(_2692_),
    .A(_2686_),
    .Y(_2694_));
 sg13g2_a21oi_1 _3103_ (.A1(_2691_),
    .A2(_2692_),
    .Y(_2695_),
    .B1(_2686_));
 sg13g2_or3_1 _3104_ (.A(_2685_),
    .B(_2693_),
    .C(_2695_),
    .X(_2696_));
 sg13g2_o21ai_1 _3105_ (.B1(_2685_),
    .Y(_2697_),
    .A1(_2693_),
    .A2(_2695_));
 sg13g2_nand3_1 _3106_ (.B(_2696_),
    .C(_2697_),
    .A(_2679_),
    .Y(_2698_));
 sg13g2_a21o_1 _3107_ (.A2(_2697_),
    .A1(_2696_),
    .B1(_2679_),
    .X(_2699_));
 sg13g2_nand3_1 _3108_ (.B(_2698_),
    .C(_2699_),
    .A(_2660_),
    .Y(_2700_));
 sg13g2_a21o_1 _3109_ (.A2(_2699_),
    .A1(_2698_),
    .B1(_2660_),
    .X(_2701_));
 sg13g2_and2_1 _3110_ (.A(_2700_),
    .B(_2701_),
    .X(_2702_));
 sg13g2_nand3_1 _3111_ (.B(_2700_),
    .C(_2701_),
    .A(_2676_),
    .Y(_2703_));
 sg13g2_a21oi_1 _3112_ (.A1(_2700_),
    .A2(_2701_),
    .Y(_2704_),
    .B1(_2676_));
 sg13g2_xor2_1 _3113_ (.B(_2702_),
    .A(_2676_),
    .X(_2705_));
 sg13g2_xnor2_1 _3114_ (.Y(_0094_),
    .A(_2678_),
    .B(_2705_));
 sg13g2_nand2_1 _3115_ (.Y(_2706_),
    .A(_2698_),
    .B(_2700_));
 sg13g2_o21ai_1 _3116_ (.B1(_2684_),
    .Y(_2707_),
    .A1(_2659_),
    .A2(_2682_));
 sg13g2_nand2_1 _3117_ (.Y(_2708_),
    .A(net1004),
    .B(net928));
 sg13g2_nand2b_2 _3118_ (.Y(_2709_),
    .B(_2707_),
    .A_N(_2708_));
 sg13g2_xor2_1 _3119_ (.B(_2708_),
    .A(_2707_),
    .X(_2710_));
 sg13g2_o21ai_1 _3120_ (.B1(_2694_),
    .Y(_2711_),
    .A1(_2685_),
    .A2(_2695_));
 sg13g2_nand2_1 _3121_ (.Y(_2712_),
    .A(net1000),
    .B(net930));
 sg13g2_nand2_1 _3122_ (.Y(_2713_),
    .A(net997),
    .B(net933));
 sg13g2_nand2_1 _3123_ (.Y(_2714_),
    .A(net997),
    .B(net935));
 sg13g2_xor2_1 _3124_ (.B(_2714_),
    .A(_2681_),
    .X(_2715_));
 sg13g2_nand2b_1 _3125_ (.Y(_2716_),
    .B(_2715_),
    .A_N(_2712_));
 sg13g2_xnor2_1 _3126_ (.Y(_2717_),
    .A(_2712_),
    .B(_2715_));
 sg13g2_o21ai_1 _3127_ (.B1(_2689_),
    .Y(_2718_),
    .A1(_2687_),
    .A2(_2690_));
 sg13g2_nand2_1 _3128_ (.Y(_2719_),
    .A(net937),
    .B(net995));
 sg13g2_and4_1 _3129_ (.A(net944),
    .B(net939),
    .C(net992),
    .D(net989),
    .X(_2720_));
 sg13g2_nand4_1 _3130_ (.B(net939),
    .C(net992),
    .A(net943),
    .Y(_2721_),
    .D(net989));
 sg13g2_a22oi_1 _3131_ (.Y(_2722_),
    .B1(net989),
    .B2(net943),
    .A2(net992),
    .A1(net939));
 sg13g2_or3_1 _3132_ (.A(_2719_),
    .B(_2720_),
    .C(_2722_),
    .X(_2723_));
 sg13g2_o21ai_1 _3133_ (.B1(_2719_),
    .Y(_2724_),
    .A1(_2720_),
    .A2(_2722_));
 sg13g2_and3_1 _3134_ (.X(_2725_),
    .A(_2718_),
    .B(_2723_),
    .C(_2724_));
 sg13g2_nand3_1 _3135_ (.B(_2723_),
    .C(_2724_),
    .A(_2718_),
    .Y(_2726_));
 sg13g2_a21o_1 _3136_ (.A2(_2724_),
    .A1(_2723_),
    .B1(_2718_),
    .X(_2727_));
 sg13g2_nand3_1 _3137_ (.B(_2726_),
    .C(_2727_),
    .A(_2717_),
    .Y(_2728_));
 sg13g2_a21o_1 _3138_ (.A2(_2727_),
    .A1(_2726_),
    .B1(_2717_),
    .X(_2729_));
 sg13g2_nand3_1 _3139_ (.B(_2728_),
    .C(_2729_),
    .A(_2711_),
    .Y(_2730_));
 sg13g2_a21oi_1 _3140_ (.A1(_2728_),
    .A2(_2729_),
    .Y(_2731_),
    .B1(_2711_));
 sg13g2_a21o_1 _3141_ (.A2(_2729_),
    .A1(_2728_),
    .B1(_2711_),
    .X(_2732_));
 sg13g2_nand2_1 _3142_ (.Y(_2733_),
    .A(_2730_),
    .B(_2732_));
 sg13g2_xnor2_1 _3143_ (.Y(_2734_),
    .A(_2710_),
    .B(_2733_));
 sg13g2_nor2b_1 _3144_ (.A(_2734_),
    .B_N(_2706_),
    .Y(_2735_));
 sg13g2_xnor2_1 _3145_ (.Y(_2736_),
    .A(_2706_),
    .B(_2734_));
 sg13g2_o21ai_1 _3146_ (.B1(_2703_),
    .Y(_2737_),
    .A1(_2678_),
    .A2(_2704_));
 sg13g2_xor2_1 _3147_ (.B(_2737_),
    .A(_2736_),
    .X(_0101_));
 sg13g2_o21ai_1 _3148_ (.B1(_2730_),
    .Y(_2738_),
    .A1(_2710_),
    .A2(_2731_));
 sg13g2_o21ai_1 _3149_ (.B1(_2716_),
    .Y(_2739_),
    .A1(_2681_),
    .A2(_2714_));
 sg13g2_a22oi_1 _3150_ (.Y(_2740_),
    .B1(net926),
    .B2(net1003),
    .A2(net928),
    .A1(net1000));
 sg13g2_nand4_1 _3151_ (.B(net1000),
    .C(net928),
    .A(net1003),
    .Y(_2741_),
    .D(net927));
 sg13g2_nor2b_2 _3152_ (.A(_2740_),
    .B_N(_2741_),
    .Y(_2742_));
 sg13g2_nand2_1 _3153_ (.Y(_2743_),
    .A(_2739_),
    .B(_2742_));
 sg13g2_xnor2_1 _3154_ (.Y(_2744_),
    .A(_2739_),
    .B(_2742_));
 sg13g2_a21o_1 _3155_ (.A2(_2727_),
    .A1(_2717_),
    .B1(_2725_),
    .X(_2745_));
 sg13g2_nand2_1 _3156_ (.Y(_2746_),
    .A(net998),
    .B(net930));
 sg13g2_nand2_1 _3157_ (.Y(_2747_),
    .A(net995),
    .B(net933));
 sg13g2_nand2_1 _3158_ (.Y(_2748_),
    .A(net934),
    .B(net995));
 sg13g2_or2_1 _3159_ (.X(_2749_),
    .B(_2747_),
    .A(_2714_));
 sg13g2_and2_1 _3160_ (.A(_2713_),
    .B(_2748_),
    .X(_2750_));
 sg13g2_xnor2_1 _3161_ (.Y(_2751_),
    .A(_2713_),
    .B(_2748_));
 sg13g2_xnor2_1 _3162_ (.Y(_2752_),
    .A(_2746_),
    .B(_2751_));
 sg13g2_o21ai_1 _3163_ (.B1(_2721_),
    .Y(_2753_),
    .A1(_2719_),
    .A2(_2722_));
 sg13g2_nand2_1 _3164_ (.Y(_2754_),
    .A(net936),
    .B(net991));
 sg13g2_and4_1 _3165_ (.A(net943),
    .B(net938),
    .C(\DP_1.matrix[78] ),
    .D(net986),
    .X(_2755_));
 sg13g2_nand4_1 _3166_ (.B(net938),
    .C(net990),
    .A(net943),
    .Y(_2756_),
    .D(net986));
 sg13g2_a22oi_1 _3167_ (.Y(_2757_),
    .B1(net986),
    .B2(net943),
    .A2(net990),
    .A1(net938));
 sg13g2_or3_1 _3168_ (.A(_2754_),
    .B(_2755_),
    .C(_2757_),
    .X(_2758_));
 sg13g2_o21ai_1 _3169_ (.B1(_2754_),
    .Y(_2759_),
    .A1(_2755_),
    .A2(_2757_));
 sg13g2_and3_1 _3170_ (.X(_2760_),
    .A(_2753_),
    .B(_2758_),
    .C(_2759_));
 sg13g2_nand3_1 _3171_ (.B(_2758_),
    .C(_2759_),
    .A(_2753_),
    .Y(_2761_));
 sg13g2_a21oi_1 _3172_ (.A1(_2758_),
    .A2(_2759_),
    .Y(_2762_),
    .B1(_2753_));
 sg13g2_or3_1 _3173_ (.A(_2752_),
    .B(_2760_),
    .C(_2762_),
    .X(_2763_));
 sg13g2_o21ai_1 _3174_ (.B1(_2752_),
    .Y(_2764_),
    .A1(_2760_),
    .A2(_2762_));
 sg13g2_and3_1 _3175_ (.X(_2765_),
    .A(_2745_),
    .B(_2763_),
    .C(_2764_));
 sg13g2_nand3_1 _3176_ (.B(_2763_),
    .C(_2764_),
    .A(_2745_),
    .Y(_2766_));
 sg13g2_a21oi_1 _3177_ (.A1(_2763_),
    .A2(_2764_),
    .Y(_2767_),
    .B1(_2745_));
 sg13g2_or3_1 _3178_ (.A(_2744_),
    .B(_2765_),
    .C(_2767_),
    .X(_2768_));
 sg13g2_o21ai_1 _3179_ (.B1(_2744_),
    .Y(_2769_),
    .A1(_2765_),
    .A2(_2767_));
 sg13g2_nand3_1 _3180_ (.B(_2768_),
    .C(_2769_),
    .A(_2738_),
    .Y(_2770_));
 sg13g2_a21oi_1 _3181_ (.A1(_2768_),
    .A2(_2769_),
    .Y(_2771_),
    .B1(_2738_));
 sg13g2_a21o_1 _3182_ (.A2(_2769_),
    .A1(_2768_),
    .B1(_2738_),
    .X(_2772_));
 sg13g2_nand2_1 _3183_ (.Y(_2773_),
    .A(_2770_),
    .B(_2772_));
 sg13g2_xor2_1 _3184_ (.B(_2773_),
    .A(_2709_),
    .X(_2774_));
 sg13g2_a21o_2 _3185_ (.A2(_2737_),
    .A1(_2736_),
    .B1(_2735_),
    .X(_2775_));
 sg13g2_nand2_1 _3186_ (.Y(_2776_),
    .A(_2774_),
    .B(_2775_));
 sg13g2_xor2_1 _3187_ (.B(_2775_),
    .A(_2774_),
    .X(_0102_));
 sg13g2_o21ai_1 _3188_ (.B1(_2766_),
    .Y(_2777_),
    .A1(_2744_),
    .A2(_2767_));
 sg13g2_o21ai_1 _3189_ (.B1(_2749_),
    .Y(_2778_),
    .A1(_2746_),
    .A2(_2750_));
 sg13g2_nand2_1 _3190_ (.Y(_2779_),
    .A(net1004),
    .B(net1051));
 sg13g2_nand2_1 _3191_ (.Y(_2780_),
    .A(net998),
    .B(net926));
 sg13g2_and4_1 _3192_ (.A(net1001),
    .B(net998),
    .C(net929),
    .D(net926),
    .X(_2781_));
 sg13g2_a22oi_1 _3193_ (.Y(_2782_),
    .B1(net927),
    .B2(net1000),
    .A2(net929),
    .A1(net998));
 sg13g2_or2_1 _3194_ (.X(_2783_),
    .B(_2782_),
    .A(_2781_));
 sg13g2_nor2_1 _3195_ (.A(_2779_),
    .B(_2783_),
    .Y(_2784_));
 sg13g2_xor2_1 _3196_ (.B(_2783_),
    .A(_2779_),
    .X(_2785_));
 sg13g2_nand2_1 _3197_ (.Y(_2786_),
    .A(_2778_),
    .B(_2785_));
 sg13g2_xnor2_1 _3198_ (.Y(_2787_),
    .A(_2778_),
    .B(_2785_));
 sg13g2_xnor2_1 _3199_ (.Y(_2788_),
    .A(_2741_),
    .B(_2787_));
 sg13g2_o21ai_1 _3200_ (.B1(_2761_),
    .Y(_2789_),
    .A1(_2752_),
    .A2(_2762_));
 sg13g2_nand2_1 _3201_ (.Y(_2790_),
    .A(net996),
    .B(net930));
 sg13g2_nand2_2 _3202_ (.Y(_2791_),
    .A(net932),
    .B(net991));
 sg13g2_nand2_1 _3203_ (.Y(_2792_),
    .A(net934),
    .B(net992));
 sg13g2_or2_1 _3204_ (.X(_2793_),
    .B(_2791_),
    .A(_2748_));
 sg13g2_xnor2_1 _3205_ (.Y(_2794_),
    .A(_2747_),
    .B(_2792_));
 sg13g2_xnor2_1 _3206_ (.Y(_2795_),
    .A(_2790_),
    .B(_2794_));
 sg13g2_o21ai_1 _3207_ (.B1(_2756_),
    .Y(_2796_),
    .A1(_2754_),
    .A2(_2757_));
 sg13g2_nand2_1 _3208_ (.Y(_2797_),
    .A(net936),
    .B(net989));
 sg13g2_and4_1 _3209_ (.A(net944),
    .B(net939),
    .C(net986),
    .D(net1054),
    .X(_2798_));
 sg13g2_nand4_1 _3210_ (.B(net938),
    .C(net986),
    .A(net943),
    .Y(_2799_),
    .D(net1054));
 sg13g2_a22oi_1 _3211_ (.Y(_2800_),
    .B1(net1055),
    .B2(net943),
    .A2(net986),
    .A1(net938));
 sg13g2_or3_1 _3212_ (.A(_2797_),
    .B(_2798_),
    .C(_2800_),
    .X(_2801_));
 sg13g2_o21ai_1 _3213_ (.B1(_2797_),
    .Y(_2802_),
    .A1(_2798_),
    .A2(_2800_));
 sg13g2_and3_1 _3214_ (.X(_2803_),
    .A(_2796_),
    .B(_2801_),
    .C(_2802_));
 sg13g2_nand3_1 _3215_ (.B(_2801_),
    .C(_2802_),
    .A(_2796_),
    .Y(_2804_));
 sg13g2_a21oi_1 _3216_ (.A1(_2801_),
    .A2(_2802_),
    .Y(_2805_),
    .B1(_2796_));
 sg13g2_or3_1 _3217_ (.A(_2795_),
    .B(_2803_),
    .C(_2805_),
    .X(_2806_));
 sg13g2_o21ai_1 _3218_ (.B1(_2795_),
    .Y(_2807_),
    .A1(_2803_),
    .A2(_2805_));
 sg13g2_and3_1 _3219_ (.X(_2808_),
    .A(_2789_),
    .B(_2806_),
    .C(_2807_));
 sg13g2_nand3_1 _3220_ (.B(_2806_),
    .C(_2807_),
    .A(_2789_),
    .Y(_2809_));
 sg13g2_a21oi_1 _3221_ (.A1(_2806_),
    .A2(_2807_),
    .Y(_2810_),
    .B1(_2789_));
 sg13g2_or3_1 _3222_ (.A(_2788_),
    .B(_2808_),
    .C(_2810_),
    .X(_2811_));
 sg13g2_o21ai_1 _3223_ (.B1(_2788_),
    .Y(_2812_),
    .A1(_2808_),
    .A2(_2810_));
 sg13g2_and3_1 _3224_ (.X(_2813_),
    .A(_2777_),
    .B(_2811_),
    .C(_2812_));
 sg13g2_nand3_1 _3225_ (.B(_2811_),
    .C(_2812_),
    .A(_2777_),
    .Y(_2814_));
 sg13g2_a21oi_1 _3226_ (.A1(_2811_),
    .A2(_2812_),
    .Y(_2815_),
    .B1(_2777_));
 sg13g2_or3_1 _3227_ (.A(_2743_),
    .B(_2813_),
    .C(_2815_),
    .X(_2816_));
 sg13g2_o21ai_1 _3228_ (.B1(_2743_),
    .Y(_2817_),
    .A1(_2813_),
    .A2(_2815_));
 sg13g2_o21ai_1 _3229_ (.B1(_2770_),
    .Y(_2818_),
    .A1(_2709_),
    .A2(_2771_));
 sg13g2_nand3_1 _3230_ (.B(_2817_),
    .C(_2818_),
    .A(_2816_),
    .Y(_2819_));
 sg13g2_a21o_1 _3231_ (.A2(_2817_),
    .A1(_2816_),
    .B1(_2818_),
    .X(_2820_));
 sg13g2_nand2_1 _3232_ (.Y(_2821_),
    .A(_2819_),
    .B(_2820_));
 sg13g2_and4_1 _3233_ (.A(_2774_),
    .B(_2775_),
    .C(_2819_),
    .D(_2820_),
    .X(_2822_));
 sg13g2_xor2_1 _3234_ (.B(_2821_),
    .A(_2776_),
    .X(_0103_));
 sg13g2_o21ai_1 _3235_ (.B1(_2819_),
    .Y(_2823_),
    .A1(_2776_),
    .A2(_2821_));
 sg13g2_o21ai_1 _3236_ (.B1(_2814_),
    .Y(_2824_),
    .A1(_2743_),
    .A2(_2815_));
 sg13g2_o21ai_1 _3237_ (.B1(_2786_),
    .Y(_2825_),
    .A1(_2741_),
    .A2(_2787_));
 sg13g2_o21ai_1 _3238_ (.B1(_2809_),
    .Y(_2826_),
    .A1(_2788_),
    .A2(_2810_));
 sg13g2_nor2_2 _3239_ (.A(_2781_),
    .B(_2784_),
    .Y(_2827_));
 sg13g2_o21ai_1 _3240_ (.B1(_2793_),
    .Y(_2828_),
    .A1(_2790_),
    .A2(_2794_));
 sg13g2_nand2_1 _3241_ (.Y(_2829_),
    .A(net1000),
    .B(net1051));
 sg13g2_nand2_1 _3242_ (.Y(_2830_),
    .A(net996),
    .B(net927));
 sg13g2_nand2_1 _3243_ (.Y(_2831_),
    .A(net996),
    .B(net928));
 sg13g2_xor2_1 _3244_ (.B(_2831_),
    .A(_2780_),
    .X(_2832_));
 sg13g2_nand2b_1 _3245_ (.Y(_2833_),
    .B(_2832_),
    .A_N(_2829_));
 sg13g2_xnor2_1 _3246_ (.Y(_2834_),
    .A(_2829_),
    .B(_2832_));
 sg13g2_xnor2_1 _3247_ (.Y(_2835_),
    .A(_2828_),
    .B(_2834_));
 sg13g2_nor2_1 _3248_ (.A(_2827_),
    .B(_2835_),
    .Y(_2836_));
 sg13g2_xnor2_1 _3249_ (.Y(_2837_),
    .A(_2827_),
    .B(_2835_));
 sg13g2_o21ai_1 _3250_ (.B1(_2804_),
    .Y(_2838_),
    .A1(_2795_),
    .A2(_2805_));
 sg13g2_nand2_1 _3251_ (.Y(_2839_),
    .A(net994),
    .B(net930));
 sg13g2_nand2_1 _3252_ (.Y(_2840_),
    .A(net934),
    .B(net989));
 sg13g2_or2_1 _3253_ (.X(_2841_),
    .B(_2840_),
    .A(_2791_));
 sg13g2_and2_1 _3254_ (.A(_2791_),
    .B(_2840_),
    .X(_2842_));
 sg13g2_xnor2_1 _3255_ (.Y(_2843_),
    .A(_2791_),
    .B(_2840_));
 sg13g2_xnor2_1 _3256_ (.Y(_2844_),
    .A(_2839_),
    .B(_2843_));
 sg13g2_o21ai_1 _3257_ (.B1(_2799_),
    .Y(_2845_),
    .A1(_2797_),
    .A2(_2800_));
 sg13g2_nand2_1 _3258_ (.Y(_2846_),
    .A(net936),
    .B(net1055));
 sg13g2_and4_1 _3259_ (.A(net938),
    .B(net936),
    .C(net986),
    .D(net1055),
    .X(_2847_));
 sg13g2_a22oi_1 _3260_ (.Y(_2848_),
    .B1(net1055),
    .B2(net938),
    .A2(net987),
    .A1(net936));
 sg13g2_nor2_1 _3261_ (.A(_2847_),
    .B(_2848_),
    .Y(_2849_));
 sg13g2_nand2_1 _3262_ (.Y(_2850_),
    .A(_2845_),
    .B(_2849_));
 sg13g2_xnor2_1 _3263_ (.Y(_2851_),
    .A(_2845_),
    .B(_2849_));
 sg13g2_xor2_1 _3264_ (.B(_2851_),
    .A(_2844_),
    .X(_2852_));
 sg13g2_nand2_1 _3265_ (.Y(_2853_),
    .A(_2838_),
    .B(_2852_));
 sg13g2_xnor2_1 _3266_ (.Y(_2854_),
    .A(_2838_),
    .B(_2852_));
 sg13g2_xor2_1 _3267_ (.B(_2854_),
    .A(_2837_),
    .X(_2855_));
 sg13g2_nand2_1 _3268_ (.Y(_2856_),
    .A(_2826_),
    .B(_2855_));
 sg13g2_xnor2_1 _3269_ (.Y(_2857_),
    .A(_2826_),
    .B(_2855_));
 sg13g2_nand2b_1 _3270_ (.Y(_2858_),
    .B(_2825_),
    .A_N(_2857_));
 sg13g2_xnor2_1 _3271_ (.Y(_2859_),
    .A(_2825_),
    .B(_2857_));
 sg13g2_nor2_1 _3272_ (.A(_2824_),
    .B(_2859_),
    .Y(_2860_));
 sg13g2_nand2_1 _3273_ (.Y(_2861_),
    .A(_2824_),
    .B(_2859_));
 sg13g2_nor2b_1 _3274_ (.A(_2860_),
    .B_N(_2861_),
    .Y(_2862_));
 sg13g2_xor2_1 _3275_ (.B(_2862_),
    .A(_2823_),
    .X(_0104_));
 sg13g2_a21oi_1 _3276_ (.A1(_2828_),
    .A2(_2834_),
    .Y(_2863_),
    .B1(_2836_));
 sg13g2_o21ai_1 _3277_ (.B1(_2853_),
    .Y(_2864_),
    .A1(_2837_),
    .A2(_2854_));
 sg13g2_o21ai_1 _3278_ (.B1(_2833_),
    .Y(_2865_),
    .A1(_2780_),
    .A2(_2831_));
 sg13g2_o21ai_1 _3279_ (.B1(_2841_),
    .Y(_2866_),
    .A1(_2839_),
    .A2(_2842_));
 sg13g2_nand2_1 _3280_ (.Y(_2867_),
    .A(net998),
    .B(net1051));
 sg13g2_nand2_1 _3281_ (.Y(_2868_),
    .A(net994),
    .B(net926));
 sg13g2_nand2_1 _3282_ (.Y(_2869_),
    .A(net994),
    .B(net929));
 sg13g2_or2_1 _3283_ (.X(_2870_),
    .B(_2868_),
    .A(_2831_));
 sg13g2_xnor2_1 _3284_ (.Y(_2871_),
    .A(_2830_),
    .B(_2869_));
 sg13g2_xor2_1 _3285_ (.B(_2871_),
    .A(_2867_),
    .X(_2872_));
 sg13g2_xnor2_1 _3286_ (.Y(_2873_),
    .A(_2866_),
    .B(_2872_));
 sg13g2_nor2b_1 _3287_ (.A(_2873_),
    .B_N(_2865_),
    .Y(_2874_));
 sg13g2_xor2_1 _3288_ (.B(_2873_),
    .A(_2865_),
    .X(_2875_));
 sg13g2_o21ai_1 _3289_ (.B1(_2850_),
    .Y(_2876_),
    .A1(_2844_),
    .A2(_2851_));
 sg13g2_a21oi_1 _3290_ (.A1(net938),
    .A2(net986),
    .Y(_2877_),
    .B1(_2846_));
 sg13g2_nand2_1 _3291_ (.Y(_2878_),
    .A(net991),
    .B(net931));
 sg13g2_nand2_1 _3292_ (.Y(_2879_),
    .A(net932),
    .B(net988));
 sg13g2_and4_1 _3293_ (.A(net935),
    .B(net932),
    .C(net989),
    .D(net987),
    .X(_2880_));
 sg13g2_a22oi_1 _3294_ (.Y(_2881_),
    .B1(net987),
    .B2(net935),
    .A2(net989),
    .A1(net932));
 sg13g2_nor3_1 _3295_ (.A(_2878_),
    .B(_2880_),
    .C(_2881_),
    .Y(_2882_));
 sg13g2_o21ai_1 _3296_ (.B1(_2878_),
    .Y(_2883_),
    .A1(_2880_),
    .A2(_2881_));
 sg13g2_nor2b_1 _3297_ (.A(_2882_),
    .B_N(_2883_),
    .Y(_2884_));
 sg13g2_xnor2_1 _3298_ (.Y(_2885_),
    .A(_2877_),
    .B(_2884_));
 sg13g2_nand2b_1 _3299_ (.Y(_2886_),
    .B(_2876_),
    .A_N(_2885_));
 sg13g2_xor2_1 _3300_ (.B(_2885_),
    .A(_2876_),
    .X(_2887_));
 sg13g2_xor2_1 _3301_ (.B(_2887_),
    .A(_2875_),
    .X(_2888_));
 sg13g2_nand2_1 _3302_ (.Y(_2889_),
    .A(_2864_),
    .B(_2888_));
 sg13g2_xor2_1 _3303_ (.B(_2888_),
    .A(_2864_),
    .X(_2890_));
 sg13g2_nand2b_1 _3304_ (.Y(_2891_),
    .B(_2890_),
    .A_N(_2863_));
 sg13g2_xor2_1 _3305_ (.B(_2890_),
    .A(_2863_),
    .X(_2892_));
 sg13g2_a21oi_1 _3306_ (.A1(_2856_),
    .A2(_2858_),
    .Y(_2893_),
    .B1(_2892_));
 sg13g2_nand3_1 _3307_ (.B(_2858_),
    .C(_2892_),
    .A(_2856_),
    .Y(_2894_));
 sg13g2_nand2b_1 _3308_ (.Y(_2895_),
    .B(_2894_),
    .A_N(_2893_));
 sg13g2_a21oi_1 _3309_ (.A1(_2819_),
    .A2(_2861_),
    .Y(_2896_),
    .B1(_2860_));
 sg13g2_a21oi_2 _3310_ (.B1(_2896_),
    .Y(_2897_),
    .A2(_2862_),
    .A1(_2822_));
 sg13g2_nor2_1 _3311_ (.A(_2895_),
    .B(_2897_),
    .Y(_2898_));
 sg13g2_xor2_1 _3312_ (.B(_2897_),
    .A(_2895_),
    .X(_0095_));
 sg13g2_a21o_1 _3313_ (.A2(_2872_),
    .A1(_2866_),
    .B1(_2874_),
    .X(_2899_));
 sg13g2_o21ai_1 _3314_ (.B1(_2886_),
    .Y(_2900_),
    .A1(_2875_),
    .A2(_2887_));
 sg13g2_a21o_1 _3315_ (.A2(_2884_),
    .A1(_2877_),
    .B1(_2847_),
    .X(_2901_));
 sg13g2_nand2_1 _3316_ (.Y(_2902_),
    .A(net930),
    .B(net990));
 sg13g2_nand2_1 _3317_ (.Y(_2903_),
    .A(net934),
    .B(net1054));
 sg13g2_or2_1 _3318_ (.X(_2904_),
    .B(_2903_),
    .A(_2879_));
 sg13g2_xnor2_1 _3319_ (.Y(_2905_),
    .A(_2879_),
    .B(_2903_));
 sg13g2_xor2_1 _3320_ (.B(_2905_),
    .A(_2902_),
    .X(_2906_));
 sg13g2_and2_1 _3321_ (.A(_2901_),
    .B(_2906_),
    .X(_2907_));
 sg13g2_or2_1 _3322_ (.X(_2908_),
    .B(_2906_),
    .A(_2901_));
 sg13g2_xnor2_1 _3323_ (.Y(_2909_),
    .A(_2901_),
    .B(_2906_));
 sg13g2_o21ai_1 _3324_ (.B1(_2870_),
    .Y(_2910_),
    .A1(_2867_),
    .A2(_2871_));
 sg13g2_or2_1 _3325_ (.X(_2911_),
    .B(_2882_),
    .A(_2880_));
 sg13g2_nand2_1 _3326_ (.Y(_2912_),
    .A(net996),
    .B(net1051));
 sg13g2_nand2_1 _3327_ (.Y(_2913_),
    .A(net991),
    .B(net928));
 sg13g2_or2_1 _3328_ (.X(_2914_),
    .B(_2913_),
    .A(_2868_));
 sg13g2_xnor2_1 _3329_ (.Y(_2915_),
    .A(_2868_),
    .B(_2913_));
 sg13g2_xor2_1 _3330_ (.B(_2915_),
    .A(_2912_),
    .X(_2916_));
 sg13g2_xnor2_1 _3331_ (.Y(_2917_),
    .A(_2911_),
    .B(_2916_));
 sg13g2_nor2b_1 _3332_ (.A(_2917_),
    .B_N(_2910_),
    .Y(_2918_));
 sg13g2_xnor2_1 _3333_ (.Y(_2919_),
    .A(_2910_),
    .B(_2917_));
 sg13g2_xnor2_1 _3334_ (.Y(_2920_),
    .A(_2909_),
    .B(_2919_));
 sg13g2_xnor2_1 _3335_ (.Y(_2921_),
    .A(_2900_),
    .B(_2920_));
 sg13g2_nor2b_1 _3336_ (.A(_2921_),
    .B_N(_2899_),
    .Y(_2922_));
 sg13g2_xor2_1 _3337_ (.B(_2921_),
    .A(_2899_),
    .X(_2923_));
 sg13g2_nand3_1 _3338_ (.B(_2891_),
    .C(_2923_),
    .A(_2889_),
    .Y(_2924_));
 sg13g2_inv_1 _3339_ (.Y(_2925_),
    .A(_2924_));
 sg13g2_a21oi_1 _3340_ (.A1(_2889_),
    .A2(_2891_),
    .Y(_2926_),
    .B1(_2923_));
 sg13g2_nor2_1 _3341_ (.A(_2925_),
    .B(_2926_),
    .Y(_2927_));
 sg13g2_nor2_1 _3342_ (.A(_2893_),
    .B(_2898_),
    .Y(_2928_));
 sg13g2_xnor2_1 _3343_ (.Y(_0096_),
    .A(_2927_),
    .B(_2928_));
 sg13g2_a21o_1 _3344_ (.A2(_2916_),
    .A1(_2911_),
    .B1(_2918_),
    .X(_2929_));
 sg13g2_a22oi_1 _3345_ (.Y(_2930_),
    .B1(net1054),
    .B2(net932),
    .A2(net988),
    .A1(net930));
 sg13g2_nand2_1 _3346_ (.Y(_2931_),
    .A(net930),
    .B(net1054));
 sg13g2_or2_1 _3347_ (.X(_2932_),
    .B(_2931_),
    .A(_2879_));
 sg13g2_nand2b_1 _3348_ (.Y(_2933_),
    .B(_2932_),
    .A_N(_2930_));
 sg13g2_o21ai_1 _3349_ (.B1(_2914_),
    .Y(_2934_),
    .A1(_2912_),
    .A2(_2915_));
 sg13g2_o21ai_1 _3350_ (.B1(_2904_),
    .Y(_2935_),
    .A1(_2902_),
    .A2(_2905_));
 sg13g2_nand2_1 _3351_ (.Y(_2936_),
    .A(net994),
    .B(net1051));
 sg13g2_nand2_1 _3352_ (.Y(_2937_),
    .A(net990),
    .B(net926));
 sg13g2_and4_1 _3353_ (.A(net993),
    .B(net990),
    .C(net928),
    .D(net926),
    .X(_2938_));
 sg13g2_or2_1 _3354_ (.X(_2939_),
    .B(_2937_),
    .A(_2913_));
 sg13g2_a22oi_1 _3355_ (.Y(_2940_),
    .B1(net926),
    .B2(net991),
    .A2(net928),
    .A1(net990));
 sg13g2_nor2_1 _3356_ (.A(_2938_),
    .B(_2940_),
    .Y(_2941_));
 sg13g2_xnor2_1 _3357_ (.Y(_2942_),
    .A(_2936_),
    .B(_2941_));
 sg13g2_xnor2_1 _3358_ (.Y(_2943_),
    .A(_2935_),
    .B(_2942_));
 sg13g2_nor2b_1 _3359_ (.A(_2943_),
    .B_N(_2934_),
    .Y(_2944_));
 sg13g2_xor2_1 _3360_ (.B(_2943_),
    .A(_2934_),
    .X(_2945_));
 sg13g2_or2_1 _3361_ (.X(_2946_),
    .B(_2945_),
    .A(_2933_));
 sg13g2_xor2_1 _3362_ (.B(_2945_),
    .A(_2933_),
    .X(_2947_));
 sg13g2_a21oi_1 _3363_ (.A1(_2908_),
    .A2(_2919_),
    .Y(_2948_),
    .B1(_2907_));
 sg13g2_nor2b_1 _3364_ (.A(_2948_),
    .B_N(_2947_),
    .Y(_2949_));
 sg13g2_xor2_1 _3365_ (.B(_2948_),
    .A(_2947_),
    .X(_2950_));
 sg13g2_nor2b_1 _3366_ (.A(_2950_),
    .B_N(_2929_),
    .Y(_2951_));
 sg13g2_xor2_1 _3367_ (.B(_2950_),
    .A(_2929_),
    .X(_2952_));
 sg13g2_a21oi_2 _3368_ (.B1(_2922_),
    .Y(_2953_),
    .A2(_2920_),
    .A1(_2900_));
 sg13g2_nor2_1 _3369_ (.A(_2952_),
    .B(_2953_),
    .Y(_2954_));
 sg13g2_xor2_1 _3370_ (.B(_2953_),
    .A(_2952_),
    .X(_2955_));
 sg13g2_a21oi_1 _3371_ (.A1(_2893_),
    .A2(_2924_),
    .Y(_2956_),
    .B1(_2926_));
 sg13g2_a21oi_1 _3372_ (.A1(_2894_),
    .A2(_2924_),
    .Y(_2957_),
    .B1(_2926_));
 sg13g2_a21oi_2 _3373_ (.B1(_2957_),
    .Y(_2958_),
    .A2(_2956_),
    .A1(_2897_));
 sg13g2_xor2_1 _3374_ (.B(_2958_),
    .A(_2955_),
    .X(_0097_));
 sg13g2_a21o_1 _3375_ (.A2(_2942_),
    .A1(_2935_),
    .B1(_2944_),
    .X(_2959_));
 sg13g2_o21ai_1 _3376_ (.B1(_2939_),
    .Y(_2960_),
    .A1(_2936_),
    .A2(_2940_));
 sg13g2_nand2_1 _3377_ (.Y(_2961_),
    .A(net993),
    .B(\DP_2.matrix[80] ));
 sg13g2_nand2_1 _3378_ (.Y(_2962_),
    .A(net988),
    .B(net927));
 sg13g2_nand2_1 _3379_ (.Y(_2963_),
    .A(net928),
    .B(net988));
 sg13g2_xor2_1 _3380_ (.B(_2963_),
    .A(_2937_),
    .X(_2964_));
 sg13g2_nand2b_1 _3381_ (.Y(_2965_),
    .B(_2964_),
    .A_N(_2961_));
 sg13g2_xnor2_1 _3382_ (.Y(_2966_),
    .A(_2961_),
    .B(_2964_));
 sg13g2_nor2b_1 _3383_ (.A(_2932_),
    .B_N(_2966_),
    .Y(_2967_));
 sg13g2_xnor2_1 _3384_ (.Y(_2968_),
    .A(_2932_),
    .B(_2966_));
 sg13g2_xnor2_1 _3385_ (.Y(_2969_),
    .A(_2960_),
    .B(_2968_));
 sg13g2_nor2_1 _3386_ (.A(_2931_),
    .B(_2969_),
    .Y(_2970_));
 sg13g2_xnor2_1 _3387_ (.Y(_2971_),
    .A(_2931_),
    .B(_2969_));
 sg13g2_nor2_1 _3388_ (.A(_2946_),
    .B(_2971_),
    .Y(_2972_));
 sg13g2_xor2_1 _3389_ (.B(_2971_),
    .A(_2946_),
    .X(_2973_));
 sg13g2_xor2_1 _3390_ (.B(_2973_),
    .A(_2959_),
    .X(_2974_));
 sg13g2_o21ai_1 _3391_ (.B1(_2974_),
    .Y(_2975_),
    .A1(_2949_),
    .A2(_2951_));
 sg13g2_or3_1 _3392_ (.A(_2949_),
    .B(_2951_),
    .C(_2974_),
    .X(_2976_));
 sg13g2_and2_1 _3393_ (.A(_2975_),
    .B(_2976_),
    .X(_2977_));
 sg13g2_a21oi_1 _3394_ (.A1(_2955_),
    .A2(_2958_),
    .Y(_2978_),
    .B1(_2954_));
 sg13g2_xnor2_1 _3395_ (.Y(_0098_),
    .A(_2977_),
    .B(_2978_));
 sg13g2_nand2_1 _3396_ (.Y(_2979_),
    .A(_2955_),
    .B(_2977_));
 sg13g2_inv_1 _3397_ (.Y(_2980_),
    .A(_2979_));
 sg13g2_o21ai_1 _3398_ (.B1(_2975_),
    .Y(_2981_),
    .A1(_2952_),
    .A2(_2953_));
 sg13g2_a22oi_1 _3399_ (.Y(_2982_),
    .B1(_2981_),
    .B2(_2976_),
    .A2(_2980_),
    .A1(_2958_));
 sg13g2_a21oi_1 _3400_ (.A1(_2959_),
    .A2(_2973_),
    .Y(_2983_),
    .B1(_2972_));
 sg13g2_a21o_1 _3401_ (.A2(_2968_),
    .A1(_2960_),
    .B1(_2967_),
    .X(_2984_));
 sg13g2_o21ai_1 _3402_ (.B1(_2965_),
    .Y(_2985_),
    .A1(_2937_),
    .A2(_2963_));
 sg13g2_nand2_1 _3403_ (.Y(_2986_),
    .A(net990),
    .B(net1051));
 sg13g2_nand2_1 _3404_ (.Y(_2987_),
    .A(net927),
    .B(net1054));
 sg13g2_nand2_1 _3405_ (.Y(_2988_),
    .A(net929),
    .B(net1054));
 sg13g2_xor2_1 _3406_ (.B(_2988_),
    .A(_2962_),
    .X(_2989_));
 sg13g2_nand2b_1 _3407_ (.Y(_2990_),
    .B(_2989_),
    .A_N(_2986_));
 sg13g2_xnor2_1 _3408_ (.Y(_2991_),
    .A(_2986_),
    .B(_2989_));
 sg13g2_nand2_1 _3409_ (.Y(_2992_),
    .A(_2985_),
    .B(_2991_));
 sg13g2_xor2_1 _3410_ (.B(_2991_),
    .A(_2985_),
    .X(_2993_));
 sg13g2_xnor2_1 _3411_ (.Y(_2994_),
    .A(_2970_),
    .B(_2993_));
 sg13g2_nor2b_1 _3412_ (.A(_2994_),
    .B_N(_2984_),
    .Y(_2995_));
 sg13g2_xor2_1 _3413_ (.B(_2994_),
    .A(_2984_),
    .X(_2996_));
 sg13g2_or2_1 _3414_ (.X(_2997_),
    .B(_2996_),
    .A(_2983_));
 sg13g2_xor2_1 _3415_ (.B(_2996_),
    .A(_2983_),
    .X(_2998_));
 sg13g2_inv_1 _3416_ (.Y(_2999_),
    .A(_2998_));
 sg13g2_xnor2_1 _3417_ (.Y(_0099_),
    .A(_2982_),
    .B(_2998_));
 sg13g2_o21ai_1 _3418_ (.B1(_2997_),
    .Y(_3000_),
    .A1(_2982_),
    .A2(_2999_));
 sg13g2_a21oi_1 _3419_ (.A1(_2970_),
    .A2(_2993_),
    .Y(_3001_),
    .B1(_2995_));
 sg13g2_nand2_1 _3420_ (.Y(_3002_),
    .A(net988),
    .B(net1051));
 sg13g2_xor2_1 _3421_ (.B(_3002_),
    .A(_2987_),
    .X(_3003_));
 sg13g2_o21ai_1 _3422_ (.B1(_2990_),
    .Y(_3004_),
    .A1(_2962_),
    .A2(_2988_));
 sg13g2_xnor2_1 _3423_ (.Y(_3005_),
    .A(_3003_),
    .B(_3004_));
 sg13g2_xnor2_1 _3424_ (.Y(_3006_),
    .A(_2992_),
    .B(_3005_));
 sg13g2_xnor2_1 _3425_ (.Y(_3007_),
    .A(_3001_),
    .B(_3006_));
 sg13g2_xnor2_1 _3426_ (.Y(_0100_),
    .A(_3000_),
    .B(_3007_));
 sg13g2_and2_1 _3427_ (.A(net1040),
    .B(net982),
    .X(_0069_));
 sg13g2_and3_2 _3428_ (.X(_3008_),
    .A(net1038),
    .B(net978),
    .C(_0069_));
 sg13g2_a22oi_1 _3429_ (.Y(_3009_),
    .B1(net978),
    .B2(net1040),
    .A2(net1038),
    .A1(net982));
 sg13g2_nor2_2 _3430_ (.A(_3008_),
    .B(_3009_),
    .Y(_0070_));
 sg13g2_nand2_1 _3431_ (.Y(_3010_),
    .A(net1040),
    .B(net976));
 sg13g2_and4_1 _3432_ (.A(net982),
    .B(net1038),
    .C(net978),
    .D(net1036),
    .X(_3011_));
 sg13g2_a22oi_1 _3433_ (.Y(_3012_),
    .B1(net1036),
    .B2(net982),
    .A2(net978),
    .A1(net1038));
 sg13g2_nor3_1 _3434_ (.A(_3010_),
    .B(_3011_),
    .C(_3012_),
    .Y(_3013_));
 sg13g2_o21ai_1 _3435_ (.B1(_3010_),
    .Y(_3014_),
    .A1(_3011_),
    .A2(_3012_));
 sg13g2_nor2b_1 _3436_ (.A(_3013_),
    .B_N(_3014_),
    .Y(_3015_));
 sg13g2_nand2_1 _3437_ (.Y(_3016_),
    .A(_3008_),
    .B(_3015_));
 sg13g2_xor2_1 _3438_ (.B(_3015_),
    .A(_3008_),
    .X(_0071_));
 sg13g2_nand2_1 _3439_ (.Y(_3017_),
    .A(net1040),
    .B(net974));
 sg13g2_or2_1 _3440_ (.X(_3018_),
    .B(_3013_),
    .A(_3011_));
 sg13g2_nand2_1 _3441_ (.Y(_3019_),
    .A(net1038),
    .B(net976));
 sg13g2_and4_1 _3442_ (.A(net982),
    .B(net978),
    .C(net1036),
    .D(net1034),
    .X(_3020_));
 sg13g2_nand4_1 _3443_ (.B(net978),
    .C(net1036),
    .A(net982),
    .Y(_3021_),
    .D(net1034));
 sg13g2_a22oi_1 _3444_ (.Y(_3022_),
    .B1(net1034),
    .B2(\DP_2.matrix[0] ),
    .A2(net1036),
    .A1(\DP_2.matrix[1] ));
 sg13g2_nor3_1 _3445_ (.A(_3019_),
    .B(_3020_),
    .C(_3022_),
    .Y(_3023_));
 sg13g2_o21ai_1 _3446_ (.B1(_3019_),
    .Y(_3024_),
    .A1(_3020_),
    .A2(_3022_));
 sg13g2_nor2b_1 _3447_ (.A(_3023_),
    .B_N(_3024_),
    .Y(_3025_));
 sg13g2_nand2_1 _3448_ (.Y(_3026_),
    .A(_3018_),
    .B(_3025_));
 sg13g2_xnor2_1 _3449_ (.Y(_3027_),
    .A(_3018_),
    .B(_3025_));
 sg13g2_xor2_1 _3450_ (.B(_3027_),
    .A(_3017_),
    .X(_3028_));
 sg13g2_nand2b_1 _3451_ (.Y(_3029_),
    .B(_3028_),
    .A_N(_3016_));
 sg13g2_xnor2_1 _3452_ (.Y(_0072_),
    .A(_3016_),
    .B(_3028_));
 sg13g2_a22oi_1 _3453_ (.Y(_3030_),
    .B1(net972),
    .B2(net1040),
    .A2(net974),
    .A1(net1038));
 sg13g2_nand2_1 _3454_ (.Y(_3031_),
    .A(net1039),
    .B(net972));
 sg13g2_and4_1 _3455_ (.A(net1041),
    .B(net1039),
    .C(net974),
    .D(net972),
    .X(_0268_));
 sg13g2_nor2_1 _3456_ (.A(_3030_),
    .B(_0268_),
    .Y(_0269_));
 sg13g2_inv_1 _3457_ (.Y(_0270_),
    .A(_0269_));
 sg13g2_o21ai_1 _3458_ (.B1(_3021_),
    .Y(_0271_),
    .A1(_3019_),
    .A2(_3022_));
 sg13g2_nand2_1 _3459_ (.Y(_0272_),
    .A(net1037),
    .B(net976));
 sg13g2_and4_1 _3460_ (.A(net985),
    .B(net981),
    .C(net1034),
    .D(net1033),
    .X(_0273_));
 sg13g2_nand4_1 _3461_ (.B(net979),
    .C(net1034),
    .A(net985),
    .Y(_0274_),
    .D(net1033));
 sg13g2_a22oi_1 _3462_ (.Y(_0275_),
    .B1(net1033),
    .B2(net985),
    .A2(net1034),
    .A1(net981));
 sg13g2_or3_1 _3463_ (.A(_0272_),
    .B(_0273_),
    .C(_0275_),
    .X(_0276_));
 sg13g2_o21ai_1 _3464_ (.B1(_0272_),
    .Y(_0277_),
    .A1(_0273_),
    .A2(_0275_));
 sg13g2_nand3_1 _3465_ (.B(_0276_),
    .C(_0277_),
    .A(_0271_),
    .Y(_0278_));
 sg13g2_a21oi_1 _3466_ (.A1(_0276_),
    .A2(_0277_),
    .Y(_0279_),
    .B1(_0271_));
 sg13g2_a21o_1 _3467_ (.A2(_0277_),
    .A1(_0276_),
    .B1(_0271_),
    .X(_0280_));
 sg13g2_nand2_1 _3468_ (.Y(_0281_),
    .A(_0278_),
    .B(_0280_));
 sg13g2_xnor2_1 _3469_ (.Y(_0282_),
    .A(_0270_),
    .B(_0281_));
 sg13g2_o21ai_1 _3470_ (.B1(_3026_),
    .Y(_0283_),
    .A1(_3017_),
    .A2(_3027_));
 sg13g2_nor2b_2 _3471_ (.A(_0282_),
    .B_N(_0283_),
    .Y(_0284_));
 sg13g2_xor2_1 _3472_ (.B(_0283_),
    .A(_0282_),
    .X(_0285_));
 sg13g2_or2_1 _3473_ (.X(_0286_),
    .B(_0285_),
    .A(_3029_));
 sg13g2_xor2_1 _3474_ (.B(_0285_),
    .A(_3029_),
    .X(_0073_));
 sg13g2_o21ai_1 _3475_ (.B1(_0278_),
    .Y(_0287_),
    .A1(_0270_),
    .A2(_0279_));
 sg13g2_nand2_1 _3476_ (.Y(_0288_),
    .A(net1040),
    .B(\DP_2.matrix[5] ));
 sg13g2_nand2_1 _3477_ (.Y(_0289_),
    .A(net1037),
    .B(net972));
 sg13g2_nand2_1 _3478_ (.Y(_0290_),
    .A(net1037),
    .B(net974));
 sg13g2_xor2_1 _3479_ (.B(_0290_),
    .A(_3031_),
    .X(_0291_));
 sg13g2_nand2b_1 _3480_ (.Y(_0292_),
    .B(_0291_),
    .A_N(_0288_));
 sg13g2_xor2_1 _3481_ (.B(_0291_),
    .A(_0288_),
    .X(_0293_));
 sg13g2_o21ai_1 _3482_ (.B1(_0274_),
    .Y(_0294_),
    .A1(_0272_),
    .A2(_0275_));
 sg13g2_nand2_1 _3483_ (.Y(_0295_),
    .A(net976),
    .B(net1035));
 sg13g2_and4_1 _3484_ (.A(net984),
    .B(net979),
    .C(net1032),
    .D(net1030),
    .X(_0296_));
 sg13g2_nand4_1 _3485_ (.B(net979),
    .C(net1033),
    .A(net983),
    .Y(_0297_),
    .D(net1030));
 sg13g2_a22oi_1 _3486_ (.Y(_0298_),
    .B1(net1030),
    .B2(net983),
    .A2(net1032),
    .A1(net979));
 sg13g2_or3_1 _3487_ (.A(_0295_),
    .B(_0296_),
    .C(_0298_),
    .X(_0299_));
 sg13g2_o21ai_1 _3488_ (.B1(_0295_),
    .Y(_0300_),
    .A1(_0296_),
    .A2(_0298_));
 sg13g2_and3_1 _3489_ (.X(_0301_),
    .A(_0294_),
    .B(_0299_),
    .C(_0300_));
 sg13g2_nand3_1 _3490_ (.B(_0299_),
    .C(_0300_),
    .A(_0294_),
    .Y(_0302_));
 sg13g2_a21oi_1 _3491_ (.A1(_0299_),
    .A2(_0300_),
    .Y(_0303_),
    .B1(_0294_));
 sg13g2_or3_1 _3492_ (.A(_0293_),
    .B(_0301_),
    .C(_0303_),
    .X(_0304_));
 sg13g2_o21ai_1 _3493_ (.B1(_0293_),
    .Y(_0305_),
    .A1(_0301_),
    .A2(_0303_));
 sg13g2_nand3_1 _3494_ (.B(_0304_),
    .C(_0305_),
    .A(_0287_),
    .Y(_0306_));
 sg13g2_a21o_1 _3495_ (.A2(_0305_),
    .A1(_0304_),
    .B1(_0287_),
    .X(_0307_));
 sg13g2_nand3_1 _3496_ (.B(_0306_),
    .C(_0307_),
    .A(_0268_),
    .Y(_0308_));
 sg13g2_a21o_1 _3497_ (.A2(_0307_),
    .A1(_0306_),
    .B1(_0268_),
    .X(_0309_));
 sg13g2_and2_1 _3498_ (.A(_0308_),
    .B(_0309_),
    .X(_0310_));
 sg13g2_nand3_1 _3499_ (.B(_0308_),
    .C(_0309_),
    .A(_0284_),
    .Y(_0311_));
 sg13g2_a21oi_1 _3500_ (.A1(_0308_),
    .A2(_0309_),
    .Y(_0312_),
    .B1(_0284_));
 sg13g2_xor2_1 _3501_ (.B(_0310_),
    .A(_0284_),
    .X(_0313_));
 sg13g2_xnor2_1 _3502_ (.Y(_0105_),
    .A(_0286_),
    .B(_0313_));
 sg13g2_nand2_1 _3503_ (.Y(_0314_),
    .A(_0306_),
    .B(_0308_));
 sg13g2_o21ai_1 _3504_ (.B1(_0292_),
    .Y(_0315_),
    .A1(_3031_),
    .A2(_0290_));
 sg13g2_nand2_1 _3505_ (.Y(_0316_),
    .A(net1041),
    .B(net970));
 sg13g2_nand2b_1 _3506_ (.Y(_0317_),
    .B(_0315_),
    .A_N(_0316_));
 sg13g2_xor2_1 _3507_ (.B(_0316_),
    .A(_0315_),
    .X(_0318_));
 sg13g2_o21ai_1 _3508_ (.B1(_0302_),
    .Y(_0319_),
    .A1(_0293_),
    .A2(_0303_));
 sg13g2_nand2_1 _3509_ (.Y(_0320_),
    .A(net1039),
    .B(\DP_2.matrix[5] ));
 sg13g2_nand2_1 _3510_ (.Y(_0321_),
    .A(net1035),
    .B(net972));
 sg13g2_nand2_2 _3511_ (.Y(_0322_),
    .A(net1035),
    .B(net974));
 sg13g2_xor2_1 _3512_ (.B(_0322_),
    .A(_0289_),
    .X(_0323_));
 sg13g2_nand2b_1 _3513_ (.Y(_0324_),
    .B(_0323_),
    .A_N(_0320_));
 sg13g2_xnor2_1 _3514_ (.Y(_0325_),
    .A(_0320_),
    .B(_0323_));
 sg13g2_o21ai_1 _3515_ (.B1(_0297_),
    .Y(_0326_),
    .A1(_0295_),
    .A2(_0298_));
 sg13g2_nand2_1 _3516_ (.Y(_0327_),
    .A(net976),
    .B(net1033));
 sg13g2_and4_1 _3517_ (.A(net983),
    .B(net979),
    .C(net1030),
    .D(net1029),
    .X(_0328_));
 sg13g2_nand4_1 _3518_ (.B(net979),
    .C(net1030),
    .A(net983),
    .Y(_0329_),
    .D(net1029));
 sg13g2_a22oi_1 _3519_ (.Y(_0330_),
    .B1(net1029),
    .B2(net983),
    .A2(net1030),
    .A1(net979));
 sg13g2_or3_1 _3520_ (.A(_0327_),
    .B(_0328_),
    .C(_0330_),
    .X(_0331_));
 sg13g2_o21ai_1 _3521_ (.B1(_0327_),
    .Y(_0332_),
    .A1(_0328_),
    .A2(_0330_));
 sg13g2_and3_1 _3522_ (.X(_0333_),
    .A(_0326_),
    .B(_0331_),
    .C(_0332_));
 sg13g2_nand3_1 _3523_ (.B(_0331_),
    .C(_0332_),
    .A(_0326_),
    .Y(_0334_));
 sg13g2_a21o_1 _3524_ (.A2(_0332_),
    .A1(_0331_),
    .B1(_0326_),
    .X(_0335_));
 sg13g2_nand3_1 _3525_ (.B(_0334_),
    .C(_0335_),
    .A(_0325_),
    .Y(_0336_));
 sg13g2_a21o_1 _3526_ (.A2(_0335_),
    .A1(_0334_),
    .B1(_0325_),
    .X(_0337_));
 sg13g2_nand3_1 _3527_ (.B(_0336_),
    .C(_0337_),
    .A(_0319_),
    .Y(_0338_));
 sg13g2_a21oi_1 _3528_ (.A1(_0336_),
    .A2(_0337_),
    .Y(_0339_),
    .B1(_0319_));
 sg13g2_a21o_1 _3529_ (.A2(_0337_),
    .A1(_0336_),
    .B1(_0319_),
    .X(_0340_));
 sg13g2_nand2_1 _3530_ (.Y(_0341_),
    .A(_0338_),
    .B(_0340_));
 sg13g2_xnor2_1 _3531_ (.Y(_0342_),
    .A(_0318_),
    .B(_0341_));
 sg13g2_nor2b_1 _3532_ (.A(_0342_),
    .B_N(_0314_),
    .Y(_0343_));
 sg13g2_xnor2_1 _3533_ (.Y(_0344_),
    .A(_0314_),
    .B(_0342_));
 sg13g2_o21ai_1 _3534_ (.B1(_0311_),
    .Y(_0345_),
    .A1(_0286_),
    .A2(_0312_));
 sg13g2_xor2_1 _3535_ (.B(_0345_),
    .A(_0344_),
    .X(_0112_));
 sg13g2_o21ai_1 _3536_ (.B1(_0338_),
    .Y(_0346_),
    .A1(_0318_),
    .A2(_0339_));
 sg13g2_o21ai_1 _3537_ (.B1(_0324_),
    .Y(_0347_),
    .A1(_0289_),
    .A2(_0322_));
 sg13g2_a22oi_1 _3538_ (.Y(_0348_),
    .B1(net966),
    .B2(net1041),
    .A2(net970),
    .A1(net1039));
 sg13g2_nand4_1 _3539_ (.B(\DP_1.matrix[1] ),
    .C(net970),
    .A(net1041),
    .Y(_0349_),
    .D(net966));
 sg13g2_nor2b_1 _3540_ (.A(_0348_),
    .B_N(_0349_),
    .Y(_0350_));
 sg13g2_nand2_1 _3541_ (.Y(_0351_),
    .A(_0347_),
    .B(_0350_));
 sg13g2_xnor2_1 _3542_ (.Y(_0352_),
    .A(_0347_),
    .B(_0350_));
 sg13g2_a21o_1 _3543_ (.A2(_0335_),
    .A1(_0325_),
    .B1(_0333_),
    .X(_0353_));
 sg13g2_nand2_1 _3544_ (.Y(_0354_),
    .A(net1036),
    .B(\DP_2.matrix[5] ));
 sg13g2_nand2_1 _3545_ (.Y(_0355_),
    .A(net1032),
    .B(net972));
 sg13g2_nand2_1 _3546_ (.Y(_0356_),
    .A(net974),
    .B(net1032));
 sg13g2_or2_1 _3547_ (.X(_0357_),
    .B(_0355_),
    .A(_0322_));
 sg13g2_and2_1 _3548_ (.A(_0321_),
    .B(_0356_),
    .X(_0358_));
 sg13g2_xnor2_1 _3549_ (.Y(_0359_),
    .A(_0321_),
    .B(_0356_));
 sg13g2_xnor2_1 _3550_ (.Y(_0360_),
    .A(_0354_),
    .B(_0359_));
 sg13g2_o21ai_1 _3551_ (.B1(_0329_),
    .Y(_0361_),
    .A1(_0327_),
    .A2(_0330_));
 sg13g2_nand2_1 _3552_ (.Y(_0362_),
    .A(net976),
    .B(net1030));
 sg13g2_and4_1 _3553_ (.A(net984),
    .B(net980),
    .C(net1028),
    .D(net1025),
    .X(_0363_));
 sg13g2_nand4_1 _3554_ (.B(net980),
    .C(net1028),
    .A(net983),
    .Y(_0364_),
    .D(net1025));
 sg13g2_a22oi_1 _3555_ (.Y(_0365_),
    .B1(net1025),
    .B2(net983),
    .A2(net1028),
    .A1(net980));
 sg13g2_or3_1 _3556_ (.A(_0362_),
    .B(_0363_),
    .C(_0365_),
    .X(_0366_));
 sg13g2_o21ai_1 _3557_ (.B1(_0362_),
    .Y(_0367_),
    .A1(_0363_),
    .A2(_0365_));
 sg13g2_and3_1 _3558_ (.X(_0368_),
    .A(_0361_),
    .B(_0366_),
    .C(_0367_));
 sg13g2_nand3_1 _3559_ (.B(_0366_),
    .C(_0367_),
    .A(_0361_),
    .Y(_0369_));
 sg13g2_a21oi_1 _3560_ (.A1(_0366_),
    .A2(_0367_),
    .Y(_0370_),
    .B1(_0361_));
 sg13g2_or3_1 _3561_ (.A(_0360_),
    .B(_0368_),
    .C(_0370_),
    .X(_0371_));
 sg13g2_o21ai_1 _3562_ (.B1(_0360_),
    .Y(_0372_),
    .A1(_0368_),
    .A2(_0370_));
 sg13g2_and3_1 _3563_ (.X(_0373_),
    .A(_0353_),
    .B(_0371_),
    .C(_0372_));
 sg13g2_nand3_1 _3564_ (.B(_0371_),
    .C(_0372_),
    .A(_0353_),
    .Y(_0374_));
 sg13g2_a21oi_1 _3565_ (.A1(_0371_),
    .A2(_0372_),
    .Y(_0375_),
    .B1(_0353_));
 sg13g2_or3_1 _3566_ (.A(_0352_),
    .B(_0373_),
    .C(_0375_),
    .X(_0376_));
 sg13g2_o21ai_1 _3567_ (.B1(_0352_),
    .Y(_0377_),
    .A1(_0373_),
    .A2(_0375_));
 sg13g2_nand3_1 _3568_ (.B(_0376_),
    .C(_0377_),
    .A(_0346_),
    .Y(_0378_));
 sg13g2_a21oi_1 _3569_ (.A1(_0376_),
    .A2(_0377_),
    .Y(_0379_),
    .B1(_0346_));
 sg13g2_a21o_1 _3570_ (.A2(_0377_),
    .A1(_0376_),
    .B1(_0346_),
    .X(_0380_));
 sg13g2_nand2_1 _3571_ (.Y(_0381_),
    .A(_0378_),
    .B(_0380_));
 sg13g2_xor2_1 _3572_ (.B(_0381_),
    .A(_0317_),
    .X(_0382_));
 sg13g2_a21o_2 _3573_ (.A2(_0345_),
    .A1(_0344_),
    .B1(_0343_),
    .X(_0383_));
 sg13g2_nand2_1 _3574_ (.Y(_0384_),
    .A(_0382_),
    .B(_0383_));
 sg13g2_xor2_1 _3575_ (.B(_0383_),
    .A(_0382_),
    .X(_0113_));
 sg13g2_o21ai_1 _3576_ (.B1(_0374_),
    .Y(_0385_),
    .A1(_0352_),
    .A2(_0375_));
 sg13g2_o21ai_1 _3577_ (.B1(_0357_),
    .Y(_0386_),
    .A1(_0354_),
    .A2(_0358_));
 sg13g2_nand2_1 _3578_ (.Y(_0387_),
    .A(net1041),
    .B(net1053));
 sg13g2_nand2_1 _3579_ (.Y(_0388_),
    .A(net1037),
    .B(net967));
 sg13g2_and4_1 _3580_ (.A(net1039),
    .B(net1037),
    .C(net970),
    .D(net967),
    .X(_0389_));
 sg13g2_a22oi_1 _3581_ (.Y(_0390_),
    .B1(net967),
    .B2(net1039),
    .A2(net970),
    .A1(net1037));
 sg13g2_or2_1 _3582_ (.X(_0391_),
    .B(_0390_),
    .A(_0389_));
 sg13g2_nor2_1 _3583_ (.A(_0387_),
    .B(_0391_),
    .Y(_0392_));
 sg13g2_xor2_1 _3584_ (.B(_0391_),
    .A(_0387_),
    .X(_0393_));
 sg13g2_nand2_1 _3585_ (.Y(_0394_),
    .A(_0386_),
    .B(_0393_));
 sg13g2_xnor2_1 _3586_ (.Y(_0395_),
    .A(_0386_),
    .B(_0393_));
 sg13g2_xnor2_1 _3587_ (.Y(_0396_),
    .A(_0349_),
    .B(_0395_));
 sg13g2_o21ai_1 _3588_ (.B1(_0369_),
    .Y(_0397_),
    .A1(_0360_),
    .A2(_0370_));
 sg13g2_nand2_1 _3589_ (.Y(_0398_),
    .A(net1035),
    .B(net971));
 sg13g2_nand2_2 _3590_ (.Y(_0399_),
    .A(net973),
    .B(net1030));
 sg13g2_nand2_1 _3591_ (.Y(_0400_),
    .A(net975),
    .B(net1031));
 sg13g2_or2_1 _3592_ (.X(_0401_),
    .B(_0399_),
    .A(_0356_));
 sg13g2_xnor2_1 _3593_ (.Y(_0402_),
    .A(_0355_),
    .B(_0400_));
 sg13g2_xnor2_1 _3594_ (.Y(_0403_),
    .A(_0398_),
    .B(_0402_));
 sg13g2_o21ai_1 _3595_ (.B1(_0364_),
    .Y(_0404_),
    .A1(_0362_),
    .A2(_0365_));
 sg13g2_nand2_1 _3596_ (.Y(_0405_),
    .A(net977),
    .B(net1028));
 sg13g2_and4_1 _3597_ (.A(net984),
    .B(net980),
    .C(net1025),
    .D(net1058),
    .X(_0406_));
 sg13g2_nand4_1 _3598_ (.B(net979),
    .C(net1025),
    .A(net983),
    .Y(_0407_),
    .D(net1058));
 sg13g2_a22oi_1 _3599_ (.Y(_0408_),
    .B1(net1058),
    .B2(net984),
    .A2(\DP_1.matrix[7] ),
    .A1(net980));
 sg13g2_or3_1 _3600_ (.A(_0405_),
    .B(_0406_),
    .C(_0408_),
    .X(_0409_));
 sg13g2_o21ai_1 _3601_ (.B1(_0405_),
    .Y(_0410_),
    .A1(_0406_),
    .A2(_0408_));
 sg13g2_and3_1 _3602_ (.X(_0411_),
    .A(_0404_),
    .B(_0409_),
    .C(_0410_));
 sg13g2_nand3_1 _3603_ (.B(_0409_),
    .C(_0410_),
    .A(_0404_),
    .Y(_0412_));
 sg13g2_a21oi_1 _3604_ (.A1(_0409_),
    .A2(_0410_),
    .Y(_0413_),
    .B1(_0404_));
 sg13g2_or3_1 _3605_ (.A(_0403_),
    .B(_0411_),
    .C(_0413_),
    .X(_0414_));
 sg13g2_o21ai_1 _3606_ (.B1(_0403_),
    .Y(_0415_),
    .A1(_0411_),
    .A2(_0413_));
 sg13g2_and3_1 _3607_ (.X(_0416_),
    .A(_0397_),
    .B(_0414_),
    .C(_0415_));
 sg13g2_nand3_1 _3608_ (.B(_0414_),
    .C(_0415_),
    .A(_0397_),
    .Y(_0417_));
 sg13g2_a21oi_1 _3609_ (.A1(_0414_),
    .A2(_0415_),
    .Y(_0418_),
    .B1(_0397_));
 sg13g2_or3_1 _3610_ (.A(_0396_),
    .B(_0416_),
    .C(_0418_),
    .X(_0419_));
 sg13g2_o21ai_1 _3611_ (.B1(_0396_),
    .Y(_0420_),
    .A1(_0416_),
    .A2(_0418_));
 sg13g2_and3_1 _3612_ (.X(_0421_),
    .A(_0385_),
    .B(_0419_),
    .C(_0420_));
 sg13g2_nand3_1 _3613_ (.B(_0419_),
    .C(_0420_),
    .A(_0385_),
    .Y(_0422_));
 sg13g2_a21oi_1 _3614_ (.A1(_0419_),
    .A2(_0420_),
    .Y(_0423_),
    .B1(_0385_));
 sg13g2_or3_1 _3615_ (.A(_0351_),
    .B(_0421_),
    .C(_0423_),
    .X(_0424_));
 sg13g2_o21ai_1 _3616_ (.B1(_0351_),
    .Y(_0425_),
    .A1(_0421_),
    .A2(_0423_));
 sg13g2_o21ai_1 _3617_ (.B1(_0378_),
    .Y(_0426_),
    .A1(_0317_),
    .A2(_0379_));
 sg13g2_nand3_1 _3618_ (.B(_0425_),
    .C(_0426_),
    .A(_0424_),
    .Y(_0427_));
 sg13g2_a21o_1 _3619_ (.A2(_0425_),
    .A1(_0424_),
    .B1(_0426_),
    .X(_0428_));
 sg13g2_nand2_1 _3620_ (.Y(_0429_),
    .A(_0427_),
    .B(_0428_));
 sg13g2_and4_1 _3621_ (.A(_0382_),
    .B(_0383_),
    .C(_0427_),
    .D(_0428_),
    .X(_0430_));
 sg13g2_xor2_1 _3622_ (.B(_0429_),
    .A(_0384_),
    .X(_0114_));
 sg13g2_o21ai_1 _3623_ (.B1(_0427_),
    .Y(_0431_),
    .A1(_0384_),
    .A2(_0429_));
 sg13g2_o21ai_1 _3624_ (.B1(_0422_),
    .Y(_0432_),
    .A1(_0351_),
    .A2(_0423_));
 sg13g2_o21ai_1 _3625_ (.B1(_0394_),
    .Y(_0433_),
    .A1(_0349_),
    .A2(_0395_));
 sg13g2_o21ai_1 _3626_ (.B1(_0417_),
    .Y(_0434_),
    .A1(_0396_),
    .A2(_0418_));
 sg13g2_nor2_1 _3627_ (.A(_0389_),
    .B(_0392_),
    .Y(_0435_));
 sg13g2_o21ai_1 _3628_ (.B1(_0401_),
    .Y(_0436_),
    .A1(_0398_),
    .A2(_0402_));
 sg13g2_nand2_1 _3629_ (.Y(_0437_),
    .A(net1039),
    .B(net1053));
 sg13g2_nand2_1 _3630_ (.Y(_0438_),
    .A(net1035),
    .B(net967));
 sg13g2_nand2_1 _3631_ (.Y(_0439_),
    .A(net1035),
    .B(net970));
 sg13g2_xor2_1 _3632_ (.B(_0439_),
    .A(_0388_),
    .X(_0440_));
 sg13g2_nand2b_1 _3633_ (.Y(_0441_),
    .B(_0440_),
    .A_N(_0437_));
 sg13g2_xnor2_1 _3634_ (.Y(_0442_),
    .A(_0437_),
    .B(_0440_));
 sg13g2_xnor2_1 _3635_ (.Y(_0443_),
    .A(_0436_),
    .B(_0442_));
 sg13g2_nor2_1 _3636_ (.A(_0435_),
    .B(_0443_),
    .Y(_0444_));
 sg13g2_xnor2_1 _3637_ (.Y(_0445_),
    .A(_0435_),
    .B(_0443_));
 sg13g2_o21ai_1 _3638_ (.B1(_0412_),
    .Y(_0446_),
    .A1(_0403_),
    .A2(_0413_));
 sg13g2_nand2_1 _3639_ (.Y(_0447_),
    .A(net1032),
    .B(net971));
 sg13g2_nand2_1 _3640_ (.Y(_0448_),
    .A(net975),
    .B(net1027));
 sg13g2_or2_1 _3641_ (.X(_0449_),
    .B(_0448_),
    .A(_0399_));
 sg13g2_and2_1 _3642_ (.A(_0399_),
    .B(_0448_),
    .X(_0450_));
 sg13g2_xnor2_1 _3643_ (.Y(_0451_),
    .A(_0399_),
    .B(_0448_));
 sg13g2_xnor2_1 _3644_ (.Y(_0452_),
    .A(_0447_),
    .B(_0451_));
 sg13g2_o21ai_1 _3645_ (.B1(_0407_),
    .Y(_0453_),
    .A1(_0405_),
    .A2(_0408_));
 sg13g2_nand2_1 _3646_ (.Y(_0454_),
    .A(net977),
    .B(net1059));
 sg13g2_and4_1 _3647_ (.A(net981),
    .B(net977),
    .C(net1025),
    .D(net1059),
    .X(_0455_));
 sg13g2_a22oi_1 _3648_ (.Y(_0456_),
    .B1(net1059),
    .B2(net980),
    .A2(net1025),
    .A1(net977));
 sg13g2_nor2_1 _3649_ (.A(_0455_),
    .B(_0456_),
    .Y(_0457_));
 sg13g2_nand2_1 _3650_ (.Y(_0458_),
    .A(_0453_),
    .B(_0457_));
 sg13g2_xnor2_1 _3651_ (.Y(_0459_),
    .A(_0453_),
    .B(_0457_));
 sg13g2_xor2_1 _3652_ (.B(_0459_),
    .A(_0452_),
    .X(_0460_));
 sg13g2_nand2_1 _3653_ (.Y(_0461_),
    .A(_0446_),
    .B(_0460_));
 sg13g2_xnor2_1 _3654_ (.Y(_0462_),
    .A(_0446_),
    .B(_0460_));
 sg13g2_xor2_1 _3655_ (.B(_0462_),
    .A(_0445_),
    .X(_0463_));
 sg13g2_nand2_1 _3656_ (.Y(_0464_),
    .A(_0434_),
    .B(_0463_));
 sg13g2_xnor2_1 _3657_ (.Y(_0465_),
    .A(_0434_),
    .B(_0463_));
 sg13g2_nand2b_1 _3658_ (.Y(_0466_),
    .B(_0433_),
    .A_N(_0465_));
 sg13g2_xnor2_1 _3659_ (.Y(_0467_),
    .A(_0433_),
    .B(_0465_));
 sg13g2_nor2_1 _3660_ (.A(_0432_),
    .B(_0467_),
    .Y(_0468_));
 sg13g2_nand2_1 _3661_ (.Y(_0469_),
    .A(_0432_),
    .B(_0467_));
 sg13g2_nor2b_2 _3662_ (.A(_0468_),
    .B_N(_0469_),
    .Y(_0470_));
 sg13g2_xor2_1 _3663_ (.B(_0470_),
    .A(_0431_),
    .X(_0115_));
 sg13g2_a21oi_1 _3664_ (.A1(_0436_),
    .A2(_0442_),
    .Y(_0471_),
    .B1(_0444_));
 sg13g2_o21ai_1 _3665_ (.B1(_0461_),
    .Y(_0472_),
    .A1(_0445_),
    .A2(_0462_));
 sg13g2_o21ai_1 _3666_ (.B1(_0441_),
    .Y(_0473_),
    .A1(_0388_),
    .A2(_0439_));
 sg13g2_o21ai_1 _3667_ (.B1(_0449_),
    .Y(_0474_),
    .A1(_0447_),
    .A2(_0450_));
 sg13g2_nand2_1 _3668_ (.Y(_0475_),
    .A(net1037),
    .B(net1053));
 sg13g2_nand2_1 _3669_ (.Y(_0476_),
    .A(net1032),
    .B(net966));
 sg13g2_nand2_1 _3670_ (.Y(_0477_),
    .A(net1032),
    .B(net969));
 sg13g2_or2_1 _3671_ (.X(_0478_),
    .B(_0476_),
    .A(_0439_));
 sg13g2_xnor2_1 _3672_ (.Y(_0479_),
    .A(_0438_),
    .B(_0477_));
 sg13g2_xor2_1 _3673_ (.B(_0479_),
    .A(_0475_),
    .X(_0480_));
 sg13g2_xnor2_1 _3674_ (.Y(_0481_),
    .A(_0474_),
    .B(_0480_));
 sg13g2_nor2b_1 _3675_ (.A(_0481_),
    .B_N(_0473_),
    .Y(_0482_));
 sg13g2_xor2_1 _3676_ (.B(_0481_),
    .A(_0473_),
    .X(_0483_));
 sg13g2_o21ai_1 _3677_ (.B1(_0458_),
    .Y(_0484_),
    .A1(_0452_),
    .A2(_0459_));
 sg13g2_a21oi_1 _3678_ (.A1(net981),
    .A2(net1025),
    .Y(_0485_),
    .B1(_0454_));
 sg13g2_nand2_1 _3679_ (.Y(_0486_),
    .A(net1031),
    .B(net971));
 sg13g2_nand2_1 _3680_ (.Y(_0487_),
    .A(net973),
    .B(net1026));
 sg13g2_and4_1 _3681_ (.A(net975),
    .B(net973),
    .C(net1027),
    .D(net1026),
    .X(_0488_));
 sg13g2_a22oi_1 _3682_ (.Y(_0489_),
    .B1(net1026),
    .B2(net975),
    .A2(net1027),
    .A1(net973));
 sg13g2_nor3_1 _3683_ (.A(_0486_),
    .B(_0488_),
    .C(_0489_),
    .Y(_0490_));
 sg13g2_o21ai_1 _3684_ (.B1(_0486_),
    .Y(_0491_),
    .A1(_0488_),
    .A2(_0489_));
 sg13g2_nor2b_1 _3685_ (.A(_0490_),
    .B_N(_0491_),
    .Y(_0492_));
 sg13g2_xnor2_1 _3686_ (.Y(_0493_),
    .A(_0485_),
    .B(_0492_));
 sg13g2_nand2b_1 _3687_ (.Y(_0494_),
    .B(_0484_),
    .A_N(_0493_));
 sg13g2_xor2_1 _3688_ (.B(_0493_),
    .A(_0484_),
    .X(_0495_));
 sg13g2_xor2_1 _3689_ (.B(_0495_),
    .A(_0483_),
    .X(_0496_));
 sg13g2_nand2_1 _3690_ (.Y(_0497_),
    .A(_0472_),
    .B(_0496_));
 sg13g2_xor2_1 _3691_ (.B(_0496_),
    .A(_0472_),
    .X(_0498_));
 sg13g2_nand2b_1 _3692_ (.Y(_0499_),
    .B(_0498_),
    .A_N(_0471_));
 sg13g2_xor2_1 _3693_ (.B(_0498_),
    .A(_0471_),
    .X(_0500_));
 sg13g2_a21oi_1 _3694_ (.A1(_0464_),
    .A2(_0466_),
    .Y(_0501_),
    .B1(_0500_));
 sg13g2_nand3_1 _3695_ (.B(_0466_),
    .C(_0500_),
    .A(_0464_),
    .Y(_0502_));
 sg13g2_nand2b_1 _3696_ (.Y(_0503_),
    .B(_0502_),
    .A_N(_0501_));
 sg13g2_a21oi_1 _3697_ (.A1(_0427_),
    .A2(_0469_),
    .Y(_0504_),
    .B1(_0468_));
 sg13g2_a21oi_2 _3698_ (.B1(_0504_),
    .Y(_0505_),
    .A2(_0470_),
    .A1(_0430_));
 sg13g2_nor2_1 _3699_ (.A(_0503_),
    .B(_0505_),
    .Y(_0506_));
 sg13g2_xor2_1 _3700_ (.B(_0505_),
    .A(_0503_),
    .X(_0106_));
 sg13g2_a21o_1 _3701_ (.A2(_0480_),
    .A1(_0474_),
    .B1(_0482_),
    .X(_0507_));
 sg13g2_o21ai_1 _3702_ (.B1(_0494_),
    .Y(_0508_),
    .A1(_0483_),
    .A2(_0495_));
 sg13g2_a21o_1 _3703_ (.A2(_0492_),
    .A1(_0485_),
    .B1(_0455_),
    .X(_0509_));
 sg13g2_nand2_1 _3704_ (.Y(_0510_),
    .A(net971),
    .B(net1027));
 sg13g2_nand2_1 _3705_ (.Y(_0511_),
    .A(net975),
    .B(net1058));
 sg13g2_or2_1 _3706_ (.X(_0512_),
    .B(_0511_),
    .A(_0487_));
 sg13g2_xnor2_1 _3707_ (.Y(_0513_),
    .A(_0487_),
    .B(_0511_));
 sg13g2_xor2_1 _3708_ (.B(_0513_),
    .A(_0510_),
    .X(_0514_));
 sg13g2_and2_1 _3709_ (.A(_0509_),
    .B(_0514_),
    .X(_0515_));
 sg13g2_or2_1 _3710_ (.X(_0516_),
    .B(_0514_),
    .A(_0509_));
 sg13g2_xnor2_1 _3711_ (.Y(_0517_),
    .A(_0509_),
    .B(_0514_));
 sg13g2_o21ai_1 _3712_ (.B1(_0478_),
    .Y(_0518_),
    .A1(_0475_),
    .A2(_0479_));
 sg13g2_or2_1 _3713_ (.X(_0519_),
    .B(_0490_),
    .A(_0488_));
 sg13g2_nand2_1 _3714_ (.Y(_0520_),
    .A(net1035),
    .B(net1053));
 sg13g2_nand2_1 _3715_ (.Y(_0521_),
    .A(net1031),
    .B(net969));
 sg13g2_or2_1 _3716_ (.X(_0522_),
    .B(_0521_),
    .A(_0476_));
 sg13g2_xnor2_1 _3717_ (.Y(_0523_),
    .A(_0476_),
    .B(_0521_));
 sg13g2_xor2_1 _3718_ (.B(_0523_),
    .A(_0520_),
    .X(_0524_));
 sg13g2_xnor2_1 _3719_ (.Y(_0525_),
    .A(_0519_),
    .B(_0524_));
 sg13g2_nor2b_1 _3720_ (.A(_0525_),
    .B_N(_0518_),
    .Y(_0526_));
 sg13g2_xnor2_1 _3721_ (.Y(_0527_),
    .A(_0518_),
    .B(_0525_));
 sg13g2_xnor2_1 _3722_ (.Y(_0528_),
    .A(_0517_),
    .B(_0527_));
 sg13g2_xnor2_1 _3723_ (.Y(_0529_),
    .A(_0508_),
    .B(_0528_));
 sg13g2_nor2b_1 _3724_ (.A(_0529_),
    .B_N(_0507_),
    .Y(_0530_));
 sg13g2_xor2_1 _3725_ (.B(_0529_),
    .A(_0507_),
    .X(_0531_));
 sg13g2_nand3_1 _3726_ (.B(_0499_),
    .C(_0531_),
    .A(_0497_),
    .Y(_0532_));
 sg13g2_inv_1 _3727_ (.Y(_0533_),
    .A(_0532_));
 sg13g2_a21oi_1 _3728_ (.A1(_0497_),
    .A2(_0499_),
    .Y(_0534_),
    .B1(_0531_));
 sg13g2_nor2_1 _3729_ (.A(_0533_),
    .B(_0534_),
    .Y(_0535_));
 sg13g2_nor2_1 _3730_ (.A(_0501_),
    .B(_0506_),
    .Y(_0536_));
 sg13g2_xnor2_1 _3731_ (.Y(_0107_),
    .A(_0535_),
    .B(_0536_));
 sg13g2_a21o_1 _3732_ (.A2(_0524_),
    .A1(_0519_),
    .B1(_0526_),
    .X(_0537_));
 sg13g2_a22oi_1 _3733_ (.Y(_0538_),
    .B1(net1058),
    .B2(net973),
    .A2(net1026),
    .A1(net971));
 sg13g2_nand2_1 _3734_ (.Y(_0539_),
    .A(net971),
    .B(net1058));
 sg13g2_or2_1 _3735_ (.X(_0540_),
    .B(_0539_),
    .A(_0487_));
 sg13g2_nand2b_1 _3736_ (.Y(_0541_),
    .B(_0540_),
    .A_N(_0538_));
 sg13g2_o21ai_1 _3737_ (.B1(_0522_),
    .Y(_0542_),
    .A1(_0520_),
    .A2(_0523_));
 sg13g2_o21ai_1 _3738_ (.B1(_0512_),
    .Y(_0543_),
    .A1(_0510_),
    .A2(_0513_));
 sg13g2_nand2_1 _3739_ (.Y(_0544_),
    .A(net1032),
    .B(net1053));
 sg13g2_nand2_1 _3740_ (.Y(_0545_),
    .A(net1027),
    .B(net966));
 sg13g2_and4_1 _3741_ (.A(net1031),
    .B(net1027),
    .C(net969),
    .D(net966),
    .X(_0546_));
 sg13g2_or2_1 _3742_ (.X(_0547_),
    .B(_0545_),
    .A(_0521_));
 sg13g2_a22oi_1 _3743_ (.Y(_0548_),
    .B1(net966),
    .B2(net1031),
    .A2(net969),
    .A1(net1027));
 sg13g2_nor2_1 _3744_ (.A(_0546_),
    .B(_0548_),
    .Y(_0549_));
 sg13g2_xnor2_1 _3745_ (.Y(_0550_),
    .A(_0544_),
    .B(_0549_));
 sg13g2_xnor2_1 _3746_ (.Y(_0551_),
    .A(_0543_),
    .B(_0550_));
 sg13g2_nor2b_1 _3747_ (.A(_0551_),
    .B_N(_0542_),
    .Y(_0552_));
 sg13g2_xor2_1 _3748_ (.B(_0551_),
    .A(_0542_),
    .X(_0553_));
 sg13g2_or2_1 _3749_ (.X(_0554_),
    .B(_0553_),
    .A(_0541_));
 sg13g2_xor2_1 _3750_ (.B(_0553_),
    .A(_0541_),
    .X(_0555_));
 sg13g2_a21oi_1 _3751_ (.A1(_0516_),
    .A2(_0527_),
    .Y(_0556_),
    .B1(_0515_));
 sg13g2_nor2b_1 _3752_ (.A(_0556_),
    .B_N(_0555_),
    .Y(_0557_));
 sg13g2_xor2_1 _3753_ (.B(_0556_),
    .A(_0555_),
    .X(_0558_));
 sg13g2_nor2b_1 _3754_ (.A(_0558_),
    .B_N(_0537_),
    .Y(_0559_));
 sg13g2_xor2_1 _3755_ (.B(_0558_),
    .A(_0537_),
    .X(_0560_));
 sg13g2_a21oi_1 _3756_ (.A1(_0508_),
    .A2(_0528_),
    .Y(_0561_),
    .B1(_0530_));
 sg13g2_nor2_1 _3757_ (.A(_0560_),
    .B(_0561_),
    .Y(_0562_));
 sg13g2_xor2_1 _3758_ (.B(_0561_),
    .A(_0560_),
    .X(_0563_));
 sg13g2_a21oi_1 _3759_ (.A1(_0501_),
    .A2(_0532_),
    .Y(_0564_),
    .B1(_0534_));
 sg13g2_a21oi_1 _3760_ (.A1(_0502_),
    .A2(_0532_),
    .Y(_0565_),
    .B1(_0534_));
 sg13g2_a21oi_2 _3761_ (.B1(_0565_),
    .Y(_0566_),
    .A2(_0564_),
    .A1(_0505_));
 sg13g2_xor2_1 _3762_ (.B(_0566_),
    .A(_0563_),
    .X(_0108_));
 sg13g2_a21o_1 _3763_ (.A2(_0550_),
    .A1(_0543_),
    .B1(_0552_),
    .X(_0567_));
 sg13g2_o21ai_1 _3764_ (.B1(_0547_),
    .Y(_0568_),
    .A1(_0544_),
    .A2(_0548_));
 sg13g2_nand2_1 _3765_ (.Y(_0569_),
    .A(net1031),
    .B(\DP_2.matrix[8] ));
 sg13g2_nand2_1 _3766_ (.Y(_0570_),
    .A(net1026),
    .B(net966));
 sg13g2_nand2_1 _3767_ (.Y(_0571_),
    .A(net969),
    .B(net1026));
 sg13g2_xor2_1 _3768_ (.B(_0571_),
    .A(_0545_),
    .X(_0572_));
 sg13g2_nand2b_1 _3769_ (.Y(_0573_),
    .B(_0572_),
    .A_N(_0569_));
 sg13g2_xnor2_1 _3770_ (.Y(_0574_),
    .A(_0569_),
    .B(_0572_));
 sg13g2_nor2b_1 _3771_ (.A(_0540_),
    .B_N(_0574_),
    .Y(_0575_));
 sg13g2_xnor2_1 _3772_ (.Y(_0576_),
    .A(_0540_),
    .B(_0574_));
 sg13g2_xnor2_1 _3773_ (.Y(_0577_),
    .A(_0568_),
    .B(_0576_));
 sg13g2_nor2_1 _3774_ (.A(_0539_),
    .B(_0577_),
    .Y(_0578_));
 sg13g2_xnor2_1 _3775_ (.Y(_0579_),
    .A(_0539_),
    .B(_0577_));
 sg13g2_nor2_1 _3776_ (.A(_0554_),
    .B(_0579_),
    .Y(_0580_));
 sg13g2_xor2_1 _3777_ (.B(_0579_),
    .A(_0554_),
    .X(_0581_));
 sg13g2_xor2_1 _3778_ (.B(_0581_),
    .A(_0567_),
    .X(_0582_));
 sg13g2_o21ai_1 _3779_ (.B1(_0582_),
    .Y(_0583_),
    .A1(_0557_),
    .A2(_0559_));
 sg13g2_or3_1 _3780_ (.A(_0557_),
    .B(_0559_),
    .C(_0582_),
    .X(_0584_));
 sg13g2_and2_1 _3781_ (.A(_0583_),
    .B(_0584_),
    .X(_0585_));
 sg13g2_a21oi_1 _3782_ (.A1(_0563_),
    .A2(_0566_),
    .Y(_0586_),
    .B1(_0562_));
 sg13g2_xnor2_1 _3783_ (.Y(_0109_),
    .A(_0585_),
    .B(_0586_));
 sg13g2_nand2_1 _3784_ (.Y(_0587_),
    .A(_0563_),
    .B(_0585_));
 sg13g2_inv_1 _3785_ (.Y(_0588_),
    .A(_0587_));
 sg13g2_o21ai_1 _3786_ (.B1(_0583_),
    .Y(_0589_),
    .A1(_0560_),
    .A2(_0561_));
 sg13g2_a22oi_1 _3787_ (.Y(_0590_),
    .B1(_0589_),
    .B2(_0584_),
    .A2(_0588_),
    .A1(_0566_));
 sg13g2_a21oi_1 _3788_ (.A1(_0567_),
    .A2(_0581_),
    .Y(_0591_),
    .B1(_0580_));
 sg13g2_a21o_1 _3789_ (.A2(_0576_),
    .A1(_0568_),
    .B1(_0575_),
    .X(_0592_));
 sg13g2_o21ai_1 _3790_ (.B1(_0573_),
    .Y(_0593_),
    .A1(_0545_),
    .A2(_0571_));
 sg13g2_nand2_1 _3791_ (.Y(_0594_),
    .A(net1027),
    .B(\DP_2.matrix[8] ));
 sg13g2_nand2_1 _3792_ (.Y(_0595_),
    .A(net966),
    .B(net1058));
 sg13g2_nand2_1 _3793_ (.Y(_0596_),
    .A(net969),
    .B(net1058));
 sg13g2_xor2_1 _3794_ (.B(_0596_),
    .A(_0570_),
    .X(_0597_));
 sg13g2_nand2b_1 _3795_ (.Y(_0598_),
    .B(_0597_),
    .A_N(_0594_));
 sg13g2_xnor2_1 _3796_ (.Y(_0599_),
    .A(_0594_),
    .B(_0597_));
 sg13g2_nand2_1 _3797_ (.Y(_0600_),
    .A(_0593_),
    .B(_0599_));
 sg13g2_xor2_1 _3798_ (.B(_0599_),
    .A(_0593_),
    .X(_0601_));
 sg13g2_xnor2_1 _3799_ (.Y(_0602_),
    .A(_0578_),
    .B(_0601_));
 sg13g2_nor2b_1 _3800_ (.A(_0602_),
    .B_N(_0592_),
    .Y(_0603_));
 sg13g2_xor2_1 _3801_ (.B(_0602_),
    .A(_0592_),
    .X(_0604_));
 sg13g2_or2_1 _3802_ (.X(_0605_),
    .B(_0604_),
    .A(_0591_));
 sg13g2_xor2_1 _3803_ (.B(_0604_),
    .A(_0591_),
    .X(_0606_));
 sg13g2_inv_1 _3804_ (.Y(_0607_),
    .A(_0606_));
 sg13g2_xnor2_1 _3805_ (.Y(_0110_),
    .A(_0590_),
    .B(_0606_));
 sg13g2_o21ai_1 _3806_ (.B1(_0605_),
    .Y(_0608_),
    .A1(_0590_),
    .A2(_0607_));
 sg13g2_a21oi_1 _3807_ (.A1(_0578_),
    .A2(_0601_),
    .Y(_0609_),
    .B1(_0603_));
 sg13g2_o21ai_1 _3808_ (.B1(_0598_),
    .Y(_0610_),
    .A1(_0570_),
    .A2(_0596_));
 sg13g2_nand2_1 _3809_ (.Y(_0611_),
    .A(net1026),
    .B(net1053));
 sg13g2_xor2_1 _3810_ (.B(_0611_),
    .A(_0595_),
    .X(_0612_));
 sg13g2_xnor2_1 _3811_ (.Y(_0613_),
    .A(_0610_),
    .B(_0612_));
 sg13g2_xnor2_1 _3812_ (.Y(_0614_),
    .A(_0600_),
    .B(_0613_));
 sg13g2_xnor2_1 _3813_ (.Y(_0615_),
    .A(_0609_),
    .B(_0614_));
 sg13g2_xnor2_1 _3814_ (.Y(_0111_),
    .A(_0608_),
    .B(_0615_));
 sg13g2_and2_1 _3815_ (.A(net1023),
    .B(net964),
    .X(_0074_));
 sg13g2_and3_2 _3816_ (.X(_0616_),
    .A(net1021),
    .B(net960),
    .C(_0074_));
 sg13g2_a22oi_1 _3817_ (.Y(_0617_),
    .B1(net960),
    .B2(net1023),
    .A2(net1021),
    .A1(net964));
 sg13g2_nor2_1 _3818_ (.A(_0616_),
    .B(net449),
    .Y(_0075_));
 sg13g2_nand2_1 _3819_ (.Y(_0618_),
    .A(net1023),
    .B(net956));
 sg13g2_and4_1 _3820_ (.A(net962),
    .B(net1021),
    .C(net958),
    .D(net1018),
    .X(_0619_));
 sg13g2_a22oi_1 _3821_ (.Y(_0620_),
    .B1(net1018),
    .B2(net962),
    .A2(net958),
    .A1(net1021));
 sg13g2_nor3_1 _3822_ (.A(_0618_),
    .B(_0619_),
    .C(_0620_),
    .Y(_0621_));
 sg13g2_o21ai_1 _3823_ (.B1(_0618_),
    .Y(_0622_),
    .A1(_0619_),
    .A2(_0620_));
 sg13g2_nor2b_1 _3824_ (.A(_0621_),
    .B_N(_0622_),
    .Y(_0623_));
 sg13g2_nand2_1 _3825_ (.Y(_0624_),
    .A(_0616_),
    .B(_0623_));
 sg13g2_xor2_1 _3826_ (.B(_0623_),
    .A(_0616_),
    .X(_0076_));
 sg13g2_nand2_1 _3827_ (.Y(_0625_),
    .A(net1023),
    .B(net954));
 sg13g2_or2_1 _3828_ (.X(_0626_),
    .B(_0621_),
    .A(_0619_));
 sg13g2_nand2_1 _3829_ (.Y(_0627_),
    .A(net1022),
    .B(net957));
 sg13g2_and4_1 _3830_ (.A(net962),
    .B(net958),
    .C(net1018),
    .D(net1016),
    .X(_0628_));
 sg13g2_nand4_1 _3831_ (.B(net961),
    .C(net1018),
    .A(net965),
    .Y(_0629_),
    .D(net1016));
 sg13g2_a22oi_1 _3832_ (.Y(_0630_),
    .B1(net1016),
    .B2(net962),
    .A2(net1018),
    .A1(net959));
 sg13g2_nor3_1 _3833_ (.A(_0627_),
    .B(_0628_),
    .C(_0630_),
    .Y(_0631_));
 sg13g2_o21ai_1 _3834_ (.B1(_0627_),
    .Y(_0632_),
    .A1(_0628_),
    .A2(_0630_));
 sg13g2_nor2b_1 _3835_ (.A(_0631_),
    .B_N(_0632_),
    .Y(_0633_));
 sg13g2_nand2_1 _3836_ (.Y(_0634_),
    .A(_0626_),
    .B(_0633_));
 sg13g2_xnor2_1 _3837_ (.Y(_0635_),
    .A(_0626_),
    .B(_0633_));
 sg13g2_xor2_1 _3838_ (.B(_0635_),
    .A(_0625_),
    .X(_0636_));
 sg13g2_nand2b_1 _3839_ (.Y(_0637_),
    .B(_0636_),
    .A_N(_0624_));
 sg13g2_xnor2_1 _3840_ (.Y(_0077_),
    .A(_0624_),
    .B(_0636_));
 sg13g2_a22oi_1 _3841_ (.Y(_0638_),
    .B1(net953),
    .B2(net1024),
    .A2(net955),
    .A1(net1022));
 sg13g2_nand2_1 _3842_ (.Y(_0639_),
    .A(net1022),
    .B(net953));
 sg13g2_and4_1 _3843_ (.A(net1024),
    .B(\DP_1.matrix[37] ),
    .C(net955),
    .D(net953),
    .X(_0640_));
 sg13g2_nor2_1 _3844_ (.A(_0638_),
    .B(_0640_),
    .Y(_0641_));
 sg13g2_inv_1 _3845_ (.Y(_0642_),
    .A(_0641_));
 sg13g2_o21ai_1 _3846_ (.B1(_0629_),
    .Y(_0643_),
    .A1(_0627_),
    .A2(_0630_));
 sg13g2_nand2_1 _3847_ (.Y(_0644_),
    .A(net1018),
    .B(net957));
 sg13g2_and4_1 _3848_ (.A(net965),
    .B(net961),
    .C(net1016),
    .D(net1013),
    .X(_0645_));
 sg13g2_nand4_1 _3849_ (.B(net961),
    .C(net1017),
    .A(net965),
    .Y(_0646_),
    .D(net1014));
 sg13g2_a22oi_1 _3850_ (.Y(_0647_),
    .B1(net1014),
    .B2(net965),
    .A2(net1017),
    .A1(net961));
 sg13g2_or3_1 _3851_ (.A(_0644_),
    .B(_0645_),
    .C(_0647_),
    .X(_0648_));
 sg13g2_o21ai_1 _3852_ (.B1(_0644_),
    .Y(_0649_),
    .A1(_0645_),
    .A2(_0647_));
 sg13g2_nand3_1 _3853_ (.B(_0648_),
    .C(_0649_),
    .A(_0643_),
    .Y(_0650_));
 sg13g2_a21oi_1 _3854_ (.A1(_0648_),
    .A2(_0649_),
    .Y(_0651_),
    .B1(_0643_));
 sg13g2_a21o_1 _3855_ (.A2(_0649_),
    .A1(_0648_),
    .B1(_0643_),
    .X(_0652_));
 sg13g2_nand2_1 _3856_ (.Y(_0653_),
    .A(_0650_),
    .B(_0652_));
 sg13g2_xnor2_1 _3857_ (.Y(_0654_),
    .A(_0642_),
    .B(_0653_));
 sg13g2_o21ai_1 _3858_ (.B1(_0634_),
    .Y(_0655_),
    .A1(_0625_),
    .A2(_0635_));
 sg13g2_nor2b_2 _3859_ (.A(_0654_),
    .B_N(_0655_),
    .Y(_0656_));
 sg13g2_xor2_1 _3860_ (.B(_0655_),
    .A(_0654_),
    .X(_0657_));
 sg13g2_or2_1 _3861_ (.X(_0658_),
    .B(_0657_),
    .A(_0637_));
 sg13g2_xor2_1 _3862_ (.B(_0657_),
    .A(_0637_),
    .X(_0078_));
 sg13g2_o21ai_1 _3863_ (.B1(_0650_),
    .Y(_0659_),
    .A1(_0642_),
    .A2(_0651_));
 sg13g2_nand2_1 _3864_ (.Y(_0660_),
    .A(net1023),
    .B(net951));
 sg13g2_nand2_1 _3865_ (.Y(_0661_),
    .A(net1019),
    .B(net952));
 sg13g2_nand2_1 _3866_ (.Y(_0662_),
    .A(net1020),
    .B(net955));
 sg13g2_xor2_1 _3867_ (.B(_0662_),
    .A(_0639_),
    .X(_0663_));
 sg13g2_nand2b_1 _3868_ (.Y(_0664_),
    .B(_0663_),
    .A_N(_0660_));
 sg13g2_xor2_1 _3869_ (.B(_0663_),
    .A(_0660_),
    .X(_0665_));
 sg13g2_o21ai_1 _3870_ (.B1(_0646_),
    .Y(_0666_),
    .A1(_0644_),
    .A2(_0647_));
 sg13g2_nand2_1 _3871_ (.Y(_0667_),
    .A(net956),
    .B(net1016));
 sg13g2_and4_1 _3872_ (.A(net962),
    .B(net958),
    .C(net1013),
    .D(net1010),
    .X(_0668_));
 sg13g2_nand4_1 _3873_ (.B(net958),
    .C(net1014),
    .A(net965),
    .Y(_0669_),
    .D(net1011));
 sg13g2_a22oi_1 _3874_ (.Y(_0670_),
    .B1(net1011),
    .B2(net962),
    .A2(net1014),
    .A1(net958));
 sg13g2_or3_1 _3875_ (.A(_0667_),
    .B(_0668_),
    .C(_0670_),
    .X(_0671_));
 sg13g2_o21ai_1 _3876_ (.B1(_0667_),
    .Y(_0672_),
    .A1(_0668_),
    .A2(_0670_));
 sg13g2_and3_1 _3877_ (.X(_0673_),
    .A(_0666_),
    .B(_0671_),
    .C(_0672_));
 sg13g2_nand3_1 _3878_ (.B(_0671_),
    .C(_0672_),
    .A(_0666_),
    .Y(_0674_));
 sg13g2_a21oi_1 _3879_ (.A1(_0671_),
    .A2(_0672_),
    .Y(_0675_),
    .B1(_0666_));
 sg13g2_or3_1 _3880_ (.A(_0665_),
    .B(_0673_),
    .C(_0675_),
    .X(_0676_));
 sg13g2_o21ai_1 _3881_ (.B1(_0665_),
    .Y(_0677_),
    .A1(_0673_),
    .A2(_0675_));
 sg13g2_nand3_1 _3882_ (.B(_0676_),
    .C(_0677_),
    .A(_0659_),
    .Y(_0678_));
 sg13g2_a21o_1 _3883_ (.A2(_0677_),
    .A1(_0676_),
    .B1(_0659_),
    .X(_0679_));
 sg13g2_nand3_1 _3884_ (.B(_0678_),
    .C(_0679_),
    .A(_0640_),
    .Y(_0680_));
 sg13g2_a21o_1 _3885_ (.A2(_0679_),
    .A1(_0678_),
    .B1(_0640_),
    .X(_0681_));
 sg13g2_and2_1 _3886_ (.A(_0680_),
    .B(_0681_),
    .X(_0682_));
 sg13g2_nand3_1 _3887_ (.B(_0680_),
    .C(_0681_),
    .A(_0656_),
    .Y(_0683_));
 sg13g2_a21oi_1 _3888_ (.A1(_0680_),
    .A2(_0681_),
    .Y(_0684_),
    .B1(_0656_));
 sg13g2_xor2_1 _3889_ (.B(_0682_),
    .A(_0656_),
    .X(_0685_));
 sg13g2_xnor2_1 _3890_ (.Y(_0116_),
    .A(_0658_),
    .B(_0685_));
 sg13g2_nand2_1 _3891_ (.Y(_0686_),
    .A(_0678_),
    .B(_0680_));
 sg13g2_o21ai_1 _3892_ (.B1(_0664_),
    .Y(_0687_),
    .A1(_0639_),
    .A2(_0662_));
 sg13g2_nand2_1 _3893_ (.Y(_0688_),
    .A(net1024),
    .B(net950));
 sg13g2_nand2b_1 _3894_ (.Y(_0689_),
    .B(_0687_),
    .A_N(_0688_));
 sg13g2_xor2_1 _3895_ (.B(_0688_),
    .A(_0687_),
    .X(_0690_));
 sg13g2_o21ai_1 _3896_ (.B1(_0674_),
    .Y(_0691_),
    .A1(_0665_),
    .A2(_0675_));
 sg13g2_nand2_1 _3897_ (.Y(_0692_),
    .A(net1021),
    .B(net951));
 sg13g2_nand2_1 _3898_ (.Y(_0693_),
    .A(net1017),
    .B(net952));
 sg13g2_nand2_1 _3899_ (.Y(_0694_),
    .A(net1017),
    .B(net954));
 sg13g2_xor2_1 _3900_ (.B(_0694_),
    .A(_0661_),
    .X(_0695_));
 sg13g2_nand2b_1 _3901_ (.Y(_0696_),
    .B(_0695_),
    .A_N(_0692_));
 sg13g2_xnor2_1 _3902_ (.Y(_0697_),
    .A(_0692_),
    .B(_0695_));
 sg13g2_o21ai_1 _3903_ (.B1(_0669_),
    .Y(_0698_),
    .A1(_0667_),
    .A2(_0670_));
 sg13g2_nand2_1 _3904_ (.Y(_0699_),
    .A(net956),
    .B(net1013));
 sg13g2_and4_1 _3905_ (.A(net962),
    .B(net959),
    .C(net1011),
    .D(net1009),
    .X(_0700_));
 sg13g2_nand4_1 _3906_ (.B(net958),
    .C(net1011),
    .A(net965),
    .Y(_0701_),
    .D(net1009));
 sg13g2_a22oi_1 _3907_ (.Y(_0702_),
    .B1(net1009),
    .B2(\DP_2.matrix[36] ),
    .A2(net1011),
    .A1(net958));
 sg13g2_or3_1 _3908_ (.A(_0699_),
    .B(_0700_),
    .C(_0702_),
    .X(_0703_));
 sg13g2_o21ai_1 _3909_ (.B1(_0699_),
    .Y(_0704_),
    .A1(_0700_),
    .A2(_0702_));
 sg13g2_and3_1 _3910_ (.X(_0705_),
    .A(_0698_),
    .B(_0703_),
    .C(_0704_));
 sg13g2_nand3_1 _3911_ (.B(_0703_),
    .C(_0704_),
    .A(_0698_),
    .Y(_0706_));
 sg13g2_a21o_1 _3912_ (.A2(_0704_),
    .A1(_0703_),
    .B1(_0698_),
    .X(_0707_));
 sg13g2_nand3_1 _3913_ (.B(_0706_),
    .C(_0707_),
    .A(_0697_),
    .Y(_0708_));
 sg13g2_a21o_1 _3914_ (.A2(_0707_),
    .A1(_0706_),
    .B1(_0697_),
    .X(_0709_));
 sg13g2_nand3_1 _3915_ (.B(_0708_),
    .C(_0709_),
    .A(_0691_),
    .Y(_0710_));
 sg13g2_a21oi_1 _3916_ (.A1(_0708_),
    .A2(_0709_),
    .Y(_0711_),
    .B1(_0691_));
 sg13g2_a21o_1 _3917_ (.A2(_0709_),
    .A1(_0708_),
    .B1(_0691_),
    .X(_0712_));
 sg13g2_nand2_1 _3918_ (.Y(_0713_),
    .A(_0710_),
    .B(_0712_));
 sg13g2_xnor2_1 _3919_ (.Y(_0714_),
    .A(_0690_),
    .B(_0713_));
 sg13g2_nor2b_1 _3920_ (.A(_0714_),
    .B_N(_0686_),
    .Y(_0715_));
 sg13g2_xnor2_1 _3921_ (.Y(_0716_),
    .A(_0686_),
    .B(_0714_));
 sg13g2_o21ai_1 _3922_ (.B1(_0683_),
    .Y(_0717_),
    .A1(_0658_),
    .A2(_0684_));
 sg13g2_xor2_1 _3923_ (.B(_0717_),
    .A(_0716_),
    .X(_0123_));
 sg13g2_o21ai_1 _3924_ (.B1(_0710_),
    .Y(_0718_),
    .A1(_0690_),
    .A2(_0711_));
 sg13g2_o21ai_1 _3925_ (.B1(_0696_),
    .Y(_0719_),
    .A1(_0661_),
    .A2(_0694_));
 sg13g2_a22oi_1 _3926_ (.Y(_0720_),
    .B1(net948),
    .B2(net1024),
    .A2(net950),
    .A1(net1022));
 sg13g2_nand4_1 _3927_ (.B(net1022),
    .C(net950),
    .A(net1024),
    .Y(_0721_),
    .D(net948));
 sg13g2_nor2b_1 _3928_ (.A(_0720_),
    .B_N(_0721_),
    .Y(_0722_));
 sg13g2_nand2_1 _3929_ (.Y(_0723_),
    .A(_0719_),
    .B(_0722_));
 sg13g2_xnor2_1 _3930_ (.Y(_0724_),
    .A(_0719_),
    .B(_0722_));
 sg13g2_a21o_1 _3931_ (.A2(_0707_),
    .A1(_0697_),
    .B1(_0705_),
    .X(_0725_));
 sg13g2_nand2_1 _3932_ (.Y(_0726_),
    .A(net1019),
    .B(\DP_2.matrix[41] ));
 sg13g2_nand2_1 _3933_ (.Y(_0727_),
    .A(net1014),
    .B(net952));
 sg13g2_nand2_1 _3934_ (.Y(_0728_),
    .A(net954),
    .B(net1013));
 sg13g2_or2_1 _3935_ (.X(_0729_),
    .B(_0727_),
    .A(_0694_));
 sg13g2_and2_1 _3936_ (.A(_0693_),
    .B(_0728_),
    .X(_0730_));
 sg13g2_xnor2_1 _3937_ (.Y(_0731_),
    .A(_0693_),
    .B(_0728_));
 sg13g2_xnor2_1 _3938_ (.Y(_0732_),
    .A(_0726_),
    .B(_0731_));
 sg13g2_o21ai_1 _3939_ (.B1(_0701_),
    .Y(_0733_),
    .A1(_0699_),
    .A2(_0702_));
 sg13g2_nand2_1 _3940_ (.Y(_0734_),
    .A(net956),
    .B(net1010));
 sg13g2_and4_1 _3941_ (.A(net962),
    .B(net959),
    .C(net1009),
    .D(net1005),
    .X(_0735_));
 sg13g2_nand4_1 _3942_ (.B(net959),
    .C(net1009),
    .A(net963),
    .Y(_0736_),
    .D(net1005));
 sg13g2_a22oi_1 _3943_ (.Y(_0737_),
    .B1(net1005),
    .B2(net963),
    .A2(net1009),
    .A1(net960));
 sg13g2_or3_1 _3944_ (.A(_0734_),
    .B(_0735_),
    .C(_0737_),
    .X(_0738_));
 sg13g2_o21ai_1 _3945_ (.B1(_0734_),
    .Y(_0739_),
    .A1(_0735_),
    .A2(_0737_));
 sg13g2_and3_1 _3946_ (.X(_0740_),
    .A(_0733_),
    .B(_0738_),
    .C(_0739_));
 sg13g2_nand3_1 _3947_ (.B(_0738_),
    .C(_0739_),
    .A(_0733_),
    .Y(_0741_));
 sg13g2_a21oi_1 _3948_ (.A1(_0738_),
    .A2(_0739_),
    .Y(_0742_),
    .B1(_0733_));
 sg13g2_or3_1 _3949_ (.A(_0732_),
    .B(_0740_),
    .C(_0742_),
    .X(_0743_));
 sg13g2_o21ai_1 _3950_ (.B1(_0732_),
    .Y(_0744_),
    .A1(_0740_),
    .A2(_0742_));
 sg13g2_and3_1 _3951_ (.X(_0745_),
    .A(_0725_),
    .B(_0743_),
    .C(_0744_));
 sg13g2_nand3_1 _3952_ (.B(_0743_),
    .C(_0744_),
    .A(_0725_),
    .Y(_0746_));
 sg13g2_a21oi_1 _3953_ (.A1(_0743_),
    .A2(_0744_),
    .Y(_0747_),
    .B1(_0725_));
 sg13g2_or3_1 _3954_ (.A(_0724_),
    .B(_0745_),
    .C(_0747_),
    .X(_0748_));
 sg13g2_o21ai_1 _3955_ (.B1(_0724_),
    .Y(_0749_),
    .A1(_0745_),
    .A2(_0747_));
 sg13g2_nand3_1 _3956_ (.B(_0748_),
    .C(_0749_),
    .A(_0718_),
    .Y(_0750_));
 sg13g2_a21oi_1 _3957_ (.A1(_0748_),
    .A2(_0749_),
    .Y(_0751_),
    .B1(_0718_));
 sg13g2_a21o_1 _3958_ (.A2(_0749_),
    .A1(_0748_),
    .B1(_0718_),
    .X(_0752_));
 sg13g2_nand2_1 _3959_ (.Y(_0753_),
    .A(_0750_),
    .B(_0752_));
 sg13g2_xor2_1 _3960_ (.B(_0753_),
    .A(_0689_),
    .X(_0754_));
 sg13g2_a21o_2 _3961_ (.A2(_0717_),
    .A1(_0716_),
    .B1(_0715_),
    .X(_0755_));
 sg13g2_nand2_1 _3962_ (.Y(_0756_),
    .A(_0754_),
    .B(_0755_));
 sg13g2_xor2_1 _3963_ (.B(_0755_),
    .A(_0754_),
    .X(_0124_));
 sg13g2_o21ai_1 _3964_ (.B1(_0746_),
    .Y(_0757_),
    .A1(_0724_),
    .A2(_0747_));
 sg13g2_o21ai_1 _3965_ (.B1(_0729_),
    .Y(_0758_),
    .A1(_0726_),
    .A2(_0730_));
 sg13g2_nand2_1 _3966_ (.Y(_0759_),
    .A(net1023),
    .B(\DP_2.matrix[44] ));
 sg13g2_nand2_1 _3967_ (.Y(_0760_),
    .A(net1019),
    .B(net948));
 sg13g2_and4_1 _3968_ (.A(net1021),
    .B(net1019),
    .C(net949),
    .D(net947),
    .X(_0761_));
 sg13g2_a22oi_1 _3969_ (.Y(_0762_),
    .B1(net947),
    .B2(net1022),
    .A2(net949),
    .A1(net1019));
 sg13g2_or2_1 _3970_ (.X(_0763_),
    .B(_0762_),
    .A(_0761_));
 sg13g2_nor2_1 _3971_ (.A(_0759_),
    .B(_0763_),
    .Y(_0764_));
 sg13g2_xor2_1 _3972_ (.B(_0763_),
    .A(_0759_),
    .X(_0765_));
 sg13g2_nand2_1 _3973_ (.Y(_0766_),
    .A(_0758_),
    .B(_0765_));
 sg13g2_xnor2_1 _3974_ (.Y(_0767_),
    .A(_0758_),
    .B(_0765_));
 sg13g2_xnor2_1 _3975_ (.Y(_0768_),
    .A(_0721_),
    .B(_0767_));
 sg13g2_o21ai_1 _3976_ (.B1(_0741_),
    .Y(_0769_),
    .A1(_0732_),
    .A2(_0742_));
 sg13g2_nand2_1 _3977_ (.Y(_0770_),
    .A(net1017),
    .B(\DP_2.matrix[41] ));
 sg13g2_nand2_2 _3978_ (.Y(_0771_),
    .A(net952),
    .B(net1010));
 sg13g2_nand2_1 _3979_ (.Y(_0772_),
    .A(net954),
    .B(net1010));
 sg13g2_or2_1 _3980_ (.X(_0773_),
    .B(_0771_),
    .A(_0728_));
 sg13g2_xnor2_1 _3981_ (.Y(_0774_),
    .A(_0727_),
    .B(_0772_));
 sg13g2_xnor2_1 _3982_ (.Y(_0775_),
    .A(_0770_),
    .B(_0774_));
 sg13g2_o21ai_1 _3983_ (.B1(_0736_),
    .Y(_0776_),
    .A1(_0734_),
    .A2(_0737_));
 sg13g2_nand2_1 _3984_ (.Y(_0777_),
    .A(net956),
    .B(net1009));
 sg13g2_and4_1 _3985_ (.A(net963),
    .B(net959),
    .C(net1005),
    .D(net1056),
    .X(_0778_));
 sg13g2_nand4_1 _3986_ (.B(net959),
    .C(net1005),
    .A(net963),
    .Y(_0779_),
    .D(net1057));
 sg13g2_a22oi_1 _3987_ (.Y(_0780_),
    .B1(net1057),
    .B2(net963),
    .A2(net1005),
    .A1(net959));
 sg13g2_or3_1 _3988_ (.A(_0777_),
    .B(_0778_),
    .C(_0780_),
    .X(_0781_));
 sg13g2_o21ai_1 _3989_ (.B1(_0777_),
    .Y(_0782_),
    .A1(_0778_),
    .A2(_0780_));
 sg13g2_and3_1 _3990_ (.X(_0783_),
    .A(_0776_),
    .B(_0781_),
    .C(_0782_));
 sg13g2_nand3_1 _3991_ (.B(_0781_),
    .C(_0782_),
    .A(_0776_),
    .Y(_0784_));
 sg13g2_a21oi_1 _3992_ (.A1(_0781_),
    .A2(_0782_),
    .Y(_0785_),
    .B1(_0776_));
 sg13g2_or3_1 _3993_ (.A(_0775_),
    .B(_0783_),
    .C(_0785_),
    .X(_0786_));
 sg13g2_o21ai_1 _3994_ (.B1(_0775_),
    .Y(_0787_),
    .A1(_0783_),
    .A2(_0785_));
 sg13g2_and3_1 _3995_ (.X(_0788_),
    .A(_0769_),
    .B(_0786_),
    .C(_0787_));
 sg13g2_nand3_1 _3996_ (.B(_0786_),
    .C(_0787_),
    .A(_0769_),
    .Y(_0789_));
 sg13g2_a21oi_1 _3997_ (.A1(_0786_),
    .A2(_0787_),
    .Y(_0790_),
    .B1(_0769_));
 sg13g2_or3_1 _3998_ (.A(_0768_),
    .B(_0788_),
    .C(_0790_),
    .X(_0791_));
 sg13g2_o21ai_1 _3999_ (.B1(_0768_),
    .Y(_0792_),
    .A1(_0788_),
    .A2(_0790_));
 sg13g2_and3_1 _4000_ (.X(_0793_),
    .A(_0757_),
    .B(_0791_),
    .C(_0792_));
 sg13g2_nand3_1 _4001_ (.B(_0791_),
    .C(_0792_),
    .A(_0757_),
    .Y(_0794_));
 sg13g2_a21oi_1 _4002_ (.A1(_0791_),
    .A2(_0792_),
    .Y(_0795_),
    .B1(_0757_));
 sg13g2_or3_1 _4003_ (.A(_0723_),
    .B(_0793_),
    .C(_0795_),
    .X(_0796_));
 sg13g2_o21ai_1 _4004_ (.B1(_0723_),
    .Y(_0797_),
    .A1(_0793_),
    .A2(_0795_));
 sg13g2_o21ai_1 _4005_ (.B1(_0750_),
    .Y(_0798_),
    .A1(_0689_),
    .A2(_0751_));
 sg13g2_nand3_1 _4006_ (.B(_0797_),
    .C(_0798_),
    .A(_0796_),
    .Y(_0799_));
 sg13g2_a21o_1 _4007_ (.A2(_0797_),
    .A1(_0796_),
    .B1(_0798_),
    .X(_0800_));
 sg13g2_nand2_1 _4008_ (.Y(_0801_),
    .A(_0799_),
    .B(_0800_));
 sg13g2_and4_1 _4009_ (.A(_0754_),
    .B(_0755_),
    .C(_0799_),
    .D(_0800_),
    .X(_0802_));
 sg13g2_xor2_1 _4010_ (.B(_0801_),
    .A(_0756_),
    .X(_0125_));
 sg13g2_o21ai_1 _4011_ (.B1(_0799_),
    .Y(_0803_),
    .A1(_0756_),
    .A2(_0801_));
 sg13g2_o21ai_1 _4012_ (.B1(_0794_),
    .Y(_0804_),
    .A1(_0723_),
    .A2(_0795_));
 sg13g2_o21ai_1 _4013_ (.B1(_0766_),
    .Y(_0805_),
    .A1(_0721_),
    .A2(_0767_));
 sg13g2_o21ai_1 _4014_ (.B1(_0789_),
    .Y(_0806_),
    .A1(_0768_),
    .A2(_0790_));
 sg13g2_nor2_1 _4015_ (.A(_0761_),
    .B(_0764_),
    .Y(_0807_));
 sg13g2_o21ai_1 _4016_ (.B1(_0773_),
    .Y(_0808_),
    .A1(_0770_),
    .A2(_0774_));
 sg13g2_nand2_1 _4017_ (.Y(_0809_),
    .A(net1021),
    .B(net1052));
 sg13g2_nand2_1 _4018_ (.Y(_0810_),
    .A(net1016),
    .B(net947));
 sg13g2_nand2_1 _4019_ (.Y(_0811_),
    .A(net1016),
    .B(net949));
 sg13g2_xor2_1 _4020_ (.B(_0811_),
    .A(_0760_),
    .X(_0812_));
 sg13g2_nand2b_1 _4021_ (.Y(_0813_),
    .B(_0812_),
    .A_N(_0809_));
 sg13g2_xnor2_1 _4022_ (.Y(_0814_),
    .A(_0809_),
    .B(_0812_));
 sg13g2_xnor2_1 _4023_ (.Y(_0815_),
    .A(_0808_),
    .B(_0814_));
 sg13g2_nor2_1 _4024_ (.A(_0807_),
    .B(_0815_),
    .Y(_0816_));
 sg13g2_xnor2_1 _4025_ (.Y(_0817_),
    .A(_0807_),
    .B(_0815_));
 sg13g2_o21ai_1 _4026_ (.B1(_0784_),
    .Y(_0818_),
    .A1(_0775_),
    .A2(_0785_));
 sg13g2_nand2_1 _4027_ (.Y(_0819_),
    .A(net1013),
    .B(net951));
 sg13g2_nand2_1 _4028_ (.Y(_0820_),
    .A(net954),
    .B(net1008));
 sg13g2_or2_1 _4029_ (.X(_0821_),
    .B(_0820_),
    .A(_0771_));
 sg13g2_and2_1 _4030_ (.A(_0771_),
    .B(_0820_),
    .X(_0822_));
 sg13g2_xnor2_1 _4031_ (.Y(_0823_),
    .A(_0771_),
    .B(_0820_));
 sg13g2_xnor2_1 _4032_ (.Y(_0824_),
    .A(_0819_),
    .B(_0823_));
 sg13g2_o21ai_1 _4033_ (.B1(_0779_),
    .Y(_0825_),
    .A1(_0777_),
    .A2(_0780_));
 sg13g2_nand2_1 _4034_ (.Y(_0826_),
    .A(net956),
    .B(net1056));
 sg13g2_and4_1 _4035_ (.A(net960),
    .B(net956),
    .C(net1005),
    .D(net1057),
    .X(_0827_));
 sg13g2_a22oi_1 _4036_ (.Y(_0828_),
    .B1(net1057),
    .B2(net960),
    .A2(net1005),
    .A1(net956));
 sg13g2_nor2_1 _4037_ (.A(_0827_),
    .B(_0828_),
    .Y(_0829_));
 sg13g2_nand2_1 _4038_ (.Y(_0830_),
    .A(_0825_),
    .B(_0829_));
 sg13g2_xnor2_1 _4039_ (.Y(_0831_),
    .A(_0825_),
    .B(_0829_));
 sg13g2_xor2_1 _4040_ (.B(_0831_),
    .A(_0824_),
    .X(_0832_));
 sg13g2_nand2_1 _4041_ (.Y(_0833_),
    .A(_0818_),
    .B(_0832_));
 sg13g2_xnor2_1 _4042_ (.Y(_0834_),
    .A(_0818_),
    .B(_0832_));
 sg13g2_xor2_1 _4043_ (.B(_0834_),
    .A(_0817_),
    .X(_0835_));
 sg13g2_nand2_1 _4044_ (.Y(_0836_),
    .A(_0806_),
    .B(_0835_));
 sg13g2_xnor2_1 _4045_ (.Y(_0837_),
    .A(_0806_),
    .B(_0835_));
 sg13g2_nand2b_1 _4046_ (.Y(_0838_),
    .B(_0805_),
    .A_N(_0837_));
 sg13g2_xnor2_1 _4047_ (.Y(_0839_),
    .A(_0805_),
    .B(_0837_));
 sg13g2_nor2_1 _4048_ (.A(_0804_),
    .B(_0839_),
    .Y(_0840_));
 sg13g2_nand2_1 _4049_ (.Y(_0841_),
    .A(_0804_),
    .B(_0839_));
 sg13g2_nor2b_2 _4050_ (.A(_0840_),
    .B_N(_0841_),
    .Y(_0842_));
 sg13g2_xor2_1 _4051_ (.B(_0842_),
    .A(_0803_),
    .X(_0126_));
 sg13g2_a21oi_1 _4052_ (.A1(_0808_),
    .A2(_0814_),
    .Y(_0843_),
    .B1(_0816_));
 sg13g2_o21ai_1 _4053_ (.B1(_0833_),
    .Y(_0844_),
    .A1(_0817_),
    .A2(_0834_));
 sg13g2_o21ai_1 _4054_ (.B1(_0813_),
    .Y(_0845_),
    .A1(_0760_),
    .A2(_0811_));
 sg13g2_o21ai_1 _4055_ (.B1(_0821_),
    .Y(_0846_),
    .A1(_0819_),
    .A2(_0822_));
 sg13g2_nand2_1 _4056_ (.Y(_0847_),
    .A(net1018),
    .B(net1052));
 sg13g2_nand2_1 _4057_ (.Y(_0848_),
    .A(net1013),
    .B(net947));
 sg13g2_nand2_1 _4058_ (.Y(_0849_),
    .A(net1013),
    .B(net949));
 sg13g2_or2_1 _4059_ (.X(_0850_),
    .B(_0848_),
    .A(_0811_));
 sg13g2_xnor2_1 _4060_ (.Y(_0851_),
    .A(_0810_),
    .B(_0849_));
 sg13g2_xor2_1 _4061_ (.B(_0851_),
    .A(_0847_),
    .X(_0852_));
 sg13g2_xnor2_1 _4062_ (.Y(_0853_),
    .A(_0846_),
    .B(_0852_));
 sg13g2_nor2b_1 _4063_ (.A(_0853_),
    .B_N(_0845_),
    .Y(_0854_));
 sg13g2_xor2_1 _4064_ (.B(_0853_),
    .A(_0845_),
    .X(_0855_));
 sg13g2_o21ai_1 _4065_ (.B1(_0830_),
    .Y(_0856_),
    .A1(_0824_),
    .A2(_0831_));
 sg13g2_a21oi_1 _4066_ (.A1(net960),
    .A2(net1006),
    .Y(_0857_),
    .B1(_0826_));
 sg13g2_nand2_1 _4067_ (.Y(_0858_),
    .A(net1010),
    .B(net951));
 sg13g2_nand2_1 _4068_ (.Y(_0859_),
    .A(net952),
    .B(net1007));
 sg13g2_and4_1 _4069_ (.A(net954),
    .B(net952),
    .C(net1008),
    .D(net1006),
    .X(_0860_));
 sg13g2_a22oi_1 _4070_ (.Y(_0861_),
    .B1(net1006),
    .B2(net954),
    .A2(net1008),
    .A1(net952));
 sg13g2_nor3_1 _4071_ (.A(_0858_),
    .B(_0860_),
    .C(_0861_),
    .Y(_0862_));
 sg13g2_o21ai_1 _4072_ (.B1(_0858_),
    .Y(_0863_),
    .A1(_0860_),
    .A2(_0861_));
 sg13g2_nor2b_1 _4073_ (.A(_0862_),
    .B_N(_0863_),
    .Y(_0864_));
 sg13g2_xnor2_1 _4074_ (.Y(_0865_),
    .A(_0857_),
    .B(_0864_));
 sg13g2_nand2b_1 _4075_ (.Y(_0866_),
    .B(_0856_),
    .A_N(_0865_));
 sg13g2_xor2_1 _4076_ (.B(_0865_),
    .A(_0856_),
    .X(_0867_));
 sg13g2_xor2_1 _4077_ (.B(_0867_),
    .A(_0855_),
    .X(_0868_));
 sg13g2_nand2_1 _4078_ (.Y(_0869_),
    .A(_0844_),
    .B(_0868_));
 sg13g2_xor2_1 _4079_ (.B(_0868_),
    .A(_0844_),
    .X(_0870_));
 sg13g2_nand2b_1 _4080_ (.Y(_0871_),
    .B(_0870_),
    .A_N(_0843_));
 sg13g2_xor2_1 _4081_ (.B(_0870_),
    .A(_0843_),
    .X(_0872_));
 sg13g2_a21oi_1 _4082_ (.A1(_0836_),
    .A2(_0838_),
    .Y(_0873_),
    .B1(_0872_));
 sg13g2_nand3_1 _4083_ (.B(_0838_),
    .C(_0872_),
    .A(_0836_),
    .Y(_0874_));
 sg13g2_nand2b_1 _4084_ (.Y(_0875_),
    .B(_0874_),
    .A_N(_0873_));
 sg13g2_a21oi_1 _4085_ (.A1(_0799_),
    .A2(_0841_),
    .Y(_0876_),
    .B1(_0840_));
 sg13g2_a21oi_2 _4086_ (.B1(_0876_),
    .Y(_0877_),
    .A2(_0842_),
    .A1(_0802_));
 sg13g2_nor2_1 _4087_ (.A(_0875_),
    .B(_0877_),
    .Y(_0878_));
 sg13g2_xor2_1 _4088_ (.B(_0877_),
    .A(_0875_),
    .X(_0117_));
 sg13g2_a21o_1 _4089_ (.A2(_0852_),
    .A1(_0846_),
    .B1(_0854_),
    .X(_0879_));
 sg13g2_o21ai_1 _4090_ (.B1(_0866_),
    .Y(_0880_),
    .A1(_0855_),
    .A2(_0867_));
 sg13g2_a21o_1 _4091_ (.A2(_0864_),
    .A1(_0857_),
    .B1(_0827_),
    .X(_0881_));
 sg13g2_nand2_1 _4092_ (.Y(_0882_),
    .A(net951),
    .B(net1008));
 sg13g2_nand2_1 _4093_ (.Y(_0883_),
    .A(net954),
    .B(net1056));
 sg13g2_or2_1 _4094_ (.X(_0884_),
    .B(_0883_),
    .A(_0859_));
 sg13g2_xnor2_1 _4095_ (.Y(_0885_),
    .A(_0859_),
    .B(_0883_));
 sg13g2_xor2_1 _4096_ (.B(_0885_),
    .A(_0882_),
    .X(_0886_));
 sg13g2_xnor2_1 _4097_ (.Y(_0887_),
    .A(_0881_),
    .B(_0886_));
 sg13g2_o21ai_1 _4098_ (.B1(_0850_),
    .Y(_0888_),
    .A1(_0847_),
    .A2(_0851_));
 sg13g2_or2_1 _4099_ (.X(_0889_),
    .B(_0862_),
    .A(_0860_));
 sg13g2_nand2_1 _4100_ (.Y(_0890_),
    .A(net1016),
    .B(net1052));
 sg13g2_nand2_2 _4101_ (.Y(_0891_),
    .A(net1010),
    .B(net949));
 sg13g2_or2_1 _4102_ (.X(_0892_),
    .B(_0891_),
    .A(_0848_));
 sg13g2_xnor2_1 _4103_ (.Y(_0893_),
    .A(_0848_),
    .B(_0891_));
 sg13g2_xor2_1 _4104_ (.B(_0893_),
    .A(_0890_),
    .X(_0894_));
 sg13g2_xnor2_1 _4105_ (.Y(_0895_),
    .A(_0889_),
    .B(_0894_));
 sg13g2_nor2b_1 _4106_ (.A(_0895_),
    .B_N(_0888_),
    .Y(_0896_));
 sg13g2_xor2_1 _4107_ (.B(_0895_),
    .A(_0888_),
    .X(_0897_));
 sg13g2_nor2_1 _4108_ (.A(_0887_),
    .B(_0897_),
    .Y(_0898_));
 sg13g2_xor2_1 _4109_ (.B(_0897_),
    .A(_0887_),
    .X(_0899_));
 sg13g2_xnor2_1 _4110_ (.Y(_0900_),
    .A(_0880_),
    .B(_0899_));
 sg13g2_nor2b_1 _4111_ (.A(_0900_),
    .B_N(_0879_),
    .Y(_0901_));
 sg13g2_xor2_1 _4112_ (.B(_0900_),
    .A(_0879_),
    .X(_0902_));
 sg13g2_nand3_1 _4113_ (.B(_0871_),
    .C(_0902_),
    .A(_0869_),
    .Y(_0903_));
 sg13g2_inv_1 _4114_ (.Y(_0904_),
    .A(_0903_));
 sg13g2_a21oi_1 _4115_ (.A1(_0869_),
    .A2(_0871_),
    .Y(_0905_),
    .B1(_0902_));
 sg13g2_nor2_1 _4116_ (.A(_0904_),
    .B(_0905_),
    .Y(_0906_));
 sg13g2_nor2_1 _4117_ (.A(_0873_),
    .B(_0878_),
    .Y(_0907_));
 sg13g2_xnor2_1 _4118_ (.Y(_0118_),
    .A(_0906_),
    .B(_0907_));
 sg13g2_a21o_1 _4119_ (.A2(_0894_),
    .A1(_0889_),
    .B1(_0896_),
    .X(_0908_));
 sg13g2_a22oi_1 _4120_ (.Y(_0909_),
    .B1(net1056),
    .B2(net952),
    .A2(net1007),
    .A1(net951));
 sg13g2_nand2_1 _4121_ (.Y(_0910_),
    .A(net951),
    .B(net1056));
 sg13g2_or2_1 _4122_ (.X(_0911_),
    .B(_0910_),
    .A(_0859_));
 sg13g2_nand2b_1 _4123_ (.Y(_0912_),
    .B(_0911_),
    .A_N(_0909_));
 sg13g2_o21ai_1 _4124_ (.B1(_0892_),
    .Y(_0913_),
    .A1(_0890_),
    .A2(_0893_));
 sg13g2_o21ai_1 _4125_ (.B1(_0884_),
    .Y(_0914_),
    .A1(_0882_),
    .A2(_0885_));
 sg13g2_nand2_1 _4126_ (.Y(_0915_),
    .A(net1013),
    .B(net1052));
 sg13g2_nand2_2 _4127_ (.Y(_0916_),
    .A(net1008),
    .B(net947));
 sg13g2_nor2_1 _4128_ (.A(_0891_),
    .B(_0916_),
    .Y(_0917_));
 sg13g2_or2_1 _4129_ (.X(_0918_),
    .B(_0916_),
    .A(_0891_));
 sg13g2_a22oi_1 _4130_ (.Y(_0919_),
    .B1(net947),
    .B2(net1010),
    .A2(net949),
    .A1(net1008));
 sg13g2_nor2_1 _4131_ (.A(_0917_),
    .B(_0919_),
    .Y(_0920_));
 sg13g2_xnor2_1 _4132_ (.Y(_0921_),
    .A(_0915_),
    .B(_0920_));
 sg13g2_xnor2_1 _4133_ (.Y(_0922_),
    .A(_0914_),
    .B(_0921_));
 sg13g2_nor2b_1 _4134_ (.A(_0922_),
    .B_N(_0913_),
    .Y(_0923_));
 sg13g2_xor2_1 _4135_ (.B(_0922_),
    .A(_0913_),
    .X(_0924_));
 sg13g2_or2_1 _4136_ (.X(_0925_),
    .B(_0924_),
    .A(_0912_));
 sg13g2_xor2_1 _4137_ (.B(_0924_),
    .A(_0912_),
    .X(_0926_));
 sg13g2_a21oi_1 _4138_ (.A1(_0881_),
    .A2(_0886_),
    .Y(_0927_),
    .B1(_0898_));
 sg13g2_nor2b_1 _4139_ (.A(_0927_),
    .B_N(_0926_),
    .Y(_0928_));
 sg13g2_xor2_1 _4140_ (.B(_0927_),
    .A(_0926_),
    .X(_0929_));
 sg13g2_nor2b_1 _4141_ (.A(_0929_),
    .B_N(_0908_),
    .Y(_0930_));
 sg13g2_xor2_1 _4142_ (.B(_0929_),
    .A(_0908_),
    .X(_0931_));
 sg13g2_a21oi_1 _4143_ (.A1(_0880_),
    .A2(_0899_),
    .Y(_0932_),
    .B1(_0901_));
 sg13g2_nor2_1 _4144_ (.A(_0931_),
    .B(_0932_),
    .Y(_0933_));
 sg13g2_xor2_1 _4145_ (.B(_0932_),
    .A(_0931_),
    .X(_0934_));
 sg13g2_a21oi_1 _4146_ (.A1(_0873_),
    .A2(_0903_),
    .Y(_0935_),
    .B1(_0905_));
 sg13g2_a21oi_1 _4147_ (.A1(_0874_),
    .A2(_0903_),
    .Y(_0936_),
    .B1(_0905_));
 sg13g2_a21oi_1 _4148_ (.A1(_0877_),
    .A2(_0935_),
    .Y(_0937_),
    .B1(_0936_));
 sg13g2_xor2_1 _4149_ (.B(_0937_),
    .A(_0934_),
    .X(_0119_));
 sg13g2_a21o_1 _4150_ (.A2(_0921_),
    .A1(_0914_),
    .B1(_0923_),
    .X(_0938_));
 sg13g2_o21ai_1 _4151_ (.B1(_0918_),
    .Y(_0939_),
    .A1(_0915_),
    .A2(_0919_));
 sg13g2_nand2_1 _4152_ (.Y(_0940_),
    .A(net1010),
    .B(net1052));
 sg13g2_nand2_1 _4153_ (.Y(_0941_),
    .A(net1007),
    .B(net947));
 sg13g2_nand2_1 _4154_ (.Y(_0942_),
    .A(net949),
    .B(net1007));
 sg13g2_xor2_1 _4155_ (.B(_0942_),
    .A(_0916_),
    .X(_0943_));
 sg13g2_nand2b_1 _4156_ (.Y(_0944_),
    .B(_0943_),
    .A_N(_0940_));
 sg13g2_xnor2_1 _4157_ (.Y(_0945_),
    .A(_0940_),
    .B(_0943_));
 sg13g2_nor2b_1 _4158_ (.A(_0911_),
    .B_N(_0945_),
    .Y(_0946_));
 sg13g2_xnor2_1 _4159_ (.Y(_0947_),
    .A(_0911_),
    .B(_0945_));
 sg13g2_xnor2_1 _4160_ (.Y(_0948_),
    .A(_0939_),
    .B(_0947_));
 sg13g2_nor2_1 _4161_ (.A(_0910_),
    .B(_0948_),
    .Y(_0949_));
 sg13g2_xor2_1 _4162_ (.B(_0948_),
    .A(_0910_),
    .X(_0950_));
 sg13g2_nand2b_1 _4163_ (.Y(_0951_),
    .B(_0950_),
    .A_N(_0925_));
 sg13g2_xnor2_1 _4164_ (.Y(_0952_),
    .A(_0925_),
    .B(_0950_));
 sg13g2_nand2_1 _4165_ (.Y(_0953_),
    .A(_0938_),
    .B(_0952_));
 sg13g2_xor2_1 _4166_ (.B(_0952_),
    .A(_0938_),
    .X(_0954_));
 sg13g2_o21ai_1 _4167_ (.B1(_0954_),
    .Y(_0955_),
    .A1(_0928_),
    .A2(_0930_));
 sg13g2_or3_1 _4168_ (.A(_0928_),
    .B(_0930_),
    .C(_0954_),
    .X(_0956_));
 sg13g2_and2_1 _4169_ (.A(_0955_),
    .B(_0956_),
    .X(_0957_));
 sg13g2_a21oi_1 _4170_ (.A1(_0934_),
    .A2(_0937_),
    .Y(_0958_),
    .B1(_0933_));
 sg13g2_xnor2_1 _4171_ (.Y(_0120_),
    .A(_0957_),
    .B(_0958_));
 sg13g2_and2_1 _4172_ (.A(_0934_),
    .B(_0957_),
    .X(_0959_));
 sg13g2_nand2_1 _4173_ (.Y(_0960_),
    .A(_0933_),
    .B(_0956_));
 sg13g2_nand2_1 _4174_ (.Y(_0961_),
    .A(_0955_),
    .B(_0960_));
 sg13g2_a21o_1 _4175_ (.A2(_0959_),
    .A1(_0937_),
    .B1(_0961_),
    .X(_0962_));
 sg13g2_and2_1 _4176_ (.A(_0951_),
    .B(_0953_),
    .X(_0963_));
 sg13g2_a21o_1 _4177_ (.A2(_0947_),
    .A1(_0939_),
    .B1(_0946_),
    .X(_0964_));
 sg13g2_o21ai_1 _4178_ (.B1(_0944_),
    .Y(_0965_),
    .A1(_0916_),
    .A2(_0942_));
 sg13g2_nand2_1 _4179_ (.Y(_0966_),
    .A(net1008),
    .B(net1052));
 sg13g2_nand2_1 _4180_ (.Y(_0967_),
    .A(net947),
    .B(net1056));
 sg13g2_nand2_1 _4181_ (.Y(_0968_),
    .A(net949),
    .B(net1056));
 sg13g2_xor2_1 _4182_ (.B(_0968_),
    .A(_0941_),
    .X(_0969_));
 sg13g2_nand2b_1 _4183_ (.Y(_0970_),
    .B(_0969_),
    .A_N(_0966_));
 sg13g2_xnor2_1 _4184_ (.Y(_0971_),
    .A(_0966_),
    .B(_0969_));
 sg13g2_nand2_1 _4185_ (.Y(_0972_),
    .A(_0965_),
    .B(_0971_));
 sg13g2_xor2_1 _4186_ (.B(_0971_),
    .A(_0965_),
    .X(_0973_));
 sg13g2_xnor2_1 _4187_ (.Y(_0974_),
    .A(_0949_),
    .B(_0973_));
 sg13g2_nor2b_1 _4188_ (.A(_0974_),
    .B_N(_0964_),
    .Y(_0975_));
 sg13g2_xor2_1 _4189_ (.B(_0974_),
    .A(_0964_),
    .X(_0976_));
 sg13g2_nor2_1 _4190_ (.A(_0963_),
    .B(_0976_),
    .Y(_0977_));
 sg13g2_xor2_1 _4191_ (.B(_0976_),
    .A(_0963_),
    .X(_0978_));
 sg13g2_xor2_1 _4192_ (.B(_0978_),
    .A(_0962_),
    .X(_0121_));
 sg13g2_a21oi_1 _4193_ (.A1(_0962_),
    .A2(_0978_),
    .Y(_0979_),
    .B1(_0977_));
 sg13g2_a21oi_1 _4194_ (.A1(_0949_),
    .A2(_0973_),
    .Y(_0980_),
    .B1(_0975_));
 sg13g2_o21ai_1 _4195_ (.B1(_0970_),
    .Y(_0981_),
    .A1(_0941_),
    .A2(_0968_));
 sg13g2_nand2_1 _4196_ (.Y(_0982_),
    .A(net1007),
    .B(net1052));
 sg13g2_xnor2_1 _4197_ (.Y(_0983_),
    .A(_0967_),
    .B(_0982_));
 sg13g2_xnor2_1 _4198_ (.Y(_0984_),
    .A(_0981_),
    .B(_0983_));
 sg13g2_xnor2_1 _4199_ (.Y(_0985_),
    .A(_0972_),
    .B(_0984_));
 sg13g2_xnor2_1 _4200_ (.Y(_0986_),
    .A(_0980_),
    .B(_0985_));
 sg13g2_xnor2_1 _4201_ (.Y(_0122_),
    .A(_0979_),
    .B(_0986_));
 sg13g2_nor2_1 _4202_ (.A(_2634_),
    .B(_2635_),
    .Y(_0079_));
 sg13g2_and3_2 _4203_ (.X(_0987_),
    .A(net905),
    .B(net847),
    .C(_0079_));
 sg13g2_a22oi_1 _4204_ (.Y(_0988_),
    .B1(net847),
    .B2(net906),
    .A2(net905),
    .A1(net850));
 sg13g2_nor2_1 _4205_ (.A(_0987_),
    .B(_0988_),
    .Y(_0080_));
 sg13g2_nand2_1 _4206_ (.Y(_0989_),
    .A(net906),
    .B(net842));
 sg13g2_and4_1 _4207_ (.A(net850),
    .B(net905),
    .C(net847),
    .D(net902),
    .X(_0990_));
 sg13g2_a22oi_1 _4208_ (.Y(_0991_),
    .B1(net902),
    .B2(net850),
    .A2(net847),
    .A1(net905));
 sg13g2_nor3_1 _4209_ (.A(_0989_),
    .B(_0990_),
    .C(_0991_),
    .Y(_0992_));
 sg13g2_o21ai_1 _4210_ (.B1(_0989_),
    .Y(_0993_),
    .A1(_0990_),
    .A2(_0991_));
 sg13g2_nor2b_1 _4211_ (.A(_0992_),
    .B_N(_0993_),
    .Y(_0994_));
 sg13g2_nand2_1 _4212_ (.Y(_0995_),
    .A(_0987_),
    .B(_0994_));
 sg13g2_xor2_1 _4213_ (.B(_0994_),
    .A(_0987_),
    .X(_0081_));
 sg13g2_nand2_1 _4214_ (.Y(_0996_),
    .A(net906),
    .B(net840));
 sg13g2_or2_1 _4215_ (.X(_0997_),
    .B(_0992_),
    .A(_0990_));
 sg13g2_nand2_1 _4216_ (.Y(_0998_),
    .A(net905),
    .B(net842));
 sg13g2_and4_1 _4217_ (.A(net850),
    .B(net847),
    .C(net902),
    .D(net900),
    .X(_0999_));
 sg13g2_nand4_1 _4218_ (.B(net846),
    .C(net902),
    .A(net850),
    .Y(_1000_),
    .D(net900));
 sg13g2_a22oi_1 _4219_ (.Y(_1001_),
    .B1(net900),
    .B2(net850),
    .A2(net902),
    .A1(net847));
 sg13g2_nor3_1 _4220_ (.A(_0998_),
    .B(_0999_),
    .C(_1001_),
    .Y(_1002_));
 sg13g2_o21ai_1 _4221_ (.B1(_0998_),
    .Y(_1003_),
    .A1(_0999_),
    .A2(_1001_));
 sg13g2_nor2b_1 _4222_ (.A(_1002_),
    .B_N(_1003_),
    .Y(_1004_));
 sg13g2_nand2_1 _4223_ (.Y(_1005_),
    .A(_0997_),
    .B(_1004_));
 sg13g2_xnor2_1 _4224_ (.Y(_1006_),
    .A(_0997_),
    .B(_1004_));
 sg13g2_xor2_1 _4225_ (.B(_1006_),
    .A(_0996_),
    .X(_1007_));
 sg13g2_nand2b_1 _4226_ (.Y(_1008_),
    .B(_1007_),
    .A_N(_0995_));
 sg13g2_xnor2_1 _4227_ (.Y(_0082_),
    .A(_0995_),
    .B(_1007_));
 sg13g2_a22oi_1 _4228_ (.Y(_1009_),
    .B1(net838),
    .B2(net906),
    .A2(net840),
    .A1(net904));
 sg13g2_nand2_1 _4229_ (.Y(_1010_),
    .A(net904),
    .B(net838));
 sg13g2_and4_1 _4230_ (.A(net906),
    .B(net904),
    .C(net840),
    .D(net838),
    .X(_1011_));
 sg13g2_nor2_1 _4231_ (.A(_1009_),
    .B(_1011_),
    .Y(_1012_));
 sg13g2_inv_1 _4232_ (.Y(_1013_),
    .A(_1012_));
 sg13g2_o21ai_1 _4233_ (.B1(_1000_),
    .Y(_1014_),
    .A1(_0998_),
    .A2(_1001_));
 sg13g2_nand2_1 _4234_ (.Y(_1015_),
    .A(net902),
    .B(net842));
 sg13g2_and4_1 _4235_ (.A(net849),
    .B(net846),
    .C(net900),
    .D(net898),
    .X(_1016_));
 sg13g2_nand4_1 _4236_ (.B(net846),
    .C(net900),
    .A(net849),
    .Y(_1017_),
    .D(net898));
 sg13g2_a22oi_1 _4237_ (.Y(_1018_),
    .B1(net898),
    .B2(net849),
    .A2(net900),
    .A1(net846));
 sg13g2_or3_1 _4238_ (.A(_1015_),
    .B(_1016_),
    .C(_1018_),
    .X(_1019_));
 sg13g2_o21ai_1 _4239_ (.B1(_1015_),
    .Y(_1020_),
    .A1(_1016_),
    .A2(_1018_));
 sg13g2_nand3_1 _4240_ (.B(_1019_),
    .C(_1020_),
    .A(_1014_),
    .Y(_1021_));
 sg13g2_a21oi_1 _4241_ (.A1(_1019_),
    .A2(_1020_),
    .Y(_1022_),
    .B1(_1014_));
 sg13g2_a21o_1 _4242_ (.A2(_1020_),
    .A1(_1019_),
    .B1(_1014_),
    .X(_1023_));
 sg13g2_nand2_1 _4243_ (.Y(_1024_),
    .A(_1021_),
    .B(_1023_));
 sg13g2_xnor2_1 _4244_ (.Y(_1025_),
    .A(_1013_),
    .B(_1024_));
 sg13g2_o21ai_1 _4245_ (.B1(_1005_),
    .Y(_1026_),
    .A1(_0996_),
    .A2(_1006_));
 sg13g2_nor2b_2 _4246_ (.A(_1025_),
    .B_N(_1026_),
    .Y(_1027_));
 sg13g2_xor2_1 _4247_ (.B(_1026_),
    .A(_1025_),
    .X(_1028_));
 sg13g2_or2_1 _4248_ (.X(_1029_),
    .B(_1028_),
    .A(_1008_));
 sg13g2_xor2_1 _4249_ (.B(_1028_),
    .A(_1008_),
    .X(_0083_));
 sg13g2_o21ai_1 _4250_ (.B1(_1021_),
    .Y(_1030_),
    .A1(_1013_),
    .A2(_1022_));
 sg13g2_nand2_1 _4251_ (.Y(_1031_),
    .A(net906),
    .B(net837));
 sg13g2_nand2_1 _4252_ (.Y(_1032_),
    .A(net903),
    .B(net838));
 sg13g2_nand2_1 _4253_ (.Y(_1033_),
    .A(net903),
    .B(net840));
 sg13g2_xor2_1 _4254_ (.B(_1033_),
    .A(_1010_),
    .X(_1034_));
 sg13g2_nand2b_1 _4255_ (.Y(_1035_),
    .B(_1034_),
    .A_N(_1031_));
 sg13g2_xor2_1 _4256_ (.B(_1034_),
    .A(_1031_),
    .X(_1036_));
 sg13g2_o21ai_1 _4257_ (.B1(_1017_),
    .Y(_1037_),
    .A1(_1015_),
    .A2(_1018_));
 sg13g2_nand2_1 _4258_ (.Y(_1038_),
    .A(net843),
    .B(net901));
 sg13g2_and4_1 _4259_ (.A(net849),
    .B(net846),
    .C(net898),
    .D(net896),
    .X(_1039_));
 sg13g2_nand4_1 _4260_ (.B(net846),
    .C(net898),
    .A(net848),
    .Y(_1040_),
    .D(net896));
 sg13g2_a22oi_1 _4261_ (.Y(_1041_),
    .B1(net896),
    .B2(net849),
    .A2(net898),
    .A1(net846));
 sg13g2_or3_1 _4262_ (.A(_1038_),
    .B(_1039_),
    .C(_1041_),
    .X(_1042_));
 sg13g2_o21ai_1 _4263_ (.B1(_1038_),
    .Y(_1043_),
    .A1(_1039_),
    .A2(_1041_));
 sg13g2_and3_1 _4264_ (.X(_1044_),
    .A(_1037_),
    .B(_1042_),
    .C(_1043_));
 sg13g2_nand3_1 _4265_ (.B(_1042_),
    .C(_1043_),
    .A(_1037_),
    .Y(_1045_));
 sg13g2_a21oi_1 _4266_ (.A1(_1042_),
    .A2(_1043_),
    .Y(_1046_),
    .B1(_1037_));
 sg13g2_or3_1 _4267_ (.A(_1036_),
    .B(_1044_),
    .C(_1046_),
    .X(_1047_));
 sg13g2_o21ai_1 _4268_ (.B1(_1036_),
    .Y(_1048_),
    .A1(_1044_),
    .A2(_1046_));
 sg13g2_nand3_1 _4269_ (.B(_1047_),
    .C(_1048_),
    .A(_1030_),
    .Y(_1049_));
 sg13g2_a21o_1 _4270_ (.A2(_1048_),
    .A1(_1047_),
    .B1(_1030_),
    .X(_1050_));
 sg13g2_nand3_1 _4271_ (.B(_1049_),
    .C(_1050_),
    .A(_1011_),
    .Y(_1051_));
 sg13g2_a21o_1 _4272_ (.A2(_1050_),
    .A1(_1049_),
    .B1(_1011_),
    .X(_1052_));
 sg13g2_and2_1 _4273_ (.A(_1051_),
    .B(_1052_),
    .X(_1053_));
 sg13g2_nand3_1 _4274_ (.B(_1051_),
    .C(_1052_),
    .A(_1027_),
    .Y(_1054_));
 sg13g2_a21oi_1 _4275_ (.A1(_1051_),
    .A2(_1052_),
    .Y(_1055_),
    .B1(_1027_));
 sg13g2_xor2_1 _4276_ (.B(_1053_),
    .A(_1027_),
    .X(_1056_));
 sg13g2_xnor2_1 _4277_ (.Y(_0127_),
    .A(_1029_),
    .B(_1056_));
 sg13g2_nand2_1 _4278_ (.Y(_1057_),
    .A(_1049_),
    .B(_1051_));
 sg13g2_o21ai_1 _4279_ (.B1(_1035_),
    .Y(_1058_),
    .A1(_1010_),
    .A2(_1033_));
 sg13g2_nand2_1 _4280_ (.Y(_1059_),
    .A(net907),
    .B(net835));
 sg13g2_nand2b_1 _4281_ (.Y(_1060_),
    .B(_1058_),
    .A_N(_1059_));
 sg13g2_xor2_1 _4282_ (.B(_1059_),
    .A(_1058_),
    .X(_1061_));
 sg13g2_o21ai_1 _4283_ (.B1(_1045_),
    .Y(_1062_),
    .A1(_1036_),
    .A2(_1046_));
 sg13g2_nand2_1 _4284_ (.Y(_1063_),
    .A(net904),
    .B(net837));
 sg13g2_nand2_1 _4285_ (.Y(_1064_),
    .A(net901),
    .B(net839));
 sg13g2_nand2_2 _4286_ (.Y(_1065_),
    .A(net901),
    .B(net840));
 sg13g2_xor2_1 _4287_ (.B(_1065_),
    .A(_1032_),
    .X(_1066_));
 sg13g2_nand2b_1 _4288_ (.Y(_1067_),
    .B(_1066_),
    .A_N(_1063_));
 sg13g2_xnor2_1 _4289_ (.Y(_1068_),
    .A(_1063_),
    .B(_1066_));
 sg13g2_o21ai_1 _4290_ (.B1(_1040_),
    .Y(_1069_),
    .A1(_1038_),
    .A2(_1041_));
 sg13g2_nand2_1 _4291_ (.Y(_1070_),
    .A(net843),
    .B(net898));
 sg13g2_and4_1 _4292_ (.A(net848),
    .B(net844),
    .C(net896),
    .D(net894),
    .X(_1071_));
 sg13g2_nand4_1 _4293_ (.B(net844),
    .C(net896),
    .A(net848),
    .Y(_1072_),
    .D(net894));
 sg13g2_a22oi_1 _4294_ (.Y(_1073_),
    .B1(net894),
    .B2(net848),
    .A2(net896),
    .A1(net844));
 sg13g2_or3_1 _4295_ (.A(_1070_),
    .B(_1071_),
    .C(_1073_),
    .X(_1074_));
 sg13g2_o21ai_1 _4296_ (.B1(_1070_),
    .Y(_1075_),
    .A1(_1071_),
    .A2(_1073_));
 sg13g2_and3_1 _4297_ (.X(_1076_),
    .A(_1069_),
    .B(_1074_),
    .C(_1075_));
 sg13g2_nand3_1 _4298_ (.B(_1074_),
    .C(_1075_),
    .A(_1069_),
    .Y(_1077_));
 sg13g2_a21o_1 _4299_ (.A2(_1075_),
    .A1(_1074_),
    .B1(_1069_),
    .X(_1078_));
 sg13g2_nand3_1 _4300_ (.B(_1077_),
    .C(_1078_),
    .A(_1068_),
    .Y(_1079_));
 sg13g2_a21o_1 _4301_ (.A2(_1078_),
    .A1(_1077_),
    .B1(_1068_),
    .X(_1080_));
 sg13g2_nand3_1 _4302_ (.B(_1079_),
    .C(_1080_),
    .A(_1062_),
    .Y(_1081_));
 sg13g2_a21oi_1 _4303_ (.A1(_1079_),
    .A2(_1080_),
    .Y(_1082_),
    .B1(_1062_));
 sg13g2_a21o_1 _4304_ (.A2(_1080_),
    .A1(_1079_),
    .B1(_1062_),
    .X(_1083_));
 sg13g2_nand2_1 _4305_ (.Y(_1084_),
    .A(_1081_),
    .B(_1083_));
 sg13g2_xnor2_1 _4306_ (.Y(_1085_),
    .A(_1061_),
    .B(_1084_));
 sg13g2_nor2b_1 _4307_ (.A(_1085_),
    .B_N(_1057_),
    .Y(_1086_));
 sg13g2_xnor2_1 _4308_ (.Y(_1087_),
    .A(_1057_),
    .B(_1085_));
 sg13g2_o21ai_1 _4309_ (.B1(_1054_),
    .Y(_1088_),
    .A1(_1029_),
    .A2(_1055_));
 sg13g2_xor2_1 _4310_ (.B(_1088_),
    .A(_1087_),
    .X(_0134_));
 sg13g2_o21ai_1 _4311_ (.B1(_1081_),
    .Y(_1089_),
    .A1(_1061_),
    .A2(_1082_));
 sg13g2_o21ai_1 _4312_ (.B1(_1067_),
    .Y(_1090_),
    .A1(_1032_),
    .A2(_1065_));
 sg13g2_a22oi_1 _4313_ (.Y(_1091_),
    .B1(net833),
    .B2(net907),
    .A2(net835),
    .A1(net904));
 sg13g2_nand4_1 _4314_ (.B(\DP_3.matrix[37] ),
    .C(net835),
    .A(net907),
    .Y(_1092_),
    .D(net833));
 sg13g2_nor2b_1 _4315_ (.A(_1091_),
    .B_N(_1092_),
    .Y(_1093_));
 sg13g2_nand2_1 _4316_ (.Y(_1094_),
    .A(_1090_),
    .B(_1093_));
 sg13g2_xnor2_1 _4317_ (.Y(_1095_),
    .A(_1090_),
    .B(_1093_));
 sg13g2_a21o_1 _4318_ (.A2(_1078_),
    .A1(_1068_),
    .B1(_1076_),
    .X(_1096_));
 sg13g2_nand2_1 _4319_ (.Y(_1097_),
    .A(net903),
    .B(net837));
 sg13g2_nand2_1 _4320_ (.Y(_1098_),
    .A(net899),
    .B(net838));
 sg13g2_nand2_1 _4321_ (.Y(_1099_),
    .A(net840),
    .B(net899));
 sg13g2_or2_1 _4322_ (.X(_1100_),
    .B(_1098_),
    .A(_1065_));
 sg13g2_and2_1 _4323_ (.A(_1064_),
    .B(_1099_),
    .X(_1101_));
 sg13g2_xnor2_1 _4324_ (.Y(_1102_),
    .A(_1064_),
    .B(_1099_));
 sg13g2_xnor2_1 _4325_ (.Y(_1103_),
    .A(_1097_),
    .B(_1102_));
 sg13g2_o21ai_1 _4326_ (.B1(_1072_),
    .Y(_1104_),
    .A1(_1070_),
    .A2(_1073_));
 sg13g2_nand2_1 _4327_ (.Y(_1105_),
    .A(net842),
    .B(net896));
 sg13g2_and4_1 _4328_ (.A(net849),
    .B(net844),
    .C(net894),
    .D(net891),
    .X(_1106_));
 sg13g2_nand4_1 _4329_ (.B(net844),
    .C(net894),
    .A(net848),
    .Y(_1107_),
    .D(net891));
 sg13g2_a22oi_1 _4330_ (.Y(_1108_),
    .B1(net891),
    .B2(net848),
    .A2(net894),
    .A1(net845));
 sg13g2_or3_1 _4331_ (.A(_1105_),
    .B(_1106_),
    .C(_1108_),
    .X(_1109_));
 sg13g2_o21ai_1 _4332_ (.B1(_1105_),
    .Y(_1110_),
    .A1(_1106_),
    .A2(_1108_));
 sg13g2_and3_1 _4333_ (.X(_1111_),
    .A(_1104_),
    .B(_1109_),
    .C(_1110_));
 sg13g2_nand3_1 _4334_ (.B(_1109_),
    .C(_1110_),
    .A(_1104_),
    .Y(_1112_));
 sg13g2_a21oi_1 _4335_ (.A1(_1109_),
    .A2(_1110_),
    .Y(_1113_),
    .B1(_1104_));
 sg13g2_or3_1 _4336_ (.A(_1103_),
    .B(_1111_),
    .C(_1113_),
    .X(_1114_));
 sg13g2_o21ai_1 _4337_ (.B1(_1103_),
    .Y(_1115_),
    .A1(_1111_),
    .A2(_1113_));
 sg13g2_and3_1 _4338_ (.X(_1116_),
    .A(_1096_),
    .B(_1114_),
    .C(_1115_));
 sg13g2_nand3_1 _4339_ (.B(_1114_),
    .C(_1115_),
    .A(_1096_),
    .Y(_1117_));
 sg13g2_a21oi_1 _4340_ (.A1(_1114_),
    .A2(_1115_),
    .Y(_1118_),
    .B1(_1096_));
 sg13g2_or3_1 _4341_ (.A(_1095_),
    .B(_1116_),
    .C(_1118_),
    .X(_1119_));
 sg13g2_o21ai_1 _4342_ (.B1(_1095_),
    .Y(_1120_),
    .A1(_1116_),
    .A2(_1118_));
 sg13g2_nand3_1 _4343_ (.B(_1119_),
    .C(_1120_),
    .A(_1089_),
    .Y(_1121_));
 sg13g2_a21oi_1 _4344_ (.A1(_1119_),
    .A2(_1120_),
    .Y(_1122_),
    .B1(_1089_));
 sg13g2_a21o_1 _4345_ (.A2(_1120_),
    .A1(_1119_),
    .B1(_1089_),
    .X(_1123_));
 sg13g2_nand2_1 _4346_ (.Y(_1124_),
    .A(_1121_),
    .B(_1123_));
 sg13g2_xor2_1 _4347_ (.B(_1124_),
    .A(_1060_),
    .X(_1125_));
 sg13g2_a21o_2 _4348_ (.A2(_1088_),
    .A1(_1087_),
    .B1(_1086_),
    .X(_1126_));
 sg13g2_nand2_1 _4349_ (.Y(_1127_),
    .A(_1125_),
    .B(_1126_));
 sg13g2_xor2_1 _4350_ (.B(_1126_),
    .A(_1125_),
    .X(_0135_));
 sg13g2_o21ai_1 _4351_ (.B1(_1117_),
    .Y(_1128_),
    .A1(_1095_),
    .A2(_1118_));
 sg13g2_o21ai_1 _4352_ (.B1(_1100_),
    .Y(_1129_),
    .A1(_1097_),
    .A2(_1101_));
 sg13g2_nand2_1 _4353_ (.Y(_1130_),
    .A(net907),
    .B(net1043));
 sg13g2_nand2_1 _4354_ (.Y(_1131_),
    .A(net903),
    .B(net833));
 sg13g2_and4_1 _4355_ (.A(net904),
    .B(net903),
    .C(net835),
    .D(net833),
    .X(_1132_));
 sg13g2_a22oi_1 _4356_ (.Y(_1133_),
    .B1(net833),
    .B2(net904),
    .A2(net835),
    .A1(net903));
 sg13g2_or2_1 _4357_ (.X(_1134_),
    .B(_1133_),
    .A(_1132_));
 sg13g2_nor2_1 _4358_ (.A(_1130_),
    .B(_1134_),
    .Y(_1135_));
 sg13g2_xor2_1 _4359_ (.B(_1134_),
    .A(_1130_),
    .X(_1136_));
 sg13g2_nand2_1 _4360_ (.Y(_1137_),
    .A(_1129_),
    .B(_1136_));
 sg13g2_xnor2_1 _4361_ (.Y(_1138_),
    .A(_1129_),
    .B(_1136_));
 sg13g2_xnor2_1 _4362_ (.Y(_1139_),
    .A(_1092_),
    .B(_1138_));
 sg13g2_o21ai_1 _4363_ (.B1(_1112_),
    .Y(_1140_),
    .A1(_1103_),
    .A2(_1113_));
 sg13g2_nand2_1 _4364_ (.Y(_1141_),
    .A(net901),
    .B(net837));
 sg13g2_nand2_2 _4365_ (.Y(_1142_),
    .A(net839),
    .B(net897));
 sg13g2_nand2_1 _4366_ (.Y(_1143_),
    .A(net840),
    .B(net897));
 sg13g2_or2_1 _4367_ (.X(_1144_),
    .B(_1142_),
    .A(_1099_));
 sg13g2_xnor2_1 _4368_ (.Y(_1145_),
    .A(_1098_),
    .B(_1143_));
 sg13g2_xnor2_1 _4369_ (.Y(_1146_),
    .A(_1141_),
    .B(_1145_));
 sg13g2_o21ai_1 _4370_ (.B1(_1107_),
    .Y(_1147_),
    .A1(_1105_),
    .A2(_1108_));
 sg13g2_nand2_1 _4371_ (.Y(_1148_),
    .A(net842),
    .B(net894));
 sg13g2_and4_1 _4372_ (.A(net849),
    .B(net844),
    .C(net891),
    .D(net1047),
    .X(_1149_));
 sg13g2_nand4_1 _4373_ (.B(net845),
    .C(net891),
    .A(net848),
    .Y(_1150_),
    .D(net1047));
 sg13g2_a22oi_1 _4374_ (.Y(_1151_),
    .B1(net1047),
    .B2(net848),
    .A2(net891),
    .A1(net845));
 sg13g2_or3_1 _4375_ (.A(_1148_),
    .B(_1149_),
    .C(_1151_),
    .X(_1152_));
 sg13g2_o21ai_1 _4376_ (.B1(_1148_),
    .Y(_1153_),
    .A1(_1149_),
    .A2(_1151_));
 sg13g2_and3_1 _4377_ (.X(_1154_),
    .A(_1147_),
    .B(_1152_),
    .C(_1153_));
 sg13g2_nand3_1 _4378_ (.B(_1152_),
    .C(_1153_),
    .A(_1147_),
    .Y(_1155_));
 sg13g2_a21oi_1 _4379_ (.A1(_1152_),
    .A2(_1153_),
    .Y(_1156_),
    .B1(_1147_));
 sg13g2_or3_1 _4380_ (.A(_1146_),
    .B(_1154_),
    .C(_1156_),
    .X(_1157_));
 sg13g2_o21ai_1 _4381_ (.B1(_1146_),
    .Y(_1158_),
    .A1(_1154_),
    .A2(_1156_));
 sg13g2_and3_1 _4382_ (.X(_1159_),
    .A(_1140_),
    .B(_1157_),
    .C(_1158_));
 sg13g2_nand3_1 _4383_ (.B(_1157_),
    .C(_1158_),
    .A(_1140_),
    .Y(_1160_));
 sg13g2_a21oi_1 _4384_ (.A1(_1157_),
    .A2(_1158_),
    .Y(_1161_),
    .B1(_1140_));
 sg13g2_or3_1 _4385_ (.A(_1139_),
    .B(_1159_),
    .C(_1161_),
    .X(_1162_));
 sg13g2_o21ai_1 _4386_ (.B1(_1139_),
    .Y(_1163_),
    .A1(_1159_),
    .A2(_1161_));
 sg13g2_and3_1 _4387_ (.X(_1164_),
    .A(_1128_),
    .B(_1162_),
    .C(_1163_));
 sg13g2_nand3_1 _4388_ (.B(_1162_),
    .C(_1163_),
    .A(_1128_),
    .Y(_1165_));
 sg13g2_a21oi_1 _4389_ (.A1(_1162_),
    .A2(_1163_),
    .Y(_1166_),
    .B1(_1128_));
 sg13g2_or3_1 _4390_ (.A(_1094_),
    .B(_1164_),
    .C(_1166_),
    .X(_1167_));
 sg13g2_o21ai_1 _4391_ (.B1(_1094_),
    .Y(_1168_),
    .A1(_1164_),
    .A2(_1166_));
 sg13g2_o21ai_1 _4392_ (.B1(_1121_),
    .Y(_1169_),
    .A1(_1060_),
    .A2(_1122_));
 sg13g2_nand3_1 _4393_ (.B(_1168_),
    .C(_1169_),
    .A(_1167_),
    .Y(_1170_));
 sg13g2_a21o_1 _4394_ (.A2(_1168_),
    .A1(_1167_),
    .B1(_1169_),
    .X(_1171_));
 sg13g2_nand2_1 _4395_ (.Y(_1172_),
    .A(_1170_),
    .B(_1171_));
 sg13g2_and4_1 _4396_ (.A(_1125_),
    .B(_1126_),
    .C(_1170_),
    .D(_1171_),
    .X(_1173_));
 sg13g2_xor2_1 _4397_ (.B(_1172_),
    .A(_1127_),
    .X(_0136_));
 sg13g2_o21ai_1 _4398_ (.B1(_1170_),
    .Y(_1174_),
    .A1(_1127_),
    .A2(_1172_));
 sg13g2_o21ai_1 _4399_ (.B1(_1165_),
    .Y(_1175_),
    .A1(_1094_),
    .A2(_1166_));
 sg13g2_o21ai_1 _4400_ (.B1(_1137_),
    .Y(_1176_),
    .A1(_1092_),
    .A2(_1138_));
 sg13g2_o21ai_1 _4401_ (.B1(_1160_),
    .Y(_1177_),
    .A1(_1139_),
    .A2(_1161_));
 sg13g2_nor2_1 _4402_ (.A(_1132_),
    .B(_1135_),
    .Y(_1178_));
 sg13g2_o21ai_1 _4403_ (.B1(_1144_),
    .Y(_1179_),
    .A1(_1141_),
    .A2(_1145_));
 sg13g2_nand2_1 _4404_ (.Y(_1180_),
    .A(net904),
    .B(net1043));
 sg13g2_nand2_1 _4405_ (.Y(_1181_),
    .A(net901),
    .B(net834));
 sg13g2_nand2_1 _4406_ (.Y(_1182_),
    .A(net901),
    .B(net836));
 sg13g2_xor2_1 _4407_ (.B(_1182_),
    .A(_1131_),
    .X(_1183_));
 sg13g2_nand2b_1 _4408_ (.Y(_1184_),
    .B(_1183_),
    .A_N(_1180_));
 sg13g2_xnor2_1 _4409_ (.Y(_1185_),
    .A(_1180_),
    .B(_1183_));
 sg13g2_xnor2_1 _4410_ (.Y(_1186_),
    .A(_1179_),
    .B(_1185_));
 sg13g2_nor2_1 _4411_ (.A(_1178_),
    .B(_1186_),
    .Y(_1187_));
 sg13g2_xnor2_1 _4412_ (.Y(_1188_),
    .A(_1178_),
    .B(_1186_));
 sg13g2_o21ai_1 _4413_ (.B1(_1155_),
    .Y(_1189_),
    .A1(_1146_),
    .A2(_1156_));
 sg13g2_nand2_1 _4414_ (.Y(_1190_),
    .A(net899),
    .B(\DP_4.matrix[41] ));
 sg13g2_nand2_1 _4415_ (.Y(_1191_),
    .A(net841),
    .B(net895));
 sg13g2_or2_1 _4416_ (.X(_1192_),
    .B(_1191_),
    .A(_1142_));
 sg13g2_and2_1 _4417_ (.A(_1142_),
    .B(_1191_),
    .X(_1193_));
 sg13g2_xnor2_1 _4418_ (.Y(_1194_),
    .A(_1142_),
    .B(_1191_));
 sg13g2_xnor2_1 _4419_ (.Y(_1195_),
    .A(_1190_),
    .B(_1194_));
 sg13g2_o21ai_1 _4420_ (.B1(_1150_),
    .Y(_1196_),
    .A1(_1148_),
    .A2(_1151_));
 sg13g2_nand2_1 _4421_ (.Y(_1197_),
    .A(net843),
    .B(net1047));
 sg13g2_and4_1 _4422_ (.A(net844),
    .B(net842),
    .C(net892),
    .D(net1047),
    .X(_1198_));
 sg13g2_a22oi_1 _4423_ (.Y(_1199_),
    .B1(net1047),
    .B2(net845),
    .A2(net891),
    .A1(net843));
 sg13g2_nor2_1 _4424_ (.A(_1198_),
    .B(_1199_),
    .Y(_1200_));
 sg13g2_nand2_1 _4425_ (.Y(_1201_),
    .A(_1196_),
    .B(_1200_));
 sg13g2_xnor2_1 _4426_ (.Y(_1202_),
    .A(_1196_),
    .B(_1200_));
 sg13g2_xor2_1 _4427_ (.B(_1202_),
    .A(_1195_),
    .X(_1203_));
 sg13g2_nand2_1 _4428_ (.Y(_1204_),
    .A(_1189_),
    .B(_1203_));
 sg13g2_xnor2_1 _4429_ (.Y(_1205_),
    .A(_1189_),
    .B(_1203_));
 sg13g2_xor2_1 _4430_ (.B(_1205_),
    .A(_1188_),
    .X(_1206_));
 sg13g2_nand2_1 _4431_ (.Y(_1207_),
    .A(_1177_),
    .B(_1206_));
 sg13g2_xnor2_1 _4432_ (.Y(_1208_),
    .A(_1177_),
    .B(_1206_));
 sg13g2_nand2b_1 _4433_ (.Y(_1209_),
    .B(_1176_),
    .A_N(_1208_));
 sg13g2_xnor2_1 _4434_ (.Y(_1210_),
    .A(_1176_),
    .B(_1208_));
 sg13g2_nor2_1 _4435_ (.A(_1175_),
    .B(_1210_),
    .Y(_1211_));
 sg13g2_nand2_1 _4436_ (.Y(_1212_),
    .A(_1175_),
    .B(_1210_));
 sg13g2_nor2b_1 _4437_ (.A(_1211_),
    .B_N(_1212_),
    .Y(_1213_));
 sg13g2_xor2_1 _4438_ (.B(_1213_),
    .A(_1174_),
    .X(_0137_));
 sg13g2_a21oi_1 _4439_ (.A1(_1179_),
    .A2(_1185_),
    .Y(_1214_),
    .B1(_1187_));
 sg13g2_o21ai_1 _4440_ (.B1(_1204_),
    .Y(_1215_),
    .A1(_1188_),
    .A2(_1205_));
 sg13g2_o21ai_1 _4441_ (.B1(_1184_),
    .Y(_1216_),
    .A1(_1131_),
    .A2(_1182_));
 sg13g2_o21ai_1 _4442_ (.B1(_1192_),
    .Y(_1217_),
    .A1(_1190_),
    .A2(_1193_));
 sg13g2_nand2_1 _4443_ (.Y(_1218_),
    .A(net903),
    .B(net1043));
 sg13g2_nand2_1 _4444_ (.Y(_1219_),
    .A(net899),
    .B(net834));
 sg13g2_nand2_1 _4445_ (.Y(_1220_),
    .A(net899),
    .B(net836));
 sg13g2_or2_1 _4446_ (.X(_1221_),
    .B(_1219_),
    .A(_1182_));
 sg13g2_xnor2_1 _4447_ (.Y(_1222_),
    .A(_1181_),
    .B(_1220_));
 sg13g2_xor2_1 _4448_ (.B(_1222_),
    .A(_1218_),
    .X(_1223_));
 sg13g2_xnor2_1 _4449_ (.Y(_1224_),
    .A(_1217_),
    .B(_1223_));
 sg13g2_nor2b_1 _4450_ (.A(_1224_),
    .B_N(_1216_),
    .Y(_1225_));
 sg13g2_xor2_1 _4451_ (.B(_1224_),
    .A(_1216_),
    .X(_1226_));
 sg13g2_o21ai_1 _4452_ (.B1(_1201_),
    .Y(_1227_),
    .A1(_1195_),
    .A2(_1202_));
 sg13g2_a21oi_1 _4453_ (.A1(net844),
    .A2(net891),
    .Y(_1228_),
    .B1(_1197_));
 sg13g2_nand2_1 _4454_ (.Y(_1229_),
    .A(net897),
    .B(\DP_4.matrix[41] ));
 sg13g2_nand2_1 _4455_ (.Y(_1230_),
    .A(net839),
    .B(net893));
 sg13g2_and4_1 _4456_ (.A(net841),
    .B(net839),
    .C(net895),
    .D(net893),
    .X(_1231_));
 sg13g2_a22oi_1 _4457_ (.Y(_1232_),
    .B1(net893),
    .B2(net841),
    .A2(net895),
    .A1(net838));
 sg13g2_nor3_1 _4458_ (.A(_1229_),
    .B(_1231_),
    .C(_1232_),
    .Y(_1233_));
 sg13g2_o21ai_1 _4459_ (.B1(_1229_),
    .Y(_1234_),
    .A1(_1231_),
    .A2(_1232_));
 sg13g2_nor2b_1 _4460_ (.A(_1233_),
    .B_N(_1234_),
    .Y(_1235_));
 sg13g2_xnor2_1 _4461_ (.Y(_1236_),
    .A(_1228_),
    .B(_1235_));
 sg13g2_nand2b_1 _4462_ (.Y(_1237_),
    .B(_1227_),
    .A_N(_1236_));
 sg13g2_xor2_1 _4463_ (.B(_1236_),
    .A(_1227_),
    .X(_1238_));
 sg13g2_xor2_1 _4464_ (.B(_1238_),
    .A(_1226_),
    .X(_1239_));
 sg13g2_nand2_1 _4465_ (.Y(_1240_),
    .A(_1215_),
    .B(_1239_));
 sg13g2_xor2_1 _4466_ (.B(_1239_),
    .A(_1215_),
    .X(_1241_));
 sg13g2_nand2b_1 _4467_ (.Y(_1242_),
    .B(_1241_),
    .A_N(_1214_));
 sg13g2_xor2_1 _4468_ (.B(_1241_),
    .A(_1214_),
    .X(_1243_));
 sg13g2_a21oi_1 _4469_ (.A1(_1207_),
    .A2(_1209_),
    .Y(_1244_),
    .B1(_1243_));
 sg13g2_nand3_1 _4470_ (.B(_1209_),
    .C(_1243_),
    .A(_1207_),
    .Y(_1245_));
 sg13g2_nand2b_1 _4471_ (.Y(_1246_),
    .B(_1245_),
    .A_N(_1244_));
 sg13g2_a21oi_1 _4472_ (.A1(_1170_),
    .A2(_1212_),
    .Y(_1247_),
    .B1(_1211_));
 sg13g2_a21oi_2 _4473_ (.B1(_1247_),
    .Y(_1248_),
    .A2(_1213_),
    .A1(_1173_));
 sg13g2_nor2_1 _4474_ (.A(_1246_),
    .B(_1248_),
    .Y(_1249_));
 sg13g2_xor2_1 _4475_ (.B(_1248_),
    .A(_1246_),
    .X(_0128_));
 sg13g2_a21o_1 _4476_ (.A2(_1223_),
    .A1(_1217_),
    .B1(_1225_),
    .X(_1250_));
 sg13g2_o21ai_1 _4477_ (.B1(_1237_),
    .Y(_1251_),
    .A1(_1226_),
    .A2(_1238_));
 sg13g2_a21o_1 _4478_ (.A2(_1235_),
    .A1(_1228_),
    .B1(_1198_),
    .X(_1252_));
 sg13g2_nand2_2 _4479_ (.Y(_1253_),
    .A(net837),
    .B(\DP_3.matrix[42] ));
 sg13g2_nand2_1 _4480_ (.Y(_1254_),
    .A(net841),
    .B(net1048));
 sg13g2_or2_1 _4481_ (.X(_1255_),
    .B(_1254_),
    .A(_1230_));
 sg13g2_xnor2_1 _4482_ (.Y(_1256_),
    .A(_1230_),
    .B(_1254_));
 sg13g2_xor2_1 _4483_ (.B(_1256_),
    .A(_1253_),
    .X(_1257_));
 sg13g2_xnor2_1 _4484_ (.Y(_1258_),
    .A(_1252_),
    .B(_1257_));
 sg13g2_o21ai_1 _4485_ (.B1(_1221_),
    .Y(_1259_),
    .A1(_1218_),
    .A2(_1222_));
 sg13g2_or2_1 _4486_ (.X(_1260_),
    .B(_1233_),
    .A(_1231_));
 sg13g2_nand2_1 _4487_ (.Y(_1261_),
    .A(net901),
    .B(net1043));
 sg13g2_nand2_2 _4488_ (.Y(_1262_),
    .A(net897),
    .B(net836));
 sg13g2_or2_1 _4489_ (.X(_1263_),
    .B(_1262_),
    .A(_1219_));
 sg13g2_xnor2_1 _4490_ (.Y(_1264_),
    .A(_1219_),
    .B(_1262_));
 sg13g2_xor2_1 _4491_ (.B(_1264_),
    .A(_1261_),
    .X(_1265_));
 sg13g2_xnor2_1 _4492_ (.Y(_1266_),
    .A(_1260_),
    .B(_1265_));
 sg13g2_nor2b_1 _4493_ (.A(_1266_),
    .B_N(_1259_),
    .Y(_1267_));
 sg13g2_xor2_1 _4494_ (.B(_1266_),
    .A(_1259_),
    .X(_1268_));
 sg13g2_nor2_1 _4495_ (.A(_1258_),
    .B(_1268_),
    .Y(_1269_));
 sg13g2_xor2_1 _4496_ (.B(_1268_),
    .A(_1258_),
    .X(_1270_));
 sg13g2_xnor2_1 _4497_ (.Y(_1271_),
    .A(_1251_),
    .B(_1270_));
 sg13g2_nor2b_1 _4498_ (.A(_1271_),
    .B_N(_1250_),
    .Y(_1272_));
 sg13g2_xor2_1 _4499_ (.B(_1271_),
    .A(_1250_),
    .X(_1273_));
 sg13g2_nand3_1 _4500_ (.B(_1242_),
    .C(_1273_),
    .A(_1240_),
    .Y(_1274_));
 sg13g2_inv_1 _4501_ (.Y(_1275_),
    .A(_1274_));
 sg13g2_a21oi_1 _4502_ (.A1(_1240_),
    .A2(_1242_),
    .Y(_1276_),
    .B1(_1273_));
 sg13g2_nor2_1 _4503_ (.A(_1275_),
    .B(_1276_),
    .Y(_1277_));
 sg13g2_nor2_1 _4504_ (.A(_1244_),
    .B(_1249_),
    .Y(_1278_));
 sg13g2_xnor2_1 _4505_ (.Y(_0129_),
    .A(_1277_),
    .B(_1278_));
 sg13g2_a21o_1 _4506_ (.A2(_1265_),
    .A1(_1260_),
    .B1(_1267_),
    .X(_1279_));
 sg13g2_a22oi_1 _4507_ (.Y(_1280_),
    .B1(net1048),
    .B2(net839),
    .A2(net893),
    .A1(\DP_4.matrix[41] ));
 sg13g2_nand2_2 _4508_ (.Y(_1281_),
    .A(net837),
    .B(net1048));
 sg13g2_or2_1 _4509_ (.X(_1282_),
    .B(_1281_),
    .A(_1230_));
 sg13g2_nand2b_1 _4510_ (.Y(_1283_),
    .B(_1282_),
    .A_N(_1280_));
 sg13g2_o21ai_1 _4511_ (.B1(_1263_),
    .Y(_1284_),
    .A1(_1261_),
    .A2(_1264_));
 sg13g2_o21ai_1 _4512_ (.B1(_1255_),
    .Y(_1285_),
    .A1(_1253_),
    .A2(_1256_));
 sg13g2_nand2_1 _4513_ (.Y(_1286_),
    .A(net899),
    .B(net1043));
 sg13g2_nand2_2 _4514_ (.Y(_1287_),
    .A(net895),
    .B(net834));
 sg13g2_nor2_1 _4515_ (.A(_1262_),
    .B(_1287_),
    .Y(_1288_));
 sg13g2_or2_1 _4516_ (.X(_1289_),
    .B(_1287_),
    .A(_1262_));
 sg13g2_a22oi_1 _4517_ (.Y(_1290_),
    .B1(net834),
    .B2(net897),
    .A2(net836),
    .A1(net895));
 sg13g2_nor2_1 _4518_ (.A(_1288_),
    .B(_1290_),
    .Y(_1291_));
 sg13g2_xnor2_1 _4519_ (.Y(_1292_),
    .A(_1286_),
    .B(_1291_));
 sg13g2_xnor2_1 _4520_ (.Y(_1293_),
    .A(_1285_),
    .B(_1292_));
 sg13g2_nor2b_1 _4521_ (.A(_1293_),
    .B_N(_1284_),
    .Y(_1294_));
 sg13g2_xor2_1 _4522_ (.B(_1293_),
    .A(_1284_),
    .X(_1295_));
 sg13g2_or2_1 _4523_ (.X(_1296_),
    .B(_1295_),
    .A(_1283_));
 sg13g2_xor2_1 _4524_ (.B(_1295_),
    .A(_1283_),
    .X(_1297_));
 sg13g2_a21oi_1 _4525_ (.A1(_1252_),
    .A2(_1257_),
    .Y(_1298_),
    .B1(_1269_));
 sg13g2_nor2b_1 _4526_ (.A(_1298_),
    .B_N(_1297_),
    .Y(_1299_));
 sg13g2_xor2_1 _4527_ (.B(_1298_),
    .A(_1297_),
    .X(_1300_));
 sg13g2_nor2b_1 _4528_ (.A(_1300_),
    .B_N(_1279_),
    .Y(_1301_));
 sg13g2_xor2_1 _4529_ (.B(_1300_),
    .A(_1279_),
    .X(_1302_));
 sg13g2_a21oi_1 _4530_ (.A1(_1251_),
    .A2(_1270_),
    .Y(_1303_),
    .B1(_1272_));
 sg13g2_nor2_1 _4531_ (.A(_1302_),
    .B(_1303_),
    .Y(_1304_));
 sg13g2_xor2_1 _4532_ (.B(_1303_),
    .A(_1302_),
    .X(_1305_));
 sg13g2_a21oi_1 _4533_ (.A1(_1244_),
    .A2(_1274_),
    .Y(_1306_),
    .B1(_1276_));
 sg13g2_a21oi_1 _4534_ (.A1(_1245_),
    .A2(_1274_),
    .Y(_1307_),
    .B1(_1276_));
 sg13g2_a21oi_2 _4535_ (.B1(_1307_),
    .Y(_1308_),
    .A2(_1306_),
    .A1(_1248_));
 sg13g2_xor2_1 _4536_ (.B(_1308_),
    .A(_1305_),
    .X(_0130_));
 sg13g2_a21o_1 _4537_ (.A2(_1292_),
    .A1(_1285_),
    .B1(_1294_),
    .X(_1309_));
 sg13g2_o21ai_1 _4538_ (.B1(_1289_),
    .Y(_1310_),
    .A1(_1286_),
    .A2(_1290_));
 sg13g2_nand2_1 _4539_ (.Y(_1311_),
    .A(net897),
    .B(\DP_4.matrix[44] ));
 sg13g2_nand2_1 _4540_ (.Y(_1312_),
    .A(net893),
    .B(net834));
 sg13g2_nand2_1 _4541_ (.Y(_1313_),
    .A(net836),
    .B(net893));
 sg13g2_xor2_1 _4542_ (.B(_1313_),
    .A(_1287_),
    .X(_1314_));
 sg13g2_nand2b_1 _4543_ (.Y(_1315_),
    .B(_1314_),
    .A_N(_1311_));
 sg13g2_xnor2_1 _4544_ (.Y(_1316_),
    .A(_1311_),
    .B(_1314_));
 sg13g2_nor2b_1 _4545_ (.A(_1282_),
    .B_N(_1316_),
    .Y(_1317_));
 sg13g2_xnor2_1 _4546_ (.Y(_1318_),
    .A(_1282_),
    .B(_1316_));
 sg13g2_xnor2_1 _4547_ (.Y(_1319_),
    .A(_1310_),
    .B(_1318_));
 sg13g2_nor2_1 _4548_ (.A(_1281_),
    .B(_1319_),
    .Y(_1320_));
 sg13g2_xor2_1 _4549_ (.B(_1319_),
    .A(_1281_),
    .X(_1321_));
 sg13g2_nand2b_1 _4550_ (.Y(_1322_),
    .B(_1321_),
    .A_N(_1296_));
 sg13g2_xnor2_1 _4551_ (.Y(_1323_),
    .A(_1296_),
    .B(_1321_));
 sg13g2_nand2_1 _4552_ (.Y(_1324_),
    .A(_1309_),
    .B(_1323_));
 sg13g2_xor2_1 _4553_ (.B(_1323_),
    .A(_1309_),
    .X(_1325_));
 sg13g2_o21ai_1 _4554_ (.B1(_1325_),
    .Y(_1326_),
    .A1(_1299_),
    .A2(_1301_));
 sg13g2_or3_1 _4555_ (.A(_1299_),
    .B(_1301_),
    .C(_1325_),
    .X(_1327_));
 sg13g2_and2_1 _4556_ (.A(_1326_),
    .B(_1327_),
    .X(_1328_));
 sg13g2_a21oi_1 _4557_ (.A1(_1305_),
    .A2(_1308_),
    .Y(_1329_),
    .B1(_1304_));
 sg13g2_xnor2_1 _4558_ (.Y(_0131_),
    .A(_1328_),
    .B(_1329_));
 sg13g2_and2_1 _4559_ (.A(_1305_),
    .B(_1328_),
    .X(_1330_));
 sg13g2_nand2_1 _4560_ (.Y(_1331_),
    .A(_1304_),
    .B(_1327_));
 sg13g2_nand2_1 _4561_ (.Y(_1332_),
    .A(_1326_),
    .B(_1331_));
 sg13g2_a21o_1 _4562_ (.A2(_1330_),
    .A1(_1308_),
    .B1(_1332_),
    .X(_1333_));
 sg13g2_and2_1 _4563_ (.A(_1322_),
    .B(_1324_),
    .X(_1334_));
 sg13g2_a21o_1 _4564_ (.A2(_1318_),
    .A1(_1310_),
    .B1(_1317_),
    .X(_1335_));
 sg13g2_o21ai_1 _4565_ (.B1(_1315_),
    .Y(_1336_),
    .A1(_1287_),
    .A2(_1313_));
 sg13g2_nand2_1 _4566_ (.Y(_1337_),
    .A(net895),
    .B(\DP_4.matrix[44] ));
 sg13g2_nand2_1 _4567_ (.Y(_1338_),
    .A(net833),
    .B(net1048));
 sg13g2_nand2_1 _4568_ (.Y(_1339_),
    .A(net835),
    .B(net1048));
 sg13g2_xor2_1 _4569_ (.B(_1339_),
    .A(_1312_),
    .X(_1340_));
 sg13g2_nand2b_1 _4570_ (.Y(_1341_),
    .B(_1340_),
    .A_N(_1337_));
 sg13g2_xnor2_1 _4571_ (.Y(_1342_),
    .A(_1337_),
    .B(_1340_));
 sg13g2_nand2_1 _4572_ (.Y(_1343_),
    .A(_1336_),
    .B(_1342_));
 sg13g2_xor2_1 _4573_ (.B(_1342_),
    .A(_1336_),
    .X(_1344_));
 sg13g2_xnor2_1 _4574_ (.Y(_1345_),
    .A(_1320_),
    .B(_1344_));
 sg13g2_nor2b_1 _4575_ (.A(_1345_),
    .B_N(_1335_),
    .Y(_1346_));
 sg13g2_xor2_1 _4576_ (.B(_1345_),
    .A(_1335_),
    .X(_1347_));
 sg13g2_nor2_1 _4577_ (.A(_1334_),
    .B(_1347_),
    .Y(_1348_));
 sg13g2_xor2_1 _4578_ (.B(_1347_),
    .A(_1334_),
    .X(_1349_));
 sg13g2_xor2_1 _4579_ (.B(_1349_),
    .A(_1333_),
    .X(_0132_));
 sg13g2_a21oi_1 _4580_ (.A1(_1333_),
    .A2(_1349_),
    .Y(_1350_),
    .B1(_1348_));
 sg13g2_a21oi_1 _4581_ (.A1(_1320_),
    .A2(_1344_),
    .Y(_1351_),
    .B1(_1346_));
 sg13g2_o21ai_1 _4582_ (.B1(_1341_),
    .Y(_1352_),
    .A1(_1312_),
    .A2(_1339_));
 sg13g2_nand2_1 _4583_ (.Y(_1353_),
    .A(net893),
    .B(net1043));
 sg13g2_xnor2_1 _4584_ (.Y(_1354_),
    .A(_1338_),
    .B(_1353_));
 sg13g2_xnor2_1 _4585_ (.Y(_1355_),
    .A(_1352_),
    .B(_1354_));
 sg13g2_xnor2_1 _4586_ (.Y(_1356_),
    .A(_1343_),
    .B(_1355_));
 sg13g2_xnor2_1 _4587_ (.Y(_1357_),
    .A(_1351_),
    .B(_1356_));
 sg13g2_xnor2_1 _4588_ (.Y(_0133_),
    .A(_1350_),
    .B(_1357_));
 sg13g2_and2_1 _4589_ (.A(net924),
    .B(net869),
    .X(_0084_));
 sg13g2_and3_2 _4590_ (.X(_1358_),
    .A(net923),
    .B(net863),
    .C(_0084_));
 sg13g2_a22oi_1 _4591_ (.Y(_1359_),
    .B1(net863),
    .B2(net924),
    .A2(net923),
    .A1(net869));
 sg13g2_nor2_1 _4592_ (.A(_1358_),
    .B(_1359_),
    .Y(_0085_));
 sg13g2_nand2_1 _4593_ (.Y(_1360_),
    .A(net924),
    .B(net861));
 sg13g2_and4_1 _4594_ (.A(net869),
    .B(net923),
    .C(net863),
    .D(net920),
    .X(_1361_));
 sg13g2_a22oi_1 _4595_ (.Y(_1362_),
    .B1(net920),
    .B2(net869),
    .A2(net863),
    .A1(net923));
 sg13g2_nor3_1 _4596_ (.A(_1360_),
    .B(_1361_),
    .C(_1362_),
    .Y(_1363_));
 sg13g2_o21ai_1 _4597_ (.B1(_1360_),
    .Y(_1364_),
    .A1(_1361_),
    .A2(_1362_));
 sg13g2_nor2b_1 _4598_ (.A(_1363_),
    .B_N(_1364_),
    .Y(_1365_));
 sg13g2_nand2_1 _4599_ (.Y(_1366_),
    .A(_1358_),
    .B(_1365_));
 sg13g2_xor2_1 _4600_ (.B(_1365_),
    .A(_1358_),
    .X(_0086_));
 sg13g2_nand2_1 _4601_ (.Y(_1367_),
    .A(net924),
    .B(net859));
 sg13g2_or2_1 _4602_ (.X(_1368_),
    .B(_1363_),
    .A(_1361_));
 sg13g2_nand2_1 _4603_ (.Y(_1369_),
    .A(net923),
    .B(net861));
 sg13g2_and4_1 _4604_ (.A(net869),
    .B(net863),
    .C(net920),
    .D(net918),
    .X(_1370_));
 sg13g2_nand4_1 _4605_ (.B(net866),
    .C(net920),
    .A(net869),
    .Y(_1371_),
    .D(net918));
 sg13g2_a22oi_1 _4606_ (.Y(_1372_),
    .B1(net918),
    .B2(net869),
    .A2(net920),
    .A1(net863));
 sg13g2_nor3_1 _4607_ (.A(_1369_),
    .B(_1370_),
    .C(_1372_),
    .Y(_1373_));
 sg13g2_o21ai_1 _4608_ (.B1(_1369_),
    .Y(_1374_),
    .A1(_1370_),
    .A2(_1372_));
 sg13g2_nor2b_1 _4609_ (.A(_1373_),
    .B_N(_1374_),
    .Y(_1375_));
 sg13g2_nand2_1 _4610_ (.Y(_1376_),
    .A(_1368_),
    .B(_1375_));
 sg13g2_xnor2_1 _4611_ (.Y(_1377_),
    .A(_1368_),
    .B(_1375_));
 sg13g2_xor2_1 _4612_ (.B(_1377_),
    .A(_1367_),
    .X(_1378_));
 sg13g2_nand2b_1 _4613_ (.Y(_1379_),
    .B(_1378_),
    .A_N(_1366_));
 sg13g2_xnor2_1 _4614_ (.Y(_0087_),
    .A(_1366_),
    .B(_1378_));
 sg13g2_a22oi_1 _4615_ (.Y(_1380_),
    .B1(net857),
    .B2(net924),
    .A2(net859),
    .A1(net922));
 sg13g2_nand2_1 _4616_ (.Y(_1381_),
    .A(net922),
    .B(net857));
 sg13g2_and4_1 _4617_ (.A(net924),
    .B(net922),
    .C(net859),
    .D(net857),
    .X(_1382_));
 sg13g2_nor2_1 _4618_ (.A(_1380_),
    .B(_1382_),
    .Y(_1383_));
 sg13g2_inv_1 _4619_ (.Y(_1384_),
    .A(_1383_));
 sg13g2_o21ai_1 _4620_ (.B1(_1371_),
    .Y(_1385_),
    .A1(_1369_),
    .A2(_1372_));
 sg13g2_nand2_1 _4621_ (.Y(_1386_),
    .A(net920),
    .B(net862));
 sg13g2_and4_1 _4622_ (.A(net868),
    .B(net865),
    .C(net918),
    .D(net916),
    .X(_1387_));
 sg13g2_nand4_1 _4623_ (.B(net865),
    .C(net918),
    .A(net868),
    .Y(_1388_),
    .D(net916));
 sg13g2_a22oi_1 _4624_ (.Y(_1389_),
    .B1(net916),
    .B2(net868),
    .A2(net918),
    .A1(net865));
 sg13g2_or3_1 _4625_ (.A(_1386_),
    .B(_1387_),
    .C(_1389_),
    .X(_1390_));
 sg13g2_o21ai_1 _4626_ (.B1(_1386_),
    .Y(_1391_),
    .A1(_1387_),
    .A2(_1389_));
 sg13g2_nand3_1 _4627_ (.B(_1390_),
    .C(_1391_),
    .A(_1385_),
    .Y(_1392_));
 sg13g2_a21oi_1 _4628_ (.A1(_1390_),
    .A2(_1391_),
    .Y(_1393_),
    .B1(_1385_));
 sg13g2_a21o_1 _4629_ (.A2(_1391_),
    .A1(_1390_),
    .B1(_1385_),
    .X(_1394_));
 sg13g2_nand2_1 _4630_ (.Y(_1395_),
    .A(_1392_),
    .B(_1394_));
 sg13g2_xnor2_1 _4631_ (.Y(_1396_),
    .A(_1384_),
    .B(_1395_));
 sg13g2_o21ai_1 _4632_ (.B1(_1376_),
    .Y(_1397_),
    .A1(_1367_),
    .A2(_1377_));
 sg13g2_nor2b_2 _4633_ (.A(_1396_),
    .B_N(_1397_),
    .Y(_1398_));
 sg13g2_xor2_1 _4634_ (.B(_1397_),
    .A(_1396_),
    .X(_1399_));
 sg13g2_or2_1 _4635_ (.X(_1400_),
    .B(_1399_),
    .A(_1379_));
 sg13g2_xor2_1 _4636_ (.B(_1399_),
    .A(_1379_),
    .X(_0088_));
 sg13g2_o21ai_1 _4637_ (.B1(_1392_),
    .Y(_1401_),
    .A1(_1384_),
    .A2(_1393_));
 sg13g2_nand2_1 _4638_ (.Y(_1402_),
    .A(net925),
    .B(net856));
 sg13g2_nand2_1 _4639_ (.Y(_1403_),
    .A(net921),
    .B(net858));
 sg13g2_nand2_1 _4640_ (.Y(_1404_),
    .A(net921),
    .B(net860));
 sg13g2_xor2_1 _4641_ (.B(_1404_),
    .A(_1381_),
    .X(_1405_));
 sg13g2_nand2b_1 _4642_ (.Y(_1406_),
    .B(_1405_),
    .A_N(_1402_));
 sg13g2_xor2_1 _4643_ (.B(_1405_),
    .A(_1402_),
    .X(_1407_));
 sg13g2_o21ai_1 _4644_ (.B1(_1388_),
    .Y(_1408_),
    .A1(_1386_),
    .A2(_1389_));
 sg13g2_nand2_1 _4645_ (.Y(_1409_),
    .A(net862),
    .B(net919));
 sg13g2_and4_1 _4646_ (.A(net868),
    .B(net865),
    .C(net916),
    .D(net915),
    .X(_1410_));
 sg13g2_nand4_1 _4647_ (.B(net865),
    .C(net916),
    .A(net868),
    .Y(_1411_),
    .D(net915));
 sg13g2_a22oi_1 _4648_ (.Y(_1412_),
    .B1(net915),
    .B2(net868),
    .A2(net916),
    .A1(net865));
 sg13g2_or3_1 _4649_ (.A(_1409_),
    .B(_1410_),
    .C(_1412_),
    .X(_1413_));
 sg13g2_o21ai_1 _4650_ (.B1(_1409_),
    .Y(_1414_),
    .A1(_1410_),
    .A2(_1412_));
 sg13g2_and3_1 _4651_ (.X(_1415_),
    .A(_1408_),
    .B(_1413_),
    .C(_1414_));
 sg13g2_nand3_1 _4652_ (.B(_1413_),
    .C(_1414_),
    .A(_1408_),
    .Y(_1416_));
 sg13g2_a21oi_1 _4653_ (.A1(_1413_),
    .A2(_1414_),
    .Y(_1417_),
    .B1(_1408_));
 sg13g2_or3_1 _4654_ (.A(_1407_),
    .B(_1415_),
    .C(_1417_),
    .X(_1418_));
 sg13g2_o21ai_1 _4655_ (.B1(_1407_),
    .Y(_1419_),
    .A1(_1415_),
    .A2(_1417_));
 sg13g2_nand3_1 _4656_ (.B(_1418_),
    .C(_1419_),
    .A(_1401_),
    .Y(_1420_));
 sg13g2_a21o_1 _4657_ (.A2(_1419_),
    .A1(_1418_),
    .B1(_1401_),
    .X(_1421_));
 sg13g2_nand3_1 _4658_ (.B(_1420_),
    .C(_1421_),
    .A(_1382_),
    .Y(_1422_));
 sg13g2_a21o_1 _4659_ (.A2(_1421_),
    .A1(_1420_),
    .B1(_1382_),
    .X(_1423_));
 sg13g2_and2_1 _4660_ (.A(_1422_),
    .B(_1423_),
    .X(_1424_));
 sg13g2_nand3_1 _4661_ (.B(_1422_),
    .C(_1423_),
    .A(_1398_),
    .Y(_1425_));
 sg13g2_a21oi_1 _4662_ (.A1(_1422_),
    .A2(_1423_),
    .Y(_1426_),
    .B1(_1398_));
 sg13g2_xor2_1 _4663_ (.B(_1424_),
    .A(_1398_),
    .X(_1427_));
 sg13g2_xnor2_1 _4664_ (.Y(_0138_),
    .A(_1400_),
    .B(_1427_));
 sg13g2_nand2_1 _4665_ (.Y(_1428_),
    .A(_1420_),
    .B(_1422_));
 sg13g2_o21ai_1 _4666_ (.B1(_1406_),
    .Y(_1429_),
    .A1(_1381_),
    .A2(_1404_));
 sg13g2_nand2_1 _4667_ (.Y(_1430_),
    .A(net925),
    .B(net855));
 sg13g2_nand2b_2 _4668_ (.Y(_1431_),
    .B(_1429_),
    .A_N(_1430_));
 sg13g2_xor2_1 _4669_ (.B(_1430_),
    .A(_1429_),
    .X(_1432_));
 sg13g2_o21ai_1 _4670_ (.B1(_1416_),
    .Y(_1433_),
    .A1(_1407_),
    .A2(_1417_));
 sg13g2_nand2_1 _4671_ (.Y(_1434_),
    .A(net922),
    .B(\DP_4.matrix[5] ));
 sg13g2_nand2_1 _4672_ (.Y(_1435_),
    .A(net919),
    .B(net857));
 sg13g2_nand2_1 _4673_ (.Y(_1436_),
    .A(net919),
    .B(net859));
 sg13g2_xor2_1 _4674_ (.B(_1436_),
    .A(_1403_),
    .X(_1437_));
 sg13g2_nand2b_1 _4675_ (.Y(_1438_),
    .B(_1437_),
    .A_N(_1434_));
 sg13g2_xnor2_1 _4676_ (.Y(_1439_),
    .A(_1434_),
    .B(_1437_));
 sg13g2_o21ai_1 _4677_ (.B1(_1411_),
    .Y(_1440_),
    .A1(_1409_),
    .A2(_1412_));
 sg13g2_nand2_1 _4678_ (.Y(_1441_),
    .A(net861),
    .B(net917));
 sg13g2_and4_1 _4679_ (.A(net867),
    .B(net865),
    .C(net914),
    .D(net913),
    .X(_1442_));
 sg13g2_nand4_1 _4680_ (.B(net864),
    .C(net914),
    .A(net867),
    .Y(_1443_),
    .D(net913));
 sg13g2_a22oi_1 _4681_ (.Y(_1444_),
    .B1(net913),
    .B2(net867),
    .A2(net914),
    .A1(net864));
 sg13g2_or3_1 _4682_ (.A(_1441_),
    .B(_1442_),
    .C(_1444_),
    .X(_1445_));
 sg13g2_o21ai_1 _4683_ (.B1(_1441_),
    .Y(_1446_),
    .A1(_1442_),
    .A2(_1444_));
 sg13g2_and3_1 _4684_ (.X(_1447_),
    .A(_1440_),
    .B(_1445_),
    .C(_1446_));
 sg13g2_nand3_1 _4685_ (.B(_1445_),
    .C(_1446_),
    .A(_1440_),
    .Y(_1448_));
 sg13g2_a21o_1 _4686_ (.A2(_1446_),
    .A1(_1445_),
    .B1(_1440_),
    .X(_1449_));
 sg13g2_nand3_1 _4687_ (.B(_1448_),
    .C(_1449_),
    .A(_1439_),
    .Y(_1450_));
 sg13g2_a21o_1 _4688_ (.A2(_1449_),
    .A1(_1448_),
    .B1(_1439_),
    .X(_1451_));
 sg13g2_nand3_1 _4689_ (.B(_1450_),
    .C(_1451_),
    .A(_1433_),
    .Y(_1452_));
 sg13g2_a21oi_1 _4690_ (.A1(_1450_),
    .A2(_1451_),
    .Y(_1453_),
    .B1(_1433_));
 sg13g2_a21o_1 _4691_ (.A2(_1451_),
    .A1(_1450_),
    .B1(_1433_),
    .X(_1454_));
 sg13g2_nand2_1 _4692_ (.Y(_1455_),
    .A(_1452_),
    .B(_1454_));
 sg13g2_xnor2_1 _4693_ (.Y(_1456_),
    .A(_1432_),
    .B(_1455_));
 sg13g2_nor2b_1 _4694_ (.A(_1456_),
    .B_N(_1428_),
    .Y(_1457_));
 sg13g2_xnor2_1 _4695_ (.Y(_1458_),
    .A(_1428_),
    .B(_1456_));
 sg13g2_o21ai_1 _4696_ (.B1(_1425_),
    .Y(_1459_),
    .A1(_1400_),
    .A2(_1426_));
 sg13g2_xor2_1 _4697_ (.B(_1459_),
    .A(_1458_),
    .X(_0145_));
 sg13g2_o21ai_1 _4698_ (.B1(_1452_),
    .Y(_1460_),
    .A1(_1432_),
    .A2(_1453_));
 sg13g2_o21ai_1 _4699_ (.B1(_1438_),
    .Y(_1461_),
    .A1(_1403_),
    .A2(_1436_));
 sg13g2_a22oi_1 _4700_ (.Y(_1462_),
    .B1(net851),
    .B2(net925),
    .A2(net854),
    .A1(net922));
 sg13g2_nand4_1 _4701_ (.B(\DP_3.matrix[1] ),
    .C(net854),
    .A(net925),
    .Y(_1463_),
    .D(net851));
 sg13g2_nor2b_1 _4702_ (.A(_1462_),
    .B_N(_1463_),
    .Y(_1464_));
 sg13g2_nand2_1 _4703_ (.Y(_1465_),
    .A(_1461_),
    .B(_1464_));
 sg13g2_xnor2_1 _4704_ (.Y(_1466_),
    .A(_1461_),
    .B(_1464_));
 sg13g2_a21o_1 _4705_ (.A2(_1449_),
    .A1(_1439_),
    .B1(_1447_),
    .X(_1467_));
 sg13g2_nand2_1 _4706_ (.Y(_1468_),
    .A(net921),
    .B(\DP_4.matrix[5] ));
 sg13g2_nand2_1 _4707_ (.Y(_1469_),
    .A(net917),
    .B(net857));
 sg13g2_nand2_1 _4708_ (.Y(_1470_),
    .A(net859),
    .B(net917));
 sg13g2_or2_1 _4709_ (.X(_1471_),
    .B(_1469_),
    .A(_1436_));
 sg13g2_and2_1 _4710_ (.A(_1435_),
    .B(_1470_),
    .X(_1472_));
 sg13g2_xnor2_1 _4711_ (.Y(_1473_),
    .A(_1435_),
    .B(_1470_));
 sg13g2_xnor2_1 _4712_ (.Y(_1474_),
    .A(_1468_),
    .B(_1473_));
 sg13g2_o21ai_1 _4713_ (.B1(_1443_),
    .Y(_1475_),
    .A1(_1441_),
    .A2(_1444_));
 sg13g2_nand2_1 _4714_ (.Y(_1476_),
    .A(net861),
    .B(net914));
 sg13g2_and4_1 _4715_ (.A(net867),
    .B(net864),
    .C(net911),
    .D(net909),
    .X(_1477_));
 sg13g2_nand4_1 _4716_ (.B(net864),
    .C(net911),
    .A(\DP_4.matrix[0] ),
    .Y(_1478_),
    .D(net909));
 sg13g2_a22oi_1 _4717_ (.Y(_1479_),
    .B1(net909),
    .B2(net867),
    .A2(net911),
    .A1(net864));
 sg13g2_or3_1 _4718_ (.A(_1476_),
    .B(_1477_),
    .C(_1479_),
    .X(_1480_));
 sg13g2_o21ai_1 _4719_ (.B1(_1476_),
    .Y(_1481_),
    .A1(_1477_),
    .A2(_1479_));
 sg13g2_and3_1 _4720_ (.X(_1482_),
    .A(_1475_),
    .B(_1480_),
    .C(_1481_));
 sg13g2_nand3_1 _4721_ (.B(_1480_),
    .C(_1481_),
    .A(_1475_),
    .Y(_1483_));
 sg13g2_a21oi_1 _4722_ (.A1(_1480_),
    .A2(_1481_),
    .Y(_1484_),
    .B1(_1475_));
 sg13g2_or3_1 _4723_ (.A(_1474_),
    .B(_1482_),
    .C(_1484_),
    .X(_1485_));
 sg13g2_o21ai_1 _4724_ (.B1(_1474_),
    .Y(_1486_),
    .A1(_1482_),
    .A2(_1484_));
 sg13g2_and3_1 _4725_ (.X(_1487_),
    .A(_1467_),
    .B(_1485_),
    .C(_1486_));
 sg13g2_nand3_1 _4726_ (.B(_1485_),
    .C(_1486_),
    .A(_1467_),
    .Y(_1488_));
 sg13g2_a21oi_1 _4727_ (.A1(_1485_),
    .A2(_1486_),
    .Y(_1489_),
    .B1(_1467_));
 sg13g2_or3_1 _4728_ (.A(_1466_),
    .B(_1487_),
    .C(_1489_),
    .X(_1490_));
 sg13g2_o21ai_1 _4729_ (.B1(_1466_),
    .Y(_1491_),
    .A1(_1487_),
    .A2(_1489_));
 sg13g2_nand3_1 _4730_ (.B(_1490_),
    .C(_1491_),
    .A(_1460_),
    .Y(_1492_));
 sg13g2_a21oi_1 _4731_ (.A1(_1490_),
    .A2(_1491_),
    .Y(_1493_),
    .B1(_1460_));
 sg13g2_a21o_1 _4732_ (.A2(_1491_),
    .A1(_1490_),
    .B1(_1460_),
    .X(_1494_));
 sg13g2_nand2_1 _4733_ (.Y(_1495_),
    .A(_1492_),
    .B(_1494_));
 sg13g2_xor2_1 _4734_ (.B(_1495_),
    .A(_1431_),
    .X(_1496_));
 sg13g2_a21o_2 _4735_ (.A2(_1459_),
    .A1(_1458_),
    .B1(_1457_),
    .X(_1497_));
 sg13g2_nand2_1 _4736_ (.Y(_1498_),
    .A(_1496_),
    .B(_1497_));
 sg13g2_xor2_1 _4737_ (.B(_1497_),
    .A(_1496_),
    .X(_0146_));
 sg13g2_o21ai_1 _4738_ (.B1(_1488_),
    .Y(_1499_),
    .A1(_1466_),
    .A2(_1489_));
 sg13g2_o21ai_1 _4739_ (.B1(_1471_),
    .Y(_1500_),
    .A1(_1468_),
    .A2(_1472_));
 sg13g2_nand2_1 _4740_ (.Y(_1501_),
    .A(net925),
    .B(net1044));
 sg13g2_nand2_1 _4741_ (.Y(_1502_),
    .A(net921),
    .B(net851));
 sg13g2_and4_1 _4742_ (.A(net922),
    .B(net921),
    .C(net854),
    .D(net851),
    .X(_1503_));
 sg13g2_a22oi_1 _4743_ (.Y(_1504_),
    .B1(net851),
    .B2(net922),
    .A2(net854),
    .A1(net921));
 sg13g2_or2_1 _4744_ (.X(_1505_),
    .B(_1504_),
    .A(_1503_));
 sg13g2_nor2_1 _4745_ (.A(_1501_),
    .B(_1505_),
    .Y(_1506_));
 sg13g2_xor2_1 _4746_ (.B(_1505_),
    .A(_1501_),
    .X(_1507_));
 sg13g2_nand2_1 _4747_ (.Y(_1508_),
    .A(_1500_),
    .B(_1507_));
 sg13g2_xnor2_1 _4748_ (.Y(_1509_),
    .A(_1500_),
    .B(_1507_));
 sg13g2_xnor2_1 _4749_ (.Y(_1510_),
    .A(_1463_),
    .B(_1509_));
 sg13g2_o21ai_1 _4750_ (.B1(_1483_),
    .Y(_1511_),
    .A1(_1474_),
    .A2(_1484_));
 sg13g2_nand2_1 _4751_ (.Y(_1512_),
    .A(net919),
    .B(net856));
 sg13g2_nand2_2 _4752_ (.Y(_1513_),
    .A(net857),
    .B(net914));
 sg13g2_nand2_1 _4753_ (.Y(_1514_),
    .A(net859),
    .B(net915));
 sg13g2_or2_1 _4754_ (.X(_1515_),
    .B(_1513_),
    .A(_1470_));
 sg13g2_xnor2_1 _4755_ (.Y(_1516_),
    .A(_1469_),
    .B(_1514_));
 sg13g2_xnor2_1 _4756_ (.Y(_1517_),
    .A(_1512_),
    .B(_1516_));
 sg13g2_o21ai_1 _4757_ (.B1(_1478_),
    .Y(_1518_),
    .A1(_1476_),
    .A2(_1479_));
 sg13g2_nand2_1 _4758_ (.Y(_1519_),
    .A(net861),
    .B(net911));
 sg13g2_and4_1 _4759_ (.A(net867),
    .B(net866),
    .C(net909),
    .D(net1049),
    .X(_1520_));
 sg13g2_nand4_1 _4760_ (.B(net864),
    .C(net909),
    .A(net867),
    .Y(_1521_),
    .D(net1049));
 sg13g2_a22oi_1 _4761_ (.Y(_1522_),
    .B1(net1049),
    .B2(net867),
    .A2(net909),
    .A1(net864));
 sg13g2_or3_1 _4762_ (.A(_1519_),
    .B(_1520_),
    .C(_1522_),
    .X(_1523_));
 sg13g2_o21ai_1 _4763_ (.B1(_1519_),
    .Y(_1524_),
    .A1(_1520_),
    .A2(_1522_));
 sg13g2_and3_1 _4764_ (.X(_1525_),
    .A(_1518_),
    .B(_1523_),
    .C(_1524_));
 sg13g2_nand3_1 _4765_ (.B(_1523_),
    .C(_1524_),
    .A(_1518_),
    .Y(_1526_));
 sg13g2_a21oi_1 _4766_ (.A1(_1523_),
    .A2(_1524_),
    .Y(_1527_),
    .B1(_1518_));
 sg13g2_or3_1 _4767_ (.A(_1517_),
    .B(_1525_),
    .C(_1527_),
    .X(_1528_));
 sg13g2_o21ai_1 _4768_ (.B1(_1517_),
    .Y(_1529_),
    .A1(_1525_),
    .A2(_1527_));
 sg13g2_and3_1 _4769_ (.X(_1530_),
    .A(_1511_),
    .B(_1528_),
    .C(_1529_));
 sg13g2_nand3_1 _4770_ (.B(_1528_),
    .C(_1529_),
    .A(_1511_),
    .Y(_1531_));
 sg13g2_a21oi_1 _4771_ (.A1(_1528_),
    .A2(_1529_),
    .Y(_1532_),
    .B1(_1511_));
 sg13g2_or3_1 _4772_ (.A(_1510_),
    .B(_1530_),
    .C(_1532_),
    .X(_1533_));
 sg13g2_o21ai_1 _4773_ (.B1(_1510_),
    .Y(_1534_),
    .A1(_1530_),
    .A2(_1532_));
 sg13g2_and3_1 _4774_ (.X(_1535_),
    .A(_1499_),
    .B(_1533_),
    .C(_1534_));
 sg13g2_nand3_1 _4775_ (.B(_1533_),
    .C(_1534_),
    .A(_1499_),
    .Y(_1536_));
 sg13g2_a21oi_1 _4776_ (.A1(_1533_),
    .A2(_1534_),
    .Y(_1537_),
    .B1(_1499_));
 sg13g2_or3_1 _4777_ (.A(_1465_),
    .B(_1535_),
    .C(_1537_),
    .X(_1538_));
 sg13g2_o21ai_1 _4778_ (.B1(_1465_),
    .Y(_1539_),
    .A1(_1535_),
    .A2(_1537_));
 sg13g2_o21ai_1 _4779_ (.B1(_1492_),
    .Y(_1540_),
    .A1(_1431_),
    .A2(_1493_));
 sg13g2_nand3_1 _4780_ (.B(_1539_),
    .C(_1540_),
    .A(_1538_),
    .Y(_1541_));
 sg13g2_a21o_1 _4781_ (.A2(_1539_),
    .A1(_1538_),
    .B1(_1540_),
    .X(_1542_));
 sg13g2_nand2_1 _4782_ (.Y(_1543_),
    .A(_1541_),
    .B(_1542_));
 sg13g2_and4_1 _4783_ (.A(_1496_),
    .B(_1497_),
    .C(_1541_),
    .D(_1542_),
    .X(_1544_));
 sg13g2_xor2_1 _4784_ (.B(_1543_),
    .A(_1498_),
    .X(_0147_));
 sg13g2_o21ai_1 _4785_ (.B1(_1541_),
    .Y(_1545_),
    .A1(_1498_),
    .A2(_1543_));
 sg13g2_o21ai_1 _4786_ (.B1(_1536_),
    .Y(_1546_),
    .A1(_1465_),
    .A2(_1537_));
 sg13g2_o21ai_1 _4787_ (.B1(_1508_),
    .Y(_1547_),
    .A1(_1463_),
    .A2(_1509_));
 sg13g2_o21ai_1 _4788_ (.B1(_1531_),
    .Y(_1548_),
    .A1(_1510_),
    .A2(_1532_));
 sg13g2_nor2_1 _4789_ (.A(_1503_),
    .B(_1506_),
    .Y(_1549_));
 sg13g2_o21ai_1 _4790_ (.B1(_1515_),
    .Y(_1550_),
    .A1(_1512_),
    .A2(_1516_));
 sg13g2_nand2_1 _4791_ (.Y(_1551_),
    .A(net922),
    .B(net1044));
 sg13g2_nand2_1 _4792_ (.Y(_1552_),
    .A(net919),
    .B(net851));
 sg13g2_nand2_1 _4793_ (.Y(_1553_),
    .A(net919),
    .B(net854));
 sg13g2_xor2_1 _4794_ (.B(_1553_),
    .A(_1502_),
    .X(_1554_));
 sg13g2_nand2b_1 _4795_ (.Y(_1555_),
    .B(_1554_),
    .A_N(_1551_));
 sg13g2_xnor2_1 _4796_ (.Y(_1556_),
    .A(_1551_),
    .B(_1554_));
 sg13g2_xnor2_1 _4797_ (.Y(_1557_),
    .A(_1550_),
    .B(_1556_));
 sg13g2_nor2_1 _4798_ (.A(_1549_),
    .B(_1557_),
    .Y(_1558_));
 sg13g2_xnor2_1 _4799_ (.Y(_1559_),
    .A(_1549_),
    .B(_1557_));
 sg13g2_o21ai_1 _4800_ (.B1(_1526_),
    .Y(_1560_),
    .A1(_1517_),
    .A2(_1527_));
 sg13g2_nand2_1 _4801_ (.Y(_1561_),
    .A(net917),
    .B(net856));
 sg13g2_nand2_1 _4802_ (.Y(_1562_),
    .A(net860),
    .B(net911));
 sg13g2_or2_1 _4803_ (.X(_1563_),
    .B(_1562_),
    .A(_1513_));
 sg13g2_and2_1 _4804_ (.A(_1513_),
    .B(_1562_),
    .X(_1564_));
 sg13g2_xnor2_1 _4805_ (.Y(_1565_),
    .A(_1513_),
    .B(_1562_));
 sg13g2_xnor2_1 _4806_ (.Y(_1566_),
    .A(_1561_),
    .B(_1565_));
 sg13g2_o21ai_1 _4807_ (.B1(_1521_),
    .Y(_1567_),
    .A1(_1519_),
    .A2(_1522_));
 sg13g2_nand2_1 _4808_ (.Y(_1568_),
    .A(net861),
    .B(net1049));
 sg13g2_and4_1 _4809_ (.A(net866),
    .B(net862),
    .C(net908),
    .D(net1050),
    .X(_1569_));
 sg13g2_a22oi_1 _4810_ (.Y(_1570_),
    .B1(net1049),
    .B2(net866),
    .A2(net908),
    .A1(net862));
 sg13g2_nor2_1 _4811_ (.A(_1569_),
    .B(_1570_),
    .Y(_1571_));
 sg13g2_nand2_1 _4812_ (.Y(_1572_),
    .A(_1567_),
    .B(_1571_));
 sg13g2_xnor2_1 _4813_ (.Y(_1573_),
    .A(_1567_),
    .B(_1571_));
 sg13g2_xor2_1 _4814_ (.B(_1573_),
    .A(_1566_),
    .X(_1574_));
 sg13g2_nand2_1 _4815_ (.Y(_1575_),
    .A(_1560_),
    .B(_1574_));
 sg13g2_xnor2_1 _4816_ (.Y(_1576_),
    .A(_1560_),
    .B(_1574_));
 sg13g2_xor2_1 _4817_ (.B(_1576_),
    .A(_1559_),
    .X(_1577_));
 sg13g2_nand2_1 _4818_ (.Y(_1578_),
    .A(_1548_),
    .B(_1577_));
 sg13g2_xnor2_1 _4819_ (.Y(_1579_),
    .A(_1548_),
    .B(_1577_));
 sg13g2_nand2b_1 _4820_ (.Y(_1580_),
    .B(_1547_),
    .A_N(_1579_));
 sg13g2_xnor2_1 _4821_ (.Y(_1581_),
    .A(_1547_),
    .B(_1579_));
 sg13g2_nor2_1 _4822_ (.A(_1546_),
    .B(_1581_),
    .Y(_1582_));
 sg13g2_nand2_1 _4823_ (.Y(_1583_),
    .A(_1546_),
    .B(_1581_));
 sg13g2_nor2b_1 _4824_ (.A(_1582_),
    .B_N(_1583_),
    .Y(_1584_));
 sg13g2_xor2_1 _4825_ (.B(_1584_),
    .A(_1545_),
    .X(_0148_));
 sg13g2_a21oi_1 _4826_ (.A1(_1550_),
    .A2(_1556_),
    .Y(_1585_),
    .B1(_1558_));
 sg13g2_o21ai_1 _4827_ (.B1(_1575_),
    .Y(_1586_),
    .A1(_1559_),
    .A2(_1576_));
 sg13g2_o21ai_1 _4828_ (.B1(_1555_),
    .Y(_1587_),
    .A1(_1502_),
    .A2(_1553_));
 sg13g2_o21ai_1 _4829_ (.B1(_1563_),
    .Y(_1588_),
    .A1(_1561_),
    .A2(_1564_));
 sg13g2_nand2_1 _4830_ (.Y(_1589_),
    .A(net921),
    .B(net1044));
 sg13g2_nand2_1 _4831_ (.Y(_1590_),
    .A(net917),
    .B(net852));
 sg13g2_nand2_1 _4832_ (.Y(_1591_),
    .A(net917),
    .B(net854));
 sg13g2_or2_1 _4833_ (.X(_1592_),
    .B(_1590_),
    .A(_1553_));
 sg13g2_xnor2_1 _4834_ (.Y(_1593_),
    .A(_1552_),
    .B(_1591_));
 sg13g2_xor2_1 _4835_ (.B(_1593_),
    .A(_1589_),
    .X(_1594_));
 sg13g2_xnor2_1 _4836_ (.Y(_1595_),
    .A(_1588_),
    .B(_1594_));
 sg13g2_nor2b_1 _4837_ (.A(_1595_),
    .B_N(_1587_),
    .Y(_1596_));
 sg13g2_xor2_1 _4838_ (.B(_1595_),
    .A(_1587_),
    .X(_1597_));
 sg13g2_o21ai_1 _4839_ (.B1(_1572_),
    .Y(_1598_),
    .A1(_1566_),
    .A2(_1573_));
 sg13g2_a21oi_1 _4840_ (.A1(net864),
    .A2(net908),
    .Y(_1599_),
    .B1(_1568_));
 sg13g2_nand2_1 _4841_ (.Y(_1600_),
    .A(net914),
    .B(net856));
 sg13g2_nand2_1 _4842_ (.Y(_1601_),
    .A(net858),
    .B(net908));
 sg13g2_and4_1 _4843_ (.A(net860),
    .B(net858),
    .C(net911),
    .D(net908),
    .X(_1602_));
 sg13g2_a22oi_1 _4844_ (.Y(_1603_),
    .B1(net910),
    .B2(net860),
    .A2(net911),
    .A1(net858));
 sg13g2_nor3_1 _4845_ (.A(_1600_),
    .B(_1602_),
    .C(_1603_),
    .Y(_1604_));
 sg13g2_o21ai_1 _4846_ (.B1(_1600_),
    .Y(_1605_),
    .A1(_1602_),
    .A2(_1603_));
 sg13g2_nor2b_1 _4847_ (.A(_1604_),
    .B_N(_1605_),
    .Y(_1606_));
 sg13g2_xnor2_1 _4848_ (.Y(_1607_),
    .A(_1599_),
    .B(_1606_));
 sg13g2_nand2b_1 _4849_ (.Y(_1608_),
    .B(_1598_),
    .A_N(_1607_));
 sg13g2_xor2_1 _4850_ (.B(_1607_),
    .A(_1598_),
    .X(_1609_));
 sg13g2_xor2_1 _4851_ (.B(_1609_),
    .A(_1597_),
    .X(_1610_));
 sg13g2_nand2_1 _4852_ (.Y(_1611_),
    .A(_1586_),
    .B(_1610_));
 sg13g2_xor2_1 _4853_ (.B(_1610_),
    .A(_1586_),
    .X(_1612_));
 sg13g2_nand2b_1 _4854_ (.Y(_1613_),
    .B(_1612_),
    .A_N(_1585_));
 sg13g2_xor2_1 _4855_ (.B(_1612_),
    .A(_1585_),
    .X(_1614_));
 sg13g2_a21oi_1 _4856_ (.A1(_1578_),
    .A2(_1580_),
    .Y(_1615_),
    .B1(_1614_));
 sg13g2_nand3_1 _4857_ (.B(_1580_),
    .C(_1614_),
    .A(_1578_),
    .Y(_1616_));
 sg13g2_nand2b_1 _4858_ (.Y(_1617_),
    .B(_1616_),
    .A_N(_1615_));
 sg13g2_a21oi_1 _4859_ (.A1(_1541_),
    .A2(_1583_),
    .Y(_1618_),
    .B1(_1582_));
 sg13g2_a21oi_2 _4860_ (.B1(_1618_),
    .Y(_1619_),
    .A2(_1584_),
    .A1(_1544_));
 sg13g2_nor2_1 _4861_ (.A(_1617_),
    .B(_1619_),
    .Y(_1620_));
 sg13g2_xor2_1 _4862_ (.B(_1619_),
    .A(_1617_),
    .X(_0139_));
 sg13g2_a21o_1 _4863_ (.A2(_1594_),
    .A1(_1588_),
    .B1(_1596_),
    .X(_1621_));
 sg13g2_o21ai_1 _4864_ (.B1(_1608_),
    .Y(_1622_),
    .A1(_1597_),
    .A2(_1609_));
 sg13g2_a21o_2 _4865_ (.A2(_1606_),
    .A1(_1599_),
    .B1(_1569_),
    .X(_1623_));
 sg13g2_nand2_1 _4866_ (.Y(_1624_),
    .A(net856),
    .B(net912));
 sg13g2_nand2_1 _4867_ (.Y(_1625_),
    .A(net860),
    .B(net1049));
 sg13g2_or2_1 _4868_ (.X(_1626_),
    .B(_1625_),
    .A(_1601_));
 sg13g2_xnor2_1 _4869_ (.Y(_1627_),
    .A(_1601_),
    .B(_1625_));
 sg13g2_xor2_1 _4870_ (.B(_1627_),
    .A(_1624_),
    .X(_1628_));
 sg13g2_and2_1 _4871_ (.A(_1623_),
    .B(_1628_),
    .X(_1629_));
 sg13g2_or2_1 _4872_ (.X(_1630_),
    .B(_1628_),
    .A(_1623_));
 sg13g2_xnor2_1 _4873_ (.Y(_1631_),
    .A(_1623_),
    .B(_1628_));
 sg13g2_o21ai_1 _4874_ (.B1(_1592_),
    .Y(_1632_),
    .A1(_1589_),
    .A2(_1593_));
 sg13g2_or2_1 _4875_ (.X(_1633_),
    .B(_1604_),
    .A(_1602_));
 sg13g2_nand2_1 _4876_ (.Y(_1634_),
    .A(net919),
    .B(net1044));
 sg13g2_nand2_1 _4877_ (.Y(_1635_),
    .A(net914),
    .B(net854));
 sg13g2_or2_1 _4878_ (.X(_1636_),
    .B(_1635_),
    .A(_1590_));
 sg13g2_xnor2_1 _4879_ (.Y(_1637_),
    .A(_1590_),
    .B(_1635_));
 sg13g2_xor2_1 _4880_ (.B(_1637_),
    .A(_1634_),
    .X(_1638_));
 sg13g2_xnor2_1 _4881_ (.Y(_1639_),
    .A(_1633_),
    .B(_1638_));
 sg13g2_nor2b_1 _4882_ (.A(_1639_),
    .B_N(_1632_),
    .Y(_1640_));
 sg13g2_xnor2_1 _4883_ (.Y(_1641_),
    .A(_1632_),
    .B(_1639_));
 sg13g2_xnor2_1 _4884_ (.Y(_1642_),
    .A(_1631_),
    .B(_1641_));
 sg13g2_xnor2_1 _4885_ (.Y(_1643_),
    .A(_1622_),
    .B(_1642_));
 sg13g2_nor2b_1 _4886_ (.A(_1643_),
    .B_N(_1621_),
    .Y(_1644_));
 sg13g2_xor2_1 _4887_ (.B(_1643_),
    .A(_1621_),
    .X(_1645_));
 sg13g2_nand3_1 _4888_ (.B(_1613_),
    .C(_1645_),
    .A(_1611_),
    .Y(_1646_));
 sg13g2_a21oi_1 _4889_ (.A1(_1611_),
    .A2(_1613_),
    .Y(_1647_),
    .B1(_1645_));
 sg13g2_inv_1 _4890_ (.Y(_1648_),
    .A(_1647_));
 sg13g2_nand2_1 _4891_ (.Y(_1649_),
    .A(_1646_),
    .B(_1648_));
 sg13g2_nor2_1 _4892_ (.A(_1615_),
    .B(_1620_),
    .Y(_1650_));
 sg13g2_xor2_1 _4893_ (.B(_1650_),
    .A(_1649_),
    .X(_0140_));
 sg13g2_a21o_1 _4894_ (.A2(_1638_),
    .A1(_1633_),
    .B1(_1640_),
    .X(_1651_));
 sg13g2_a22oi_1 _4895_ (.Y(_1652_),
    .B1(net1049),
    .B2(net858),
    .A2(net908),
    .A1(net856));
 sg13g2_nand2_2 _4896_ (.Y(_1653_),
    .A(\DP_4.matrix[5] ),
    .B(net1049));
 sg13g2_or2_1 _4897_ (.X(_1654_),
    .B(_1653_),
    .A(_1601_));
 sg13g2_nand2b_1 _4898_ (.Y(_1655_),
    .B(_1654_),
    .A_N(_1652_));
 sg13g2_o21ai_1 _4899_ (.B1(_1636_),
    .Y(_1656_),
    .A1(_1634_),
    .A2(_1637_));
 sg13g2_o21ai_1 _4900_ (.B1(_1626_),
    .Y(_1657_),
    .A1(_1624_),
    .A2(_1627_));
 sg13g2_nand2_1 _4901_ (.Y(_1658_),
    .A(net917),
    .B(net1044));
 sg13g2_nand2_1 _4902_ (.Y(_1659_),
    .A(net912),
    .B(net852));
 sg13g2_and4_1 _4903_ (.A(net914),
    .B(net911),
    .C(net854),
    .D(net852),
    .X(_1660_));
 sg13g2_or2_1 _4904_ (.X(_1661_),
    .B(_1659_),
    .A(_1635_));
 sg13g2_a22oi_1 _4905_ (.Y(_1662_),
    .B1(net852),
    .B2(\DP_3.matrix[5] ),
    .A2(net855),
    .A1(net912));
 sg13g2_nor2_1 _4906_ (.A(_1660_),
    .B(_1662_),
    .Y(_1663_));
 sg13g2_xnor2_1 _4907_ (.Y(_1664_),
    .A(_1658_),
    .B(_1663_));
 sg13g2_xnor2_1 _4908_ (.Y(_1665_),
    .A(_1657_),
    .B(_1664_));
 sg13g2_nor2b_1 _4909_ (.A(_1665_),
    .B_N(_1656_),
    .Y(_1666_));
 sg13g2_xor2_1 _4910_ (.B(_1665_),
    .A(_1656_),
    .X(_1667_));
 sg13g2_or2_1 _4911_ (.X(_1668_),
    .B(_1667_),
    .A(_1655_));
 sg13g2_xor2_1 _4912_ (.B(_1667_),
    .A(_1655_),
    .X(_1669_));
 sg13g2_a21oi_1 _4913_ (.A1(_1630_),
    .A2(_1641_),
    .Y(_1670_),
    .B1(_1629_));
 sg13g2_nor2b_1 _4914_ (.A(_1670_),
    .B_N(_1669_),
    .Y(_1671_));
 sg13g2_xor2_1 _4915_ (.B(_1670_),
    .A(_1669_),
    .X(_1672_));
 sg13g2_nor2b_1 _4916_ (.A(_1672_),
    .B_N(_1651_),
    .Y(_1673_));
 sg13g2_xor2_1 _4917_ (.B(_1672_),
    .A(_1651_),
    .X(_1674_));
 sg13g2_a21oi_1 _4918_ (.A1(_1622_),
    .A2(_1642_),
    .Y(_1675_),
    .B1(_1644_));
 sg13g2_nor2_1 _4919_ (.A(_1674_),
    .B(_1675_),
    .Y(_1676_));
 sg13g2_xor2_1 _4920_ (.B(_1675_),
    .A(_1674_),
    .X(_1677_));
 sg13g2_a21oi_1 _4921_ (.A1(_1615_),
    .A2(_1646_),
    .Y(_1678_),
    .B1(_1647_));
 sg13g2_nand2_1 _4922_ (.Y(_1679_),
    .A(_1616_),
    .B(_1646_));
 sg13g2_a22oi_1 _4923_ (.Y(_1680_),
    .B1(_1679_),
    .B2(_1648_),
    .A2(_1678_),
    .A1(_1619_));
 sg13g2_xor2_1 _4924_ (.B(_1680_),
    .A(_1677_),
    .X(_0141_));
 sg13g2_a21o_1 _4925_ (.A2(_1664_),
    .A1(_1657_),
    .B1(_1666_),
    .X(_1681_));
 sg13g2_o21ai_1 _4926_ (.B1(_1661_),
    .Y(_1682_),
    .A1(_1658_),
    .A2(_1662_));
 sg13g2_nand2_1 _4927_ (.Y(_1683_),
    .A(net915),
    .B(net1044));
 sg13g2_nand2_1 _4928_ (.Y(_1684_),
    .A(net909),
    .B(net851));
 sg13g2_nand2_1 _4929_ (.Y(_1685_),
    .A(net855),
    .B(net908));
 sg13g2_xor2_1 _4930_ (.B(_1685_),
    .A(_1659_),
    .X(_1686_));
 sg13g2_nand2b_1 _4931_ (.Y(_1687_),
    .B(_1686_),
    .A_N(_1683_));
 sg13g2_xnor2_1 _4932_ (.Y(_1688_),
    .A(_1683_),
    .B(_1686_));
 sg13g2_nor2b_1 _4933_ (.A(_1654_),
    .B_N(_1688_),
    .Y(_1689_));
 sg13g2_xnor2_1 _4934_ (.Y(_1690_),
    .A(_1654_),
    .B(_1688_));
 sg13g2_xnor2_1 _4935_ (.Y(_1691_),
    .A(_1682_),
    .B(_1690_));
 sg13g2_nor2_1 _4936_ (.A(_1653_),
    .B(_1691_),
    .Y(_1692_));
 sg13g2_xnor2_1 _4937_ (.Y(_1693_),
    .A(_1653_),
    .B(_1691_));
 sg13g2_nor2_1 _4938_ (.A(_1668_),
    .B(_1693_),
    .Y(_1694_));
 sg13g2_xor2_1 _4939_ (.B(_1693_),
    .A(_1668_),
    .X(_1695_));
 sg13g2_xor2_1 _4940_ (.B(_1695_),
    .A(_1681_),
    .X(_1696_));
 sg13g2_o21ai_1 _4941_ (.B1(_1696_),
    .Y(_1697_),
    .A1(_1671_),
    .A2(_1673_));
 sg13g2_or3_1 _4942_ (.A(_1671_),
    .B(_1673_),
    .C(_1696_),
    .X(_1698_));
 sg13g2_and2_1 _4943_ (.A(_1697_),
    .B(_1698_),
    .X(_1699_));
 sg13g2_a21oi_1 _4944_ (.A1(_1677_),
    .A2(_1680_),
    .Y(_1700_),
    .B1(_1676_));
 sg13g2_xnor2_1 _4945_ (.Y(_0142_),
    .A(_1699_),
    .B(_1700_));
 sg13g2_nand2_1 _4946_ (.Y(_1701_),
    .A(_1677_),
    .B(_1699_));
 sg13g2_a221oi_1 _4947_ (.B2(_1648_),
    .C1(_1701_),
    .B1(_1679_),
    .A1(_1619_),
    .Y(_1702_),
    .A2(_1678_));
 sg13g2_nand2_1 _4948_ (.Y(_1703_),
    .A(_1676_),
    .B(_1698_));
 sg13g2_nand2_1 _4949_ (.Y(_1704_),
    .A(_1697_),
    .B(_1703_));
 sg13g2_a21oi_1 _4950_ (.A1(_1681_),
    .A2(_1695_),
    .Y(_1705_),
    .B1(_1694_));
 sg13g2_a21o_1 _4951_ (.A2(_1690_),
    .A1(_1682_),
    .B1(_1689_),
    .X(_1706_));
 sg13g2_o21ai_1 _4952_ (.B1(_1687_),
    .Y(_1707_),
    .A1(_1659_),
    .A2(_1685_));
 sg13g2_nand2_1 _4953_ (.Y(_1708_),
    .A(net912),
    .B(\DP_4.matrix[8] ));
 sg13g2_nand2_1 _4954_ (.Y(_1709_),
    .A(net851),
    .B(net1050));
 sg13g2_nand2_1 _4955_ (.Y(_1710_),
    .A(net855),
    .B(net1050));
 sg13g2_xor2_1 _4956_ (.B(_1710_),
    .A(_1684_),
    .X(_1711_));
 sg13g2_nand2b_1 _4957_ (.Y(_1712_),
    .B(_1711_),
    .A_N(_1708_));
 sg13g2_xnor2_1 _4958_ (.Y(_1713_),
    .A(_1708_),
    .B(_1711_));
 sg13g2_nand2_1 _4959_ (.Y(_1714_),
    .A(_1707_),
    .B(_1713_));
 sg13g2_xor2_1 _4960_ (.B(_1713_),
    .A(_1707_),
    .X(_1715_));
 sg13g2_xnor2_1 _4961_ (.Y(_1716_),
    .A(_1692_),
    .B(_1715_));
 sg13g2_nor2b_1 _4962_ (.A(_1716_),
    .B_N(_1706_),
    .Y(_1717_));
 sg13g2_xor2_1 _4963_ (.B(_1716_),
    .A(_1706_),
    .X(_1718_));
 sg13g2_xor2_1 _4964_ (.B(_1718_),
    .A(_1705_),
    .X(_1719_));
 sg13g2_o21ai_1 _4965_ (.B1(_1719_),
    .Y(_1720_),
    .A1(_1702_),
    .A2(_1704_));
 sg13g2_or3_1 _4966_ (.A(_1702_),
    .B(_1704_),
    .C(_1719_),
    .X(_1721_));
 sg13g2_and2_1 _4967_ (.A(_1720_),
    .B(_1721_),
    .X(_0143_));
 sg13g2_o21ai_1 _4968_ (.B1(_1720_),
    .Y(_1722_),
    .A1(_1705_),
    .A2(_1718_));
 sg13g2_a21oi_1 _4969_ (.A1(_1692_),
    .A2(_1715_),
    .Y(_1723_),
    .B1(_1717_));
 sg13g2_o21ai_1 _4970_ (.B1(_1712_),
    .Y(_1724_),
    .A1(_1684_),
    .A2(_1710_));
 sg13g2_nand2_1 _4971_ (.Y(_1725_),
    .A(net908),
    .B(\DP_4.matrix[8] ));
 sg13g2_xor2_1 _4972_ (.B(_1725_),
    .A(_1709_),
    .X(_1726_));
 sg13g2_xnor2_1 _4973_ (.Y(_1727_),
    .A(_1724_),
    .B(_1726_));
 sg13g2_xnor2_1 _4974_ (.Y(_1728_),
    .A(_1714_),
    .B(_1727_));
 sg13g2_xnor2_1 _4975_ (.Y(_1729_),
    .A(_1723_),
    .B(_1728_));
 sg13g2_xnor2_1 _4976_ (.Y(_0144_),
    .A(_1722_),
    .B(_1729_));
 sg13g2_and2_1 _4977_ (.A(net890),
    .B(net832),
    .X(_0089_));
 sg13g2_and3_2 _4978_ (.X(_1730_),
    .A(net888),
    .B(net827),
    .C(_0089_));
 sg13g2_a22oi_1 _4979_ (.Y(_1731_),
    .B1(net827),
    .B2(net890),
    .A2(net888),
    .A1(net832));
 sg13g2_nor2_1 _4980_ (.A(_1730_),
    .B(_1731_),
    .Y(_0090_));
 sg13g2_nand2_1 _4981_ (.Y(_1732_),
    .A(net890),
    .B(net822));
 sg13g2_and4_1 _4982_ (.A(net830),
    .B(net887),
    .C(net825),
    .D(net884),
    .X(_1733_));
 sg13g2_a22oi_1 _4983_ (.Y(_1734_),
    .B1(net884),
    .B2(net831),
    .A2(net826),
    .A1(net887));
 sg13g2_nor3_1 _4984_ (.A(_1732_),
    .B(_1733_),
    .C(_1734_),
    .Y(_1735_));
 sg13g2_o21ai_1 _4985_ (.B1(_1732_),
    .Y(_1736_),
    .A1(_1733_),
    .A2(_1734_));
 sg13g2_nor2b_1 _4986_ (.A(_1735_),
    .B_N(_1736_),
    .Y(_1737_));
 sg13g2_nand2_1 _4987_ (.Y(_1738_),
    .A(_1730_),
    .B(_1737_));
 sg13g2_xor2_1 _4988_ (.B(_1737_),
    .A(_1730_),
    .X(_0091_));
 sg13g2_nand2_1 _4989_ (.Y(_1739_),
    .A(net889),
    .B(net820));
 sg13g2_or2_1 _4990_ (.X(_1740_),
    .B(_1735_),
    .A(_1733_));
 sg13g2_nand2_1 _4991_ (.Y(_1741_),
    .A(net887),
    .B(net822));
 sg13g2_and4_1 _4992_ (.A(net828),
    .B(net825),
    .C(net883),
    .D(net880),
    .X(_1742_));
 sg13g2_nand4_1 _4993_ (.B(net825),
    .C(net883),
    .A(net830),
    .Y(_1743_),
    .D(net880));
 sg13g2_a22oi_1 _4994_ (.Y(_1744_),
    .B1(net880),
    .B2(net830),
    .A2(net883),
    .A1(net825));
 sg13g2_nor3_1 _4995_ (.A(_1741_),
    .B(_1742_),
    .C(_1744_),
    .Y(_1745_));
 sg13g2_o21ai_1 _4996_ (.B1(_1741_),
    .Y(_1746_),
    .A1(_1742_),
    .A2(_1744_));
 sg13g2_nor2b_1 _4997_ (.A(_1745_),
    .B_N(_1746_),
    .Y(_1747_));
 sg13g2_nand2_1 _4998_ (.Y(_1748_),
    .A(_1740_),
    .B(_1747_));
 sg13g2_xnor2_1 _4999_ (.Y(_1749_),
    .A(_1740_),
    .B(_1747_));
 sg13g2_xor2_1 _5000_ (.B(_1749_),
    .A(_1739_),
    .X(_1750_));
 sg13g2_nand2b_1 _5001_ (.Y(_1751_),
    .B(_1750_),
    .A_N(_1738_));
 sg13g2_xnor2_1 _5002_ (.Y(_0092_),
    .A(_1738_),
    .B(_1750_));
 sg13g2_a22oi_1 _5003_ (.Y(_1752_),
    .B1(net818),
    .B2(net889),
    .A2(net820),
    .A1(net886));
 sg13g2_nand2_1 _5004_ (.Y(_1753_),
    .A(net886),
    .B(net818));
 sg13g2_and4_1 _5005_ (.A(net889),
    .B(net886),
    .C(net820),
    .D(net818),
    .X(_1754_));
 sg13g2_nor2_1 _5006_ (.A(_1752_),
    .B(_1754_),
    .Y(_1755_));
 sg13g2_inv_1 _5007_ (.Y(_1756_),
    .A(_1755_));
 sg13g2_o21ai_1 _5008_ (.B1(_1743_),
    .Y(_1757_),
    .A1(_1741_),
    .A2(_1744_));
 sg13g2_nand2_1 _5009_ (.Y(_1758_),
    .A(net883),
    .B(net822));
 sg13g2_and4_1 _5010_ (.A(net828),
    .B(net825),
    .C(net881),
    .D(net877),
    .X(_1759_));
 sg13g2_nand4_1 _5011_ (.B(net825),
    .C(net880),
    .A(net828),
    .Y(_1760_),
    .D(net877));
 sg13g2_a22oi_1 _5012_ (.Y(_1761_),
    .B1(net877),
    .B2(net828),
    .A2(net881),
    .A1(net825));
 sg13g2_or3_1 _5013_ (.A(_1758_),
    .B(_1759_),
    .C(_1761_),
    .X(_1762_));
 sg13g2_o21ai_1 _5014_ (.B1(_1758_),
    .Y(_1763_),
    .A1(_1759_),
    .A2(_1761_));
 sg13g2_nand3_1 _5015_ (.B(_1762_),
    .C(_1763_),
    .A(_1757_),
    .Y(_1764_));
 sg13g2_a21oi_1 _5016_ (.A1(_1762_),
    .A2(_1763_),
    .Y(_1765_),
    .B1(_1757_));
 sg13g2_a21o_1 _5017_ (.A2(_1763_),
    .A1(_1762_),
    .B1(_1757_),
    .X(_1766_));
 sg13g2_nand2_1 _5018_ (.Y(_1767_),
    .A(_1764_),
    .B(_1766_));
 sg13g2_xnor2_1 _5019_ (.Y(_1768_),
    .A(_1756_),
    .B(_1767_));
 sg13g2_o21ai_1 _5020_ (.B1(_1748_),
    .Y(_1769_),
    .A1(_1739_),
    .A2(_1749_));
 sg13g2_nor2b_2 _5021_ (.A(_1768_),
    .B_N(_1769_),
    .Y(_1770_));
 sg13g2_xor2_1 _5022_ (.B(_1769_),
    .A(_1768_),
    .X(_1771_));
 sg13g2_or2_1 _5023_ (.X(_1772_),
    .B(_1771_),
    .A(_1751_));
 sg13g2_xor2_1 _5024_ (.B(_1771_),
    .A(_1751_),
    .X(_0093_));
 sg13g2_o21ai_1 _5025_ (.B1(_1764_),
    .Y(_1773_),
    .A1(_1756_),
    .A2(_1765_));
 sg13g2_nand2_1 _5026_ (.Y(_1774_),
    .A(net889),
    .B(net816));
 sg13g2_nand2_1 _5027_ (.Y(_1775_),
    .A(net883),
    .B(net818));
 sg13g2_nand2_1 _5028_ (.Y(_1776_),
    .A(net883),
    .B(net820));
 sg13g2_xor2_1 _5029_ (.B(_1776_),
    .A(_1753_),
    .X(_1777_));
 sg13g2_nand2b_1 _5030_ (.Y(_1778_),
    .B(_1777_),
    .A_N(_1774_));
 sg13g2_xor2_1 _5031_ (.B(_1777_),
    .A(_1774_),
    .X(_1779_));
 sg13g2_o21ai_1 _5032_ (.B1(_1760_),
    .Y(_1780_),
    .A1(_1758_),
    .A2(_1761_));
 sg13g2_nand2_1 _5033_ (.Y(_1781_),
    .A(net822),
    .B(net880));
 sg13g2_and4_1 _5034_ (.A(net828),
    .B(net824),
    .C(net878),
    .D(net875),
    .X(_1782_));
 sg13g2_nand4_1 _5035_ (.B(net824),
    .C(net877),
    .A(net829),
    .Y(_1783_),
    .D(net875));
 sg13g2_a22oi_1 _5036_ (.Y(_1784_),
    .B1(net875),
    .B2(net828),
    .A2(net877),
    .A1(net824));
 sg13g2_or3_1 _5037_ (.A(_1781_),
    .B(_1782_),
    .C(_1784_),
    .X(_1785_));
 sg13g2_o21ai_1 _5038_ (.B1(_1781_),
    .Y(_1786_),
    .A1(_1782_),
    .A2(_1784_));
 sg13g2_and3_1 _5039_ (.X(_1787_),
    .A(_1780_),
    .B(_1785_),
    .C(_1786_));
 sg13g2_nand3_1 _5040_ (.B(_1785_),
    .C(_1786_),
    .A(_1780_),
    .Y(_1788_));
 sg13g2_a21oi_1 _5041_ (.A1(_1785_),
    .A2(_1786_),
    .Y(_1789_),
    .B1(_1780_));
 sg13g2_or3_1 _5042_ (.A(_1779_),
    .B(_1787_),
    .C(_1789_),
    .X(_1790_));
 sg13g2_o21ai_1 _5043_ (.B1(_1779_),
    .Y(_1791_),
    .A1(_1787_),
    .A2(_1789_));
 sg13g2_nand3_1 _5044_ (.B(_1790_),
    .C(_1791_),
    .A(_1773_),
    .Y(_1792_));
 sg13g2_a21o_1 _5045_ (.A2(_1791_),
    .A1(_1790_),
    .B1(_1773_),
    .X(_1793_));
 sg13g2_nand3_1 _5046_ (.B(_1792_),
    .C(_1793_),
    .A(_1754_),
    .Y(_1794_));
 sg13g2_a21o_1 _5047_ (.A2(_1793_),
    .A1(_1792_),
    .B1(_1754_),
    .X(_1795_));
 sg13g2_and2_1 _5048_ (.A(_1794_),
    .B(_1795_),
    .X(_1796_));
 sg13g2_nand3_1 _5049_ (.B(_1794_),
    .C(_1795_),
    .A(_1770_),
    .Y(_1797_));
 sg13g2_a21oi_1 _5050_ (.A1(_1794_),
    .A2(_1795_),
    .Y(_1798_),
    .B1(_1770_));
 sg13g2_xor2_1 _5051_ (.B(_1796_),
    .A(_1770_),
    .X(_1799_));
 sg13g2_xnor2_1 _5052_ (.Y(_0149_),
    .A(_1772_),
    .B(_1799_));
 sg13g2_nand2_1 _5053_ (.Y(_1800_),
    .A(_1792_),
    .B(_1794_));
 sg13g2_o21ai_1 _5054_ (.B1(_1778_),
    .Y(_1801_),
    .A1(_1753_),
    .A2(_1776_));
 sg13g2_nand2_1 _5055_ (.Y(_1802_),
    .A(net889),
    .B(net814));
 sg13g2_nand2b_1 _5056_ (.Y(_1803_),
    .B(_1801_),
    .A_N(_1802_));
 sg13g2_xor2_1 _5057_ (.B(_1802_),
    .A(_1801_),
    .X(_1804_));
 sg13g2_o21ai_1 _5058_ (.B1(_1788_),
    .Y(_1805_),
    .A1(_1779_),
    .A2(_1789_));
 sg13g2_nand2_1 _5059_ (.Y(_1806_),
    .A(net886),
    .B(net816));
 sg13g2_nand2_1 _5060_ (.Y(_1807_),
    .A(net880),
    .B(net818));
 sg13g2_nand2_1 _5061_ (.Y(_1808_),
    .A(net880),
    .B(net820));
 sg13g2_xor2_1 _5062_ (.B(_1808_),
    .A(_1775_),
    .X(_1809_));
 sg13g2_nand2b_1 _5063_ (.Y(_1810_),
    .B(_1809_),
    .A_N(_1806_));
 sg13g2_xnor2_1 _5064_ (.Y(_1811_),
    .A(_1806_),
    .B(_1809_));
 sg13g2_o21ai_1 _5065_ (.B1(_1783_),
    .Y(_1812_),
    .A1(_1781_),
    .A2(_1784_));
 sg13g2_nand2_1 _5066_ (.Y(_1813_),
    .A(net822),
    .B(net877));
 sg13g2_and4_1 _5067_ (.A(net829),
    .B(net824),
    .C(net875),
    .D(net873),
    .X(_1814_));
 sg13g2_nand4_1 _5068_ (.B(net824),
    .C(net875),
    .A(net828),
    .Y(_1815_),
    .D(net873));
 sg13g2_a22oi_1 _5069_ (.Y(_1816_),
    .B1(net873),
    .B2(net829),
    .A2(net875),
    .A1(net824));
 sg13g2_or3_1 _5070_ (.A(_1813_),
    .B(_1814_),
    .C(_1816_),
    .X(_1817_));
 sg13g2_o21ai_1 _5071_ (.B1(_1813_),
    .Y(_1818_),
    .A1(_1814_),
    .A2(_1816_));
 sg13g2_and3_1 _5072_ (.X(_1819_),
    .A(_1812_),
    .B(_1817_),
    .C(_1818_));
 sg13g2_nand3_1 _5073_ (.B(_1817_),
    .C(_1818_),
    .A(_1812_),
    .Y(_1820_));
 sg13g2_a21o_1 _5074_ (.A2(_1818_),
    .A1(_1817_),
    .B1(_1812_),
    .X(_1821_));
 sg13g2_nand3_1 _5075_ (.B(_1820_),
    .C(_1821_),
    .A(_1811_),
    .Y(_1822_));
 sg13g2_a21o_1 _5076_ (.A2(_1821_),
    .A1(_1820_),
    .B1(_1811_),
    .X(_1823_));
 sg13g2_nand3_1 _5077_ (.B(_1822_),
    .C(_1823_),
    .A(_1805_),
    .Y(_1824_));
 sg13g2_a21oi_1 _5078_ (.A1(_1822_),
    .A2(_1823_),
    .Y(_1825_),
    .B1(_1805_));
 sg13g2_a21o_1 _5079_ (.A2(_1823_),
    .A1(_1822_),
    .B1(_1805_),
    .X(_1826_));
 sg13g2_nand2_1 _5080_ (.Y(_1827_),
    .A(_1824_),
    .B(_1826_));
 sg13g2_xnor2_1 _5081_ (.Y(_1828_),
    .A(_1804_),
    .B(_1827_));
 sg13g2_nor2b_1 _5082_ (.A(_1828_),
    .B_N(_1800_),
    .Y(_1829_));
 sg13g2_xnor2_1 _5083_ (.Y(_1830_),
    .A(_1800_),
    .B(_1828_));
 sg13g2_o21ai_1 _5084_ (.B1(_1797_),
    .Y(_1831_),
    .A1(_1772_),
    .A2(_1798_));
 sg13g2_xor2_1 _5085_ (.B(_1831_),
    .A(_1830_),
    .X(_0156_));
 sg13g2_o21ai_1 _5086_ (.B1(_1824_),
    .Y(_1832_),
    .A1(_1804_),
    .A2(_1825_));
 sg13g2_o21ai_1 _5087_ (.B1(_1810_),
    .Y(_1833_),
    .A1(_1775_),
    .A2(_1808_));
 sg13g2_a22oi_1 _5088_ (.Y(_1834_),
    .B1(net811),
    .B2(net889),
    .A2(net814),
    .A1(net886));
 sg13g2_nand4_1 _5089_ (.B(net886),
    .C(net814),
    .A(net889),
    .Y(_1835_),
    .D(net811));
 sg13g2_nor2b_1 _5090_ (.A(_1834_),
    .B_N(_1835_),
    .Y(_1836_));
 sg13g2_nand2_1 _5091_ (.Y(_1837_),
    .A(_1833_),
    .B(_1836_));
 sg13g2_xnor2_1 _5092_ (.Y(_1838_),
    .A(_1833_),
    .B(_1836_));
 sg13g2_a21o_1 _5093_ (.A2(_1821_),
    .A1(_1811_),
    .B1(_1819_),
    .X(_1839_));
 sg13g2_nand2_1 _5094_ (.Y(_1840_),
    .A(net883),
    .B(net816));
 sg13g2_nand2_1 _5095_ (.Y(_1841_),
    .A(net877),
    .B(net818));
 sg13g2_nand2_1 _5096_ (.Y(_1842_),
    .A(net820),
    .B(net877));
 sg13g2_or2_1 _5097_ (.X(_1843_),
    .B(_1841_),
    .A(_1808_));
 sg13g2_and2_1 _5098_ (.A(_1807_),
    .B(_1842_),
    .X(_1844_));
 sg13g2_xnor2_1 _5099_ (.Y(_1845_),
    .A(_1807_),
    .B(_1842_));
 sg13g2_xnor2_1 _5100_ (.Y(_1846_),
    .A(_1840_),
    .B(_1845_));
 sg13g2_o21ai_1 _5101_ (.B1(_1815_),
    .Y(_1847_),
    .A1(_1813_),
    .A2(_1816_));
 sg13g2_nand2_1 _5102_ (.Y(_1848_),
    .A(net822),
    .B(net875));
 sg13g2_and4_1 _5103_ (.A(net829),
    .B(net824),
    .C(net873),
    .D(net870),
    .X(_1849_));
 sg13g2_nand4_1 _5104_ (.B(net824),
    .C(net873),
    .A(net828),
    .Y(_1850_),
    .D(net870));
 sg13g2_a22oi_1 _5105_ (.Y(_1851_),
    .B1(net870),
    .B2(net829),
    .A2(net873),
    .A1(net825));
 sg13g2_or3_1 _5106_ (.A(_1848_),
    .B(_1849_),
    .C(_1851_),
    .X(_1852_));
 sg13g2_o21ai_1 _5107_ (.B1(_1848_),
    .Y(_1853_),
    .A1(_1849_),
    .A2(_1851_));
 sg13g2_and3_1 _5108_ (.X(_1854_),
    .A(_1847_),
    .B(_1852_),
    .C(_1853_));
 sg13g2_nand3_1 _5109_ (.B(_1852_),
    .C(_1853_),
    .A(_1847_),
    .Y(_1855_));
 sg13g2_a21oi_1 _5110_ (.A1(_1852_),
    .A2(_1853_),
    .Y(_1856_),
    .B1(_1847_));
 sg13g2_or3_1 _5111_ (.A(_1846_),
    .B(_1854_),
    .C(_1856_),
    .X(_1857_));
 sg13g2_o21ai_1 _5112_ (.B1(_1846_),
    .Y(_1858_),
    .A1(_1854_),
    .A2(_1856_));
 sg13g2_and3_1 _5113_ (.X(_1859_),
    .A(_1839_),
    .B(_1857_),
    .C(_1858_));
 sg13g2_nand3_1 _5114_ (.B(_1857_),
    .C(_1858_),
    .A(_1839_),
    .Y(_1860_));
 sg13g2_a21oi_1 _5115_ (.A1(_1857_),
    .A2(_1858_),
    .Y(_1861_),
    .B1(_1839_));
 sg13g2_or3_1 _5116_ (.A(_1838_),
    .B(_1859_),
    .C(_1861_),
    .X(_1862_));
 sg13g2_o21ai_1 _5117_ (.B1(_1838_),
    .Y(_1863_),
    .A1(_1859_),
    .A2(_1861_));
 sg13g2_nand3_1 _5118_ (.B(_1862_),
    .C(_1863_),
    .A(_1832_),
    .Y(_1864_));
 sg13g2_a21oi_1 _5119_ (.A1(_1862_),
    .A2(_1863_),
    .Y(_1865_),
    .B1(_1832_));
 sg13g2_a21o_1 _5120_ (.A2(_1863_),
    .A1(_1862_),
    .B1(_1832_),
    .X(_1866_));
 sg13g2_nand2_1 _5121_ (.Y(_1867_),
    .A(_1864_),
    .B(_1866_));
 sg13g2_xor2_1 _5122_ (.B(_1867_),
    .A(_1803_),
    .X(_1868_));
 sg13g2_a21o_1 _5123_ (.A2(_1831_),
    .A1(_1830_),
    .B1(_1829_),
    .X(_1869_));
 sg13g2_nand2_1 _5124_ (.Y(_1870_),
    .A(_1868_),
    .B(_1869_));
 sg13g2_xor2_1 _5125_ (.B(_1869_),
    .A(_1868_),
    .X(_0157_));
 sg13g2_o21ai_1 _5126_ (.B1(_1860_),
    .Y(_1871_),
    .A1(_1838_),
    .A2(_1861_));
 sg13g2_o21ai_1 _5127_ (.B1(_1843_),
    .Y(_1872_),
    .A1(_1840_),
    .A2(_1844_));
 sg13g2_nand2_1 _5128_ (.Y(_1873_),
    .A(net889),
    .B(net1042));
 sg13g2_nand2_1 _5129_ (.Y(_1874_),
    .A(net884),
    .B(net811));
 sg13g2_and4_1 _5130_ (.A(net886),
    .B(net883),
    .C(net814),
    .D(net811),
    .X(_1875_));
 sg13g2_a22oi_1 _5131_ (.Y(_1876_),
    .B1(net811),
    .B2(net886),
    .A2(net814),
    .A1(net884));
 sg13g2_or2_1 _5132_ (.X(_1877_),
    .B(_1876_),
    .A(_1875_));
 sg13g2_nor2_1 _5133_ (.A(_1873_),
    .B(_1877_),
    .Y(_1878_));
 sg13g2_xor2_1 _5134_ (.B(_1877_),
    .A(_1873_),
    .X(_1879_));
 sg13g2_nand2_1 _5135_ (.Y(_1880_),
    .A(_1872_),
    .B(_1879_));
 sg13g2_xnor2_1 _5136_ (.Y(_1881_),
    .A(_1872_),
    .B(_1879_));
 sg13g2_xnor2_1 _5137_ (.Y(_1882_),
    .A(_1835_),
    .B(_1881_));
 sg13g2_o21ai_1 _5138_ (.B1(_1855_),
    .Y(_1883_),
    .A1(_1846_),
    .A2(_1856_));
 sg13g2_nand2_1 _5139_ (.Y(_1884_),
    .A(net880),
    .B(net816));
 sg13g2_nand2_2 _5140_ (.Y(_1885_),
    .A(net818),
    .B(net876));
 sg13g2_nand2_1 _5141_ (.Y(_1886_),
    .A(net820),
    .B(net875));
 sg13g2_or2_1 _5142_ (.X(_1887_),
    .B(_1885_),
    .A(_1842_));
 sg13g2_xnor2_1 _5143_ (.Y(_1888_),
    .A(_1841_),
    .B(_1886_));
 sg13g2_xnor2_1 _5144_ (.Y(_1889_),
    .A(_1884_),
    .B(_1888_));
 sg13g2_o21ai_1 _5145_ (.B1(_1850_),
    .Y(_1890_),
    .A1(_1848_),
    .A2(_1851_));
 sg13g2_nand2_1 _5146_ (.Y(_1891_),
    .A(net822),
    .B(net873));
 sg13g2_and4_1 _5147_ (.A(net831),
    .B(net826),
    .C(net870),
    .D(net1045),
    .X(_1892_));
 sg13g2_nand4_1 _5148_ (.B(net827),
    .C(net870),
    .A(net831),
    .Y(_1893_),
    .D(net1045));
 sg13g2_a22oi_1 _5149_ (.Y(_1894_),
    .B1(net1045),
    .B2(net831),
    .A2(net870),
    .A1(net826));
 sg13g2_or3_1 _5150_ (.A(_1891_),
    .B(_1892_),
    .C(_1894_),
    .X(_1895_));
 sg13g2_o21ai_1 _5151_ (.B1(_1891_),
    .Y(_1896_),
    .A1(_1892_),
    .A2(_1894_));
 sg13g2_and3_1 _5152_ (.X(_1897_),
    .A(_1890_),
    .B(_1895_),
    .C(_1896_));
 sg13g2_nand3_1 _5153_ (.B(_1895_),
    .C(_1896_),
    .A(_1890_),
    .Y(_1898_));
 sg13g2_a21oi_1 _5154_ (.A1(_1895_),
    .A2(_1896_),
    .Y(_1899_),
    .B1(_1890_));
 sg13g2_or3_1 _5155_ (.A(_1889_),
    .B(_1897_),
    .C(_1899_),
    .X(_1900_));
 sg13g2_o21ai_1 _5156_ (.B1(_1889_),
    .Y(_1901_),
    .A1(_1897_),
    .A2(_1899_));
 sg13g2_and3_1 _5157_ (.X(_1902_),
    .A(_1883_),
    .B(_1900_),
    .C(_1901_));
 sg13g2_nand3_1 _5158_ (.B(_1900_),
    .C(_1901_),
    .A(_1883_),
    .Y(_1903_));
 sg13g2_a21oi_1 _5159_ (.A1(_1900_),
    .A2(_1901_),
    .Y(_1904_),
    .B1(_1883_));
 sg13g2_or3_1 _5160_ (.A(_1882_),
    .B(_1902_),
    .C(_1904_),
    .X(_1905_));
 sg13g2_o21ai_1 _5161_ (.B1(_1882_),
    .Y(_1906_),
    .A1(_1902_),
    .A2(_1904_));
 sg13g2_and3_1 _5162_ (.X(_1907_),
    .A(_1871_),
    .B(_1905_),
    .C(_1906_));
 sg13g2_nand3_1 _5163_ (.B(_1905_),
    .C(_1906_),
    .A(_1871_),
    .Y(_1908_));
 sg13g2_a21oi_1 _5164_ (.A1(_1905_),
    .A2(_1906_),
    .Y(_1909_),
    .B1(_1871_));
 sg13g2_or3_1 _5165_ (.A(_1837_),
    .B(_1907_),
    .C(_1909_),
    .X(_1910_));
 sg13g2_o21ai_1 _5166_ (.B1(_1837_),
    .Y(_1911_),
    .A1(_1907_),
    .A2(_1909_));
 sg13g2_o21ai_1 _5167_ (.B1(_1864_),
    .Y(_1912_),
    .A1(_1803_),
    .A2(_1865_));
 sg13g2_nand3_1 _5168_ (.B(_1911_),
    .C(_1912_),
    .A(_1910_),
    .Y(_1913_));
 sg13g2_a21o_1 _5169_ (.A2(_1911_),
    .A1(_1910_),
    .B1(_1912_),
    .X(_1914_));
 sg13g2_nand2_1 _5170_ (.Y(_1915_),
    .A(_1913_),
    .B(_1914_));
 sg13g2_and4_1 _5171_ (.A(_1868_),
    .B(_1869_),
    .C(_1913_),
    .D(_1914_),
    .X(_1916_));
 sg13g2_xor2_1 _5172_ (.B(_1915_),
    .A(_1870_),
    .X(_0158_));
 sg13g2_o21ai_1 _5173_ (.B1(_1913_),
    .Y(_1917_),
    .A1(_1870_),
    .A2(_1915_));
 sg13g2_o21ai_1 _5174_ (.B1(_1908_),
    .Y(_1918_),
    .A1(_1837_),
    .A2(_1909_));
 sg13g2_o21ai_1 _5175_ (.B1(_1880_),
    .Y(_1919_),
    .A1(_1835_),
    .A2(_1881_));
 sg13g2_o21ai_1 _5176_ (.B1(_1903_),
    .Y(_1920_),
    .A1(_1882_),
    .A2(_1904_));
 sg13g2_nor2_1 _5177_ (.A(_1875_),
    .B(_1878_),
    .Y(_1921_));
 sg13g2_o21ai_1 _5178_ (.B1(_1887_),
    .Y(_1922_),
    .A1(_1884_),
    .A2(_1888_));
 sg13g2_nand2_1 _5179_ (.Y(_1923_),
    .A(net887),
    .B(net1042));
 sg13g2_nand2_1 _5180_ (.Y(_1924_),
    .A(net882),
    .B(net811));
 sg13g2_nand2_1 _5181_ (.Y(_1925_),
    .A(net881),
    .B(net814));
 sg13g2_xor2_1 _5182_ (.B(_1925_),
    .A(_1874_),
    .X(_1926_));
 sg13g2_nand2b_1 _5183_ (.Y(_1927_),
    .B(_1926_),
    .A_N(_1923_));
 sg13g2_xnor2_1 _5184_ (.Y(_1928_),
    .A(_1923_),
    .B(_1926_));
 sg13g2_xnor2_1 _5185_ (.Y(_1929_),
    .A(_1922_),
    .B(_1928_));
 sg13g2_nor2_1 _5186_ (.A(_1921_),
    .B(_1929_),
    .Y(_1930_));
 sg13g2_xnor2_1 _5187_ (.Y(_1931_),
    .A(_1921_),
    .B(_1929_));
 sg13g2_o21ai_1 _5188_ (.B1(_1898_),
    .Y(_1932_),
    .A1(_1889_),
    .A2(_1899_));
 sg13g2_nand2_1 _5189_ (.Y(_1933_),
    .A(net878),
    .B(net816));
 sg13g2_nand2_1 _5190_ (.Y(_1934_),
    .A(net820),
    .B(net873));
 sg13g2_or2_1 _5191_ (.X(_1935_),
    .B(_1934_),
    .A(_1885_));
 sg13g2_and2_1 _5192_ (.A(_1885_),
    .B(_1934_),
    .X(_1936_));
 sg13g2_xnor2_1 _5193_ (.Y(_1937_),
    .A(_1885_),
    .B(_1934_));
 sg13g2_xnor2_1 _5194_ (.Y(_1938_),
    .A(_1933_),
    .B(_1937_));
 sg13g2_o21ai_1 _5195_ (.B1(_1893_),
    .Y(_1939_),
    .A1(_1891_),
    .A2(_1894_));
 sg13g2_nand2_1 _5196_ (.Y(_1940_),
    .A(net823),
    .B(net1045));
 sg13g2_and4_1 _5197_ (.A(net826),
    .B(net823),
    .C(net870),
    .D(net1045),
    .X(_1941_));
 sg13g2_a22oi_1 _5198_ (.Y(_1942_),
    .B1(net1045),
    .B2(net826),
    .A2(net871),
    .A1(net822));
 sg13g2_nor2_1 _5199_ (.A(_1941_),
    .B(_1942_),
    .Y(_1943_));
 sg13g2_nand2_1 _5200_ (.Y(_1944_),
    .A(_1939_),
    .B(_1943_));
 sg13g2_xnor2_1 _5201_ (.Y(_1945_),
    .A(_1939_),
    .B(_1943_));
 sg13g2_xor2_1 _5202_ (.B(_1945_),
    .A(_1938_),
    .X(_1946_));
 sg13g2_nand2_1 _5203_ (.Y(_1947_),
    .A(_1932_),
    .B(_1946_));
 sg13g2_xnor2_1 _5204_ (.Y(_1948_),
    .A(_1932_),
    .B(_1946_));
 sg13g2_xor2_1 _5205_ (.B(_1948_),
    .A(_1931_),
    .X(_1949_));
 sg13g2_nand2_1 _5206_ (.Y(_1950_),
    .A(_1920_),
    .B(_1949_));
 sg13g2_xnor2_1 _5207_ (.Y(_1951_),
    .A(_1920_),
    .B(_1949_));
 sg13g2_nand2b_1 _5208_ (.Y(_1952_),
    .B(_1919_),
    .A_N(_1951_));
 sg13g2_xnor2_1 _5209_ (.Y(_1953_),
    .A(_1919_),
    .B(_1951_));
 sg13g2_nor2_1 _5210_ (.A(_1918_),
    .B(_1953_),
    .Y(_1954_));
 sg13g2_nand2_1 _5211_ (.Y(_1955_),
    .A(_1918_),
    .B(_1953_));
 sg13g2_nor2b_2 _5212_ (.A(_1954_),
    .B_N(_1955_),
    .Y(_1956_));
 sg13g2_xor2_1 _5213_ (.B(_1956_),
    .A(_1917_),
    .X(_0159_));
 sg13g2_a21oi_1 _5214_ (.A1(_1922_),
    .A2(_1928_),
    .Y(_1957_),
    .B1(_1930_));
 sg13g2_o21ai_1 _5215_ (.B1(_1947_),
    .Y(_1958_),
    .A1(_1931_),
    .A2(_1948_));
 sg13g2_o21ai_1 _5216_ (.B1(_1927_),
    .Y(_1959_),
    .A1(_1874_),
    .A2(_1925_));
 sg13g2_o21ai_1 _5217_ (.B1(_1935_),
    .Y(_1960_),
    .A1(_1933_),
    .A2(_1936_));
 sg13g2_nand2_1 _5218_ (.Y(_1961_),
    .A(net885),
    .B(net1042));
 sg13g2_nand2_1 _5219_ (.Y(_1962_),
    .A(net878),
    .B(net811));
 sg13g2_nand2_1 _5220_ (.Y(_1963_),
    .A(net878),
    .B(net814));
 sg13g2_or2_1 _5221_ (.X(_1964_),
    .B(_1962_),
    .A(_1925_));
 sg13g2_xnor2_1 _5222_ (.Y(_1965_),
    .A(_1924_),
    .B(_1963_));
 sg13g2_xor2_1 _5223_ (.B(_1965_),
    .A(_1961_),
    .X(_1966_));
 sg13g2_xnor2_1 _5224_ (.Y(_1967_),
    .A(_1960_),
    .B(_1966_));
 sg13g2_nor2b_1 _5225_ (.A(_1967_),
    .B_N(_1959_),
    .Y(_1968_));
 sg13g2_xor2_1 _5226_ (.B(_1967_),
    .A(_1959_),
    .X(_1969_));
 sg13g2_o21ai_1 _5227_ (.B1(_1944_),
    .Y(_1970_),
    .A1(_1938_),
    .A2(_1945_));
 sg13g2_a21oi_1 _5228_ (.A1(net827),
    .A2(net871),
    .Y(_1971_),
    .B1(_1940_));
 sg13g2_nand2_1 _5229_ (.Y(_1972_),
    .A(net876),
    .B(net816));
 sg13g2_nand2_1 _5230_ (.Y(_1973_),
    .A(net819),
    .B(net871));
 sg13g2_and4_1 _5231_ (.A(net821),
    .B(net818),
    .C(net874),
    .D(net871),
    .X(_1974_));
 sg13g2_a22oi_1 _5232_ (.Y(_1975_),
    .B1(net871),
    .B2(net821),
    .A2(net874),
    .A1(net819));
 sg13g2_nor3_1 _5233_ (.A(_1972_),
    .B(_1974_),
    .C(_1975_),
    .Y(_1976_));
 sg13g2_o21ai_1 _5234_ (.B1(_1972_),
    .Y(_1977_),
    .A1(_1974_),
    .A2(_1975_));
 sg13g2_nor2b_1 _5235_ (.A(_1976_),
    .B_N(_1977_),
    .Y(_1978_));
 sg13g2_xnor2_1 _5236_ (.Y(_1979_),
    .A(_1971_),
    .B(_1978_));
 sg13g2_nand2b_1 _5237_ (.Y(_1980_),
    .B(_1970_),
    .A_N(_1979_));
 sg13g2_xor2_1 _5238_ (.B(_1979_),
    .A(_1970_),
    .X(_1981_));
 sg13g2_xor2_1 _5239_ (.B(_1981_),
    .A(_1969_),
    .X(_1982_));
 sg13g2_nand2_1 _5240_ (.Y(_1983_),
    .A(_1958_),
    .B(_1982_));
 sg13g2_xor2_1 _5241_ (.B(_1982_),
    .A(_1958_),
    .X(_1984_));
 sg13g2_nand2b_1 _5242_ (.Y(_1985_),
    .B(_1984_),
    .A_N(_1957_));
 sg13g2_xor2_1 _5243_ (.B(_1984_),
    .A(_1957_),
    .X(_1986_));
 sg13g2_a21oi_1 _5244_ (.A1(_1950_),
    .A2(_1952_),
    .Y(_1987_),
    .B1(_1986_));
 sg13g2_nand3_1 _5245_ (.B(_1952_),
    .C(_1986_),
    .A(_1950_),
    .Y(_1988_));
 sg13g2_nand2b_1 _5246_ (.Y(_1989_),
    .B(_1988_),
    .A_N(_1987_));
 sg13g2_a21oi_1 _5247_ (.A1(_1913_),
    .A2(_1955_),
    .Y(_1990_),
    .B1(_1954_));
 sg13g2_a21oi_2 _5248_ (.B1(_1990_),
    .Y(_1991_),
    .A2(_1956_),
    .A1(_1916_));
 sg13g2_nor2_1 _5249_ (.A(_1989_),
    .B(_1991_),
    .Y(_1992_));
 sg13g2_xor2_1 _5250_ (.B(_1991_),
    .A(_1989_),
    .X(_0150_));
 sg13g2_a21o_1 _5251_ (.A2(_1966_),
    .A1(_1960_),
    .B1(_1968_),
    .X(_1993_));
 sg13g2_o21ai_1 _5252_ (.B1(_1980_),
    .Y(_1994_),
    .A1(_1969_),
    .A2(_1981_));
 sg13g2_a21o_1 _5253_ (.A2(_1978_),
    .A1(_1971_),
    .B1(_1941_),
    .X(_1995_));
 sg13g2_nand2_1 _5254_ (.Y(_1996_),
    .A(net816),
    .B(net874));
 sg13g2_nand2_1 _5255_ (.Y(_1997_),
    .A(net821),
    .B(net1046));
 sg13g2_or2_1 _5256_ (.X(_1998_),
    .B(_1997_),
    .A(_1973_));
 sg13g2_xnor2_1 _5257_ (.Y(_1999_),
    .A(_1973_),
    .B(_1997_));
 sg13g2_xor2_1 _5258_ (.B(_1999_),
    .A(_1996_),
    .X(_2000_));
 sg13g2_and2_1 _5259_ (.A(_1995_),
    .B(_2000_),
    .X(_2001_));
 sg13g2_or2_1 _5260_ (.X(_2002_),
    .B(_2000_),
    .A(_1995_));
 sg13g2_xnor2_1 _5261_ (.Y(_2003_),
    .A(_1995_),
    .B(_2000_));
 sg13g2_o21ai_1 _5262_ (.B1(_1964_),
    .Y(_2004_),
    .A1(_1961_),
    .A2(_1965_));
 sg13g2_or2_1 _5263_ (.X(_2005_),
    .B(_1976_),
    .A(_1974_));
 sg13g2_nand2_1 _5264_ (.Y(_2006_),
    .A(net882),
    .B(net1042));
 sg13g2_nand2_1 _5265_ (.Y(_2007_),
    .A(net876),
    .B(net815));
 sg13g2_or2_1 _5266_ (.X(_2008_),
    .B(_2007_),
    .A(_1962_));
 sg13g2_xnor2_1 _5267_ (.Y(_2009_),
    .A(_1962_),
    .B(_2007_));
 sg13g2_xor2_1 _5268_ (.B(_2009_),
    .A(_2006_),
    .X(_2010_));
 sg13g2_xnor2_1 _5269_ (.Y(_2011_),
    .A(_2005_),
    .B(_2010_));
 sg13g2_nor2b_1 _5270_ (.A(_2011_),
    .B_N(_2004_),
    .Y(_2012_));
 sg13g2_xnor2_1 _5271_ (.Y(_2013_),
    .A(_2004_),
    .B(_2011_));
 sg13g2_xnor2_1 _5272_ (.Y(_2014_),
    .A(_2003_),
    .B(_2013_));
 sg13g2_xnor2_1 _5273_ (.Y(_2015_),
    .A(_1994_),
    .B(_2014_));
 sg13g2_nor2b_1 _5274_ (.A(_2015_),
    .B_N(_1993_),
    .Y(_2016_));
 sg13g2_xor2_1 _5275_ (.B(_2015_),
    .A(_1993_),
    .X(_2017_));
 sg13g2_nand3_1 _5276_ (.B(_1985_),
    .C(_2017_),
    .A(_1983_),
    .Y(_2018_));
 sg13g2_inv_1 _5277_ (.Y(_2019_),
    .A(_2018_));
 sg13g2_a21oi_1 _5278_ (.A1(_1983_),
    .A2(_1985_),
    .Y(_2020_),
    .B1(_2017_));
 sg13g2_nor2_1 _5279_ (.A(_2019_),
    .B(_2020_),
    .Y(_2021_));
 sg13g2_nor2_1 _5280_ (.A(_1987_),
    .B(_1992_),
    .Y(_2022_));
 sg13g2_xnor2_1 _5281_ (.Y(_0151_),
    .A(_2021_),
    .B(_2022_));
 sg13g2_a21o_1 _5282_ (.A2(_2010_),
    .A1(_2005_),
    .B1(_2012_),
    .X(_2023_));
 sg13g2_a22oi_1 _5283_ (.Y(_2024_),
    .B1(net1045),
    .B2(net819),
    .A2(net870),
    .A1(net816));
 sg13g2_nand2_1 _5284_ (.Y(_2025_),
    .A(net817),
    .B(net1045));
 sg13g2_or2_1 _5285_ (.X(_2026_),
    .B(_2025_),
    .A(_1973_));
 sg13g2_nand2b_1 _5286_ (.Y(_2027_),
    .B(_2026_),
    .A_N(_2024_));
 sg13g2_o21ai_1 _5287_ (.B1(_2008_),
    .Y(_2028_),
    .A1(_2006_),
    .A2(_2009_));
 sg13g2_o21ai_1 _5288_ (.B1(_1998_),
    .Y(_2029_),
    .A1(_1996_),
    .A2(_1999_));
 sg13g2_nand2_1 _5289_ (.Y(_2030_),
    .A(net879),
    .B(net1042));
 sg13g2_nand2_1 _5290_ (.Y(_2031_),
    .A(net874),
    .B(net812));
 sg13g2_and4_1 _5291_ (.A(net876),
    .B(net874),
    .C(net815),
    .D(net812),
    .X(_2032_));
 sg13g2_or2_1 _5292_ (.X(_2033_),
    .B(_2031_),
    .A(_2007_));
 sg13g2_a22oi_1 _5293_ (.Y(_2034_),
    .B1(net812),
    .B2(net876),
    .A2(net814),
    .A1(net874));
 sg13g2_nor2_1 _5294_ (.A(_2032_),
    .B(_2034_),
    .Y(_2035_));
 sg13g2_xnor2_1 _5295_ (.Y(_2036_),
    .A(_2030_),
    .B(_2035_));
 sg13g2_xnor2_1 _5296_ (.Y(_2037_),
    .A(_2029_),
    .B(_2036_));
 sg13g2_nor2b_1 _5297_ (.A(_2037_),
    .B_N(_2028_),
    .Y(_2038_));
 sg13g2_xor2_1 _5298_ (.B(_2037_),
    .A(_2028_),
    .X(_2039_));
 sg13g2_or2_1 _5299_ (.X(_2040_),
    .B(_2039_),
    .A(_2027_));
 sg13g2_xor2_1 _5300_ (.B(_2039_),
    .A(_2027_),
    .X(_2041_));
 sg13g2_a21oi_1 _5301_ (.A1(_2002_),
    .A2(_2013_),
    .Y(_2042_),
    .B1(_2001_));
 sg13g2_nor2b_1 _5302_ (.A(_2042_),
    .B_N(_2041_),
    .Y(_2043_));
 sg13g2_xor2_1 _5303_ (.B(_2042_),
    .A(_2041_),
    .X(_2044_));
 sg13g2_nor2b_1 _5304_ (.A(_2044_),
    .B_N(_2023_),
    .Y(_2045_));
 sg13g2_xor2_1 _5305_ (.B(_2044_),
    .A(_2023_),
    .X(_2046_));
 sg13g2_a21oi_1 _5306_ (.A1(_1994_),
    .A2(_2014_),
    .Y(_2047_),
    .B1(_2016_));
 sg13g2_nor2_1 _5307_ (.A(_2046_),
    .B(_2047_),
    .Y(_2048_));
 sg13g2_xor2_1 _5308_ (.B(_2047_),
    .A(_2046_),
    .X(_2049_));
 sg13g2_a21oi_1 _5309_ (.A1(_1987_),
    .A2(_2018_),
    .Y(_2050_),
    .B1(_2020_));
 sg13g2_a21oi_1 _5310_ (.A1(_1988_),
    .A2(_2018_),
    .Y(_2051_),
    .B1(_2020_));
 sg13g2_a21oi_2 _5311_ (.B1(_2051_),
    .Y(_2052_),
    .A2(_2050_),
    .A1(_1991_));
 sg13g2_xor2_1 _5312_ (.B(_2052_),
    .A(_2049_),
    .X(_0152_));
 sg13g2_a21o_1 _5313_ (.A2(_2036_),
    .A1(_2029_),
    .B1(_2038_),
    .X(_2053_));
 sg13g2_o21ai_1 _5314_ (.B1(_2033_),
    .Y(_2054_),
    .A1(_2030_),
    .A2(_2034_));
 sg13g2_nand2_1 _5315_ (.Y(_2055_),
    .A(net876),
    .B(net1042));
 sg13g2_nand2_1 _5316_ (.Y(_2056_),
    .A(net872),
    .B(net811));
 sg13g2_nand2_1 _5317_ (.Y(_2057_),
    .A(net815),
    .B(net872));
 sg13g2_xor2_1 _5318_ (.B(_2057_),
    .A(_2031_),
    .X(_2058_));
 sg13g2_nand2b_1 _5319_ (.Y(_2059_),
    .B(_2058_),
    .A_N(_2055_));
 sg13g2_xnor2_1 _5320_ (.Y(_2060_),
    .A(_2055_),
    .B(_2058_));
 sg13g2_nor2b_1 _5321_ (.A(_2026_),
    .B_N(_2060_),
    .Y(_2061_));
 sg13g2_xnor2_1 _5322_ (.Y(_2062_),
    .A(_2026_),
    .B(_2060_));
 sg13g2_xnor2_1 _5323_ (.Y(_2063_),
    .A(_2054_),
    .B(_2062_));
 sg13g2_nor2_1 _5324_ (.A(_2025_),
    .B(_2063_),
    .Y(_2064_));
 sg13g2_xnor2_1 _5325_ (.Y(_2065_),
    .A(_2025_),
    .B(_2063_));
 sg13g2_nor2_1 _5326_ (.A(_2040_),
    .B(_2065_),
    .Y(_2066_));
 sg13g2_xor2_1 _5327_ (.B(_2065_),
    .A(_2040_),
    .X(_2067_));
 sg13g2_xor2_1 _5328_ (.B(_2067_),
    .A(_2053_),
    .X(_2068_));
 sg13g2_o21ai_1 _5329_ (.B1(_2068_),
    .Y(_2069_),
    .A1(_2043_),
    .A2(_2045_));
 sg13g2_or3_1 _5330_ (.A(_2043_),
    .B(_2045_),
    .C(_2068_),
    .X(_2070_));
 sg13g2_and2_1 _5331_ (.A(_2069_),
    .B(_2070_),
    .X(_2071_));
 sg13g2_a21oi_1 _5332_ (.A1(_2049_),
    .A2(_2052_),
    .Y(_2072_),
    .B1(_2048_));
 sg13g2_xnor2_1 _5333_ (.Y(_0153_),
    .A(_2071_),
    .B(_2072_));
 sg13g2_nand2_1 _5334_ (.Y(_2073_),
    .A(_2049_),
    .B(_2071_));
 sg13g2_inv_1 _5335_ (.Y(_2074_),
    .A(_2073_));
 sg13g2_o21ai_1 _5336_ (.B1(_2069_),
    .Y(_2075_),
    .A1(_2046_),
    .A2(_2047_));
 sg13g2_a22oi_1 _5337_ (.Y(_2076_),
    .B1(_2075_),
    .B2(_2070_),
    .A2(_2074_),
    .A1(_2052_));
 sg13g2_a21oi_1 _5338_ (.A1(_2053_),
    .A2(_2067_),
    .Y(_2077_),
    .B1(_2066_));
 sg13g2_a21o_1 _5339_ (.A2(_2062_),
    .A1(_2054_),
    .B1(_2061_),
    .X(_2078_));
 sg13g2_o21ai_1 _5340_ (.B1(_2059_),
    .Y(_2079_),
    .A1(_2031_),
    .A2(_2057_));
 sg13g2_nand2_1 _5341_ (.Y(_2080_),
    .A(net874),
    .B(net1042));
 sg13g2_nand2_1 _5342_ (.Y(_2081_),
    .A(net812),
    .B(net1046));
 sg13g2_nand2_1 _5343_ (.Y(_2082_),
    .A(net815),
    .B(net1046));
 sg13g2_xor2_1 _5344_ (.B(_2082_),
    .A(_2056_),
    .X(_2083_));
 sg13g2_nand2b_1 _5345_ (.Y(_2084_),
    .B(_2083_),
    .A_N(_2080_));
 sg13g2_xnor2_1 _5346_ (.Y(_2085_),
    .A(_2080_),
    .B(_2083_));
 sg13g2_nand2_1 _5347_ (.Y(_2086_),
    .A(_2079_),
    .B(_2085_));
 sg13g2_xor2_1 _5348_ (.B(_2085_),
    .A(_2079_),
    .X(_2087_));
 sg13g2_xnor2_1 _5349_ (.Y(_2088_),
    .A(_2064_),
    .B(_2087_));
 sg13g2_nor2b_1 _5350_ (.A(_2088_),
    .B_N(_2078_),
    .Y(_2089_));
 sg13g2_xor2_1 _5351_ (.B(_2088_),
    .A(_2078_),
    .X(_2090_));
 sg13g2_or2_1 _5352_ (.X(_2091_),
    .B(_2090_),
    .A(_2077_));
 sg13g2_xor2_1 _5353_ (.B(_2090_),
    .A(_2077_),
    .X(_2092_));
 sg13g2_inv_1 _5354_ (.Y(_2093_),
    .A(_2092_));
 sg13g2_xnor2_1 _5355_ (.Y(_0154_),
    .A(_2076_),
    .B(_2092_));
 sg13g2_o21ai_1 _5356_ (.B1(_2091_),
    .Y(_2094_),
    .A1(_2076_),
    .A2(_2093_));
 sg13g2_a21oi_1 _5357_ (.A1(_2064_),
    .A2(_2087_),
    .Y(_2095_),
    .B1(_2089_));
 sg13g2_o21ai_1 _5358_ (.B1(_2084_),
    .Y(_2096_),
    .A1(_2056_),
    .A2(_2082_));
 sg13g2_nand2_1 _5359_ (.Y(_2097_),
    .A(net872),
    .B(net1042));
 sg13g2_xor2_1 _5360_ (.B(_2097_),
    .A(_2081_),
    .X(_2098_));
 sg13g2_xnor2_1 _5361_ (.Y(_2099_),
    .A(_2096_),
    .B(_2098_));
 sg13g2_xnor2_1 _5362_ (.Y(_2100_),
    .A(_2086_),
    .B(_2099_));
 sg13g2_xnor2_1 _5363_ (.Y(_2101_),
    .A(_2095_),
    .B(_2100_));
 sg13g2_xnor2_1 _5364_ (.Y(_0155_),
    .A(_2094_),
    .B(_2101_));
 sg13g2_nand2_1 _5365_ (.Y(_2102_),
    .A(net287),
    .B(net267));
 sg13g2_nand2_1 _5366_ (.Y(_2103_),
    .A(\mac1.sum_lvl2_ff[20] ),
    .B(\mac1.sum_lvl2_ff[1] ));
 sg13g2_nor2_1 _5367_ (.A(\mac1.sum_lvl2_ff[20] ),
    .B(\mac1.sum_lvl2_ff[1] ),
    .Y(_2104_));
 sg13g2_xor2_1 _5368_ (.B(\mac1.sum_lvl2_ff[1] ),
    .A(\mac1.sum_lvl2_ff[20] ),
    .X(_2105_));
 sg13g2_xnor2_1 _5369_ (.Y(_0007_),
    .A(_2102_),
    .B(_2105_));
 sg13g2_o21ai_1 _5370_ (.B1(_2103_),
    .Y(_2106_),
    .A1(_2102_),
    .A2(_2104_));
 sg13g2_and2_1 _5371_ (.A(\mac1.sum_lvl2_ff[21] ),
    .B(net389),
    .X(_2107_));
 sg13g2_xor2_1 _5372_ (.B(net389),
    .A(\mac1.sum_lvl2_ff[21] ),
    .X(_2108_));
 sg13g2_xor2_1 _5373_ (.B(net390),
    .A(_2106_),
    .X(_0008_));
 sg13g2_a21oi_2 _5374_ (.B1(_2107_),
    .Y(_2109_),
    .A2(net390),
    .A1(_2106_));
 sg13g2_nand2_1 _5375_ (.Y(_2110_),
    .A(\mac1.sum_lvl2_ff[22] ),
    .B(\mac1.sum_lvl2_ff[3] ));
 sg13g2_xnor2_1 _5376_ (.Y(_2111_),
    .A(\mac1.sum_lvl2_ff[22] ),
    .B(net475));
 sg13g2_xor2_1 _5377_ (.B(net476),
    .A(_2109_),
    .X(_0009_));
 sg13g2_o21ai_1 _5378_ (.B1(_2110_),
    .Y(_2112_),
    .A1(_2109_),
    .A2(_2111_));
 sg13g2_and2_1 _5379_ (.A(\mac1.sum_lvl2_ff[23] ),
    .B(net340),
    .X(_2113_));
 sg13g2_xor2_1 _5380_ (.B(net340),
    .A(\mac1.sum_lvl2_ff[23] ),
    .X(_2114_));
 sg13g2_xor2_1 _5381_ (.B(net341),
    .A(_2112_),
    .X(_0010_));
 sg13g2_a21oi_1 _5382_ (.A1(_2112_),
    .A2(_2114_),
    .Y(_2115_),
    .B1(_2113_));
 sg13g2_nor2_1 _5383_ (.A(\mac1.sum_lvl2_ff[24] ),
    .B(net294),
    .Y(_2116_));
 sg13g2_xor2_1 _5384_ (.B(net294),
    .A(\mac1.sum_lvl2_ff[24] ),
    .X(_2117_));
 sg13g2_xnor2_1 _5385_ (.Y(_0011_),
    .A(_2115_),
    .B(net295));
 sg13g2_and2_1 _5386_ (.A(\mac1.sum_lvl2_ff[25] ),
    .B(net461),
    .X(_2118_));
 sg13g2_xnor2_1 _5387_ (.Y(_2119_),
    .A(\mac1.sum_lvl2_ff[25] ),
    .B(net461));
 sg13g2_a221oi_1 _5388_ (.B2(_2114_),
    .C1(_2113_),
    .B1(_2112_),
    .A1(\mac1.sum_lvl2_ff[24] ),
    .Y(_2120_),
    .A2(net294));
 sg13g2_nor3_1 _5389_ (.A(_2116_),
    .B(net462),
    .C(_2120_),
    .Y(_2121_));
 sg13g2_o21ai_1 _5390_ (.B1(net462),
    .Y(_2122_),
    .A1(_2116_),
    .A2(_2120_));
 sg13g2_nor2b_1 _5391_ (.A(_2121_),
    .B_N(net463),
    .Y(_0012_));
 sg13g2_nand2_1 _5392_ (.Y(_2123_),
    .A(\mac1.sum_lvl2_ff[26] ),
    .B(\mac1.sum_lvl2_ff[7] ));
 sg13g2_xor2_1 _5393_ (.B(net535),
    .A(\mac1.sum_lvl2_ff[26] ),
    .X(_2124_));
 sg13g2_o21ai_1 _5394_ (.B1(net536),
    .Y(_2125_),
    .A1(_2118_),
    .A2(_2121_));
 sg13g2_or3_1 _5395_ (.A(_2118_),
    .B(_2121_),
    .C(net536),
    .X(_2126_));
 sg13g2_and2_1 _5396_ (.A(net537),
    .B(_2126_),
    .X(_0013_));
 sg13g2_xnor2_1 _5397_ (.Y(_2127_),
    .A(\mac1.sum_lvl2_ff[27] ),
    .B(net392));
 sg13g2_a21oi_1 _5398_ (.A1(_2123_),
    .A2(_2125_),
    .Y(_2128_),
    .B1(net393));
 sg13g2_nand3_1 _5399_ (.B(_2125_),
    .C(net393),
    .A(_2123_),
    .Y(_2129_));
 sg13g2_nor2b_1 _5400_ (.A(net394),
    .B_N(_2129_),
    .Y(_0014_));
 sg13g2_a21o_1 _5401_ (.A2(net392),
    .A1(net458),
    .B1(net394),
    .X(_2130_));
 sg13g2_and2_1 _5402_ (.A(\mac1.sum_lvl2_ff[28] ),
    .B(\mac1.sum_lvl2_ff[9] ),
    .X(_2131_));
 sg13g2_or2_1 _5403_ (.X(_2132_),
    .B(\mac1.sum_lvl2_ff[9] ),
    .A(\mac1.sum_lvl2_ff[28] ));
 sg13g2_nand2b_1 _5404_ (.Y(_2133_),
    .B(_2132_),
    .A_N(_2131_));
 sg13g2_xnor2_1 _5405_ (.Y(_0015_),
    .A(_2130_),
    .B(_2133_));
 sg13g2_nand2_1 _5406_ (.Y(_2134_),
    .A(net365),
    .B(\mac1.sum_lvl2_ff[10] ));
 sg13g2_xor2_1 _5407_ (.B(net478),
    .A(net365),
    .X(_2135_));
 sg13g2_inv_1 _5408_ (.Y(_2136_),
    .A(_2135_));
 sg13g2_a21o_2 _5409_ (.A2(_2132_),
    .A1(_2130_),
    .B1(_2131_),
    .X(_2137_));
 sg13g2_nand2_1 _5410_ (.Y(_2138_),
    .A(_2135_),
    .B(_2137_));
 sg13g2_xnor2_1 _5411_ (.Y(_0001_),
    .A(_2136_),
    .B(_2137_));
 sg13g2_nor2_1 _5412_ (.A(\mac1.sum_lvl2_ff[30] ),
    .B(\mac1.sum_lvl2_ff[11] ),
    .Y(_2139_));
 sg13g2_xnor2_1 _5413_ (.Y(_2140_),
    .A(\mac1.sum_lvl2_ff[30] ),
    .B(\mac1.sum_lvl2_ff[11] ));
 sg13g2_nand2_1 _5414_ (.Y(_2141_),
    .A(net366),
    .B(_2138_));
 sg13g2_xnor2_1 _5415_ (.Y(_0002_),
    .A(_2140_),
    .B(net367));
 sg13g2_nand2_1 _5416_ (.Y(_2142_),
    .A(\mac1.sum_lvl2_ff[31] ),
    .B(net319));
 sg13g2_nor2_1 _5417_ (.A(\mac1.sum_lvl2_ff[31] ),
    .B(net319),
    .Y(_2143_));
 sg13g2_xor2_1 _5418_ (.B(net319),
    .A(\mac1.sum_lvl2_ff[31] ),
    .X(_2144_));
 sg13g2_nor2_1 _5419_ (.A(_2134_),
    .B(_2139_),
    .Y(_2145_));
 sg13g2_nor2_1 _5420_ (.A(_2136_),
    .B(_2140_),
    .Y(_2146_));
 sg13g2_a221oi_1 _5421_ (.B2(_2146_),
    .C1(_2145_),
    .B1(_2137_),
    .A1(\mac1.sum_lvl2_ff[30] ),
    .Y(_2147_),
    .A2(\mac1.sum_lvl2_ff[11] ));
 sg13g2_xnor2_1 _5422_ (.Y(_0003_),
    .A(net320),
    .B(_2147_));
 sg13g2_o21ai_1 _5423_ (.B1(_2142_),
    .Y(_2148_),
    .A1(_2143_),
    .A2(_2147_));
 sg13g2_and2_1 _5424_ (.A(\mac1.sum_lvl2_ff[32] ),
    .B(net465),
    .X(_2149_));
 sg13g2_or2_1 _5425_ (.X(_2150_),
    .B(net465),
    .A(\mac1.sum_lvl2_ff[32] ));
 sg13g2_nand2b_1 _5426_ (.Y(_2151_),
    .B(net466),
    .A_N(_2149_));
 sg13g2_xnor2_1 _5427_ (.Y(_0004_),
    .A(_2148_),
    .B(net467));
 sg13g2_a21oi_1 _5428_ (.A1(_2148_),
    .A2(_2150_),
    .Y(_2152_),
    .B1(_2149_));
 sg13g2_nand2_1 _5429_ (.Y(_2153_),
    .A(\mac1.sum_lvl2_ff[33] ),
    .B(\mac1.sum_lvl2_ff[14] ));
 sg13g2_nor2_1 _5430_ (.A(\mac1.sum_lvl2_ff[33] ),
    .B(\mac1.sum_lvl2_ff[14] ),
    .Y(_2154_));
 sg13g2_xor2_1 _5431_ (.B(net303),
    .A(\mac1.sum_lvl2_ff[33] ),
    .X(_2155_));
 sg13g2_xnor2_1 _5432_ (.Y(_0005_),
    .A(_2152_),
    .B(net304));
 sg13g2_o21ai_1 _5433_ (.B1(_2153_),
    .Y(_2156_),
    .A1(_2152_),
    .A2(_2154_));
 sg13g2_xnor2_1 _5434_ (.Y(_2157_),
    .A(\mac1.sum_lvl2_ff[34] ),
    .B(net284));
 sg13g2_xnor2_1 _5435_ (.Y(_0006_),
    .A(_2156_),
    .B(net285));
 sg13g2_xor2_1 _5436_ (.B(net267),
    .A(\mac1.sum_lvl2_ff[19] ),
    .X(_0000_));
 sg13g2_nand2_1 _5437_ (.Y(_2158_),
    .A(net292),
    .B(net265));
 sg13g2_nand2_1 _5438_ (.Y(_2159_),
    .A(\mac1.sum_lvl3_ff[21] ),
    .B(\mac1.sum_lvl3_ff[1] ));
 sg13g2_nor2_1 _5439_ (.A(\mac1.sum_lvl3_ff[21] ),
    .B(\mac1.sum_lvl3_ff[1] ),
    .Y(_2160_));
 sg13g2_xor2_1 _5440_ (.B(\mac1.sum_lvl3_ff[1] ),
    .A(\mac1.sum_lvl3_ff[21] ),
    .X(_2161_));
 sg13g2_xnor2_1 _5441_ (.Y(_0023_),
    .A(_2158_),
    .B(_2161_));
 sg13g2_o21ai_1 _5442_ (.B1(_2159_),
    .Y(_2162_),
    .A1(_2158_),
    .A2(_2160_));
 sg13g2_and2_1 _5443_ (.A(\mac1.sum_lvl3_ff[22] ),
    .B(net381),
    .X(_2163_));
 sg13g2_xor2_1 _5444_ (.B(net381),
    .A(\mac1.sum_lvl3_ff[22] ),
    .X(_2164_));
 sg13g2_xor2_1 _5445_ (.B(net382),
    .A(_2162_),
    .X(_0024_));
 sg13g2_a21oi_1 _5446_ (.A1(_2162_),
    .A2(_2164_),
    .Y(_2165_),
    .B1(_2163_));
 sg13g2_nand2_1 _5447_ (.Y(_2166_),
    .A(\mac1.sum_lvl3_ff[23] ),
    .B(\mac1.sum_lvl3_ff[3] ));
 sg13g2_xnor2_1 _5448_ (.Y(_2167_),
    .A(\mac1.sum_lvl3_ff[23] ),
    .B(net441));
 sg13g2_xor2_1 _5449_ (.B(net442),
    .A(_2165_),
    .X(_0025_));
 sg13g2_o21ai_1 _5450_ (.B1(_2166_),
    .Y(_2168_),
    .A1(_2165_),
    .A2(_2167_));
 sg13g2_and2_1 _5451_ (.A(\mac1.sum_lvl3_ff[24] ),
    .B(\mac1.sum_lvl3_ff[4] ),
    .X(_2169_));
 sg13g2_xor2_1 _5452_ (.B(net551),
    .A(\mac1.sum_lvl3_ff[24] ),
    .X(_2170_));
 sg13g2_xor2_1 _5453_ (.B(_2170_),
    .A(_2168_),
    .X(_0026_));
 sg13g2_a21oi_1 _5454_ (.A1(_2168_),
    .A2(_2170_),
    .Y(_2171_),
    .B1(_2169_));
 sg13g2_nor2_1 _5455_ (.A(\mac1.sum_lvl3_ff[25] ),
    .B(\mac1.sum_lvl3_ff[5] ),
    .Y(_2172_));
 sg13g2_xor2_1 _5456_ (.B(net546),
    .A(\mac1.sum_lvl3_ff[25] ),
    .X(_2173_));
 sg13g2_xnor2_1 _5457_ (.Y(_0027_),
    .A(_2171_),
    .B(net547));
 sg13g2_and2_1 _5458_ (.A(\mac1.sum_lvl3_ff[26] ),
    .B(\mac1.sum_lvl3_ff[6] ),
    .X(_2174_));
 sg13g2_xnor2_1 _5459_ (.Y(_2175_),
    .A(\mac1.sum_lvl3_ff[26] ),
    .B(net532));
 sg13g2_a221oi_1 _5460_ (.B2(_2170_),
    .C1(_2169_),
    .B1(_2168_),
    .A1(\mac1.sum_lvl3_ff[25] ),
    .Y(_2176_),
    .A2(\mac1.sum_lvl3_ff[5] ));
 sg13g2_nor3_1 _5461_ (.A(_2172_),
    .B(_2175_),
    .C(_2176_),
    .Y(_2177_));
 sg13g2_o21ai_1 _5462_ (.B1(net533),
    .Y(_2178_),
    .A1(_2172_),
    .A2(_2176_));
 sg13g2_nor2b_2 _5463_ (.A(_2177_),
    .B_N(net534),
    .Y(_0028_));
 sg13g2_nand2_1 _5464_ (.Y(_2179_),
    .A(\mac1.sum_lvl3_ff[27] ),
    .B(\mac1.sum_lvl3_ff[7] ));
 sg13g2_xor2_1 _5465_ (.B(\mac1.sum_lvl3_ff[7] ),
    .A(\mac1.sum_lvl3_ff[27] ),
    .X(_2180_));
 sg13g2_o21ai_1 _5466_ (.B1(_2180_),
    .Y(_2181_),
    .A1(_2174_),
    .A2(_2177_));
 sg13g2_or3_1 _5467_ (.A(_2174_),
    .B(_2177_),
    .C(_2180_),
    .X(_2182_));
 sg13g2_and2_1 _5468_ (.A(_2181_),
    .B(_2182_),
    .X(_0029_));
 sg13g2_and2_1 _5469_ (.A(\mac1.sum_lvl3_ff[28] ),
    .B(\mac1.sum_lvl3_ff[8] ),
    .X(_2183_));
 sg13g2_xnor2_1 _5470_ (.Y(_2184_),
    .A(\mac1.sum_lvl3_ff[28] ),
    .B(net494));
 sg13g2_a21oi_2 _5471_ (.B1(net495),
    .Y(_2185_),
    .A2(_2181_),
    .A1(_2179_));
 sg13g2_nand3_1 _5472_ (.B(_2181_),
    .C(_2184_),
    .A(_2179_),
    .Y(_2186_));
 sg13g2_nor2b_2 _5473_ (.A(net496),
    .B_N(_2186_),
    .Y(_0030_));
 sg13g2_nor2_1 _5474_ (.A(_2183_),
    .B(_2185_),
    .Y(_2187_));
 sg13g2_nand2_1 _5475_ (.Y(_2188_),
    .A(\mac1.sum_lvl3_ff[29] ),
    .B(net509));
 sg13g2_xor2_1 _5476_ (.B(net509),
    .A(\mac1.sum_lvl3_ff[29] ),
    .X(_2189_));
 sg13g2_o21ai_1 _5477_ (.B1(_2189_),
    .Y(_2190_),
    .A1(_2183_),
    .A2(_2185_));
 sg13g2_xnor2_1 _5478_ (.Y(_0031_),
    .A(_2187_),
    .B(net510));
 sg13g2_nand2_1 _5479_ (.Y(_2191_),
    .A(_2188_),
    .B(_2190_));
 sg13g2_nand2_1 _5480_ (.Y(_2192_),
    .A(net525),
    .B(net521));
 sg13g2_xor2_1 _5481_ (.B(net521),
    .A(\mac1.sum_lvl3_ff[30] ),
    .X(_2193_));
 sg13g2_nand2_1 _5482_ (.Y(_2194_),
    .A(_2191_),
    .B(_2193_));
 sg13g2_xor2_1 _5483_ (.B(net522),
    .A(_2191_),
    .X(_0017_));
 sg13g2_nor2_1 _5484_ (.A(\mac1.sum_lvl3_ff[31] ),
    .B(\mac1.sum_lvl3_ff[11] ),
    .Y(_2195_));
 sg13g2_nand2_1 _5485_ (.Y(_2196_),
    .A(\mac1.sum_lvl3_ff[31] ),
    .B(\mac1.sum_lvl3_ff[11] ));
 sg13g2_nand2b_1 _5486_ (.Y(_2197_),
    .B(_2196_),
    .A_N(_2195_));
 sg13g2_nand2_1 _5487_ (.Y(_2198_),
    .A(_2192_),
    .B(_2194_));
 sg13g2_xnor2_1 _5488_ (.Y(_0018_),
    .A(_2197_),
    .B(_2198_));
 sg13g2_nand2_1 _5489_ (.Y(_2199_),
    .A(\mac1.sum_lvl3_ff[32] ),
    .B(\mac1.sum_lvl3_ff[12] ));
 sg13g2_xor2_1 _5490_ (.B(net540),
    .A(\mac1.sum_lvl3_ff[32] ),
    .X(_2200_));
 sg13g2_o21ai_1 _5491_ (.B1(_2196_),
    .Y(_2201_),
    .A1(_2192_),
    .A2(_2195_));
 sg13g2_nand3b_1 _5492_ (.B(_2196_),
    .C(_2193_),
    .Y(_2202_),
    .A_N(_2195_));
 sg13g2_a21oi_2 _5493_ (.B1(_2202_),
    .Y(_2203_),
    .A2(_2190_),
    .A1(_2188_));
 sg13g2_o21ai_1 _5494_ (.B1(net541),
    .Y(_2204_),
    .A1(_2201_),
    .A2(_2203_));
 sg13g2_or3_1 _5495_ (.A(net541),
    .B(_2201_),
    .C(_2203_),
    .X(_2205_));
 sg13g2_and2_1 _5496_ (.A(_2204_),
    .B(_2205_),
    .X(_0019_));
 sg13g2_xnor2_1 _5497_ (.Y(_2206_),
    .A(\mac1.sum_lvl3_ff[33] ),
    .B(net427));
 sg13g2_a21oi_1 _5498_ (.A1(_2199_),
    .A2(_2204_),
    .Y(_2207_),
    .B1(net428));
 sg13g2_nand3_1 _5499_ (.B(_2204_),
    .C(net428),
    .A(_2199_),
    .Y(_2208_));
 sg13g2_nor2b_1 _5500_ (.A(net429),
    .B_N(_2208_),
    .Y(_0020_));
 sg13g2_a21oi_1 _5501_ (.A1(\mac1.sum_lvl3_ff[33] ),
    .A2(\mac1.sum_lvl3_ff[13] ),
    .Y(_2209_),
    .B1(_2207_));
 sg13g2_nand2_1 _5502_ (.Y(_2210_),
    .A(\mac1.sum_lvl3_ff[34] ),
    .B(\mac1.sum_lvl3_ff[14] ));
 sg13g2_nor2_1 _5503_ (.A(\mac1.sum_lvl3_ff[34] ),
    .B(\mac1.sum_lvl3_ff[14] ),
    .Y(_2211_));
 sg13g2_xor2_1 _5504_ (.B(net331),
    .A(\mac1.sum_lvl3_ff[34] ),
    .X(_2212_));
 sg13g2_xnor2_1 _5505_ (.Y(_0021_),
    .A(_2209_),
    .B(net332));
 sg13g2_o21ai_1 _5506_ (.B1(_2210_),
    .Y(_2213_),
    .A1(_2209_),
    .A2(_2211_));
 sg13g2_xnor2_1 _5507_ (.Y(_2214_),
    .A(\mac1.sum_lvl3_ff[35] ),
    .B(net289));
 sg13g2_xnor2_1 _5508_ (.Y(_0022_),
    .A(_2213_),
    .B(net290));
 sg13g2_xor2_1 _5509_ (.B(net265),
    .A(\mac1.sum_lvl3_ff[20] ),
    .X(_0016_));
 sg13g2_nand2_1 _5510_ (.Y(_2215_),
    .A(net308),
    .B(net271));
 sg13g2_nand2_1 _5511_ (.Y(_2216_),
    .A(\mac2.sum_lvl2_ff[20] ),
    .B(\mac2.sum_lvl2_ff[1] ));
 sg13g2_nor2_1 _5512_ (.A(\mac2.sum_lvl2_ff[20] ),
    .B(\mac2.sum_lvl2_ff[1] ),
    .Y(_2217_));
 sg13g2_xor2_1 _5513_ (.B(\mac2.sum_lvl2_ff[1] ),
    .A(\mac2.sum_lvl2_ff[20] ),
    .X(_2218_));
 sg13g2_xnor2_1 _5514_ (.Y(_0039_),
    .A(_2215_),
    .B(_2218_));
 sg13g2_o21ai_1 _5515_ (.B1(_2216_),
    .Y(_2219_),
    .A1(_2215_),
    .A2(_2217_));
 sg13g2_and2_1 _5516_ (.A(\mac2.sum_lvl2_ff[21] ),
    .B(net350),
    .X(_2220_));
 sg13g2_xor2_1 _5517_ (.B(net350),
    .A(\mac2.sum_lvl2_ff[21] ),
    .X(_2221_));
 sg13g2_xor2_1 _5518_ (.B(net351),
    .A(_2219_),
    .X(_0040_));
 sg13g2_a21oi_1 _5519_ (.A1(_2219_),
    .A2(_2221_),
    .Y(_2222_),
    .B1(_2220_));
 sg13g2_nand2_1 _5520_ (.Y(_2223_),
    .A(\mac2.sum_lvl2_ff[22] ),
    .B(net432));
 sg13g2_xnor2_1 _5521_ (.Y(_2224_),
    .A(\mac2.sum_lvl2_ff[22] ),
    .B(net432));
 sg13g2_xor2_1 _5522_ (.B(net433),
    .A(_2222_),
    .X(_0041_));
 sg13g2_o21ai_1 _5523_ (.B1(_2223_),
    .Y(_2225_),
    .A1(_2222_),
    .A2(_2224_));
 sg13g2_and2_1 _5524_ (.A(\mac2.sum_lvl2_ff[23] ),
    .B(\mac2.sum_lvl2_ff[4] ),
    .X(_2226_));
 sg13g2_xor2_1 _5525_ (.B(net512),
    .A(\mac2.sum_lvl2_ff[23] ),
    .X(_2227_));
 sg13g2_xor2_1 _5526_ (.B(net513),
    .A(_2225_),
    .X(_0042_));
 sg13g2_a21oi_1 _5527_ (.A1(_2225_),
    .A2(_2227_),
    .Y(_2228_),
    .B1(_2226_));
 sg13g2_nor2_1 _5528_ (.A(net548),
    .B(net469),
    .Y(_2229_));
 sg13g2_xor2_1 _5529_ (.B(net469),
    .A(\mac2.sum_lvl2_ff[24] ),
    .X(_2230_));
 sg13g2_xnor2_1 _5530_ (.Y(_0043_),
    .A(_2228_),
    .B(net470));
 sg13g2_and2_1 _5531_ (.A(\mac2.sum_lvl2_ff[25] ),
    .B(\mac2.sum_lvl2_ff[6] ),
    .X(_2231_));
 sg13g2_xnor2_1 _5532_ (.Y(_2232_),
    .A(\mac2.sum_lvl2_ff[25] ),
    .B(\mac2.sum_lvl2_ff[6] ));
 sg13g2_a221oi_1 _5533_ (.B2(_2227_),
    .C1(_2226_),
    .B1(_2225_),
    .A1(\mac2.sum_lvl2_ff[24] ),
    .Y(_2233_),
    .A2(\mac2.sum_lvl2_ff[5] ));
 sg13g2_nor3_2 _5534_ (.A(_2229_),
    .B(_2232_),
    .C(_2233_),
    .Y(_2234_));
 sg13g2_o21ai_1 _5535_ (.B1(_2232_),
    .Y(_2235_),
    .A1(_2229_),
    .A2(_2233_));
 sg13g2_nor2b_2 _5536_ (.A(_2234_),
    .B_N(net549),
    .Y(_0044_));
 sg13g2_nand2_1 _5537_ (.Y(_2236_),
    .A(\mac2.sum_lvl2_ff[26] ),
    .B(\mac2.sum_lvl2_ff[7] ));
 sg13g2_xor2_1 _5538_ (.B(\mac2.sum_lvl2_ff[7] ),
    .A(\mac2.sum_lvl2_ff[26] ),
    .X(_2237_));
 sg13g2_o21ai_1 _5539_ (.B1(_2237_),
    .Y(_2238_),
    .A1(_2231_),
    .A2(_2234_));
 sg13g2_or3_1 _5540_ (.A(_2231_),
    .B(_2234_),
    .C(_2237_),
    .X(_2239_));
 sg13g2_and2_1 _5541_ (.A(_2238_),
    .B(_2239_),
    .X(_0045_));
 sg13g2_xnor2_1 _5542_ (.Y(_2240_),
    .A(\mac2.sum_lvl2_ff[27] ),
    .B(net517));
 sg13g2_a21oi_1 _5543_ (.A1(_2236_),
    .A2(_2238_),
    .Y(_2241_),
    .B1(net518));
 sg13g2_nand3_1 _5544_ (.B(_2238_),
    .C(_2240_),
    .A(_2236_),
    .Y(_2242_));
 sg13g2_nor2b_2 _5545_ (.A(net519),
    .B_N(_2242_),
    .Y(_0046_));
 sg13g2_a21o_1 _5546_ (.A2(\mac2.sum_lvl2_ff[8] ),
    .A1(\mac2.sum_lvl2_ff[27] ),
    .B1(_2241_),
    .X(_2243_));
 sg13g2_and2_1 _5547_ (.A(\mac2.sum_lvl2_ff[28] ),
    .B(\mac2.sum_lvl2_ff[9] ),
    .X(_2244_));
 sg13g2_or2_1 _5548_ (.X(_2245_),
    .B(\mac2.sum_lvl2_ff[9] ),
    .A(\mac2.sum_lvl2_ff[28] ));
 sg13g2_nand2b_1 _5549_ (.Y(_2246_),
    .B(_2245_),
    .A_N(_2244_));
 sg13g2_xnor2_1 _5550_ (.Y(_0047_),
    .A(_2243_),
    .B(_2246_));
 sg13g2_nand2_1 _5551_ (.Y(_2247_),
    .A(\mac2.sum_lvl2_ff[29] ),
    .B(\mac2.sum_lvl2_ff[10] ));
 sg13g2_xor2_1 _5552_ (.B(\mac2.sum_lvl2_ff[10] ),
    .A(\mac2.sum_lvl2_ff[29] ),
    .X(_2248_));
 sg13g2_inv_1 _5553_ (.Y(_2249_),
    .A(_2248_));
 sg13g2_a21o_2 _5554_ (.A2(_2245_),
    .A1(_2243_),
    .B1(_2244_),
    .X(_2250_));
 sg13g2_nand2_1 _5555_ (.Y(_2251_),
    .A(_2248_),
    .B(_2250_));
 sg13g2_xnor2_1 _5556_ (.Y(_0033_),
    .A(_2249_),
    .B(_2250_));
 sg13g2_nor2_1 _5557_ (.A(\mac2.sum_lvl2_ff[30] ),
    .B(\mac2.sum_lvl2_ff[11] ),
    .Y(_2252_));
 sg13g2_xnor2_1 _5558_ (.Y(_2253_),
    .A(\mac2.sum_lvl2_ff[30] ),
    .B(\mac2.sum_lvl2_ff[11] ));
 sg13g2_nand2_1 _5559_ (.Y(_2254_),
    .A(_2247_),
    .B(_2251_));
 sg13g2_xnor2_1 _5560_ (.Y(_0034_),
    .A(_2253_),
    .B(_2254_));
 sg13g2_nand2_1 _5561_ (.Y(_2255_),
    .A(\mac2.sum_lvl2_ff[31] ),
    .B(\mac2.sum_lvl2_ff[12] ));
 sg13g2_nor2_1 _5562_ (.A(\mac2.sum_lvl2_ff[31] ),
    .B(\mac2.sum_lvl2_ff[12] ),
    .Y(_2256_));
 sg13g2_xor2_1 _5563_ (.B(\mac2.sum_lvl2_ff[12] ),
    .A(\mac2.sum_lvl2_ff[31] ),
    .X(_2257_));
 sg13g2_nor2_1 _5564_ (.A(_2247_),
    .B(_2252_),
    .Y(_2258_));
 sg13g2_nor2_1 _5565_ (.A(_2249_),
    .B(_2253_),
    .Y(_2259_));
 sg13g2_a221oi_1 _5566_ (.B2(_2259_),
    .C1(_2258_),
    .B1(_2250_),
    .A1(\mac2.sum_lvl2_ff[30] ),
    .Y(_2260_),
    .A2(\mac2.sum_lvl2_ff[11] ));
 sg13g2_xnor2_1 _5567_ (.Y(_0035_),
    .A(_2257_),
    .B(_2260_));
 sg13g2_o21ai_1 _5568_ (.B1(_2255_),
    .Y(_2261_),
    .A1(_2256_),
    .A2(_2260_));
 sg13g2_and2_1 _5569_ (.A(\mac2.sum_lvl2_ff[32] ),
    .B(\mac2.sum_lvl2_ff[13] ),
    .X(_2262_));
 sg13g2_or2_1 _5570_ (.X(_2263_),
    .B(\mac2.sum_lvl2_ff[13] ),
    .A(\mac2.sum_lvl2_ff[32] ));
 sg13g2_nand2b_1 _5571_ (.Y(_2264_),
    .B(_2263_),
    .A_N(_2262_));
 sg13g2_xnor2_1 _5572_ (.Y(_0036_),
    .A(_2261_),
    .B(_2264_));
 sg13g2_a21oi_1 _5573_ (.A1(_2261_),
    .A2(_2263_),
    .Y(_2265_),
    .B1(_2262_));
 sg13g2_nand2_1 _5574_ (.Y(_2266_),
    .A(\mac2.sum_lvl2_ff[33] ),
    .B(\mac2.sum_lvl2_ff[14] ));
 sg13g2_nor2_1 _5575_ (.A(\mac2.sum_lvl2_ff[33] ),
    .B(\mac2.sum_lvl2_ff[14] ),
    .Y(_2267_));
 sg13g2_xor2_1 _5576_ (.B(net552),
    .A(\mac2.sum_lvl2_ff[33] ),
    .X(_2268_));
 sg13g2_xnor2_1 _5577_ (.Y(_0037_),
    .A(_2265_),
    .B(_2268_));
 sg13g2_o21ai_1 _5578_ (.B1(_2266_),
    .Y(_2269_),
    .A1(_2265_),
    .A2(_2267_));
 sg13g2_xnor2_1 _5579_ (.Y(_2270_),
    .A(\mac2.sum_lvl2_ff[34] ),
    .B(net484));
 sg13g2_xnor2_1 _5580_ (.Y(_0038_),
    .A(_2269_),
    .B(net485));
 sg13g2_xor2_1 _5581_ (.B(net271),
    .A(\mac2.sum_lvl2_ff[19] ),
    .X(_0032_));
 sg13g2_nand2_1 _5582_ (.Y(_2271_),
    .A(net480),
    .B(net325));
 sg13g2_nand2_1 _5583_ (.Y(_2272_),
    .A(\mac2.sum_lvl3_ff[21] ),
    .B(\mac2.sum_lvl3_ff[1] ));
 sg13g2_nor2_1 _5584_ (.A(\mac2.sum_lvl3_ff[21] ),
    .B(\mac2.sum_lvl3_ff[1] ),
    .Y(_2273_));
 sg13g2_xor2_1 _5585_ (.B(\mac2.sum_lvl3_ff[1] ),
    .A(\mac2.sum_lvl3_ff[21] ),
    .X(_2274_));
 sg13g2_xnor2_1 _5586_ (.Y(_0055_),
    .A(_2271_),
    .B(_2274_));
 sg13g2_o21ai_1 _5587_ (.B1(_2272_),
    .Y(_2275_),
    .A1(_2271_),
    .A2(_2273_));
 sg13g2_and2_1 _5588_ (.A(\mac2.sum_lvl3_ff[22] ),
    .B(net498),
    .X(_2276_));
 sg13g2_xor2_1 _5589_ (.B(net498),
    .A(\mac2.sum_lvl3_ff[22] ),
    .X(_2277_));
 sg13g2_xor2_1 _5590_ (.B(net499),
    .A(_2275_),
    .X(_0056_));
 sg13g2_a21oi_1 _5591_ (.A1(_2275_),
    .A2(_2277_),
    .Y(_2278_),
    .B1(_2276_));
 sg13g2_nand2_1 _5592_ (.Y(_2279_),
    .A(\mac2.sum_lvl3_ff[23] ),
    .B(\mac2.sum_lvl3_ff[3] ));
 sg13g2_xnor2_1 _5593_ (.Y(_2280_),
    .A(\mac2.sum_lvl3_ff[23] ),
    .B(net501));
 sg13g2_xor2_1 _5594_ (.B(net502),
    .A(_2278_),
    .X(_0057_));
 sg13g2_o21ai_1 _5595_ (.B1(_2279_),
    .Y(_2281_),
    .A1(_2278_),
    .A2(_2280_));
 sg13g2_and2_1 _5596_ (.A(\mac2.sum_lvl3_ff[24] ),
    .B(net444),
    .X(_2282_));
 sg13g2_xor2_1 _5597_ (.B(net444),
    .A(\mac2.sum_lvl3_ff[24] ),
    .X(_2283_));
 sg13g2_xor2_1 _5598_ (.B(net445),
    .A(_2281_),
    .X(_0058_));
 sg13g2_a21oi_1 _5599_ (.A1(_2281_),
    .A2(_2283_),
    .Y(_2284_),
    .B1(_2282_));
 sg13g2_nor2_1 _5600_ (.A(\mac2.sum_lvl3_ff[25] ),
    .B(net359),
    .Y(_2285_));
 sg13g2_xor2_1 _5601_ (.B(net359),
    .A(\mac2.sum_lvl3_ff[25] ),
    .X(_2286_));
 sg13g2_xnor2_1 _5602_ (.Y(_0059_),
    .A(_2284_),
    .B(net360));
 sg13g2_and2_1 _5603_ (.A(net487),
    .B(\mac2.sum_lvl3_ff[6] ),
    .X(_2287_));
 sg13g2_xnor2_1 _5604_ (.Y(_2288_),
    .A(net487),
    .B(\mac2.sum_lvl3_ff[6] ));
 sg13g2_a221oi_1 _5605_ (.B2(_2283_),
    .C1(_2282_),
    .B1(_2281_),
    .A1(\mac2.sum_lvl3_ff[25] ),
    .Y(_2289_),
    .A2(net359));
 sg13g2_nor3_1 _5606_ (.A(_2285_),
    .B(net488),
    .C(_2289_),
    .Y(_2290_));
 sg13g2_o21ai_1 _5607_ (.B1(net488),
    .Y(_2291_),
    .A1(_2285_),
    .A2(_2289_));
 sg13g2_nor2b_1 _5608_ (.A(_2290_),
    .B_N(net489),
    .Y(_0060_));
 sg13g2_nand2_1 _5609_ (.Y(_2292_),
    .A(net454),
    .B(\mac2.sum_lvl3_ff[7] ));
 sg13g2_xor2_1 _5610_ (.B(net545),
    .A(net454),
    .X(_2293_));
 sg13g2_o21ai_1 _5611_ (.B1(_2293_),
    .Y(_2294_),
    .A1(_2287_),
    .A2(_2290_));
 sg13g2_or3_1 _5612_ (.A(_2287_),
    .B(_2290_),
    .C(_2293_),
    .X(_2295_));
 sg13g2_and2_1 _5613_ (.A(_2294_),
    .B(_2295_),
    .X(_0061_));
 sg13g2_and2_1 _5614_ (.A(\mac2.sum_lvl3_ff[28] ),
    .B(\mac2.sum_lvl3_ff[8] ),
    .X(_2296_));
 sg13g2_xnor2_1 _5615_ (.Y(_2297_),
    .A(\mac2.sum_lvl3_ff[28] ),
    .B(\mac2.sum_lvl3_ff[8] ));
 sg13g2_a21oi_1 _5616_ (.A1(net455),
    .A2(_2294_),
    .Y(_2298_),
    .B1(_2297_));
 sg13g2_nand3_1 _5617_ (.B(_2294_),
    .C(_2297_),
    .A(net455),
    .Y(_2299_));
 sg13g2_nor2b_1 _5618_ (.A(_2298_),
    .B_N(net456),
    .Y(_0062_));
 sg13g2_nor2_1 _5619_ (.A(_2296_),
    .B(_2298_),
    .Y(_2300_));
 sg13g2_nand2_1 _5620_ (.Y(_2301_),
    .A(\mac2.sum_lvl3_ff[29] ),
    .B(net315));
 sg13g2_xor2_1 _5621_ (.B(net315),
    .A(\mac2.sum_lvl3_ff[29] ),
    .X(_2302_));
 sg13g2_o21ai_1 _5622_ (.B1(_2302_),
    .Y(_2303_),
    .A1(_2296_),
    .A2(_2298_));
 sg13g2_xnor2_1 _5623_ (.Y(_0063_),
    .A(_2300_),
    .B(net316));
 sg13g2_nand2_1 _5624_ (.Y(_2304_),
    .A(_2301_),
    .B(_2303_));
 sg13g2_nand2_1 _5625_ (.Y(_2305_),
    .A(net401),
    .B(net346));
 sg13g2_xor2_1 _5626_ (.B(net346),
    .A(\mac2.sum_lvl3_ff[30] ),
    .X(_2306_));
 sg13g2_nand2_1 _5627_ (.Y(_2307_),
    .A(_2304_),
    .B(net347));
 sg13g2_xor2_1 _5628_ (.B(net347),
    .A(_2304_),
    .X(_0049_));
 sg13g2_nor2_1 _5629_ (.A(\mac2.sum_lvl3_ff[31] ),
    .B(\mac2.sum_lvl3_ff[11] ),
    .Y(_2308_));
 sg13g2_nand2_1 _5630_ (.Y(_2309_),
    .A(\mac2.sum_lvl3_ff[31] ),
    .B(\mac2.sum_lvl3_ff[11] ));
 sg13g2_nand2b_1 _5631_ (.Y(_2310_),
    .B(_2309_),
    .A_N(_2308_));
 sg13g2_nand2_1 _5632_ (.Y(_2311_),
    .A(_2305_),
    .B(_2307_));
 sg13g2_xnor2_1 _5633_ (.Y(_0050_),
    .A(_2310_),
    .B(net402));
 sg13g2_nand2_1 _5634_ (.Y(_2312_),
    .A(\mac2.sum_lvl3_ff[32] ),
    .B(\mac2.sum_lvl3_ff[12] ));
 sg13g2_xor2_1 _5635_ (.B(net530),
    .A(\mac2.sum_lvl3_ff[32] ),
    .X(_2313_));
 sg13g2_o21ai_1 _5636_ (.B1(_2309_),
    .Y(_2314_),
    .A1(_2305_),
    .A2(_2308_));
 sg13g2_nand3b_1 _5637_ (.B(_2309_),
    .C(_2306_),
    .Y(_2315_),
    .A_N(_2308_));
 sg13g2_a21oi_1 _5638_ (.A1(_2301_),
    .A2(_2303_),
    .Y(_2316_),
    .B1(_2315_));
 sg13g2_o21ai_1 _5639_ (.B1(net531),
    .Y(_2317_),
    .A1(_2314_),
    .A2(_2316_));
 sg13g2_or3_1 _5640_ (.A(net531),
    .B(_2314_),
    .C(_2316_),
    .X(_2318_));
 sg13g2_and2_1 _5641_ (.A(_2317_),
    .B(_2318_),
    .X(_0051_));
 sg13g2_xnor2_1 _5642_ (.Y(_2319_),
    .A(\mac2.sum_lvl3_ff[33] ),
    .B(net410));
 sg13g2_a21oi_1 _5643_ (.A1(_2312_),
    .A2(_2317_),
    .Y(_2320_),
    .B1(net411));
 sg13g2_nand3_1 _5644_ (.B(_2317_),
    .C(net411),
    .A(_2312_),
    .Y(_2321_));
 sg13g2_nor2b_1 _5645_ (.A(net412),
    .B_N(_2321_),
    .Y(_0052_));
 sg13g2_a21oi_1 _5646_ (.A1(\mac2.sum_lvl3_ff[33] ),
    .A2(net410),
    .Y(_2322_),
    .B1(_2320_));
 sg13g2_nand2_1 _5647_ (.Y(_2323_),
    .A(\mac2.sum_lvl3_ff[34] ),
    .B(net297));
 sg13g2_nor2_1 _5648_ (.A(\mac2.sum_lvl3_ff[34] ),
    .B(net297),
    .Y(_2324_));
 sg13g2_xor2_1 _5649_ (.B(net297),
    .A(\mac2.sum_lvl3_ff[34] ),
    .X(_2325_));
 sg13g2_xnor2_1 _5650_ (.Y(_0053_),
    .A(_2322_),
    .B(net298));
 sg13g2_o21ai_1 _5651_ (.B1(_2323_),
    .Y(_2326_),
    .A1(_2322_),
    .A2(_2324_));
 sg13g2_xnor2_1 _5652_ (.Y(_2327_),
    .A(net437),
    .B(\mac2.sum_lvl3_ff[15] ));
 sg13g2_xnor2_1 _5653_ (.Y(_0054_),
    .A(_2326_),
    .B(net438));
 sg13g2_xor2_1 _5654_ (.B(net325),
    .A(\mac2.sum_lvl3_ff[20] ),
    .X(_0048_));
 sg13g2_nand2_1 _5655_ (.Y(_2328_),
    .A(\mac1.total_sum[0] ),
    .B(\mac2.total_sum[0] ));
 sg13g2_nand2_1 _5656_ (.Y(_2329_),
    .A(\mac1.total_sum[1] ),
    .B(\mac2.total_sum[1] ));
 sg13g2_nor2_1 _5657_ (.A(\mac1.total_sum[1] ),
    .B(\mac2.total_sum[1] ),
    .Y(_2330_));
 sg13g2_xor2_1 _5658_ (.B(\mac2.total_sum[1] ),
    .A(\mac1.total_sum[1] ),
    .X(_2331_));
 sg13g2_xnor2_1 _5659_ (.Y(net26),
    .A(_2328_),
    .B(_2331_));
 sg13g2_o21ai_1 _5660_ (.B1(_2329_),
    .Y(_2332_),
    .A1(_2328_),
    .A2(_2330_));
 sg13g2_and2_1 _5661_ (.A(\mac1.total_sum[2] ),
    .B(\mac2.total_sum[2] ),
    .X(_2333_));
 sg13g2_xor2_1 _5662_ (.B(\mac2.total_sum[2] ),
    .A(\mac1.total_sum[2] ),
    .X(_2334_));
 sg13g2_xor2_1 _5663_ (.B(_2334_),
    .A(_2332_),
    .X(net27));
 sg13g2_a21oi_1 _5664_ (.A1(_2332_),
    .A2(_2334_),
    .Y(_2335_),
    .B1(_2333_));
 sg13g2_nand2_1 _5665_ (.Y(_2336_),
    .A(\mac1.total_sum[3] ),
    .B(\mac2.total_sum[3] ));
 sg13g2_xnor2_1 _5666_ (.Y(_2337_),
    .A(\mac1.total_sum[3] ),
    .B(\mac2.total_sum[3] ));
 sg13g2_xor2_1 _5667_ (.B(_2337_),
    .A(_2335_),
    .X(net28));
 sg13g2_o21ai_1 _5668_ (.B1(_2336_),
    .Y(_2338_),
    .A1(_2335_),
    .A2(_2337_));
 sg13g2_and2_1 _5669_ (.A(\mac1.total_sum[4] ),
    .B(\mac2.total_sum[4] ),
    .X(_2339_));
 sg13g2_xor2_1 _5670_ (.B(\mac2.total_sum[4] ),
    .A(\mac1.total_sum[4] ),
    .X(_2340_));
 sg13g2_xor2_1 _5671_ (.B(_2340_),
    .A(_2338_),
    .X(net29));
 sg13g2_a21oi_1 _5672_ (.A1(_2338_),
    .A2(_2340_),
    .Y(_2341_),
    .B1(_2339_));
 sg13g2_nor2_1 _5673_ (.A(\mac1.total_sum[5] ),
    .B(\mac2.total_sum[5] ),
    .Y(_2342_));
 sg13g2_xor2_1 _5674_ (.B(\mac2.total_sum[5] ),
    .A(\mac1.total_sum[5] ),
    .X(_2343_));
 sg13g2_xnor2_1 _5675_ (.Y(net30),
    .A(_2341_),
    .B(_2343_));
 sg13g2_and2_1 _5676_ (.A(\mac1.total_sum[6] ),
    .B(\mac2.total_sum[6] ),
    .X(_2344_));
 sg13g2_xnor2_1 _5677_ (.Y(_2345_),
    .A(\mac1.total_sum[6] ),
    .B(\mac2.total_sum[6] ));
 sg13g2_a221oi_1 _5678_ (.B2(_2340_),
    .C1(_2339_),
    .B1(_2338_),
    .A1(\mac1.total_sum[5] ),
    .Y(_2346_),
    .A2(\mac2.total_sum[5] ));
 sg13g2_nor3_1 _5679_ (.A(_2342_),
    .B(_2345_),
    .C(_2346_),
    .Y(_2347_));
 sg13g2_o21ai_1 _5680_ (.B1(_2345_),
    .Y(_2348_),
    .A1(_2342_),
    .A2(_2346_));
 sg13g2_nor2b_2 _5681_ (.A(_2347_),
    .B_N(_2348_),
    .Y(net31));
 sg13g2_nand2_1 _5682_ (.Y(_2349_),
    .A(\mac1.total_sum[7] ),
    .B(\mac2.total_sum[7] ));
 sg13g2_xor2_1 _5683_ (.B(\mac2.total_sum[7] ),
    .A(\mac1.total_sum[7] ),
    .X(_2350_));
 sg13g2_o21ai_1 _5684_ (.B1(_2350_),
    .Y(_2351_),
    .A1(_2344_),
    .A2(_2347_));
 sg13g2_or3_1 _5685_ (.A(_2344_),
    .B(_2347_),
    .C(_2350_),
    .X(_2352_));
 sg13g2_and2_1 _5686_ (.A(_2351_),
    .B(_2352_),
    .X(net32));
 sg13g2_xnor2_1 _5687_ (.Y(_2353_),
    .A(\mac1.total_sum[8] ),
    .B(\mac2.total_sum[8] ));
 sg13g2_a21oi_1 _5688_ (.A1(_2349_),
    .A2(_2351_),
    .Y(_2354_),
    .B1(_2353_));
 sg13g2_nand3_1 _5689_ (.B(_2351_),
    .C(_2353_),
    .A(_2349_),
    .Y(_2355_));
 sg13g2_nor2b_2 _5690_ (.A(_2354_),
    .B_N(_2355_),
    .Y(net17));
 sg13g2_a21o_1 _5691_ (.A2(\mac2.total_sum[8] ),
    .A1(\mac1.total_sum[8] ),
    .B1(_2354_),
    .X(_2356_));
 sg13g2_and2_1 _5692_ (.A(\mac1.total_sum[9] ),
    .B(\mac2.total_sum[9] ),
    .X(_2357_));
 sg13g2_or2_1 _5693_ (.X(_2358_),
    .B(\mac2.total_sum[9] ),
    .A(\mac1.total_sum[9] ));
 sg13g2_nand2b_1 _5694_ (.Y(_2359_),
    .B(_2358_),
    .A_N(_2357_));
 sg13g2_xnor2_1 _5695_ (.Y(net18),
    .A(_2356_),
    .B(_2359_));
 sg13g2_nand2_1 _5696_ (.Y(_2360_),
    .A(\mac1.total_sum[10] ),
    .B(\mac2.total_sum[10] ));
 sg13g2_xor2_1 _5697_ (.B(\mac2.total_sum[10] ),
    .A(\mac1.total_sum[10] ),
    .X(_2361_));
 sg13g2_inv_1 _5698_ (.Y(_2362_),
    .A(_2361_));
 sg13g2_a21o_1 _5699_ (.A2(_2358_),
    .A1(_2356_),
    .B1(_2357_),
    .X(_2363_));
 sg13g2_nand2_1 _5700_ (.Y(_2364_),
    .A(_2361_),
    .B(_2363_));
 sg13g2_xnor2_1 _5701_ (.Y(net19),
    .A(_2362_),
    .B(_2363_));
 sg13g2_nor2_1 _5702_ (.A(\mac1.total_sum[11] ),
    .B(\mac2.total_sum[11] ),
    .Y(_2365_));
 sg13g2_xnor2_1 _5703_ (.Y(_2366_),
    .A(\mac1.total_sum[11] ),
    .B(\mac2.total_sum[11] ));
 sg13g2_nand2_1 _5704_ (.Y(_2367_),
    .A(_2360_),
    .B(_2364_));
 sg13g2_xnor2_1 _5705_ (.Y(net20),
    .A(_2366_),
    .B(_2367_));
 sg13g2_nand2_1 _5706_ (.Y(_2368_),
    .A(\mac1.total_sum[12] ),
    .B(\mac2.total_sum[12] ));
 sg13g2_nor2_1 _5707_ (.A(\mac1.total_sum[12] ),
    .B(\mac2.total_sum[12] ),
    .Y(_2369_));
 sg13g2_xor2_1 _5708_ (.B(\mac2.total_sum[12] ),
    .A(\mac1.total_sum[12] ),
    .X(_2370_));
 sg13g2_nor2_1 _5709_ (.A(_2360_),
    .B(_2365_),
    .Y(_2371_));
 sg13g2_nor2_1 _5710_ (.A(_2362_),
    .B(_2366_),
    .Y(_2372_));
 sg13g2_a221oi_1 _5711_ (.B2(_2372_),
    .C1(_2371_),
    .B1(_2363_),
    .A1(\mac1.total_sum[11] ),
    .Y(_2373_),
    .A2(\mac2.total_sum[11] ));
 sg13g2_xnor2_1 _5712_ (.Y(net21),
    .A(_2370_),
    .B(_2373_));
 sg13g2_o21ai_1 _5713_ (.B1(_2368_),
    .Y(_2374_),
    .A1(_2369_),
    .A2(_2373_));
 sg13g2_and2_1 _5714_ (.A(\mac1.total_sum[13] ),
    .B(\mac2.total_sum[13] ),
    .X(_2375_));
 sg13g2_or2_1 _5715_ (.X(_2376_),
    .B(\mac2.total_sum[13] ),
    .A(\mac1.total_sum[13] ));
 sg13g2_nand2b_1 _5716_ (.Y(_2377_),
    .B(_2376_),
    .A_N(_2375_));
 sg13g2_xnor2_1 _5717_ (.Y(net22),
    .A(_2374_),
    .B(_2377_));
 sg13g2_a21oi_1 _5718_ (.A1(_2374_),
    .A2(_2376_),
    .Y(_2378_),
    .B1(_2375_));
 sg13g2_nand2_1 _5719_ (.Y(_2379_),
    .A(\mac1.total_sum[14] ),
    .B(\mac2.total_sum[14] ));
 sg13g2_nor2_1 _5720_ (.A(\mac1.total_sum[14] ),
    .B(\mac2.total_sum[14] ),
    .Y(_2380_));
 sg13g2_xor2_1 _5721_ (.B(\mac2.total_sum[14] ),
    .A(\mac1.total_sum[14] ),
    .X(_2381_));
 sg13g2_xnor2_1 _5722_ (.Y(net23),
    .A(_2378_),
    .B(_2381_));
 sg13g2_o21ai_1 _5723_ (.B1(_2379_),
    .Y(_2382_),
    .A1(_2378_),
    .A2(_2380_));
 sg13g2_xnor2_1 _5724_ (.Y(_2383_),
    .A(\mac1.total_sum[15] ),
    .B(\mac2.total_sum[15] ));
 sg13g2_xnor2_1 _5725_ (.Y(net24),
    .A(_2382_),
    .B(_2383_));
 sg13g2_xor2_1 _5726_ (.B(\mac2.total_sum[0] ),
    .A(\mac1.total_sum[0] ),
    .X(net25));
 sg13g2_nor2b_1 _5727_ (.A(\DP_1.Q_range.out_data[4] ),
    .B_N(\DP_1.I_range.out_data[5] ),
    .Y(_2384_));
 sg13g2_o21ai_1 _5728_ (.B1(_2384_),
    .Y(_2385_),
    .A1(\DP_1.I_range.out_data[3] ),
    .A2(\DP_1.Q_range.out_data[5] ));
 sg13g2_nand2_1 _5729_ (.Y(_2386_),
    .A(\DP_1.I_range.out_data[2] ),
    .B(\DP_1.Q_range.out_data[2] ));
 sg13g2_nand3b_1 _5730_ (.B(\DP_1.Q_range.out_data[3] ),
    .C(\DP_1.Q_range.out_data[5] ),
    .Y(_2387_),
    .A_N(\DP_1.I_range.out_data[3] ));
 sg13g2_nor2b_1 _5731_ (.A(\DP_1.Q_range.out_data[3] ),
    .B_N(\DP_1.I_range.out_data[3] ),
    .Y(_2388_));
 sg13g2_o21ai_1 _5732_ (.B1(\DP_1.I_range.out_data[4] ),
    .Y(_2389_),
    .A1(_2386_),
    .A2(_2388_));
 sg13g2_nor3_1 _5733_ (.A(\DP_1.I_range.out_data[4] ),
    .B(_2386_),
    .C(_2388_),
    .Y(_2390_));
 sg13g2_a21oi_1 _5734_ (.A1(_2386_),
    .A2(_2387_),
    .Y(_2391_),
    .B1(_2390_));
 sg13g2_nand2_1 _5735_ (.Y(_2392_),
    .A(_2389_),
    .B(_2391_));
 sg13g2_nor4_2 _5736_ (.A(\DP_1.I_range.out_data[2] ),
    .B(\DP_1.Q_range.out_data[2] ),
    .C(_2385_),
    .Y(_2393_),
    .D(_2392_));
 sg13g2_nor2_1 _5737_ (.A(net1059),
    .B(net786),
    .Y(_2394_));
 sg13g2_xor2_1 _5738_ (.B(\DP_1.Q_range.out_data[3] ),
    .A(\DP_1.I_range.out_data[3] ),
    .X(_2395_));
 sg13g2_xor2_1 _5739_ (.B(\DP_1.Q_range.out_data[2] ),
    .A(\DP_1.I_range.out_data[2] ),
    .X(_2396_));
 sg13g2_xnor2_1 _5740_ (.Y(_2397_),
    .A(\DP_1.I_range.out_data[2] ),
    .B(\DP_1.Q_range.out_data[2] ));
 sg13g2_nor2_1 _5741_ (.A(_2395_),
    .B(net809),
    .Y(_2398_));
 sg13g2_nand2_1 _5742_ (.Y(_2399_),
    .A(net418),
    .B(net801));
 sg13g2_nor2b_2 _5743_ (.A(\DP_1.Q_range.out_data[2] ),
    .B_N(\DP_1.I_range.out_data[2] ),
    .Y(_2400_));
 sg13g2_xor2_1 _5744_ (.B(_2400_),
    .A(_2395_),
    .X(_2401_));
 sg13g2_xnor2_1 _5745_ (.Y(_2402_),
    .A(_2395_),
    .B(_2400_));
 sg13g2_nor2_1 _5746_ (.A(net1059),
    .B(net810),
    .Y(_2403_));
 sg13g2_o21ai_1 _5747_ (.B1(net799),
    .Y(_2404_),
    .A1(\DP_1.matrix[44] ),
    .A2(net808));
 sg13g2_o21ai_1 _5748_ (.B1(_2399_),
    .Y(_2405_),
    .A1(_2403_),
    .A2(_2404_));
 sg13g2_a21oi_1 _5749_ (.A1(net787),
    .A2(_2405_),
    .Y(_2406_),
    .B1(_2394_));
 sg13g2_mux2_1 _5750_ (.A0(\DP_1.matrix[5] ),
    .A1(net1012),
    .S(net810),
    .X(_2407_));
 sg13g2_a22oi_1 _5751_ (.Y(_2408_),
    .B1(net800),
    .B2(_2407_),
    .A2(net802),
    .A1(\DP_1.matrix[77] ));
 sg13g2_and2_1 _5752_ (.A(net1034),
    .B(_2397_),
    .X(_2409_));
 sg13g2_a21oi_1 _5753_ (.A1(net1017),
    .A2(net809),
    .Y(_2410_),
    .B1(_2409_));
 sg13g2_nand3_1 _5754_ (.B(net808),
    .C(_2402_),
    .A(net997),
    .Y(_2411_));
 sg13g2_o21ai_1 _5755_ (.B1(_2411_),
    .Y(_2412_),
    .A1(_2402_),
    .A2(_2410_));
 sg13g2_nand2_1 _5756_ (.Y(_2413_),
    .A(net1003),
    .B(net801));
 sg13g2_nor2_1 _5757_ (.A(net1040),
    .B(net809),
    .Y(_2414_));
 sg13g2_o21ai_1 _5758_ (.B1(net799),
    .Y(_2415_),
    .A1(net1023),
    .A2(net808));
 sg13g2_o21ai_1 _5759_ (.B1(_2413_),
    .Y(_2416_),
    .A1(_2414_),
    .A2(_2415_));
 sg13g2_nand2_1 _5760_ (.Y(_2417_),
    .A(_2395_),
    .B(net808));
 sg13g2_a22oi_1 _5761_ (.Y(_2418_),
    .B1(net799),
    .B2(net1022),
    .A2(net808),
    .A1(net1002));
 sg13g2_nor2_1 _5762_ (.A(net1038),
    .B(_2417_),
    .Y(_2419_));
 sg13g2_a21oi_1 _5763_ (.A1(_2417_),
    .A2(_2418_),
    .Y(_2420_),
    .B1(_2419_));
 sg13g2_and2_1 _5764_ (.A(_2416_),
    .B(_2420_),
    .X(_2421_));
 sg13g2_mux2_1 _5765_ (.A0(net1036),
    .A1(net1020),
    .S(net809),
    .X(_2422_));
 sg13g2_a22oi_1 _5766_ (.Y(_2423_),
    .B1(net800),
    .B2(_2422_),
    .A2(net801),
    .A1(net999));
 sg13g2_nor2b_1 _5767_ (.A(_2423_),
    .B_N(_2421_),
    .Y(_2424_));
 sg13g2_nand2_1 _5768_ (.Y(_2425_),
    .A(_2412_),
    .B(_2424_));
 sg13g2_mux2_1 _5769_ (.A0(net1033),
    .A1(net1015),
    .S(net810),
    .X(_2426_));
 sg13g2_a22oi_1 _5770_ (.Y(_2427_),
    .B1(net800),
    .B2(_2426_),
    .A2(net802),
    .A1(\DP_1.matrix[76] ));
 sg13g2_or2_1 _5771_ (.X(_2428_),
    .B(_2427_),
    .A(_2425_));
 sg13g2_or2_1 _5772_ (.X(_2429_),
    .B(_2428_),
    .A(_2408_));
 sg13g2_mux2_1 _5773_ (.A0(net1029),
    .A1(\DP_1.matrix[42] ),
    .S(net810),
    .X(_2430_));
 sg13g2_a22oi_1 _5774_ (.Y(_2431_),
    .B1(net800),
    .B2(_2430_),
    .A2(net802),
    .A1(\DP_1.matrix[78] ));
 sg13g2_nor2_1 _5775_ (.A(_2429_),
    .B(_2431_),
    .Y(_2432_));
 sg13g2_inv_1 _5776_ (.Y(_2433_),
    .A(_2432_));
 sg13g2_mux2_1 _5777_ (.A0(net1026),
    .A1(\DP_1.matrix[43] ),
    .S(net810),
    .X(_2434_));
 sg13g2_a22oi_1 _5778_ (.Y(_2435_),
    .B1(net800),
    .B2(_2434_),
    .A2(net802),
    .A1(\DP_1.matrix[79] ));
 sg13g2_o21ai_1 _5779_ (.B1(net786),
    .Y(_2436_),
    .A1(_2433_),
    .A2(_2435_));
 sg13g2_mux2_1 _5780_ (.A0(_2405_),
    .A1(_2406_),
    .S(_2436_),
    .X(_0160_));
 sg13g2_nor2_1 _5781_ (.A(net1053),
    .B(net784),
    .Y(_2437_));
 sg13g2_nand2_1 _5782_ (.Y(_2438_),
    .A(net386),
    .B(net802));
 sg13g2_nor2_1 _5783_ (.A(net1053),
    .B(net809),
    .Y(_2439_));
 sg13g2_o21ai_1 _5784_ (.B1(net799),
    .Y(_2440_),
    .A1(net1052),
    .A2(_2397_));
 sg13g2_o21ai_1 _5785_ (.B1(_2438_),
    .Y(_2441_),
    .A1(_2439_),
    .A2(_2440_));
 sg13g2_a21oi_1 _5786_ (.A1(net784),
    .A2(_2441_),
    .Y(_2442_),
    .B1(_2437_));
 sg13g2_mux2_1 _5787_ (.A0(net971),
    .A1(\DP_2.matrix[41] ),
    .S(net809),
    .X(_2443_));
 sg13g2_a22oi_1 _5788_ (.Y(_2444_),
    .B1(net799),
    .B2(_2443_),
    .A2(net801),
    .A1(net931));
 sg13g2_and2_1 _5789_ (.A(net974),
    .B(_2397_),
    .X(_2445_));
 sg13g2_a21oi_1 _5790_ (.A1(net955),
    .A2(net809),
    .Y(_2446_),
    .B1(_2445_));
 sg13g2_nand3_1 _5791_ (.B(net808),
    .C(_2402_),
    .A(\DP_2.matrix[75] ),
    .Y(_2447_));
 sg13g2_o21ai_1 _5792_ (.B1(_2447_),
    .Y(_2448_),
    .A1(_2402_),
    .A2(_2446_));
 sg13g2_nand2_1 _5793_ (.Y(_2449_),
    .A(net946),
    .B(net801));
 sg13g2_nor2_1 _5794_ (.A(net982),
    .B(net809),
    .Y(_2450_));
 sg13g2_o21ai_1 _5795_ (.B1(net799),
    .Y(_2451_),
    .A1(net965),
    .A2(net808));
 sg13g2_o21ai_1 _5796_ (.B1(_2449_),
    .Y(_2452_),
    .A1(_2450_),
    .A2(_2451_));
 sg13g2_a22oi_1 _5797_ (.Y(_2453_),
    .B1(net799),
    .B2(net961),
    .A2(net808),
    .A1(net942));
 sg13g2_nor2_1 _5798_ (.A(net978),
    .B(_2417_),
    .Y(_2454_));
 sg13g2_a21oi_1 _5799_ (.A1(_2417_),
    .A2(_2453_),
    .Y(_2455_),
    .B1(_2454_));
 sg13g2_and2_1 _5800_ (.A(_2452_),
    .B(_2455_),
    .X(_2456_));
 sg13g2_mux2_1 _5801_ (.A0(net976),
    .A1(net957),
    .S(net810),
    .X(_2457_));
 sg13g2_a22oi_1 _5802_ (.Y(_2458_),
    .B1(net800),
    .B2(_2457_),
    .A2(net801),
    .A1(net937));
 sg13g2_nor2b_1 _5803_ (.A(_2458_),
    .B_N(_2456_),
    .Y(_2459_));
 sg13g2_nand2_1 _5804_ (.Y(_2460_),
    .A(_2448_),
    .B(_2459_));
 sg13g2_mux2_1 _5805_ (.A0(net972),
    .A1(net953),
    .S(net810),
    .X(_2461_));
 sg13g2_a22oi_1 _5806_ (.Y(_2462_),
    .B1(net799),
    .B2(_2461_),
    .A2(net801),
    .A1(net404));
 sg13g2_or2_1 _5807_ (.X(_2463_),
    .B(_2462_),
    .A(_2460_));
 sg13g2_or2_1 _5808_ (.X(_2464_),
    .B(_2463_),
    .A(_2444_));
 sg13g2_mux2_1 _5809_ (.A0(net969),
    .A1(net950),
    .S(_2396_),
    .X(_2465_));
 sg13g2_a22oi_1 _5810_ (.Y(_2466_),
    .B1(net800),
    .B2(_2465_),
    .A2(net801),
    .A1(\DP_2.matrix[78] ));
 sg13g2_nor2_1 _5811_ (.A(_2464_),
    .B(_2466_),
    .Y(_2467_));
 sg13g2_inv_1 _5812_ (.Y(_2468_),
    .A(_2467_));
 sg13g2_mux2_1 _5813_ (.A0(net968),
    .A1(net948),
    .S(_2396_),
    .X(_2469_));
 sg13g2_a22oi_1 _5814_ (.Y(_2470_),
    .B1(net800),
    .B2(_2469_),
    .A2(net802),
    .A1(\DP_2.matrix[79] ));
 sg13g2_o21ai_1 _5815_ (.B1(net784),
    .Y(_2471_),
    .A1(_2468_),
    .A2(_2470_));
 sg13g2_mux2_1 _5816_ (.A0(_2441_),
    .A1(_2442_),
    .S(_2471_),
    .X(_0163_));
 sg13g2_nand2_1 _5817_ (.Y(_2472_),
    .A(\DP_3.Q_range.out_data[3] ),
    .B(\DP_3.Q_range.out_data[5] ));
 sg13g2_nor3_1 _5818_ (.A(\DP_3.Q_range.out_data[2] ),
    .B(net505),
    .C(_2472_),
    .Y(_2473_));
 sg13g2_nor4_1 _5819_ (.A(\DP_3.I_range.out_data[2] ),
    .B(\DP_3.I_range.out_data[3] ),
    .C(_2633_),
    .D(\DP_3.I_range.out_data[4] ),
    .Y(_2474_));
 sg13g2_nand2_2 _5820_ (.Y(_2475_),
    .A(net506),
    .B(_2474_));
 sg13g2_xor2_1 _5821_ (.B(\DP_3.Q_range.out_data[3] ),
    .A(\DP_3.I_range.out_data[3] ),
    .X(_2476_));
 sg13g2_nor2b_1 _5822_ (.A(\DP_3.Q_range.out_data[2] ),
    .B_N(\DP_3.I_range.out_data[2] ),
    .Y(_2477_));
 sg13g2_xnor2_1 _5823_ (.Y(_2478_),
    .A(\DP_3.I_range.out_data[2] ),
    .B(\DP_3.Q_range.out_data[2] ));
 sg13g2_xor2_1 _5824_ (.B(\DP_3.Q_range.out_data[2] ),
    .A(\DP_3.I_range.out_data[2] ),
    .X(_2479_));
 sg13g2_nor2_1 _5825_ (.A(_2476_),
    .B(net805),
    .Y(_2480_));
 sg13g2_xnor2_1 _5826_ (.Y(_2481_),
    .A(_2476_),
    .B(_2477_));
 sg13g2_nor2_1 _5827_ (.A(net896),
    .B(net807),
    .Y(_2482_));
 sg13g2_nor2_1 _5828_ (.A(net915),
    .B(net804),
    .Y(_2483_));
 sg13g2_nor3_1 _5829_ (.A(net794),
    .B(_2482_),
    .C(_2483_),
    .Y(_2484_));
 sg13g2_a21oi_1 _5830_ (.A1(net277),
    .A2(net797),
    .Y(_2485_),
    .B1(_2484_));
 sg13g2_and2_1 _5831_ (.A(net900),
    .B(net805),
    .X(_2486_));
 sg13g2_a21oi_1 _5832_ (.A1(net918),
    .A2(net806),
    .Y(_2487_),
    .B1(_2486_));
 sg13g2_nand3_1 _5833_ (.B(net806),
    .C(net795),
    .A(net882),
    .Y(_2488_));
 sg13g2_o21ai_1 _5834_ (.B1(_2488_),
    .Y(_2489_),
    .A1(net795),
    .A2(_2487_));
 sg13g2_nand2_1 _5835_ (.Y(_2490_),
    .A(net275),
    .B(net798));
 sg13g2_a21oi_1 _5836_ (.A1(_2634_),
    .A2(net805),
    .Y(_2491_),
    .B1(net795));
 sg13g2_o21ai_1 _5837_ (.B1(_2491_),
    .Y(_2492_),
    .A1(net924),
    .A2(net805));
 sg13g2_nand2_1 _5838_ (.Y(_2493_),
    .A(_2490_),
    .B(_2492_));
 sg13g2_nand2b_1 _5839_ (.Y(_2494_),
    .B(net905),
    .A_N(net795));
 sg13g2_nand2_1 _5840_ (.Y(_2495_),
    .A(_2476_),
    .B(net806));
 sg13g2_o21ai_1 _5841_ (.B1(net806),
    .Y(_2496_),
    .A1(net888),
    .A2(_2476_));
 sg13g2_nor2_1 _5842_ (.A(net923),
    .B(_2495_),
    .Y(_2497_));
 sg13g2_a21oi_1 _5843_ (.A1(_2494_),
    .A2(_2496_),
    .Y(_2498_),
    .B1(_2497_));
 sg13g2_and2_1 _5844_ (.A(_2493_),
    .B(_2498_),
    .X(_2499_));
 sg13g2_nor2_1 _5845_ (.A(net920),
    .B(net805),
    .Y(_2500_));
 sg13g2_nor2_1 _5846_ (.A(net902),
    .B(net806),
    .Y(_2501_));
 sg13g2_nor3_1 _5847_ (.A(net795),
    .B(_2500_),
    .C(_2501_),
    .Y(_2502_));
 sg13g2_a21oi_1 _5848_ (.A1(net885),
    .A2(net798),
    .Y(_2503_),
    .B1(_2502_));
 sg13g2_nor2b_1 _5849_ (.A(_2503_),
    .B_N(_2499_),
    .Y(_2504_));
 sg13g2_nand2_1 _5850_ (.Y(_2505_),
    .A(_2489_),
    .B(_2504_));
 sg13g2_nor2_1 _5851_ (.A(net916),
    .B(net804),
    .Y(_2506_));
 sg13g2_nor2_1 _5852_ (.A(net898),
    .B(net807),
    .Y(_2507_));
 sg13g2_nor3_1 _5853_ (.A(net794),
    .B(_2506_),
    .C(_2507_),
    .Y(_2508_));
 sg13g2_a21oi_1 _5854_ (.A1(net879),
    .A2(net797),
    .Y(_2509_),
    .B1(_2508_));
 sg13g2_or2_1 _5855_ (.X(_2510_),
    .B(_2509_),
    .A(_2505_));
 sg13g2_or2_1 _5856_ (.X(_2511_),
    .B(_2510_),
    .A(_2485_));
 sg13g2_nand2_1 _5857_ (.Y(_2512_),
    .A(net279),
    .B(net797));
 sg13g2_nand2b_1 _5858_ (.Y(_2513_),
    .B(net803),
    .A_N(net895));
 sg13g2_o21ai_1 _5859_ (.B1(_2513_),
    .Y(_2514_),
    .A1(net913),
    .A2(net803));
 sg13g2_o21ai_1 _5860_ (.B1(_2512_),
    .Y(_2515_),
    .A1(net794),
    .A2(_2514_));
 sg13g2_nor2b_1 _5861_ (.A(_2511_),
    .B_N(_2515_),
    .Y(_2516_));
 sg13g2_nor2_1 _5862_ (.A(net910),
    .B(net803),
    .Y(_2517_));
 sg13g2_nor2_1 _5863_ (.A(net892),
    .B(net807),
    .Y(_2518_));
 sg13g2_nor3_1 _5864_ (.A(net796),
    .B(_2517_),
    .C(_2518_),
    .Y(_2519_));
 sg13g2_a21oi_1 _5865_ (.A1(net276),
    .A2(net798),
    .Y(_2520_),
    .B1(_2519_));
 sg13g2_inv_1 _5866_ (.Y(_2521_),
    .A(_2520_));
 sg13g2_a21oi_1 _5867_ (.A1(_2516_),
    .A2(_2521_),
    .Y(_2522_),
    .B1(net792));
 sg13g2_nand2_1 _5868_ (.Y(_2523_),
    .A(net1050),
    .B(net791));
 sg13g2_nor2_1 _5869_ (.A(net1050),
    .B(net804),
    .Y(_2524_));
 sg13g2_nor2_1 _5870_ (.A(net1047),
    .B(net807),
    .Y(_2525_));
 sg13g2_nor3_1 _5871_ (.A(net794),
    .B(_2524_),
    .C(_2525_),
    .Y(_2526_));
 sg13g2_a21oi_1 _5872_ (.A1(net273),
    .A2(net797),
    .Y(_2527_),
    .B1(_2526_));
 sg13g2_o21ai_1 _5873_ (.B1(_2523_),
    .Y(_2528_),
    .A1(net791),
    .A2(_2526_));
 sg13g2_nor2_1 _5874_ (.A(_2522_),
    .B(_2528_),
    .Y(_2529_));
 sg13g2_a21oi_1 _5875_ (.A1(_2522_),
    .A2(_2527_),
    .Y(_0166_),
    .B1(_2529_));
 sg13g2_nand2_1 _5876_ (.Y(_2530_),
    .A(net817),
    .B(net797));
 sg13g2_nand2b_1 _5877_ (.Y(_2531_),
    .B(net804),
    .A_N(net837));
 sg13g2_o21ai_1 _5878_ (.B1(_2531_),
    .Y(_2532_),
    .A1(net856),
    .A2(net803));
 sg13g2_o21ai_1 _5879_ (.B1(_2530_),
    .Y(_2533_),
    .A1(net794),
    .A2(_2532_));
 sg13g2_nor2_1 _5880_ (.A(net859),
    .B(net804),
    .Y(_2534_));
 sg13g2_nor2_1 _5881_ (.A(net840),
    .B(net807),
    .Y(_2535_));
 sg13g2_nor3_1 _5882_ (.A(net794),
    .B(_2534_),
    .C(_2535_),
    .Y(_2536_));
 sg13g2_a21oi_1 _5883_ (.A1(net270),
    .A2(net797),
    .Y(_2537_),
    .B1(_2536_));
 sg13g2_nand2_1 _5884_ (.Y(_2538_),
    .A(net376),
    .B(net798));
 sg13g2_a21oi_1 _5885_ (.A1(_2635_),
    .A2(net805),
    .Y(_2539_),
    .B1(net795));
 sg13g2_o21ai_1 _5886_ (.B1(_2539_),
    .Y(_2540_),
    .A1(net869),
    .A2(net805));
 sg13g2_nand2_1 _5887_ (.Y(_2541_),
    .A(_2538_),
    .B(_2540_));
 sg13g2_nand2b_1 _5888_ (.Y(_2542_),
    .B(net847),
    .A_N(net795));
 sg13g2_o21ai_1 _5889_ (.B1(net806),
    .Y(_2543_),
    .A1(\DP_4.matrix[73] ),
    .A2(_2476_));
 sg13g2_nor2_1 _5890_ (.A(net863),
    .B(_2495_),
    .Y(_2544_));
 sg13g2_a21oi_1 _5891_ (.A1(_2542_),
    .A2(_2543_),
    .Y(_2545_),
    .B1(_2544_));
 sg13g2_and2_1 _5892_ (.A(_2541_),
    .B(_2545_),
    .X(_2546_));
 sg13g2_nor2_1 _5893_ (.A(net861),
    .B(net805),
    .Y(_2547_));
 sg13g2_nor2_1 _5894_ (.A(net842),
    .B(net806),
    .Y(_2548_));
 sg13g2_nor3_1 _5895_ (.A(net795),
    .B(_2547_),
    .C(_2548_),
    .Y(_2549_));
 sg13g2_a21oi_1 _5896_ (.A1(net370),
    .A2(net798),
    .Y(_2550_),
    .B1(_2549_));
 sg13g2_nor2b_1 _5897_ (.A(_2550_),
    .B_N(_2546_),
    .Y(_2551_));
 sg13g2_nand2b_1 _5898_ (.Y(_2552_),
    .B(_2551_),
    .A_N(_2537_));
 sg13g2_nand2_1 _5899_ (.Y(_2553_),
    .A(net269),
    .B(net797));
 sg13g2_nand2b_1 _5900_ (.Y(_2554_),
    .B(net803),
    .A_N(net838));
 sg13g2_o21ai_1 _5901_ (.B1(_2554_),
    .Y(_2555_),
    .A1(net857),
    .A2(net804));
 sg13g2_o21ai_1 _5902_ (.B1(_2553_),
    .Y(_2556_),
    .A1(net794),
    .A2(_2555_));
 sg13g2_nand2b_1 _5903_ (.Y(_2557_),
    .B(_2556_),
    .A_N(_2552_));
 sg13g2_nand2b_1 _5904_ (.Y(_2558_),
    .B(_2533_),
    .A_N(_2557_));
 sg13g2_nand2_1 _5905_ (.Y(_2559_),
    .A(\DP_4.matrix[78] ),
    .B(net797));
 sg13g2_nand2b_1 _5906_ (.Y(_2560_),
    .B(net803),
    .A_N(net835));
 sg13g2_o21ai_1 _5907_ (.B1(_2560_),
    .Y(_2561_),
    .A1(net855),
    .A2(net804));
 sg13g2_o21ai_1 _5908_ (.B1(_2559_),
    .Y(_2562_),
    .A1(net794),
    .A2(_2561_));
 sg13g2_nor2b_1 _5909_ (.A(_2558_),
    .B_N(_2562_),
    .Y(_2563_));
 sg13g2_nor2_1 _5910_ (.A(net853),
    .B(net803),
    .Y(_2564_));
 sg13g2_nor2_1 _5911_ (.A(net833),
    .B(net807),
    .Y(_2565_));
 sg13g2_nor3_1 _5912_ (.A(net796),
    .B(_2564_),
    .C(_2565_),
    .Y(_2566_));
 sg13g2_a21oi_1 _5913_ (.A1(net813),
    .A2(net798),
    .Y(_2567_),
    .B1(_2566_));
 sg13g2_inv_1 _5914_ (.Y(_2568_),
    .A(_2567_));
 sg13g2_nor2_1 _5915_ (.A(net1044),
    .B(net803),
    .Y(_2569_));
 sg13g2_nor2_1 _5916_ (.A(net1043),
    .B(net806),
    .Y(_2570_));
 sg13g2_nor3_1 _5917_ (.A(net796),
    .B(_2569_),
    .C(_2570_),
    .Y(_2571_));
 sg13g2_a21oi_1 _5918_ (.A1(net278),
    .A2(net798),
    .Y(_2572_),
    .B1(_2571_));
 sg13g2_a21oi_1 _5919_ (.A1(_2563_),
    .A2(_2568_),
    .Y(_2573_),
    .B1(net791));
 sg13g2_nand2_1 _5920_ (.Y(_2574_),
    .A(net1044),
    .B(net791));
 sg13g2_o21ai_1 _5921_ (.B1(_2574_),
    .Y(_2575_),
    .A1(net791),
    .A2(_2571_));
 sg13g2_nor2_1 _5922_ (.A(_2573_),
    .B(_2575_),
    .Y(_2576_));
 sg13g2_a21oi_1 _5923_ (.A1(_2572_),
    .A2(_2573_),
    .Y(_0169_),
    .B1(_2576_));
 sg13g2_xor2_1 _5924_ (.B(net786),
    .A(net1040),
    .X(_0172_));
 sg13g2_nor2_1 _5925_ (.A(net1038),
    .B(net785),
    .Y(_2577_));
 sg13g2_xnor2_1 _5926_ (.Y(_2578_),
    .A(_2416_),
    .B(_2420_));
 sg13g2_a21oi_1 _5927_ (.A1(net785),
    .A2(_2578_),
    .Y(_0173_),
    .B1(_2577_));
 sg13g2_nor2_1 _5928_ (.A(net1036),
    .B(net785),
    .Y(_2579_));
 sg13g2_xor2_1 _5929_ (.B(_2423_),
    .A(_2421_),
    .X(_2580_));
 sg13g2_a21oi_1 _5930_ (.A1(net785),
    .A2(_2580_),
    .Y(_0174_),
    .B1(_2579_));
 sg13g2_nor2_1 _5931_ (.A(net1034),
    .B(net784),
    .Y(_2581_));
 sg13g2_xnor2_1 _5932_ (.Y(_2582_),
    .A(_2412_),
    .B(_2424_));
 sg13g2_a21oi_1 _5933_ (.A1(net784),
    .A2(_2582_),
    .Y(_0175_),
    .B1(_2581_));
 sg13g2_nor2_1 _5934_ (.A(net1033),
    .B(net786),
    .Y(_2583_));
 sg13g2_xnor2_1 _5935_ (.Y(_2584_),
    .A(_2425_),
    .B(_2427_));
 sg13g2_a21oi_1 _5936_ (.A1(net786),
    .A2(_2584_),
    .Y(_0176_),
    .B1(_2583_));
 sg13g2_nor2_1 _5937_ (.A(net282),
    .B(net786),
    .Y(_2585_));
 sg13g2_xnor2_1 _5938_ (.Y(_2586_),
    .A(_2408_),
    .B(_2428_));
 sg13g2_a21oi_1 _5939_ (.A1(net787),
    .A2(_2586_),
    .Y(_0177_),
    .B1(_2585_));
 sg13g2_nor2_1 _5940_ (.A(net1029),
    .B(net787),
    .Y(_2587_));
 sg13g2_xnor2_1 _5941_ (.Y(_2588_),
    .A(_2429_),
    .B(_2431_));
 sg13g2_a21oi_1 _5942_ (.A1(net787),
    .A2(_2588_),
    .Y(_0178_),
    .B1(_2587_));
 sg13g2_nand2b_1 _5943_ (.Y(_2589_),
    .B(net280),
    .A_N(net787));
 sg13g2_nor2b_1 _5944_ (.A(_2432_),
    .B_N(_2435_),
    .Y(_2590_));
 sg13g2_o21ai_1 _5945_ (.B1(_2589_),
    .Y(_0179_),
    .A1(_2436_),
    .A2(_2590_));
 sg13g2_xor2_1 _5946_ (.B(net785),
    .A(net982),
    .X(_0196_));
 sg13g2_nor2_1 _5947_ (.A(net978),
    .B(net785),
    .Y(_2591_));
 sg13g2_xnor2_1 _5948_ (.Y(_2592_),
    .A(_2452_),
    .B(_2455_));
 sg13g2_a21oi_1 _5949_ (.A1(net785),
    .A2(_2592_),
    .Y(_0197_),
    .B1(_2591_));
 sg13g2_nor2_1 _5950_ (.A(net976),
    .B(net786),
    .Y(_2593_));
 sg13g2_xor2_1 _5951_ (.B(_2458_),
    .A(_2456_),
    .X(_2594_));
 sg13g2_a21oi_1 _5952_ (.A1(net786),
    .A2(_2594_),
    .Y(_0198_),
    .B1(_2593_));
 sg13g2_nor2_1 _5953_ (.A(net974),
    .B(net783),
    .Y(_2595_));
 sg13g2_xnor2_1 _5954_ (.Y(_2596_),
    .A(_2448_),
    .B(_2459_));
 sg13g2_a21oi_1 _5955_ (.A1(net783),
    .A2(_2596_),
    .Y(_0199_),
    .B1(_2595_));
 sg13g2_nor2_1 _5956_ (.A(net972),
    .B(net783),
    .Y(_2597_));
 sg13g2_xnor2_1 _5957_ (.Y(_2598_),
    .A(_2460_),
    .B(_2462_));
 sg13g2_a21oi_1 _5958_ (.A1(net783),
    .A2(_2598_),
    .Y(_0200_),
    .B1(_2597_));
 sg13g2_nor2_1 _5959_ (.A(net971),
    .B(net783),
    .Y(_2599_));
 sg13g2_xnor2_1 _5960_ (.Y(_2600_),
    .A(_2444_),
    .B(_2463_));
 sg13g2_a21oi_1 _5961_ (.A1(net783),
    .A2(_2600_),
    .Y(_0201_),
    .B1(_2599_));
 sg13g2_nor2_1 _5962_ (.A(net969),
    .B(net783),
    .Y(_2601_));
 sg13g2_xnor2_1 _5963_ (.Y(_2602_),
    .A(_2464_),
    .B(_2466_));
 sg13g2_a21oi_1 _5964_ (.A1(net783),
    .A2(_2602_),
    .Y(_0202_),
    .B1(_2601_));
 sg13g2_nand2b_1 _5965_ (.Y(_2603_),
    .B(net968),
    .A_N(net784));
 sg13g2_nor2b_1 _5966_ (.A(_2467_),
    .B_N(_2470_),
    .Y(_2604_));
 sg13g2_o21ai_1 _5967_ (.B1(_2603_),
    .Y(_0203_),
    .A1(_2471_),
    .A2(_2604_));
 sg13g2_xnor2_1 _5968_ (.Y(_0220_),
    .A(net924),
    .B(net792));
 sg13g2_xnor2_1 _5969_ (.Y(_2605_),
    .A(_2493_),
    .B(_2498_));
 sg13g2_nand2_1 _5970_ (.Y(_2606_),
    .A(net923),
    .B(net789));
 sg13g2_o21ai_1 _5971_ (.B1(_2606_),
    .Y(_0221_),
    .A1(net789),
    .A2(_2605_));
 sg13g2_xor2_1 _5972_ (.B(_2503_),
    .A(_2499_),
    .X(_2607_));
 sg13g2_nand2_1 _5973_ (.Y(_2608_),
    .A(net920),
    .B(net789));
 sg13g2_o21ai_1 _5974_ (.B1(_2608_),
    .Y(_0222_),
    .A1(net789),
    .A2(_2607_));
 sg13g2_xnor2_1 _5975_ (.Y(_2609_),
    .A(_2489_),
    .B(_2504_));
 sg13g2_nand2_1 _5976_ (.Y(_2610_),
    .A(net918),
    .B(net790));
 sg13g2_o21ai_1 _5977_ (.B1(_2610_),
    .Y(_0223_),
    .A1(net790),
    .A2(_2609_));
 sg13g2_nand2_1 _5978_ (.Y(_2611_),
    .A(net916),
    .B(net793));
 sg13g2_xnor2_1 _5979_ (.Y(_2612_),
    .A(_2505_),
    .B(_2509_));
 sg13g2_o21ai_1 _5980_ (.B1(_2611_),
    .Y(_0224_),
    .A1(net793),
    .A2(_2612_));
 sg13g2_nand2b_1 _5981_ (.Y(_2613_),
    .B(_2511_),
    .A_N(net793));
 sg13g2_a21oi_1 _5982_ (.A1(_2485_),
    .A2(_2510_),
    .Y(_2614_),
    .B1(_2613_));
 sg13g2_a21o_1 _5983_ (.A2(net793),
    .A1(net915),
    .B1(_2614_),
    .X(_0225_));
 sg13g2_nand2_1 _5984_ (.Y(_2615_),
    .A(net913),
    .B(net792));
 sg13g2_xor2_1 _5985_ (.B(_2515_),
    .A(_2511_),
    .X(_2616_));
 sg13g2_o21ai_1 _5986_ (.B1(_2615_),
    .Y(_0226_),
    .A1(net792),
    .A2(_2616_));
 sg13g2_nand2b_1 _5987_ (.Y(_2617_),
    .B(_2520_),
    .A_N(_2516_));
 sg13g2_a22oi_1 _5988_ (.Y(_2618_),
    .B1(_2522_),
    .B2(_2617_),
    .A2(net792),
    .A1(net910));
 sg13g2_inv_1 _5989_ (.Y(_0227_),
    .A(_2618_));
 sg13g2_xnor2_1 _5990_ (.Y(_0244_),
    .A(net868),
    .B(net793));
 sg13g2_xnor2_1 _5991_ (.Y(_2619_),
    .A(_2541_),
    .B(_2545_));
 sg13g2_nand2_1 _5992_ (.Y(_2620_),
    .A(net863),
    .B(net789));
 sg13g2_o21ai_1 _5993_ (.B1(_2620_),
    .Y(_0245_),
    .A1(net789),
    .A2(_2619_));
 sg13g2_xor2_1 _5994_ (.B(_2550_),
    .A(_2546_),
    .X(_2621_));
 sg13g2_nand2_1 _5995_ (.Y(_2622_),
    .A(net861),
    .B(net789));
 sg13g2_o21ai_1 _5996_ (.B1(_2622_),
    .Y(_0246_),
    .A1(net789),
    .A2(_2621_));
 sg13g2_xor2_1 _5997_ (.B(_2551_),
    .A(_2537_),
    .X(_2623_));
 sg13g2_nand2_1 _5998_ (.Y(_2624_),
    .A(net859),
    .B(net790));
 sg13g2_o21ai_1 _5999_ (.B1(_2624_),
    .Y(_0247_),
    .A1(net790),
    .A2(_2623_));
 sg13g2_nand2_1 _6000_ (.Y(_2625_),
    .A(net857),
    .B(net793));
 sg13g2_xor2_1 _6001_ (.B(_2556_),
    .A(_2552_),
    .X(_2626_));
 sg13g2_o21ai_1 _6002_ (.B1(_2625_),
    .Y(_0248_),
    .A1(net793),
    .A2(_2626_));
 sg13g2_nand2_1 _6003_ (.Y(_2627_),
    .A(net856),
    .B(net792));
 sg13g2_xor2_1 _6004_ (.B(_2557_),
    .A(_2533_),
    .X(_2628_));
 sg13g2_o21ai_1 _6005_ (.B1(_2627_),
    .Y(_0249_),
    .A1(net792),
    .A2(_2628_));
 sg13g2_nand2_1 _6006_ (.Y(_2629_),
    .A(net855),
    .B(net791));
 sg13g2_xor2_1 _6007_ (.B(_2562_),
    .A(_2558_),
    .X(_2630_));
 sg13g2_o21ai_1 _6008_ (.B1(_2629_),
    .Y(_0250_),
    .A1(net791),
    .A2(_2630_));
 sg13g2_nand2b_1 _6009_ (.Y(_2631_),
    .B(_2567_),
    .A_N(_2563_));
 sg13g2_a22oi_1 _6010_ (.Y(_2632_),
    .B1(_2573_),
    .B2(_2631_),
    .A2(net791),
    .A1(net853));
 sg13g2_inv_1 _6011_ (.Y(_0251_),
    .A(_2632_));
 sg13g2_buf_1 _6012_ (.A(net1056),
    .X(_0161_));
 sg13g2_buf_1 _6013_ (.A(net1054),
    .X(_0162_));
 sg13g2_buf_1 _6014_ (.A(net274),
    .X(_0164_));
 sg13g2_buf_1 _6015_ (.A(net1051),
    .X(_0165_));
 sg13g2_buf_1 _6016_ (.A(net1047),
    .X(_0167_));
 sg13g2_buf_1 _6017_ (.A(net273),
    .X(_0168_));
 sg13g2_buf_1 _6018_ (.A(net1043),
    .X(_0170_));
 sg13g2_buf_1 _6019_ (.A(net278),
    .X(_0171_));
 sg13g2_buf_1 _6020_ (.A(net1023),
    .X(_0180_));
 sg13g2_buf_1 _6021_ (.A(net1021),
    .X(_0181_));
 sg13g2_buf_1 _6022_ (.A(net1018),
    .X(_0182_));
 sg13g2_buf_1 _6023_ (.A(net1017),
    .X(_0183_));
 sg13g2_buf_1 _6024_ (.A(net1015),
    .X(_0184_));
 sg13g2_buf_1 _6025_ (.A(net1012),
    .X(_0185_));
 sg13g2_buf_1 _6026_ (.A(net1008),
    .X(_0186_));
 sg13g2_buf_1 _6027_ (.A(net1007),
    .X(_0187_));
 sg13g2_buf_1 _6028_ (.A(net1004),
    .X(_0188_));
 sg13g2_buf_1 _6029_ (.A(net1001),
    .X(_0189_));
 sg13g2_buf_1 _6030_ (.A(net998),
    .X(_0190_));
 sg13g2_buf_1 _6031_ (.A(net997),
    .X(_0191_));
 sg13g2_buf_1 _6032_ (.A(net994),
    .X(_0192_));
 sg13g2_buf_1 _6033_ (.A(net991),
    .X(_0193_));
 sg13g2_buf_1 _6034_ (.A(net989),
    .X(_0194_));
 sg13g2_buf_1 _6035_ (.A(net987),
    .X(_0195_));
 sg13g2_buf_1 _6036_ (.A(net964),
    .X(_0204_));
 sg13g2_buf_1 _6037_ (.A(net960),
    .X(_0205_));
 sg13g2_buf_1 _6038_ (.A(net957),
    .X(_0206_));
 sg13g2_buf_1 _6039_ (.A(net955),
    .X(_0207_));
 sg13g2_buf_1 _6040_ (.A(net953),
    .X(_0208_));
 sg13g2_buf_1 _6041_ (.A(net951),
    .X(_0209_));
 sg13g2_buf_1 _6042_ (.A(net950),
    .X(_0210_));
 sg13g2_buf_1 _6043_ (.A(net948),
    .X(_0211_));
 sg13g2_buf_1 _6044_ (.A(net943),
    .X(_0212_));
 sg13g2_buf_1 _6045_ (.A(net940),
    .X(_0213_));
 sg13g2_buf_1 _6046_ (.A(net936),
    .X(_0214_));
 sg13g2_buf_1 _6047_ (.A(net934),
    .X(_0215_));
 sg13g2_buf_1 _6048_ (.A(net933),
    .X(_0216_));
 sg13g2_buf_1 _6049_ (.A(net931),
    .X(_0217_));
 sg13g2_buf_1 _6050_ (.A(net929),
    .X(_0218_));
 sg13g2_buf_1 _6051_ (.A(net926),
    .X(_0219_));
 sg13g2_buf_1 _6052_ (.A(net906),
    .X(_0228_));
 sg13g2_buf_1 _6053_ (.A(net905),
    .X(_0229_));
 sg13g2_buf_1 _6054_ (.A(net902),
    .X(_0230_));
 sg13g2_buf_1 _6055_ (.A(net900),
    .X(_0231_));
 sg13g2_buf_1 _6056_ (.A(net899),
    .X(_0232_));
 sg13g2_buf_1 _6057_ (.A(net897),
    .X(_0233_));
 sg13g2_buf_1 _6058_ (.A(net894),
    .X(_0234_));
 sg13g2_buf_1 _6059_ (.A(net892),
    .X(_0235_));
 sg13g2_buf_1 _6060_ (.A(net275),
    .X(_0236_));
 sg13g2_buf_1 _6061_ (.A(net888),
    .X(_0237_));
 sg13g2_buf_1 _6062_ (.A(net885),
    .X(_0238_));
 sg13g2_buf_1 _6063_ (.A(net882),
    .X(_0239_));
 sg13g2_buf_1 _6064_ (.A(net879),
    .X(_0240_));
 sg13g2_buf_1 _6065_ (.A(net277),
    .X(_0241_));
 sg13g2_buf_1 _6066_ (.A(net279),
    .X(_0242_));
 sg13g2_buf_1 _6067_ (.A(net276),
    .X(_0243_));
 sg13g2_buf_1 _6068_ (.A(net850),
    .X(_0252_));
 sg13g2_buf_1 _6069_ (.A(net847),
    .X(_0253_));
 sg13g2_buf_1 _6070_ (.A(net842),
    .X(_0254_));
 sg13g2_buf_1 _6071_ (.A(net841),
    .X(_0255_));
 sg13g2_buf_1 _6072_ (.A(net838),
    .X(_0256_));
 sg13g2_buf_1 _6073_ (.A(net837),
    .X(_0257_));
 sg13g2_buf_1 _6074_ (.A(net835),
    .X(_0258_));
 sg13g2_buf_1 _6075_ (.A(net833),
    .X(_0259_));
 sg13g2_buf_1 _6076_ (.A(net832),
    .X(_0260_));
 sg13g2_buf_1 _6077_ (.A(net826),
    .X(_0261_));
 sg13g2_buf_1 _6078_ (.A(net823),
    .X(_0262_));
 sg13g2_buf_1 _6079_ (.A(net270),
    .X(_0263_));
 sg13g2_buf_1 _6080_ (.A(net269),
    .X(_0264_));
 sg13g2_buf_1 _6081_ (.A(net817),
    .X(_0265_));
 sg13g2_buf_1 _6082_ (.A(net815),
    .X(_0266_));
 sg13g2_buf_1 _6083_ (.A(net813),
    .X(_0267_));
 sg13g2_dfrbpq_2 _6084_ (.RESET_B(net1080),
    .D(net9),
    .Q(\DP_3.Q_range.out_data[2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6085_ (.RESET_B(net1080),
    .D(net10),
    .Q(\DP_3.Q_range.out_data[3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6086_ (.RESET_B(net1080),
    .D(net11),
    .Q(\DP_3.Q_range.out_data[4] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6087_ (.RESET_B(net1080),
    .D(\DP_3.Q_range.data_plus_4[6] ),
    .Q(\DP_3.Q_range.out_data[5] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6088_ (.RESET_B(net1063),
    .D(_0069_),
    .Q(\mac1.products_ff[0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6089_ (.RESET_B(net1063),
    .D(_0070_),
    .Q(\mac1.products_ff[1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6090_ (.RESET_B(net1070),
    .D(_0071_),
    .Q(\mac1.products_ff[2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6091_ (.RESET_B(net1071),
    .D(_0072_),
    .Q(\mac1.products_ff[3] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6092_ (.RESET_B(net1092),
    .D(_0073_),
    .Q(\mac1.products_ff[4] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6093_ (.RESET_B(net1109),
    .D(_0105_),
    .Q(\mac1.products_ff[5] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6094_ (.RESET_B(net1109),
    .D(_0112_),
    .Q(\mac1.products_ff[6] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6095_ (.RESET_B(net1115),
    .D(_0113_),
    .Q(\mac1.products_ff[7] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6096_ (.RESET_B(net1114),
    .D(_0114_),
    .Q(\mac1.products_ff[8] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6097_ (.RESET_B(net1115),
    .D(_0115_),
    .Q(\mac1.products_ff[9] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6098_ (.RESET_B(net1121),
    .D(_0106_),
    .Q(\mac1.products_ff[10] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6099_ (.RESET_B(net1121),
    .D(_0107_),
    .Q(\mac1.products_ff[11] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6100_ (.RESET_B(net1098),
    .D(_0108_),
    .Q(\mac1.products_ff[12] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6101_ (.RESET_B(net1098),
    .D(_0109_),
    .Q(\mac1.products_ff[13] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6102_ (.RESET_B(net1097),
    .D(_0110_),
    .Q(\mac1.products_ff[14] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6103_ (.RESET_B(net1084),
    .D(_0111_),
    .Q(\mac1.products_ff[15] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6104_ (.RESET_B(net1070),
    .D(_0074_),
    .Q(\mac1.products_ff[68] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6105_ (.RESET_B(net1063),
    .D(_0075_),
    .Q(\mac1.products_ff[69] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6106_ (.RESET_B(net1069),
    .D(_0076_),
    .Q(\mac1.products_ff[70] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _6107_ (.RESET_B(net1088),
    .D(_0077_),
    .Q(\mac1.products_ff[71] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6108_ (.RESET_B(net1090),
    .D(_0078_),
    .Q(\mac1.products_ff[72] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6109_ (.RESET_B(net1090),
    .D(_0116_),
    .Q(\mac1.products_ff[73] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6110_ (.RESET_B(net1090),
    .D(_0123_),
    .Q(\mac1.products_ff[74] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6111_ (.RESET_B(net1090),
    .D(_0124_),
    .Q(\mac1.products_ff[75] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6112_ (.RESET_B(net1092),
    .D(_0125_),
    .Q(\mac1.products_ff[76] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6113_ (.RESET_B(net1092),
    .D(_0126_),
    .Q(\mac1.products_ff[77] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6114_ (.RESET_B(net1089),
    .D(_0117_),
    .Q(\mac1.products_ff[78] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6115_ (.RESET_B(net1098),
    .D(_0118_),
    .Q(\mac1.products_ff[79] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6116_ (.RESET_B(net1089),
    .D(_0119_),
    .Q(\mac1.products_ff[80] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6117_ (.RESET_B(net1096),
    .D(_0120_),
    .Q(\mac1.products_ff[81] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6118_ (.RESET_B(net1083),
    .D(_0121_),
    .Q(\mac1.products_ff[82] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6119_ (.RESET_B(net1083),
    .D(_0122_),
    .Q(\mac1.products_ff[83] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6120_ (.RESET_B(net1095),
    .D(_0160_),
    .Q(\DP_1.matrix[8] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _6121_ (.RESET_B(net1073),
    .D(_0161_),
    .Q(\DP_1.matrix[44] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _6122_ (.RESET_B(net1135),
    .D(_0162_),
    .Q(\DP_1.matrix[80] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _6123_ (.RESET_B(net1094),
    .D(_0163_),
    .Q(\DP_2.matrix[8] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _6124_ (.RESET_B(net1089),
    .D(_0164_),
    .Q(\DP_2.matrix[44] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _6125_ (.RESET_B(net1118),
    .D(_0165_),
    .Q(\DP_2.matrix[80] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6126_ (.RESET_B(net1127),
    .D(_0166_),
    .Q(\DP_3.matrix[8] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6127_ (.RESET_B(net1127),
    .D(_0167_),
    .Q(\DP_3.matrix[44] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6128_ (.RESET_B(net1106),
    .D(_0168_),
    .Q(\DP_3.matrix[80] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6129_ (.RESET_B(net1127),
    .D(_0169_),
    .Q(\DP_4.matrix[8] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6130_ (.RESET_B(net1129),
    .D(_0170_),
    .Q(\DP_4.matrix[44] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _6131_ (.RESET_B(net1124),
    .D(_0171_),
    .Q(\DP_4.matrix[80] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6132_ (.RESET_B(net1062),
    .D(_0064_),
    .Q(\mac1.products_ff[136] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6133_ (.RESET_B(net1093),
    .D(_0172_),
    .Q(\DP_1.matrix[0] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _6134_ (.RESET_B(net1091),
    .D(_0173_),
    .Q(\DP_1.matrix[1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6135_ (.RESET_B(net1062),
    .D(_0065_),
    .Q(\mac1.products_ff[137] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _6136_ (.RESET_B(net1091),
    .D(_0174_),
    .Q(\DP_1.matrix[2] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _6137_ (.RESET_B(net1094),
    .D(_0175_),
    .Q(\DP_1.matrix[3] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6138_ (.RESET_B(net1062),
    .D(_0066_),
    .Q(\mac1.products_ff[138] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _6139_ (.RESET_B(net1094),
    .D(net397),
    .Q(\DP_1.matrix[4] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _6140_ (.RESET_B(net1094),
    .D(net283),
    .Q(\DP_1.matrix[5] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6141_ (.RESET_B(net1071),
    .D(_0067_),
    .Q(\mac1.products_ff[139] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6142_ (.RESET_B(net1095),
    .D(net409),
    .Q(\DP_1.matrix[6] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6143_ (.RESET_B(net1095),
    .D(net281),
    .Q(\DP_1.matrix[7] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6144_ (.RESET_B(net1116),
    .D(_0068_),
    .Q(\mac1.products_ff[140] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6145_ (.RESET_B(net1072),
    .D(_0180_),
    .Q(\DP_1.matrix[36] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6146_ (.RESET_B(net1071),
    .D(_0181_),
    .Q(\DP_1.matrix[37] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6147_ (.RESET_B(net1116),
    .D(_0094_),
    .Q(\mac1.products_ff[141] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6148_ (.RESET_B(net1088),
    .D(_0182_),
    .Q(\DP_1.matrix[38] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6149_ (.RESET_B(net1088),
    .D(_0183_),
    .Q(\DP_1.matrix[39] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6150_ (.RESET_B(net1116),
    .D(_0101_),
    .Q(\mac1.products_ff[142] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6151_ (.RESET_B(net1090),
    .D(_0184_),
    .Q(\DP_1.matrix[40] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6152_ (.RESET_B(net1090),
    .D(_0185_),
    .Q(\DP_1.matrix[41] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6153_ (.RESET_B(net1131),
    .D(_0102_),
    .Q(\mac1.products_ff[143] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _6154_ (.RESET_B(net1072),
    .D(_0186_),
    .Q(\DP_1.matrix[42] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _6155_ (.RESET_B(net1070),
    .D(_0187_),
    .Q(\DP_1.matrix[43] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6156_ (.RESET_B(net1111),
    .D(_0103_),
    .Q(\mac1.products_ff[144] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6157_ (.RESET_B(net1112),
    .D(_0188_),
    .Q(\DP_1.matrix[72] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6158_ (.RESET_B(net1116),
    .D(_0189_),
    .Q(\DP_1.matrix[73] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6159_ (.RESET_B(net1132),
    .D(_0104_),
    .Q(\mac1.products_ff[145] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6160_ (.RESET_B(net1112),
    .D(_0190_),
    .Q(\DP_1.matrix[74] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6161_ (.RESET_B(net1112),
    .D(_0191_),
    .Q(\DP_1.matrix[75] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6162_ (.RESET_B(net1133),
    .D(_0095_),
    .Q(\mac1.products_ff[146] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _6163_ (.RESET_B(net1117),
    .D(_0192_),
    .Q(\DP_1.matrix[76] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _6164_ (.RESET_B(net1117),
    .D(_0193_),
    .Q(\DP_1.matrix[77] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6165_ (.RESET_B(net1133),
    .D(_0096_),
    .Q(\mac1.products_ff[147] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _6166_ (.RESET_B(net1132),
    .D(_0194_),
    .Q(\DP_1.matrix[78] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _6167_ (.RESET_B(net1135),
    .D(_0195_),
    .Q(\DP_1.matrix[79] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _6168_ (.RESET_B(net1119),
    .D(_0097_),
    .Q(\mac1.products_ff[148] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _6169_ (.RESET_B(net1091),
    .D(_0196_),
    .Q(\DP_2.matrix[0] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6170_ (.RESET_B(net1091),
    .D(_0197_),
    .Q(\DP_2.matrix[1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6171_ (.RESET_B(net1067),
    .D(_0098_),
    .Q(\mac1.products_ff[149] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6172_ (.RESET_B(net1093),
    .D(_0198_),
    .Q(\DP_2.matrix[2] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6173_ (.RESET_B(net1094),
    .D(net407),
    .Q(\DP_2.matrix[3] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6174_ (.RESET_B(net1067),
    .D(_0099_),
    .Q(\mac1.products_ff[150] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6175_ (.RESET_B(net1094),
    .D(_0200_),
    .Q(\DP_2.matrix[4] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _6176_ (.RESET_B(net1089),
    .D(_0201_),
    .Q(\DP_2.matrix[5] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _6177_ (.RESET_B(net1118),
    .D(_0100_),
    .Q(\mac1.products_ff[151] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6178_ (.RESET_B(net1094),
    .D(net417),
    .Q(\DP_2.matrix[6] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6179_ (.RESET_B(net1094),
    .D(net378),
    .Q(\DP_2.matrix[7] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6180_ (.RESET_B(net1063),
    .D(net107),
    .Q(\mac1.sum_lvl1_ff[0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6181_ (.RESET_B(net1071),
    .D(_0204_),
    .Q(\DP_2.matrix[36] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6182_ (.RESET_B(net1072),
    .D(_0205_),
    .Q(\DP_2.matrix[37] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6183_ (.RESET_B(net1063),
    .D(net219),
    .Q(\mac1.sum_lvl1_ff[1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6184_ (.RESET_B(net1090),
    .D(_0206_),
    .Q(\DP_2.matrix[38] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6185_ (.RESET_B(net1090),
    .D(_0207_),
    .Q(\DP_2.matrix[39] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6186_ (.RESET_B(net1070),
    .D(net103),
    .Q(\mac1.sum_lvl1_ff[2] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6187_ (.RESET_B(net1088),
    .D(_0208_),
    .Q(\DP_2.matrix[40] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _6188_ (.RESET_B(net1070),
    .D(_0209_),
    .Q(\DP_2.matrix[41] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6189_ (.RESET_B(net1088),
    .D(net96),
    .Q(\mac1.sum_lvl1_ff[3] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6190_ (.RESET_B(net1091),
    .D(_0210_),
    .Q(\DP_2.matrix[42] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6191_ (.RESET_B(net1091),
    .D(_0211_),
    .Q(\DP_2.matrix[43] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6192_ (.RESET_B(net1109),
    .D(net183),
    .Q(\mac1.sum_lvl1_ff[4] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6193_ (.RESET_B(net1131),
    .D(_0212_),
    .Q(\DP_2.matrix[72] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6194_ (.RESET_B(net1131),
    .D(_0213_),
    .Q(\DP_2.matrix[73] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6195_ (.RESET_B(net1109),
    .D(net86),
    .Q(\mac1.sum_lvl1_ff[5] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6196_ (.RESET_B(net1131),
    .D(_0214_),
    .Q(\DP_2.matrix[74] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _6197_ (.RESET_B(net1117),
    .D(_0215_),
    .Q(\DP_2.matrix[75] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6198_ (.RESET_B(net1110),
    .D(net149),
    .Q(\mac1.sum_lvl1_ff[6] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _6199_ (.RESET_B(net1112),
    .D(_0216_),
    .Q(\DP_2.matrix[76] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6200_ (.RESET_B(net1114),
    .D(_0217_),
    .Q(\DP_2.matrix[77] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6201_ (.RESET_B(net1115),
    .D(net81),
    .Q(\mac1.sum_lvl1_ff[7] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _6202_ (.RESET_B(net1116),
    .D(_0218_),
    .Q(\DP_2.matrix[78] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _6203_ (.RESET_B(net1116),
    .D(_0219_),
    .Q(\DP_2.matrix[79] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6204_ (.RESET_B(net1114),
    .D(net77),
    .Q(\mac1.sum_lvl1_ff[8] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6205_ (.RESET_B(net1127),
    .D(_0220_),
    .Q(\DP_3.matrix[0] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6206_ (.RESET_B(net1105),
    .D(net423),
    .Q(\DP_3.matrix[1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6207_ (.RESET_B(net1114),
    .D(net74),
    .Q(\mac1.sum_lvl1_ff[9] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _6208_ (.RESET_B(net1122),
    .D(net436),
    .Q(\DP_3.matrix[2] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6209_ (.RESET_B(net1122),
    .D(net388),
    .Q(\DP_3.matrix[3] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6210_ (.RESET_B(net1120),
    .D(net246),
    .Q(\mac1.sum_lvl1_ff[10] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _6211_ (.RESET_B(net1124),
    .D(net421),
    .Q(\DP_3.matrix[4] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6212_ (.RESET_B(net1128),
    .D(_0225_),
    .Q(\DP_3.matrix[5] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6213_ (.RESET_B(net1121),
    .D(net134),
    .Q(\mac1.sum_lvl1_ff[11] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6214_ (.RESET_B(net1126),
    .D(_0226_),
    .Q(\DP_3.matrix[6] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6215_ (.RESET_B(net1126),
    .D(_0227_),
    .Q(\DP_3.matrix[7] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6216_ (.RESET_B(net1098),
    .D(net71),
    .Q(\mac1.sum_lvl1_ff[12] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6217_ (.RESET_B(net1121),
    .D(_0228_),
    .Q(\DP_3.matrix[36] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _6218_ (.RESET_B(net1122),
    .D(_0229_),
    .Q(\DP_3.matrix[37] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6219_ (.RESET_B(net1098),
    .D(net151),
    .Q(\mac1.sum_lvl1_ff[13] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6220_ (.RESET_B(net1126),
    .D(_0230_),
    .Q(\DP_3.matrix[38] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6221_ (.RESET_B(net1129),
    .D(_0231_),
    .Q(\DP_3.matrix[39] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6222_ (.RESET_B(net1097),
    .D(net200),
    .Q(\mac1.sum_lvl1_ff[14] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _6223_ (.RESET_B(net1139),
    .D(_0232_),
    .Q(\DP_3.matrix[40] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _6224_ (.RESET_B(net1146),
    .D(_0233_),
    .Q(\DP_3.matrix[41] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6225_ (.RESET_B(net1097),
    .D(net181),
    .Q(\mac1.sum_lvl1_ff[15] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _6226_ (.RESET_B(net1127),
    .D(_0234_),
    .Q(\DP_3.matrix[42] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6227_ (.RESET_B(net1129),
    .D(_0235_),
    .Q(\DP_3.matrix[43] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6228_ (.RESET_B(net1100),
    .D(_0236_),
    .Q(\DP_3.matrix[72] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6229_ (.RESET_B(net1104),
    .D(_0237_),
    .Q(\DP_3.matrix[73] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6230_ (.RESET_B(net1104),
    .D(_0238_),
    .Q(\DP_3.matrix[74] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6231_ (.RESET_B(net1104),
    .D(_0239_),
    .Q(\DP_3.matrix[75] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6232_ (.RESET_B(net1123),
    .D(_0240_),
    .Q(\DP_3.matrix[76] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6233_ (.RESET_B(net1124),
    .D(_0241_),
    .Q(\DP_3.matrix[77] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6234_ (.RESET_B(net1104),
    .D(_0242_),
    .Q(\DP_3.matrix[78] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6235_ (.RESET_B(net1123),
    .D(_0243_),
    .Q(\DP_3.matrix[79] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6236_ (.RESET_B(net1127),
    .D(net375),
    .Q(\DP_4.matrix[0] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6237_ (.RESET_B(net1105),
    .D(net508),
    .Q(\DP_4.matrix[1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6238_ (.RESET_B(net1122),
    .D(net380),
    .Q(\DP_4.matrix[2] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6239_ (.RESET_B(net1124),
    .D(net385),
    .Q(\DP_4.matrix[3] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6240_ (.RESET_B(net1126),
    .D(net372),
    .Q(\DP_4.matrix[4] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _6241_ (.RESET_B(net1126),
    .D(_0249_),
    .Q(\DP_4.matrix[5] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6242_ (.RESET_B(net1128),
    .D(net358),
    .Q(\DP_4.matrix[6] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6243_ (.RESET_B(net1126),
    .D(_0251_),
    .Q(\DP_4.matrix[7] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6244_ (.RESET_B(net1121),
    .D(_0252_),
    .Q(\DP_4.matrix[36] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6245_ (.RESET_B(net1105),
    .D(_0253_),
    .Q(\DP_4.matrix[37] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6246_ (.RESET_B(net1120),
    .D(_0254_),
    .Q(\DP_4.matrix[38] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6247_ (.RESET_B(net1129),
    .D(_0255_),
    .Q(\DP_4.matrix[39] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6248_ (.RESET_B(net1139),
    .D(_0256_),
    .Q(\DP_4.matrix[40] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _6249_ (.RESET_B(net1139),
    .D(_0257_),
    .Q(\DP_4.matrix[41] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6250_ (.RESET_B(net1139),
    .D(_0258_),
    .Q(\DP_4.matrix[42] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6251_ (.RESET_B(net1139),
    .D(_0259_),
    .Q(\DP_4.matrix[43] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6252_ (.RESET_B(net1085),
    .D(_0260_),
    .Q(\DP_4.matrix[72] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6253_ (.RESET_B(net1085),
    .D(_0261_),
    .Q(\DP_4.matrix[73] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6254_ (.RESET_B(net1101),
    .D(_0262_),
    .Q(\DP_4.matrix[74] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6255_ (.RESET_B(net1104),
    .D(_0263_),
    .Q(\DP_4.matrix[75] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6256_ (.RESET_B(net1123),
    .D(_0264_),
    .Q(\DP_4.matrix[76] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6257_ (.RESET_B(net1123),
    .D(_0265_),
    .Q(\DP_4.matrix[77] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6258_ (.RESET_B(net1100),
    .D(_0266_),
    .Q(\DP_4.matrix[78] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6259_ (.RESET_B(net1125),
    .D(_0267_),
    .Q(\DP_4.matrix[79] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6260_ (.RESET_B(net1064),
    .D(net239),
    .Q(\mac1.sum_lvl1_ff[36] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6261_ (.RESET_B(net1063),
    .D(net217),
    .Q(\mac1.sum_lvl1_ff[37] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6262_ (.RESET_B(net1069),
    .D(net54),
    .Q(\mac1.sum_lvl1_ff[38] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _6263_ (.RESET_B(net1088),
    .D(net120),
    .Q(\mac1.sum_lvl1_ff[39] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6264_ (.RESET_B(net1092),
    .D(net72),
    .Q(\mac1.sum_lvl1_ff[40] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6265_ (.RESET_B(net1092),
    .D(net237),
    .Q(\mac1.sum_lvl1_ff[41] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6266_ (.RESET_B(net1092),
    .D(net189),
    .Q(\mac1.sum_lvl1_ff[42] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6267_ (.RESET_B(net1092),
    .D(net146),
    .Q(\mac1.sum_lvl1_ff[43] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6268_ (.RESET_B(net1110),
    .D(net175),
    .Q(\mac1.sum_lvl1_ff[44] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6269_ (.RESET_B(net1115),
    .D(net241),
    .Q(\mac1.sum_lvl1_ff[45] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6270_ (.RESET_B(net1089),
    .D(net124),
    .Q(\mac1.sum_lvl1_ff[46] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6271_ (.RESET_B(net1098),
    .D(net63),
    .Q(\mac1.sum_lvl1_ff[47] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6272_ (.RESET_B(net1096),
    .D(net230),
    .Q(\mac1.sum_lvl1_ff[48] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6273_ (.RESET_B(net1097),
    .D(net253),
    .Q(\mac1.sum_lvl1_ff[49] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6274_ (.RESET_B(net1096),
    .D(net177),
    .Q(\mac1.sum_lvl1_ff[50] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6275_ (.RESET_B(net1096),
    .D(net98),
    .Q(\mac1.sum_lvl1_ff[51] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6276_ (.RESET_B(net1064),
    .D(net142),
    .Q(\mac1.sum_lvl2_ff[0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6277_ (.RESET_B(net1063),
    .D(net59),
    .Q(\mac1.sum_lvl2_ff[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6278_ (.RESET_B(net1069),
    .D(net234),
    .Q(\mac1.sum_lvl2_ff[2] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6279_ (.RESET_B(net1088),
    .D(net62),
    .Q(\mac1.sum_lvl2_ff[3] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6280_ (.RESET_B(net1109),
    .D(net88),
    .Q(\mac1.sum_lvl2_ff[4] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6281_ (.RESET_B(net1109),
    .D(net127),
    .Q(\mac1.sum_lvl2_ff[5] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6282_ (.RESET_B(net1111),
    .D(net73),
    .Q(\mac1.sum_lvl2_ff[6] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6283_ (.RESET_B(net1114),
    .D(net168),
    .Q(\mac1.sum_lvl2_ff[7] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6284_ (.RESET_B(net1114),
    .D(net156),
    .Q(\mac1.sum_lvl2_ff[8] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6285_ (.RESET_B(net1114),
    .D(net182),
    .Q(\mac1.sum_lvl2_ff[9] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6286_ (.RESET_B(net1120),
    .D(net46),
    .Q(\mac1.sum_lvl2_ff[10] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6287_ (.RESET_B(net1120),
    .D(net226),
    .Q(\mac1.sum_lvl2_ff[11] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6288_ (.RESET_B(net1098),
    .D(net204),
    .Q(\mac1.sum_lvl2_ff[12] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6289_ (.RESET_B(net1099),
    .D(net197),
    .Q(\mac1.sum_lvl2_ff[13] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6290_ (.RESET_B(net1097),
    .D(net58),
    .Q(\mac1.sum_lvl2_ff[14] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6291_ (.RESET_B(net1097),
    .D(net56),
    .Q(\mac1.sum_lvl2_ff[15] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6292_ (.RESET_B(net1064),
    .D(net212),
    .Q(\mac1.sum_lvl2_ff[19] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6293_ (.RESET_B(net1063),
    .D(net78),
    .Q(\mac1.sum_lvl2_ff[20] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6294_ (.RESET_B(net1069),
    .D(net68),
    .Q(\mac1.sum_lvl2_ff[21] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6295_ (.RESET_B(net1088),
    .D(net147),
    .Q(\mac1.sum_lvl2_ff[22] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6296_ (.RESET_B(net1109),
    .D(net255),
    .Q(\mac1.sum_lvl2_ff[23] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6297_ (.RESET_B(net1109),
    .D(net211),
    .Q(\mac1.sum_lvl2_ff[24] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6298_ (.RESET_B(net1092),
    .D(net52),
    .Q(\mac1.sum_lvl2_ff[25] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6299_ (.RESET_B(net1110),
    .D(net260),
    .Q(\mac1.sum_lvl2_ff[26] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6300_ (.RESET_B(net1110),
    .D(net139),
    .Q(\mac1.sum_lvl2_ff[27] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6301_ (.RESET_B(net1115),
    .D(net206),
    .Q(\mac1.sum_lvl2_ff[28] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6302_ (.RESET_B(net1120),
    .D(net262),
    .Q(\mac1.sum_lvl2_ff[29] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _6303_ (.RESET_B(net1107),
    .D(net42),
    .Q(\mac1.sum_lvl2_ff[30] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6304_ (.RESET_B(net1098),
    .D(net148),
    .Q(\mac1.sum_lvl2_ff[31] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6305_ (.RESET_B(net1097),
    .D(net99),
    .Q(\mac1.sum_lvl2_ff[32] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6306_ (.RESET_B(net1096),
    .D(net188),
    .Q(\mac1.sum_lvl2_ff[33] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6307_ (.RESET_B(net1096),
    .D(net208),
    .Q(\mac1.sum_lvl2_ff[34] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6308_ (.RESET_B(net1064),
    .D(net164),
    .Q(\mac1.sum_lvl2_ff[38] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6309_ (.RESET_B(net1062),
    .D(net215),
    .Q(\mac1.sum_lvl2_ff[39] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6310_ (.RESET_B(net1069),
    .D(net150),
    .Q(\mac1.sum_lvl2_ff[40] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6311_ (.RESET_B(net1071),
    .D(net157),
    .Q(\mac1.sum_lvl2_ff[41] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6312_ (.RESET_B(net1117),
    .D(net254),
    .Q(\mac1.sum_lvl2_ff[42] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6313_ (.RESET_B(net1131),
    .D(net48),
    .Q(\mac1.sum_lvl2_ff[43] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6314_ (.RESET_B(net1131),
    .D(net159),
    .Q(\mac1.sum_lvl2_ff[44] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6315_ (.RESET_B(net1132),
    .D(net244),
    .Q(\mac1.sum_lvl2_ff[45] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6316_ (.RESET_B(net1111),
    .D(net243),
    .Q(\mac1.sum_lvl2_ff[46] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6317_ (.RESET_B(net1138),
    .D(net138),
    .Q(\mac1.sum_lvl2_ff[47] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6318_ (.RESET_B(net1133),
    .D(net109),
    .Q(\mac1.sum_lvl2_ff[48] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6319_ (.RESET_B(net1137),
    .D(net102),
    .Q(\mac1.sum_lvl2_ff[49] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6320_ (.RESET_B(net1073),
    .D(net248),
    .Q(\mac1.sum_lvl2_ff[50] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6321_ (.RESET_B(net1074),
    .D(net166),
    .Q(\mac1.sum_lvl2_ff[51] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6322_ (.RESET_B(net1073),
    .D(net229),
    .Q(\mac1.sum_lvl2_ff[52] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6323_ (.RESET_B(net1089),
    .D(net79),
    .Q(\mac1.sum_lvl2_ff[53] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6324_ (.RESET_B(net1102),
    .D(net190),
    .Q(\mac2.sum_lvl2_ff[38] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6325_ (.RESET_B(net1101),
    .D(net163),
    .Q(\mac2.sum_lvl2_ff[39] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6326_ (.RESET_B(net1100),
    .D(net152),
    .Q(\mac2.sum_lvl2_ff[40] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6327_ (.RESET_B(net1100),
    .D(net165),
    .Q(\mac2.sum_lvl2_ff[41] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6328_ (.RESET_B(net1084),
    .D(net171),
    .Q(\mac2.sum_lvl2_ff[42] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6329_ (.RESET_B(net1082),
    .D(net112),
    .Q(\mac2.sum_lvl2_ff[43] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6330_ (.RESET_B(net1081),
    .D(net47),
    .Q(\mac2.sum_lvl2_ff[44] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6331_ (.RESET_B(net1078),
    .D(net93),
    .Q(\mac2.sum_lvl2_ff[45] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6332_ (.RESET_B(net1077),
    .D(net64),
    .Q(\mac2.sum_lvl2_ff[46] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6333_ (.RESET_B(net1078),
    .D(net51),
    .Q(\mac2.sum_lvl2_ff[47] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6334_ (.RESET_B(net1077),
    .D(net106),
    .Q(\mac2.sum_lvl2_ff[48] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6335_ (.RESET_B(net1077),
    .D(net69),
    .Q(\mac2.sum_lvl2_ff[49] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6336_ (.RESET_B(net1076),
    .D(net94),
    .Q(\mac2.sum_lvl2_ff[50] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6337_ (.RESET_B(net1081),
    .D(net202),
    .Q(\mac2.sum_lvl2_ff[51] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6338_ (.RESET_B(net1084),
    .D(net194),
    .Q(\mac2.sum_lvl2_ff[52] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6339_ (.RESET_B(net1103),
    .D(net44),
    .Q(\mac2.sum_lvl2_ff[53] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6340_ (.RESET_B(net1062),
    .D(net91),
    .Q(\mac1.sum_lvl1_ff[72] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6341_ (.RESET_B(net1062),
    .D(net95),
    .Q(\mac1.sum_lvl1_ff[73] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6342_ (.RESET_B(net1069),
    .D(net43),
    .Q(\mac1.sum_lvl1_ff[74] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6343_ (.RESET_B(net1071),
    .D(net126),
    .Q(\mac1.sum_lvl1_ff[75] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6344_ (.RESET_B(net1116),
    .D(net207),
    .Q(\mac1.sum_lvl1_ff[76] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6345_ (.RESET_B(net1131),
    .D(net135),
    .Q(\mac1.sum_lvl1_ff[77] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6346_ (.RESET_B(net1116),
    .D(net201),
    .Q(\mac1.sum_lvl1_ff[78] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6347_ (.RESET_B(net1132),
    .D(net90),
    .Q(\mac1.sum_lvl1_ff[79] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6348_ (.RESET_B(net1111),
    .D(net176),
    .Q(\mac1.sum_lvl1_ff[80] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6349_ (.RESET_B(net1132),
    .D(net228),
    .Q(\mac1.sum_lvl1_ff[81] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6350_ (.RESET_B(net1133),
    .D(net155),
    .Q(\mac1.sum_lvl1_ff[82] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6351_ (.RESET_B(net1133),
    .D(net57),
    .Q(\mac1.sum_lvl1_ff[83] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6352_ (.RESET_B(net1073),
    .D(net263),
    .Q(\mac1.sum_lvl1_ff[84] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6353_ (.RESET_B(net1073),
    .D(net192),
    .Q(\mac1.sum_lvl1_ff[85] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6354_ (.RESET_B(net1067),
    .D(net223),
    .Q(\mac1.sum_lvl1_ff[86] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6355_ (.RESET_B(net1089),
    .D(net264),
    .Q(\mac1.sum_lvl1_ff[87] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6356_ (.RESET_B(net1102),
    .D(net145),
    .Q(\mac2.sum_lvl1_ff[72] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6357_ (.RESET_B(net1102),
    .D(net61),
    .Q(\mac2.sum_lvl1_ff[73] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6358_ (.RESET_B(net1100),
    .D(net67),
    .Q(\mac2.sum_lvl1_ff[74] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6359_ (.RESET_B(net1086),
    .D(net144),
    .Q(\mac2.sum_lvl1_ff[75] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6360_ (.RESET_B(net1081),
    .D(net153),
    .Q(\mac2.sum_lvl1_ff[76] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6361_ (.RESET_B(net1081),
    .D(net128),
    .Q(\mac2.sum_lvl1_ff[77] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6362_ (.RESET_B(net1079),
    .D(net60),
    .Q(\mac2.sum_lvl1_ff[78] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6363_ (.RESET_B(net1079),
    .D(net196),
    .Q(\mac2.sum_lvl1_ff[79] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6364_ (.RESET_B(net1076),
    .D(net140),
    .Q(\mac2.sum_lvl1_ff[80] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6365_ (.RESET_B(net1079),
    .D(net121),
    .Q(\mac2.sum_lvl1_ff[81] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6366_ (.RESET_B(net1077),
    .D(net236),
    .Q(\mac2.sum_lvl1_ff[82] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6367_ (.RESET_B(net1077),
    .D(net108),
    .Q(\mac2.sum_lvl1_ff[83] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6368_ (.RESET_B(net1076),
    .D(net232),
    .Q(\mac2.sum_lvl1_ff[84] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6369_ (.RESET_B(net1081),
    .D(net258),
    .Q(\mac2.sum_lvl1_ff[85] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6370_ (.RESET_B(net1085),
    .D(net233),
    .Q(\mac2.sum_lvl1_ff[86] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6371_ (.RESET_B(net1101),
    .D(net172),
    .Q(\mac2.sum_lvl1_ff[87] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6372_ (.RESET_B(net1062),
    .D(net170),
    .Q(\mac1.sum_lvl3_ff[20] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6373_ (.RESET_B(net1064),
    .D(net119),
    .Q(\mac1.sum_lvl3_ff[21] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6374_ (.RESET_B(net1069),
    .D(net129),
    .Q(\mac1.sum_lvl3_ff[22] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6375_ (.RESET_B(net1071),
    .D(net161),
    .Q(\mac1.sum_lvl3_ff[23] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6376_ (.RESET_B(net1117),
    .D(net136),
    .Q(\mac1.sum_lvl3_ff[24] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _6377_ (.RESET_B(net1132),
    .D(net193),
    .Q(\mac1.sum_lvl3_ff[25] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _6378_ (.RESET_B(net1131),
    .D(net216),
    .Q(\mac1.sum_lvl3_ff[26] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _6379_ (.RESET_B(net1138),
    .D(net209),
    .Q(\mac1.sum_lvl3_ff[27] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6380_ (.RESET_B(net1111),
    .D(net174),
    .Q(\mac1.sum_lvl3_ff[28] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _6381_ (.RESET_B(net1138),
    .D(net186),
    .Q(\mac1.sum_lvl3_ff[29] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _6382_ (.RESET_B(net1133),
    .D(net187),
    .Q(\mac1.sum_lvl3_ff[30] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _6383_ (.RESET_B(net1137),
    .D(net125),
    .Q(\mac1.sum_lvl3_ff[31] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6384_ (.RESET_B(net1073),
    .D(net104),
    .Q(\mac1.sum_lvl3_ff[32] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6385_ (.RESET_B(net1074),
    .D(net213),
    .Q(\mac1.sum_lvl3_ff[33] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6386_ (.RESET_B(net1073),
    .D(net87),
    .Q(\mac1.sum_lvl3_ff[34] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6387_ (.RESET_B(net1089),
    .D(net143),
    .Q(\mac1.sum_lvl3_ff[35] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6388_ (.RESET_B(net1064),
    .D(net268),
    .Q(\mac1.sum_lvl3_ff[0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6389_ (.RESET_B(net1062),
    .D(net288),
    .Q(\mac1.sum_lvl3_ff[1] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6390_ (.RESET_B(net1069),
    .D(net391),
    .Q(\mac1.sum_lvl3_ff[2] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6391_ (.RESET_B(net1071),
    .D(net477),
    .Q(\mac1.sum_lvl3_ff[3] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6392_ (.RESET_B(net1111),
    .D(net342),
    .Q(\mac1.sum_lvl3_ff[4] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6393_ (.RESET_B(net1111),
    .D(net296),
    .Q(\mac1.sum_lvl3_ff[5] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6394_ (.RESET_B(net1111),
    .D(net464),
    .Q(\mac1.sum_lvl3_ff[6] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6395_ (.RESET_B(net1112),
    .D(net538),
    .Q(\mac1.sum_lvl3_ff[7] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6396_ (.RESET_B(net1112),
    .D(net395),
    .Q(\mac1.sum_lvl3_ff[8] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6397_ (.RESET_B(net1114),
    .D(net459),
    .Q(\mac1.sum_lvl3_ff[9] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6398_ (.RESET_B(net1118),
    .D(net479),
    .Q(\mac1.sum_lvl3_ff[10] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6399_ (.RESET_B(net1118),
    .D(net368),
    .Q(\mac1.sum_lvl3_ff[11] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6400_ (.RESET_B(net1083),
    .D(net321),
    .Q(\mac1.sum_lvl3_ff[12] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6401_ (.RESET_B(net1083),
    .D(net468),
    .Q(\mac1.sum_lvl3_ff[13] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6402_ (.RESET_B(net1083),
    .D(net305),
    .Q(\mac1.sum_lvl3_ff[14] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6403_ (.RESET_B(net1096),
    .D(net286),
    .Q(\mac1.sum_lvl3_ff[15] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6404_ (.RESET_B(net1102),
    .D(net116),
    .Q(\mac2.sum_lvl3_ff[20] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6405_ (.RESET_B(net1101),
    .D(net123),
    .Q(\mac2.sum_lvl3_ff[21] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6406_ (.RESET_B(net1101),
    .D(net195),
    .Q(\mac2.sum_lvl3_ff[22] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6407_ (.RESET_B(net1100),
    .D(net76),
    .Q(\mac2.sum_lvl3_ff[23] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6408_ (.RESET_B(net1084),
    .D(net97),
    .Q(\mac2.sum_lvl3_ff[24] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6409_ (.RESET_B(net1084),
    .D(net115),
    .Q(\mac2.sum_lvl3_ff[25] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6410_ (.RESET_B(net1082),
    .D(net113),
    .Q(\mac2.sum_lvl3_ff[26] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6411_ (.RESET_B(net1082),
    .D(net85),
    .Q(\mac2.sum_lvl3_ff[27] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6412_ (.RESET_B(net1078),
    .D(net205),
    .Q(\mac2.sum_lvl3_ff[28] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6413_ (.RESET_B(net1078),
    .D(net162),
    .Q(\mac2.sum_lvl3_ff[29] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6414_ (.RESET_B(net1067),
    .D(net101),
    .Q(\mac2.sum_lvl3_ff[30] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6415_ (.RESET_B(net1077),
    .D(net118),
    .Q(\mac2.sum_lvl3_ff[31] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6416_ (.RESET_B(net1077),
    .D(net50),
    .Q(\mac2.sum_lvl3_ff[32] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6417_ (.RESET_B(net1081),
    .D(net105),
    .Q(\mac2.sum_lvl3_ff[33] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6418_ (.RESET_B(net1084),
    .D(net92),
    .Q(\mac2.sum_lvl3_ff[34] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6419_ (.RESET_B(net1103),
    .D(net167),
    .Q(\mac2.sum_lvl3_ff[35] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6420_ (.RESET_B(net1061),
    .D(net266),
    .Q(\mac1.total_sum[0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6421_ (.RESET_B(net1061),
    .D(net293),
    .Q(\mac1.total_sum[1] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6422_ (.RESET_B(net1061),
    .D(net383),
    .Q(\mac1.total_sum[2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6423_ (.RESET_B(net1061),
    .D(net443),
    .Q(\mac1.total_sum[3] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6424_ (.RESET_B(net1060),
    .D(_0026_),
    .Q(\mac1.total_sum[4] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6425_ (.RESET_B(net1060),
    .D(_0027_),
    .Q(\mac1.total_sum[5] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6426_ (.RESET_B(net1060),
    .D(_0028_),
    .Q(\mac1.total_sum[6] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6427_ (.RESET_B(net1060),
    .D(_0029_),
    .Q(\mac1.total_sum[7] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6428_ (.RESET_B(net1060),
    .D(net497),
    .Q(\mac1.total_sum[8] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6429_ (.RESET_B(net1065),
    .D(net511),
    .Q(\mac1.total_sum[9] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6430_ (.RESET_B(net1065),
    .D(_0017_),
    .Q(\mac1.total_sum[10] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6431_ (.RESET_B(net1065),
    .D(net526),
    .Q(\mac1.total_sum[11] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6432_ (.RESET_B(net1065),
    .D(_0019_),
    .Q(\mac1.total_sum[12] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6433_ (.RESET_B(net1066),
    .D(net430),
    .Q(\mac1.total_sum[13] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6434_ (.RESET_B(net1066),
    .D(net333),
    .Q(\mac1.total_sum[14] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6435_ (.RESET_B(net1074),
    .D(net291),
    .Q(\mac1.total_sum[15] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6436_ (.RESET_B(net1103),
    .D(_0084_),
    .Q(\mac2.products_ff[0] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6437_ (.RESET_B(net1106),
    .D(_0085_),
    .Q(\mac2.products_ff[1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6438_ (.RESET_B(net1122),
    .D(_0086_),
    .Q(\mac2.products_ff[2] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6439_ (.RESET_B(net1124),
    .D(_0087_),
    .Q(\mac2.products_ff[3] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6440_ (.RESET_B(net1126),
    .D(_0088_),
    .Q(\mac2.products_ff[4] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6441_ (.RESET_B(net1127),
    .D(_0138_),
    .Q(\mac2.products_ff[5] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6442_ (.RESET_B(net1139),
    .D(_0145_),
    .Q(\mac2.products_ff[6] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6443_ (.RESET_B(net1140),
    .D(_0146_),
    .Q(\mac2.products_ff[7] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6444_ (.RESET_B(net1140),
    .D(_0147_),
    .Q(\mac2.products_ff[8] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6445_ (.RESET_B(net1140),
    .D(_0148_),
    .Q(\mac2.products_ff[9] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6446_ (.RESET_B(net1140),
    .D(_0139_),
    .Q(\mac2.products_ff[10] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6447_ (.RESET_B(net1140),
    .D(_0140_),
    .Q(\mac2.products_ff[11] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6448_ (.RESET_B(net1145),
    .D(_0141_),
    .Q(\mac2.products_ff[12] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6449_ (.RESET_B(net1145),
    .D(_0142_),
    .Q(\mac2.products_ff[13] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6450_ (.RESET_B(net1145),
    .D(_0143_),
    .Q(\mac2.products_ff[14] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6451_ (.RESET_B(net1146),
    .D(_0144_),
    .Q(\mac2.products_ff[15] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6452_ (.RESET_B(net1103),
    .D(_0079_),
    .Q(\mac2.products_ff[68] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6453_ (.RESET_B(net1105),
    .D(_0080_),
    .Q(\mac2.products_ff[69] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6454_ (.RESET_B(net1122),
    .D(_0081_),
    .Q(\mac2.products_ff[70] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6455_ (.RESET_B(net1120),
    .D(_0082_),
    .Q(\mac2.products_ff[71] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6456_ (.RESET_B(net1129),
    .D(_0083_),
    .Q(\mac2.products_ff[72] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6457_ (.RESET_B(net1118),
    .D(_0127_),
    .Q(\mac2.products_ff[73] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6458_ (.RESET_B(net1134),
    .D(_0134_),
    .Q(\mac2.products_ff[74] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6459_ (.RESET_B(net1134),
    .D(_0135_),
    .Q(\mac2.products_ff[75] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6460_ (.RESET_B(net1134),
    .D(_0136_),
    .Q(\mac2.products_ff[76] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6461_ (.RESET_B(net1133),
    .D(_0137_),
    .Q(\mac2.products_ff[77] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6462_ (.RESET_B(net1133),
    .D(_0128_),
    .Q(\mac2.products_ff[78] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6463_ (.RESET_B(net1134),
    .D(_0129_),
    .Q(\mac2.products_ff[79] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6464_ (.RESET_B(net1141),
    .D(_0130_),
    .Q(\mac2.products_ff[80] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6465_ (.RESET_B(net1141),
    .D(_0131_),
    .Q(\mac2.products_ff[81] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6466_ (.RESET_B(net1140),
    .D(_0132_),
    .Q(\mac2.products_ff[82] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6467_ (.RESET_B(net1140),
    .D(_0133_),
    .Q(\mac2.products_ff[83] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6468_ (.RESET_B(net1100),
    .D(_0089_),
    .Q(\mac2.products_ff[136] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6469_ (.RESET_B(net1100),
    .D(_0090_),
    .Q(\mac2.products_ff[137] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6470_ (.RESET_B(net1086),
    .D(_0091_),
    .Q(\mac2.products_ff[138] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6471_ (.RESET_B(net1086),
    .D(_0092_),
    .Q(\mac2.products_ff[139] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6472_ (.RESET_B(net1081),
    .D(_0093_),
    .Q(\mac2.products_ff[140] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6473_ (.RESET_B(net1081),
    .D(_0149_),
    .Q(\mac2.products_ff[141] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6474_ (.RESET_B(net1079),
    .D(_0156_),
    .Q(\mac2.products_ff[142] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6475_ (.RESET_B(net1075),
    .D(_0157_),
    .Q(\mac2.products_ff[143] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6476_ (.RESET_B(net1075),
    .D(_0158_),
    .Q(\mac2.products_ff[144] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6477_ (.RESET_B(net1075),
    .D(_0159_),
    .Q(\mac2.products_ff[145] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6478_ (.RESET_B(net1079),
    .D(_0150_),
    .Q(\mac2.products_ff[146] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6479_ (.RESET_B(net1079),
    .D(_0151_),
    .Q(\mac2.products_ff[147] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6480_ (.RESET_B(net1075),
    .D(_0152_),
    .Q(\mac2.products_ff[148] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6481_ (.RESET_B(net1085),
    .D(_0153_),
    .Q(\mac2.products_ff[149] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6482_ (.RESET_B(net1085),
    .D(_0154_),
    .Q(\mac2.products_ff[150] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6483_ (.RESET_B(net1101),
    .D(_0155_),
    .Q(\mac2.products_ff[151] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6484_ (.RESET_B(net1103),
    .D(net185),
    .Q(\mac2.sum_lvl1_ff[0] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6485_ (.RESET_B(net1105),
    .D(net220),
    .Q(\mac2.sum_lvl1_ff[1] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6486_ (.RESET_B(net1122),
    .D(net169),
    .Q(\mac2.sum_lvl1_ff[2] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6487_ (.RESET_B(net1124),
    .D(net179),
    .Q(\mac2.sum_lvl1_ff[3] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6488_ (.RESET_B(net1127),
    .D(net133),
    .Q(\mac2.sum_lvl1_ff[4] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6489_ (.RESET_B(net1139),
    .D(net249),
    .Q(\mac2.sum_lvl1_ff[5] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6490_ (.RESET_B(net1141),
    .D(net261),
    .Q(\mac2.sum_lvl1_ff[6] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6491_ (.RESET_B(net1141),
    .D(net160),
    .Q(\mac2.sum_lvl1_ff[7] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6492_ (.RESET_B(net1144),
    .D(net235),
    .Q(\mac2.sum_lvl1_ff[8] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6493_ (.RESET_B(net1140),
    .D(net83),
    .Q(\mac2.sum_lvl1_ff[9] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6494_ (.RESET_B(net1142),
    .D(net80),
    .Q(\mac2.sum_lvl1_ff[10] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6495_ (.RESET_B(net1142),
    .D(net84),
    .Q(\mac2.sum_lvl1_ff[11] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6496_ (.RESET_B(net1142),
    .D(net225),
    .Q(\mac2.sum_lvl1_ff[12] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6497_ (.RESET_B(net1142),
    .D(net242),
    .Q(\mac2.sum_lvl1_ff[13] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6498_ (.RESET_B(net1145),
    .D(net130),
    .Q(\mac2.sum_lvl1_ff[14] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6499_ (.RESET_B(net1145),
    .D(net70),
    .Q(\mac2.sum_lvl1_ff[15] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6500_ (.RESET_B(net1103),
    .D(net49),
    .Q(\mac2.sum_lvl1_ff[36] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6501_ (.RESET_B(net1105),
    .D(net218),
    .Q(\mac2.sum_lvl1_ff[37] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6502_ (.RESET_B(net1122),
    .D(net154),
    .Q(\mac2.sum_lvl1_ff[38] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6503_ (.RESET_B(net1120),
    .D(net238),
    .Q(\mac2.sum_lvl1_ff[39] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6504_ (.RESET_B(net1118),
    .D(net214),
    .Q(\mac2.sum_lvl1_ff[40] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6505_ (.RESET_B(net1118),
    .D(net184),
    .Q(\mac2.sum_lvl1_ff[41] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6506_ (.RESET_B(net1136),
    .D(net131),
    .Q(\mac2.sum_lvl1_ff[42] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6507_ (.RESET_B(net1136),
    .D(net114),
    .Q(\mac2.sum_lvl1_ff[43] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6508_ (.RESET_B(net1136),
    .D(net199),
    .Q(\mac2.sum_lvl1_ff[44] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6509_ (.RESET_B(net1136),
    .D(net252),
    .Q(\mac2.sum_lvl1_ff[45] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6510_ (.RESET_B(net1136),
    .D(net245),
    .Q(\mac2.sum_lvl1_ff[46] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6511_ (.RESET_B(net1136),
    .D(net224),
    .Q(\mac2.sum_lvl1_ff[47] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6512_ (.RESET_B(net1141),
    .D(net110),
    .Q(\mac2.sum_lvl1_ff[48] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6513_ (.RESET_B(net1141),
    .D(net178),
    .Q(\mac2.sum_lvl1_ff[49] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6514_ (.RESET_B(net1142),
    .D(net45),
    .Q(\mac2.sum_lvl1_ff[50] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6515_ (.RESET_B(net1142),
    .D(net240),
    .Q(\mac2.sum_lvl1_ff[51] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6516_ (.RESET_B(net1103),
    .D(net100),
    .Q(\mac2.sum_lvl2_ff[0] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6517_ (.RESET_B(net1105),
    .D(net65),
    .Q(\mac2.sum_lvl2_ff[1] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6518_ (.RESET_B(net1124),
    .D(net158),
    .Q(\mac2.sum_lvl2_ff[2] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6519_ (.RESET_B(net1126),
    .D(net222),
    .Q(\mac2.sum_lvl2_ff[3] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6520_ (.RESET_B(net1129),
    .D(net198),
    .Q(\mac2.sum_lvl2_ff[4] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6521_ (.RESET_B(net1139),
    .D(net227),
    .Q(\mac2.sum_lvl2_ff[5] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6522_ (.RESET_B(net1141),
    .D(net82),
    .Q(\mac2.sum_lvl2_ff[6] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6523_ (.RESET_B(net1143),
    .D(net221),
    .Q(\mac2.sum_lvl2_ff[7] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6524_ (.RESET_B(net1143),
    .D(net247),
    .Q(\mac2.sum_lvl2_ff[8] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6525_ (.RESET_B(net1143),
    .D(net259),
    .Q(\mac2.sum_lvl2_ff[9] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6526_ (.RESET_B(net1143),
    .D(net257),
    .Q(\mac2.sum_lvl2_ff[10] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6527_ (.RESET_B(net1143),
    .D(net256),
    .Q(\mac2.sum_lvl2_ff[11] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6528_ (.RESET_B(net1143),
    .D(net251),
    .Q(\mac2.sum_lvl2_ff[12] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6529_ (.RESET_B(net1144),
    .D(net250),
    .Q(\mac2.sum_lvl2_ff[13] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _6530_ (.RESET_B(net1145),
    .D(net117),
    .Q(\mac2.sum_lvl2_ff[14] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6531_ (.RESET_B(net1145),
    .D(net137),
    .Q(\mac2.sum_lvl2_ff[15] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6532_ (.RESET_B(net1103),
    .D(net66),
    .Q(\mac2.sum_lvl2_ff[19] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6533_ (.RESET_B(net1105),
    .D(net122),
    .Q(\mac2.sum_lvl2_ff[20] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6534_ (.RESET_B(net1124),
    .D(net210),
    .Q(\mac2.sum_lvl2_ff[21] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6535_ (.RESET_B(net1120),
    .D(net203),
    .Q(\mac2.sum_lvl2_ff[22] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6536_ (.RESET_B(net1118),
    .D(net173),
    .Q(\mac2.sum_lvl2_ff[23] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _6537_ (.RESET_B(net1135),
    .D(net231),
    .Q(\mac2.sum_lvl2_ff[24] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6538_ (.RESET_B(net1136),
    .D(net180),
    .Q(\mac2.sum_lvl2_ff[25] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6539_ (.RESET_B(net1137),
    .D(net53),
    .Q(\mac2.sum_lvl2_ff[26] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6540_ (.RESET_B(net1137),
    .D(net191),
    .Q(\mac2.sum_lvl2_ff[27] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6541_ (.RESET_B(net1137),
    .D(net55),
    .Q(\mac2.sum_lvl2_ff[28] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6542_ (.RESET_B(net1141),
    .D(net41),
    .Q(\mac2.sum_lvl2_ff[29] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6543_ (.RESET_B(net1136),
    .D(net111),
    .Q(\mac2.sum_lvl2_ff[30] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6544_ (.RESET_B(net1143),
    .D(net89),
    .Q(\mac2.sum_lvl2_ff[31] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6545_ (.RESET_B(net1142),
    .D(net132),
    .Q(\mac2.sum_lvl2_ff[32] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6546_ (.RESET_B(net1142),
    .D(net141),
    .Q(\mac2.sum_lvl2_ff[33] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6547_ (.RESET_B(net1145),
    .D(net75),
    .Q(\mac2.sum_lvl2_ff[34] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _6548_ (.RESET_B(net1076),
    .D(net1),
    .Q(\DP_1.I_range.out_data[2] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6549_ (.RESET_B(net1076),
    .D(net2),
    .Q(\DP_1.I_range.out_data[3] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6550_ (.RESET_B(net1076),
    .D(net3),
    .Q(\DP_1.I_range.out_data[4] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6551_ (.RESET_B(net1075),
    .D(\DP_1.I_range.data_plus_4[6] ),
    .Q(\DP_1.I_range.out_data[5] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6552_ (.RESET_B(net1102),
    .D(net272),
    .Q(\mac2.sum_lvl3_ff[0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6553_ (.RESET_B(net1101),
    .D(net309),
    .Q(\mac2.sum_lvl3_ff[1] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6554_ (.RESET_B(net1101),
    .D(net352),
    .Q(\mac2.sum_lvl3_ff[2] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6555_ (.RESET_B(net1096),
    .D(net434),
    .Q(\mac2.sum_lvl3_ff[3] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6556_ (.RESET_B(net1083),
    .D(net514),
    .Q(\mac2.sum_lvl3_ff[4] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _6557_ (.RESET_B(net1083),
    .D(net471),
    .Q(\mac2.sum_lvl3_ff[5] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6558_ (.RESET_B(net1083),
    .D(_0044_),
    .Q(\mac2.sum_lvl3_ff[6] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6559_ (.RESET_B(net1082),
    .D(_0045_),
    .Q(\mac2.sum_lvl3_ff[7] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6560_ (.RESET_B(net1073),
    .D(net520),
    .Q(\mac2.sum_lvl3_ff[8] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6561_ (.RESET_B(net1067),
    .D(_0047_),
    .Q(\mac2.sum_lvl3_ff[9] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6562_ (.RESET_B(net1067),
    .D(_0033_),
    .Q(\mac2.sum_lvl3_ff[10] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6563_ (.RESET_B(net1077),
    .D(_0034_),
    .Q(\mac2.sum_lvl3_ff[11] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6564_ (.RESET_B(net1082),
    .D(_0035_),
    .Q(\mac2.sum_lvl3_ff[12] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6565_ (.RESET_B(net1084),
    .D(_0036_),
    .Q(\mac2.sum_lvl3_ff[13] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6566_ (.RESET_B(net1084),
    .D(_0037_),
    .Q(\mac2.sum_lvl3_ff[14] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6567_ (.RESET_B(net1129),
    .D(net486),
    .Q(\mac2.sum_lvl3_ff[15] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6568_ (.RESET_B(net1061),
    .D(net326),
    .Q(\mac2.total_sum[0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6569_ (.RESET_B(net1061),
    .D(net481),
    .Q(\mac2.total_sum[1] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6570_ (.RESET_B(net1061),
    .D(net500),
    .Q(\mac2.total_sum[2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6571_ (.RESET_B(net1060),
    .D(net503),
    .Q(\mac2.total_sum[3] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6572_ (.RESET_B(net1060),
    .D(net446),
    .Q(\mac2.total_sum[4] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6573_ (.RESET_B(net1060),
    .D(net361),
    .Q(\mac2.total_sum[5] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6574_ (.RESET_B(net1061),
    .D(net490),
    .Q(\mac2.total_sum[6] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6575_ (.RESET_B(net1065),
    .D(_0061_),
    .Q(\mac2.total_sum[7] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6576_ (.RESET_B(net1065),
    .D(net457),
    .Q(\mac2.total_sum[8] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6577_ (.RESET_B(net1066),
    .D(net317),
    .Q(\mac2.total_sum[9] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6578_ (.RESET_B(net1065),
    .D(net348),
    .Q(\mac2.total_sum[10] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6579_ (.RESET_B(net1065),
    .D(net403),
    .Q(\mac2.total_sum[11] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6580_ (.RESET_B(net1066),
    .D(_0051_),
    .Q(\mac2.total_sum[12] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6581_ (.RESET_B(net1066),
    .D(net413),
    .Q(\mac2.total_sum[13] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6582_ (.RESET_B(net1066),
    .D(net299),
    .Q(\mac2.total_sum[14] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6583_ (.RESET_B(net1074),
    .D(net439),
    .Q(\mac2.total_sum[15] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _6584_ (.RESET_B(net1076),
    .D(net5),
    .Q(\DP_1.Q_range.out_data[2] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6585_ (.RESET_B(net1075),
    .D(net6),
    .Q(\DP_1.Q_range.out_data[3] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6586_ (.RESET_B(net1075),
    .D(net7),
    .Q(\DP_1.Q_range.out_data[4] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6587_ (.RESET_B(net1075),
    .D(\DP_1.Q_range.data_plus_4[6] ),
    .Q(\DP_1.Q_range.out_data[5] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _6588_ (.RESET_B(net1080),
    .D(net13),
    .Q(\DP_3.I_range.out_data[2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6589_ (.RESET_B(net1080),
    .D(net14),
    .Q(\DP_3.I_range.out_data[3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6590_ (.RESET_B(net1086),
    .D(net15),
    .Q(\DP_3.I_range.out_data[4] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6591_ (.RESET_B(net1086),
    .D(\DP_3.I_range.data_plus_4[6] ),
    .Q(\DP_3.I_range.out_data[5] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_tiehi heichips25_template_34 (.L_HI(net34));
 sg13g2_tiehi heichips25_template_35 (.L_HI(net35));
 sg13g2_tiehi heichips25_template_36 (.L_HI(net36));
 sg13g2_tiehi heichips25_template_37 (.L_HI(net37));
 sg13g2_tiehi heichips25_template_38 (.L_HI(net38));
 sg13g2_tiehi heichips25_template_39 (.L_HI(net39));
 sg13g2_tiehi heichips25_template_40 (.L_HI(net40));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_2 fanout783 (.A(net788),
    .X(net783));
 sg13g2_buf_1 fanout784 (.A(net785),
    .X(net784));
 sg13g2_buf_8 fanout785 (.A(net788),
    .X(net785));
 sg13g2_buf_8 fanout786 (.A(net788),
    .X(net786));
 sg13g2_buf_1 fanout787 (.A(net788),
    .X(net787));
 sg13g2_buf_2 fanout788 (.A(_2393_),
    .X(net788));
 sg13g2_buf_8 fanout789 (.A(net507),
    .X(net789));
 sg13g2_buf_1 fanout790 (.A(_2475_),
    .X(net790));
 sg13g2_buf_8 fanout791 (.A(net792),
    .X(net791));
 sg13g2_buf_8 fanout792 (.A(net793),
    .X(net792));
 sg13g2_buf_8 fanout793 (.A(_2475_),
    .X(net793));
 sg13g2_buf_8 fanout794 (.A(net796),
    .X(net794));
 sg13g2_buf_8 fanout795 (.A(_2481_),
    .X(net795));
 sg13g2_buf_1 fanout796 (.A(_2481_),
    .X(net796));
 sg13g2_buf_8 fanout797 (.A(net798),
    .X(net797));
 sg13g2_buf_8 fanout798 (.A(_2480_),
    .X(net798));
 sg13g2_buf_8 fanout799 (.A(_2401_),
    .X(net799));
 sg13g2_buf_8 fanout800 (.A(_2401_),
    .X(net800));
 sg13g2_buf_8 fanout801 (.A(_2398_),
    .X(net801));
 sg13g2_buf_2 fanout802 (.A(_2398_),
    .X(net802));
 sg13g2_buf_8 fanout803 (.A(net804),
    .X(net803));
 sg13g2_buf_8 fanout804 (.A(_2479_),
    .X(net804));
 sg13g2_buf_8 fanout805 (.A(_2479_),
    .X(net805));
 sg13g2_buf_8 fanout806 (.A(_2478_),
    .X(net806));
 sg13g2_buf_1 fanout807 (.A(_2478_),
    .X(net807));
 sg13g2_buf_8 fanout808 (.A(_2397_),
    .X(net808));
 sg13g2_buf_8 fanout809 (.A(net810),
    .X(net809));
 sg13g2_buf_8 fanout810 (.A(_2396_),
    .X(net810));
 sg13g2_buf_8 fanout811 (.A(net813),
    .X(net811));
 sg13g2_buf_1 fanout812 (.A(net813),
    .X(net812));
 sg13g2_buf_2 fanout813 (.A(net324),
    .X(net813));
 sg13g2_buf_8 fanout814 (.A(\DP_4.matrix[78] ),
    .X(net814));
 sg13g2_buf_1 fanout815 (.A(net419),
    .X(net815));
 sg13g2_buf_8 fanout816 (.A(net817),
    .X(net816));
 sg13g2_buf_2 fanout817 (.A(net318),
    .X(net817));
 sg13g2_buf_8 fanout818 (.A(net819),
    .X(net818));
 sg13g2_buf_1 fanout819 (.A(\DP_4.matrix[76] ),
    .X(net819));
 sg13g2_buf_8 fanout820 (.A(net821),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(\DP_4.matrix[75] ),
    .X(net821));
 sg13g2_buf_8 fanout822 (.A(net823),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(net370),
    .X(net823));
 sg13g2_buf_8 fanout824 (.A(net826),
    .X(net824));
 sg13g2_buf_8 fanout825 (.A(net826),
    .X(net825));
 sg13g2_buf_8 fanout826 (.A(net827),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(net473),
    .X(net827));
 sg13g2_buf_8 fanout828 (.A(net830),
    .X(net828));
 sg13g2_buf_1 fanout829 (.A(net830),
    .X(net829));
 sg13g2_buf_1 fanout830 (.A(net831),
    .X(net830));
 sg13g2_buf_1 fanout831 (.A(net832),
    .X(net831));
 sg13g2_buf_1 fanout832 (.A(net376),
    .X(net832));
 sg13g2_buf_8 fanout833 (.A(net334),
    .X(net833));
 sg13g2_buf_1 fanout834 (.A(\DP_4.matrix[43] ),
    .X(net834));
 sg13g2_buf_8 fanout835 (.A(net335),
    .X(net835));
 sg13g2_buf_1 fanout836 (.A(\DP_4.matrix[42] ),
    .X(net836));
 sg13g2_buf_8 fanout837 (.A(net364),
    .X(net837));
 sg13g2_buf_8 fanout838 (.A(net330),
    .X(net838));
 sg13g2_buf_1 fanout839 (.A(\DP_4.matrix[40] ),
    .X(net839));
 sg13g2_buf_8 fanout840 (.A(net398),
    .X(net840));
 sg13g2_buf_1 fanout841 (.A(net398),
    .X(net841));
 sg13g2_buf_8 fanout842 (.A(net329),
    .X(net842));
 sg13g2_buf_1 fanout843 (.A(\DP_4.matrix[38] ),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(net846),
    .X(net844));
 sg13g2_buf_1 fanout845 (.A(\DP_4.matrix[37] ),
    .X(net845));
 sg13g2_buf_8 fanout846 (.A(\DP_4.matrix[37] ),
    .X(net846));
 sg13g2_buf_8 fanout847 (.A(net373),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(net849),
    .X(net848));
 sg13g2_buf_8 fanout849 (.A(\DP_4.matrix[36] ),
    .X(net849));
 sg13g2_buf_8 fanout850 (.A(net343),
    .X(net850));
 sg13g2_buf_8 fanout851 (.A(net853),
    .X(net851));
 sg13g2_buf_1 fanout852 (.A(net853),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(net405),
    .X(net853));
 sg13g2_buf_8 fanout854 (.A(net855),
    .X(net854));
 sg13g2_buf_8 fanout855 (.A(net357),
    .X(net855));
 sg13g2_buf_8 fanout856 (.A(net450),
    .X(net856));
 sg13g2_buf_8 fanout857 (.A(net371),
    .X(net857));
 sg13g2_buf_1 fanout858 (.A(\DP_4.matrix[4] ),
    .X(net858));
 sg13g2_buf_8 fanout859 (.A(net384),
    .X(net859));
 sg13g2_buf_1 fanout860 (.A(\DP_4.matrix[3] ),
    .X(net860));
 sg13g2_buf_8 fanout861 (.A(net379),
    .X(net861));
 sg13g2_buf_1 fanout862 (.A(\DP_4.matrix[2] ),
    .X(net862));
 sg13g2_buf_8 fanout863 (.A(net866),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(net865),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(net866),
    .X(net865));
 sg13g2_buf_8 fanout866 (.A(net474),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(net868),
    .X(net867));
 sg13g2_buf_8 fanout868 (.A(net374),
    .X(net868));
 sg13g2_buf_8 fanout869 (.A(net374),
    .X(net869));
 sg13g2_buf_8 fanout870 (.A(net872),
    .X(net870));
 sg13g2_buf_1 fanout871 (.A(net872),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(\DP_3.matrix[79] ),
    .X(net872));
 sg13g2_buf_8 fanout873 (.A(net874),
    .X(net873));
 sg13g2_buf_8 fanout874 (.A(\DP_3.matrix[78] ),
    .X(net874));
 sg13g2_buf_8 fanout875 (.A(net876),
    .X(net875));
 sg13g2_buf_8 fanout876 (.A(\DP_3.matrix[77] ),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(net878),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(net879),
    .X(net878));
 sg13g2_buf_1 fanout879 (.A(net353),
    .X(net879));
 sg13g2_buf_8 fanout880 (.A(net881),
    .X(net880));
 sg13g2_buf_1 fanout881 (.A(net882),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(net301),
    .X(net882));
 sg13g2_buf_8 fanout883 (.A(net884),
    .X(net883));
 sg13g2_buf_1 fanout884 (.A(net885),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(net307),
    .X(net885));
 sg13g2_buf_8 fanout886 (.A(net887),
    .X(net886));
 sg13g2_buf_1 fanout887 (.A(net888),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(net310),
    .X(net888));
 sg13g2_buf_8 fanout889 (.A(net890),
    .X(net889));
 sg13g2_buf_1 fanout890 (.A(net275),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(net892),
    .X(net891));
 sg13g2_buf_1 fanout892 (.A(net893),
    .X(net892));
 sg13g2_buf_8 fanout893 (.A(net529),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(net895),
    .X(net894));
 sg13g2_buf_8 fanout895 (.A(net539),
    .X(net895));
 sg13g2_buf_8 fanout896 (.A(\DP_3.matrix[41] ),
    .X(net896));
 sg13g2_buf_8 fanout897 (.A(net356),
    .X(net897));
 sg13g2_buf_8 fanout898 (.A(\DP_3.matrix[40] ),
    .X(net898));
 sg13g2_buf_8 fanout899 (.A(net337),
    .X(net899));
 sg13g2_buf_8 fanout900 (.A(net901),
    .X(net900));
 sg13g2_buf_8 fanout901 (.A(net483),
    .X(net901));
 sg13g2_buf_8 fanout902 (.A(net339),
    .X(net902));
 sg13g2_buf_8 fanout903 (.A(\DP_3.matrix[38] ),
    .X(net903));
 sg13g2_buf_8 fanout904 (.A(net905),
    .X(net904));
 sg13g2_buf_8 fanout905 (.A(net338),
    .X(net905));
 sg13g2_buf_8 fanout906 (.A(net349),
    .X(net906));
 sg13g2_buf_1 fanout907 (.A(\DP_3.matrix[36] ),
    .X(net907));
 sg13g2_buf_8 fanout908 (.A(net909),
    .X(net908));
 sg13g2_buf_8 fanout909 (.A(net910),
    .X(net909));
 sg13g2_buf_2 fanout910 (.A(net451),
    .X(net910));
 sg13g2_buf_8 fanout911 (.A(net913),
    .X(net911));
 sg13g2_buf_1 fanout912 (.A(net913),
    .X(net912));
 sg13g2_buf_8 fanout913 (.A(net345),
    .X(net913));
 sg13g2_buf_8 fanout914 (.A(net915),
    .X(net914));
 sg13g2_buf_8 fanout915 (.A(net447),
    .X(net915));
 sg13g2_buf_8 fanout916 (.A(net420),
    .X(net916));
 sg13g2_buf_8 fanout917 (.A(\DP_3.matrix[4] ),
    .X(net917));
 sg13g2_buf_8 fanout918 (.A(net387),
    .X(net918));
 sg13g2_buf_8 fanout919 (.A(\DP_3.matrix[3] ),
    .X(net919));
 sg13g2_buf_8 fanout920 (.A(net435),
    .X(net920));
 sg13g2_buf_8 fanout921 (.A(\DP_3.matrix[2] ),
    .X(net921));
 sg13g2_buf_8 fanout922 (.A(net923),
    .X(net922));
 sg13g2_buf_8 fanout923 (.A(net422),
    .X(net923));
 sg13g2_buf_8 fanout924 (.A(net355),
    .X(net924));
 sg13g2_buf_1 fanout925 (.A(\DP_3.matrix[0] ),
    .X(net925));
 sg13g2_buf_8 fanout926 (.A(net927),
    .X(net926));
 sg13g2_buf_8 fanout927 (.A(net523),
    .X(net927));
 sg13g2_buf_8 fanout928 (.A(net929),
    .X(net928));
 sg13g2_buf_2 fanout929 (.A(net426),
    .X(net929));
 sg13g2_buf_8 fanout930 (.A(net931),
    .X(net930));
 sg13g2_buf_8 fanout931 (.A(net311),
    .X(net931));
 sg13g2_buf_8 fanout932 (.A(net933),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(net404),
    .X(net933));
 sg13g2_buf_8 fanout934 (.A(net935),
    .X(net934));
 sg13g2_buf_1 fanout935 (.A(net550),
    .X(net935));
 sg13g2_buf_8 fanout936 (.A(net937),
    .X(net936));
 sg13g2_buf_8 fanout937 (.A(net482),
    .X(net937));
 sg13g2_buf_2 fanout938 (.A(net939),
    .X(net938));
 sg13g2_buf_1 fanout939 (.A(net940),
    .X(net939));
 sg13g2_buf_1 fanout940 (.A(net941),
    .X(net940));
 sg13g2_buf_1 fanout941 (.A(net543),
    .X(net941));
 sg13g2_buf_8 fanout942 (.A(\DP_2.matrix[73] ),
    .X(net942));
 sg13g2_buf_8 fanout943 (.A(net944),
    .X(net943));
 sg13g2_buf_1 fanout944 (.A(net945),
    .X(net944));
 sg13g2_buf_1 fanout945 (.A(\DP_2.matrix[72] ),
    .X(net945));
 sg13g2_buf_8 fanout946 (.A(net491),
    .X(net946));
 sg13g2_buf_8 fanout947 (.A(net948),
    .X(net947));
 sg13g2_buf_8 fanout948 (.A(net300),
    .X(net948));
 sg13g2_buf_8 fanout949 (.A(\DP_2.matrix[42] ),
    .X(net949));
 sg13g2_buf_1 fanout950 (.A(net415),
    .X(net950));
 sg13g2_buf_8 fanout951 (.A(net400),
    .X(net951));
 sg13g2_buf_8 fanout952 (.A(\DP_2.matrix[40] ),
    .X(net952));
 sg13g2_buf_1 fanout953 (.A(net452),
    .X(net953));
 sg13g2_buf_8 fanout954 (.A(\DP_2.matrix[39] ),
    .X(net954));
 sg13g2_buf_1 fanout955 (.A(net431),
    .X(net955));
 sg13g2_buf_8 fanout956 (.A(net957),
    .X(net956));
 sg13g2_buf_8 fanout957 (.A(net306),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(net959),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(net960),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(net961),
    .X(net960));
 sg13g2_buf_8 fanout961 (.A(net524),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(net964),
    .X(net962));
 sg13g2_buf_1 fanout963 (.A(net964),
    .X(net963));
 sg13g2_buf_1 fanout964 (.A(net965),
    .X(net964));
 sg13g2_buf_8 fanout965 (.A(net363),
    .X(net965));
 sg13g2_buf_8 fanout966 (.A(net968),
    .X(net966));
 sg13g2_buf_1 fanout967 (.A(net968),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(net377),
    .X(net968));
 sg13g2_buf_8 fanout969 (.A(net416),
    .X(net969));
 sg13g2_buf_1 fanout970 (.A(\DP_2.matrix[6] ),
    .X(net970));
 sg13g2_buf_8 fanout971 (.A(net460),
    .X(net971));
 sg13g2_buf_8 fanout972 (.A(net414),
    .X(net972));
 sg13g2_buf_1 fanout973 (.A(\DP_2.matrix[4] ),
    .X(net973));
 sg13g2_buf_8 fanout974 (.A(net406),
    .X(net974));
 sg13g2_buf_1 fanout975 (.A(\DP_2.matrix[3] ),
    .X(net975));
 sg13g2_buf_8 fanout976 (.A(net440),
    .X(net976));
 sg13g2_buf_1 fanout977 (.A(\DP_2.matrix[2] ),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(net472),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(net981),
    .X(net979));
 sg13g2_buf_1 fanout980 (.A(net981),
    .X(net980));
 sg13g2_buf_1 fanout981 (.A(\DP_2.matrix[1] ),
    .X(net981));
 sg13g2_buf_8 fanout982 (.A(net322),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(net984),
    .X(net983));
 sg13g2_buf_1 fanout984 (.A(net985),
    .X(net984));
 sg13g2_buf_1 fanout985 (.A(\DP_2.matrix[0] ),
    .X(net985));
 sg13g2_buf_2 fanout986 (.A(net987),
    .X(net986));
 sg13g2_buf_1 fanout987 (.A(net988),
    .X(net987));
 sg13g2_buf_1 fanout988 (.A(\DP_1.matrix[79] ),
    .X(net988));
 sg13g2_buf_8 fanout989 (.A(net990),
    .X(net989));
 sg13g2_buf_8 fanout990 (.A(net544),
    .X(net990));
 sg13g2_buf_8 fanout991 (.A(net993),
    .X(net991));
 sg13g2_buf_1 fanout992 (.A(net993),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(net542),
    .X(net993));
 sg13g2_buf_8 fanout994 (.A(net995),
    .X(net994));
 sg13g2_buf_8 fanout995 (.A(net528),
    .X(net995));
 sg13g2_buf_8 fanout996 (.A(net997),
    .X(net996));
 sg13g2_buf_8 fanout997 (.A(net314),
    .X(net997));
 sg13g2_buf_8 fanout998 (.A(net999),
    .X(net998));
 sg13g2_buf_8 fanout999 (.A(net492),
    .X(net999));
 sg13g2_buf_8 fanout1000 (.A(net1001),
    .X(net1000));
 sg13g2_buf_1 fanout1001 (.A(net1002),
    .X(net1001));
 sg13g2_buf_8 fanout1002 (.A(net515),
    .X(net1002));
 sg13g2_buf_8 fanout1003 (.A(net424),
    .X(net1003));
 sg13g2_buf_1 fanout1004 (.A(net424),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(net1006),
    .X(net1005));
 sg13g2_buf_1 fanout1006 (.A(net1007),
    .X(net1006));
 sg13g2_buf_2 fanout1007 (.A(net399),
    .X(net1007));
 sg13g2_buf_8 fanout1008 (.A(net369),
    .X(net1008));
 sg13g2_buf_1 fanout1009 (.A(\DP_1.matrix[42] ),
    .X(net1009));
 sg13g2_buf_8 fanout1010 (.A(net1012),
    .X(net1010));
 sg13g2_buf_1 fanout1011 (.A(net1012),
    .X(net1011));
 sg13g2_buf_2 fanout1012 (.A(net323),
    .X(net1012));
 sg13g2_buf_8 fanout1013 (.A(net1015),
    .X(net1013));
 sg13g2_buf_1 fanout1014 (.A(net1015),
    .X(net1014));
 sg13g2_buf_2 fanout1015 (.A(net313),
    .X(net1015));
 sg13g2_buf_8 fanout1016 (.A(net1017),
    .X(net1016));
 sg13g2_buf_8 fanout1017 (.A(net312),
    .X(net1017));
 sg13g2_buf_8 fanout1018 (.A(net1020),
    .X(net1018));
 sg13g2_buf_1 fanout1019 (.A(net1020),
    .X(net1019));
 sg13g2_buf_2 fanout1020 (.A(net493),
    .X(net1020));
 sg13g2_buf_8 fanout1021 (.A(net1022),
    .X(net1021));
 sg13g2_buf_8 fanout1022 (.A(net448),
    .X(net1022));
 sg13g2_buf_8 fanout1023 (.A(net328),
    .X(net1023));
 sg13g2_buf_1 fanout1024 (.A(\DP_1.matrix[36] ),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(\DP_1.matrix[7] ),
    .X(net1025));
 sg13g2_buf_8 fanout1026 (.A(\DP_1.matrix[7] ),
    .X(net1026));
 sg13g2_buf_8 fanout1027 (.A(net1029),
    .X(net1027));
 sg13g2_buf_1 fanout1028 (.A(net1029),
    .X(net1028));
 sg13g2_buf_8 fanout1029 (.A(net408),
    .X(net1029));
 sg13g2_buf_8 fanout1030 (.A(net1031),
    .X(net1030));
 sg13g2_buf_8 fanout1031 (.A(\DP_1.matrix[5] ),
    .X(net1031));
 sg13g2_buf_8 fanout1032 (.A(net1033),
    .X(net1032));
 sg13g2_buf_8 fanout1033 (.A(net396),
    .X(net1033));
 sg13g2_buf_8 fanout1034 (.A(net453),
    .X(net1034));
 sg13g2_buf_8 fanout1035 (.A(\DP_1.matrix[3] ),
    .X(net1035));
 sg13g2_buf_8 fanout1036 (.A(net425),
    .X(net1036));
 sg13g2_buf_8 fanout1037 (.A(\DP_1.matrix[2] ),
    .X(net1037));
 sg13g2_buf_8 fanout1038 (.A(net1039),
    .X(net1038));
 sg13g2_buf_8 fanout1039 (.A(net504),
    .X(net1039));
 sg13g2_buf_8 fanout1040 (.A(net336),
    .X(net1040));
 sg13g2_buf_1 fanout1041 (.A(\DP_1.matrix[0] ),
    .X(net1041));
 sg13g2_buf_8 fanout1042 (.A(\DP_4.matrix[80] ),
    .X(net1042));
 sg13g2_buf_8 fanout1043 (.A(net344),
    .X(net1043));
 sg13g2_buf_8 fanout1044 (.A(net327),
    .X(net1044));
 sg13g2_buf_8 fanout1045 (.A(net1046),
    .X(net1045));
 sg13g2_buf_1 fanout1046 (.A(\DP_3.matrix[80] ),
    .X(net1046));
 sg13g2_buf_8 fanout1047 (.A(net354),
    .X(net1047));
 sg13g2_buf_1 fanout1048 (.A(\DP_3.matrix[44] ),
    .X(net1048));
 sg13g2_buf_8 fanout1049 (.A(net1050),
    .X(net1049));
 sg13g2_buf_8 fanout1050 (.A(net302),
    .X(net1050));
 sg13g2_buf_8 fanout1051 (.A(net386),
    .X(net1051));
 sg13g2_buf_8 fanout1052 (.A(\DP_2.matrix[44] ),
    .X(net1052));
 sg13g2_buf_8 fanout1053 (.A(net527),
    .X(net1053));
 sg13g2_buf_8 fanout1054 (.A(net418),
    .X(net1054));
 sg13g2_buf_1 fanout1055 (.A(\DP_1.matrix[80] ),
    .X(net1055));
 sg13g2_buf_8 fanout1056 (.A(net362),
    .X(net1056));
 sg13g2_buf_1 fanout1057 (.A(\DP_1.matrix[44] ),
    .X(net1057));
 sg13g2_buf_8 fanout1058 (.A(\DP_1.matrix[8] ),
    .X(net1058));
 sg13g2_buf_1 fanout1059 (.A(\DP_1.matrix[8] ),
    .X(net1059));
 sg13g2_buf_8 fanout1060 (.A(net1068),
    .X(net1060));
 sg13g2_buf_8 fanout1061 (.A(net1068),
    .X(net1061));
 sg13g2_buf_8 fanout1062 (.A(net1064),
    .X(net1062));
 sg13g2_buf_8 fanout1063 (.A(net1064),
    .X(net1063));
 sg13g2_buf_8 fanout1064 (.A(net1068),
    .X(net1064));
 sg13g2_buf_8 fanout1065 (.A(net1066),
    .X(net1065));
 sg13g2_buf_8 fanout1066 (.A(net1067),
    .X(net1066));
 sg13g2_buf_8 fanout1067 (.A(net1068),
    .X(net1067));
 sg13g2_buf_8 fanout1068 (.A(net1087),
    .X(net1068));
 sg13g2_buf_8 fanout1069 (.A(net1072),
    .X(net1069));
 sg13g2_buf_8 fanout1070 (.A(net1072),
    .X(net1070));
 sg13g2_buf_8 fanout1071 (.A(net1072),
    .X(net1071));
 sg13g2_buf_8 fanout1072 (.A(net1087),
    .X(net1072));
 sg13g2_buf_8 fanout1073 (.A(net1074),
    .X(net1073));
 sg13g2_buf_8 fanout1074 (.A(net1087),
    .X(net1074));
 sg13g2_buf_8 fanout1075 (.A(net1076),
    .X(net1075));
 sg13g2_buf_8 fanout1076 (.A(net1080),
    .X(net1076));
 sg13g2_buf_8 fanout1077 (.A(net1079),
    .X(net1077));
 sg13g2_buf_2 fanout1078 (.A(net1079),
    .X(net1078));
 sg13g2_buf_8 fanout1079 (.A(net1080),
    .X(net1079));
 sg13g2_buf_8 fanout1080 (.A(net1086),
    .X(net1080));
 sg13g2_buf_8 fanout1081 (.A(net1082),
    .X(net1081));
 sg13g2_buf_8 fanout1082 (.A(net1085),
    .X(net1082));
 sg13g2_buf_8 fanout1083 (.A(net1085),
    .X(net1083));
 sg13g2_buf_8 fanout1084 (.A(net1085),
    .X(net1084));
 sg13g2_buf_8 fanout1085 (.A(net1086),
    .X(net1085));
 sg13g2_buf_8 fanout1086 (.A(net1087),
    .X(net1086));
 sg13g2_buf_8 fanout1087 (.A(net1148),
    .X(net1087));
 sg13g2_buf_8 fanout1088 (.A(net1108),
    .X(net1088));
 sg13g2_buf_8 fanout1089 (.A(net1108),
    .X(net1089));
 sg13g2_buf_8 fanout1090 (.A(net1093),
    .X(net1090));
 sg13g2_buf_8 fanout1091 (.A(net1093),
    .X(net1091));
 sg13g2_buf_8 fanout1092 (.A(net1093),
    .X(net1092));
 sg13g2_buf_8 fanout1093 (.A(net1095),
    .X(net1093));
 sg13g2_buf_8 fanout1094 (.A(net1095),
    .X(net1094));
 sg13g2_buf_8 fanout1095 (.A(net1108),
    .X(net1095));
 sg13g2_buf_8 fanout1096 (.A(net1099),
    .X(net1096));
 sg13g2_buf_8 fanout1097 (.A(net1099),
    .X(net1097));
 sg13g2_buf_8 fanout1098 (.A(net1099),
    .X(net1098));
 sg13g2_buf_8 fanout1099 (.A(net1107),
    .X(net1099));
 sg13g2_buf_8 fanout1100 (.A(net1102),
    .X(net1100));
 sg13g2_buf_8 fanout1101 (.A(net1102),
    .X(net1101));
 sg13g2_buf_8 fanout1102 (.A(net1107),
    .X(net1102));
 sg13g2_buf_8 fanout1103 (.A(net1106),
    .X(net1103));
 sg13g2_buf_8 fanout1104 (.A(net1106),
    .X(net1104));
 sg13g2_buf_8 fanout1105 (.A(net1106),
    .X(net1105));
 sg13g2_buf_8 fanout1106 (.A(net1107),
    .X(net1106));
 sg13g2_buf_8 fanout1107 (.A(net1108),
    .X(net1107));
 sg13g2_buf_8 fanout1108 (.A(net1148),
    .X(net1108));
 sg13g2_buf_8 fanout1109 (.A(net1113),
    .X(net1109));
 sg13g2_buf_1 fanout1110 (.A(net1113),
    .X(net1110));
 sg13g2_buf_8 fanout1111 (.A(net1113),
    .X(net1111));
 sg13g2_buf_8 fanout1112 (.A(net1113),
    .X(net1112));
 sg13g2_buf_8 fanout1113 (.A(net1130),
    .X(net1113));
 sg13g2_buf_8 fanout1114 (.A(net1115),
    .X(net1114));
 sg13g2_buf_8 fanout1115 (.A(net1130),
    .X(net1115));
 sg13g2_buf_8 fanout1116 (.A(net1119),
    .X(net1116));
 sg13g2_buf_8 fanout1117 (.A(net1119),
    .X(net1117));
 sg13g2_buf_8 fanout1118 (.A(net1119),
    .X(net1118));
 sg13g2_buf_8 fanout1119 (.A(net1130),
    .X(net1119));
 sg13g2_buf_8 fanout1120 (.A(net1121),
    .X(net1120));
 sg13g2_buf_8 fanout1121 (.A(net1130),
    .X(net1121));
 sg13g2_buf_8 fanout1122 (.A(net1125),
    .X(net1122));
 sg13g2_buf_1 fanout1123 (.A(net1125),
    .X(net1123));
 sg13g2_buf_8 fanout1124 (.A(net1125),
    .X(net1124));
 sg13g2_buf_8 fanout1125 (.A(net1130),
    .X(net1125));
 sg13g2_buf_8 fanout1126 (.A(net1128),
    .X(net1126));
 sg13g2_buf_8 fanout1127 (.A(net1128),
    .X(net1127));
 sg13g2_buf_8 fanout1128 (.A(net1129),
    .X(net1128));
 sg13g2_buf_8 fanout1129 (.A(net1130),
    .X(net1129));
 sg13g2_buf_8 fanout1130 (.A(net1148),
    .X(net1130));
 sg13g2_buf_8 fanout1131 (.A(net1132),
    .X(net1131));
 sg13g2_buf_8 fanout1132 (.A(net1147),
    .X(net1132));
 sg13g2_buf_8 fanout1133 (.A(net1135),
    .X(net1133));
 sg13g2_buf_1 fanout1134 (.A(net1135),
    .X(net1134));
 sg13g2_buf_8 fanout1135 (.A(net1147),
    .X(net1135));
 sg13g2_buf_8 fanout1136 (.A(net1137),
    .X(net1136));
 sg13g2_buf_8 fanout1137 (.A(net1138),
    .X(net1137));
 sg13g2_buf_8 fanout1138 (.A(net1147),
    .X(net1138));
 sg13g2_buf_8 fanout1139 (.A(net1146),
    .X(net1139));
 sg13g2_buf_8 fanout1140 (.A(net1144),
    .X(net1140));
 sg13g2_buf_8 fanout1141 (.A(net1144),
    .X(net1141));
 sg13g2_buf_8 fanout1142 (.A(net1143),
    .X(net1142));
 sg13g2_buf_8 fanout1143 (.A(net1144),
    .X(net1143));
 sg13g2_buf_8 fanout1144 (.A(net1146),
    .X(net1144));
 sg13g2_buf_8 fanout1145 (.A(net1146),
    .X(net1145));
 sg13g2_buf_8 fanout1146 (.A(net1147),
    .X(net1146));
 sg13g2_buf_8 fanout1147 (.A(net1148),
    .X(net1147));
 sg13g2_buf_8 fanout1148 (.A(rst_n),
    .X(net1148));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[7]),
    .X(net16));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[0]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[1]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_out[2]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_out[3]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uio_out[4]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uio_out[5]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uio_out[6]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uio_out[7]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[0]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[1]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uo_out[2]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uo_out[3]));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uo_out[4]));
 sg13g2_buf_1 output30 (.A(net30),
    .X(uo_out[5]));
 sg13g2_buf_1 output31 (.A(net31),
    .X(uo_out[6]));
 sg13g2_buf_1 output32 (.A(net32),
    .X(uo_out[7]));
 sg13g2_tiehi heichips25_template_33 (.L_HI(net33));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_4_5_0_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_4_6_0_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_4_7_0_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_4_9_0_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_4_10_0_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_4_11_0_clk));
 sg13g2_buf_8 clkload9 (.A(clknet_4_13_0_clk));
 sg13g2_buf_8 clkload10 (.A(clknet_4_14_0_clk));
 sg13g2_buf_8 clkload11 (.A(clknet_4_15_0_clk));
 sg13g2_inv_4 clkload12 (.A(clknet_leaf_67_clk));
 sg13g2_buf_8 clkload13 (.A(clknet_leaf_65_clk));
 sg13g2_buf_8 clkload14 (.A(clknet_leaf_24_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_47_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_60_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_51_clk));
 sg13g2_inv_4 clkload18 (.A(clknet_leaf_50_clk));
 sg13g2_inv_4 clkload19 (.A(clknet_leaf_37_clk));
 sg13g2_buf_8 clkload20 (.A(clknet_leaf_44_clk));
 sg13g2_inv_2 clkload21 (.A(clknet_leaf_45_clk));
 sg13g2_inv_2 clkload22 (.A(clknet_leaf_34_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\mac2.sum_lvl1_ff[46] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold2 (.A(\mac1.sum_lvl1_ff[47] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold3 (.A(\mac1.products_ff[138] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold4 (.A(\mac2.sum_lvl1_ff[87] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold5 (.A(\mac2.products_ff[82] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold6 (.A(\mac1.sum_lvl1_ff[10] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold7 (.A(\mac2.sum_lvl1_ff[78] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold8 (.A(\mac1.sum_lvl1_ff[77] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold9 (.A(\mac2.products_ff[68] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold10 (.A(\mac2.sum_lvl2_ff[50] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold11 (.A(\mac2.sum_lvl1_ff[81] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold12 (.A(\mac1.sum_lvl1_ff[42] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold13 (.A(\mac2.sum_lvl1_ff[43] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold14 (.A(\mac1.products_ff[70] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold15 (.A(\mac2.sum_lvl1_ff[45] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold16 (.A(\mac1.sum_lvl1_ff[15] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold17 (.A(\mac1.products_ff[147] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold18 (.A(\mac1.sum_lvl1_ff[14] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold19 (.A(\mac1.sum_lvl1_ff[1] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold20 (.A(\mac2.products_ff[142] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold21 (.A(\mac2.products_ff[137] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold22 (.A(\mac1.sum_lvl1_ff[3] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold23 (.A(\mac1.products_ff[79] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold24 (.A(\mac2.sum_lvl1_ff[80] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold25 (.A(\mac2.sum_lvl1_ff[1] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold26 (.A(\mac2.sum_lvl1_ff[36] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold27 (.A(\mac2.products_ff[138] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold28 (.A(\mac1.sum_lvl1_ff[38] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold29 (.A(\mac2.sum_lvl1_ff[83] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold30 (.A(\mac2.products_ff[15] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold31 (.A(\mac1.products_ff[12] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold32 (.A(\mac1.products_ff[72] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold33 (.A(\mac1.sum_lvl1_ff[6] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold34 (.A(\mac1.products_ff[9] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold35 (.A(\mac2.sum_lvl1_ff[51] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold36 (.A(\mac2.sum_lvl2_ff[41] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold37 (.A(\mac1.products_ff[8] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold38 (.A(\mac1.sum_lvl1_ff[37] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold39 (.A(\mac1.sum_lvl1_ff[87] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold40 (.A(\mac2.products_ff[10] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold41 (.A(\mac1.products_ff[7] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold42 (.A(\mac2.sum_lvl1_ff[6] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold43 (.A(\mac2.products_ff[9] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold44 (.A(\mac2.products_ff[11] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold45 (.A(\mac2.sum_lvl2_ff[45] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold46 (.A(\mac1.products_ff[5] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold47 (.A(\mac1.sum_lvl2_ff[52] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold48 (.A(\mac1.sum_lvl1_ff[4] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold49 (.A(\mac2.sum_lvl1_ff[48] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold50 (.A(\mac1.products_ff[143] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold51 (.A(\mac1.products_ff[136] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold52 (.A(\mac2.sum_lvl2_ff[52] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold53 (.A(\mac2.sum_lvl1_ff[79] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold54 (.A(\mac2.sum_lvl1_ff[84] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold55 (.A(\mac1.products_ff[137] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold56 (.A(\mac1.products_ff[3] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold57 (.A(\mac2.sum_lvl2_ff[42] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold58 (.A(\mac1.products_ff[83] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold59 (.A(\mac1.sum_lvl1_ff[49] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold60 (.A(\mac2.sum_lvl1_ff[0] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold61 (.A(\mac2.sum_lvl2_ff[48] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold62 (.A(\mac1.sum_lvl1_ff[83] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold63 (.A(\mac1.products_ff[2] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold64 (.A(\mac1.sum_lvl2_ff[50] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold65 (.A(\mac2.sum_lvl2_ff[51] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold66 (.A(\mac2.sum_lvl1_ff[82] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold67 (.A(\mac1.products_ff[0] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold68 (.A(\mac2.products_ff[147] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold69 (.A(\mac1.sum_lvl1_ff[82] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold70 (.A(\mac2.products_ff[80] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold71 (.A(\mac2.sum_lvl1_ff[47] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold72 (.A(\mac2.sum_lvl1_ff[77] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold73 (.A(\mac2.sum_lvl2_ff[44] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold74 (.A(\mac2.products_ff[75] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold75 (.A(\mac2.sum_lvl2_ff[43] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold76 (.A(\mac2.sum_lvl2_ff[38] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold77 (.A(\mac2.sum_lvl1_ff[14] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold78 (.A(\mac2.sum_lvl2_ff[49] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold79 (.A(\mac1.sum_lvl2_ff[39] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold80 (.A(\mac1.products_ff[71] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold81 (.A(\mac2.products_ff[145] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold82 (.A(\mac2.sum_lvl1_ff[37] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold83 (.A(\mac2.sum_lvl2_ff[39] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold84 (.A(\mac1.products_ff[78] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold85 (.A(\mac1.sum_lvl2_ff[49] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold86 (.A(\mac1.products_ff[139] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold87 (.A(\mac1.sum_lvl1_ff[5] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold88 (.A(\mac2.products_ff[141] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold89 (.A(\mac1.sum_lvl2_ff[40] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold90 (.A(\mac2.products_ff[14] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold91 (.A(\mac2.products_ff[74] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold92 (.A(\mac2.sum_lvl1_ff[49] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold93 (.A(\mac2.products_ff[4] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold94 (.A(\mac1.products_ff[11] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold95 (.A(\mac1.products_ff[141] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold96 (.A(\mac1.sum_lvl2_ff[42] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold97 (.A(\mac2.sum_lvl1_ff[15] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold98 (.A(\mac1.sum_lvl1_ff[81] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold99 (.A(\mac1.sum_lvl1_ff[44] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold100 (.A(\mac2.products_ff[144] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold101 (.A(\mac2.sum_lvl1_ff[50] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold102 (.A(\mac1.sum_lvl1_ff[0] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold103 (.A(\mac1.sum_lvl2_ff[53] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold104 (.A(\mac2.products_ff[139] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold105 (.A(\mac2.products_ff[136] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold106 (.A(\mac1.products_ff[75] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold107 (.A(\mac1.sum_lvl1_ff[39] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold108 (.A(\mac1.sum_lvl1_ff[48] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold109 (.A(\mac1.products_ff[6] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold110 (.A(\mac1.sum_lvl1_ff[74] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold111 (.A(\mac1.products_ff[13] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold112 (.A(\mac2.sum_lvl1_ff[74] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold113 (.A(\mac2.products_ff[140] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold114 (.A(\mac2.products_ff[70] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold115 (.A(\mac1.products_ff[146] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold116 (.A(\mac1.sum_lvl1_ff[8] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold117 (.A(\mac1.sum_lvl1_ff[75] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold118 (.A(\mac2.sum_lvl1_ff[2] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold119 (.A(\mac1.sum_lvl1_ff[78] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold120 (.A(\mac2.products_ff[7] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold121 (.A(\mac1.sum_lvl2_ff[41] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold122 (.A(\mac2.sum_lvl2_ff[47] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold123 (.A(\mac2.sum_lvl1_ff[73] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold124 (.A(\mac1.sum_lvl1_ff[72] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold125 (.A(\mac2.sum_lvl1_ff[75] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold126 (.A(\mac1.sum_lvl1_ff[85] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold127 (.A(\mac2.sum_lvl2_ff[53] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold128 (.A(\mac1.sum_lvl1_ff[7] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold129 (.A(\mac2.products_ff[2] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold130 (.A(\mac1.sum_lvl2_ff[38] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold131 (.A(\mac2.sum_lvl1_ff[76] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold132 (.A(\mac2.products_ff[151] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold133 (.A(\mac2.sum_lvl1_ff[40] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold134 (.A(\mac1.sum_lvl2_ff[46] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold135 (.A(\mac1.products_ff[76] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold136 (.A(\mac1.products_ff[144] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold137 (.A(\mac1.products_ff[82] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold138 (.A(\mac2.products_ff[81] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold139 (.A(\mac2.products_ff[3] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold140 (.A(\mac2.sum_lvl1_ff[42] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold141 (.A(\mac1.products_ff[15] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold142 (.A(\mac1.sum_lvl1_ff[9] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold143 (.A(\mac1.products_ff[4] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold144 (.A(\mac2.products_ff[73] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold145 (.A(\mac2.products_ff[0] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold146 (.A(\mac1.sum_lvl2_ff[47] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold147 (.A(\mac1.sum_lvl2_ff[48] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold148 (.A(\mac1.sum_lvl1_ff[50] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold149 (.A(\mac1.products_ff[74] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold150 (.A(\mac2.sum_lvl1_ff[72] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold151 (.A(\mac2.sum_lvl1_ff[44] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold152 (.A(\mac1.products_ff[149] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold153 (.A(\mac1.sum_lvl2_ff[43] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold154 (.A(\mac2.sum_lvl1_ff[86] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold155 (.A(\mac2.sum_lvl2_ff[40] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold156 (.A(\mac2.products_ff[143] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold157 (.A(\mac1.sum_lvl1_ff[13] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold158 (.A(\mac2.sum_lvl1_ff[4] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold159 (.A(\mac2.products_ff[76] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold160 (.A(\mac1.products_ff[14] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold161 (.A(\mac1.products_ff[142] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold162 (.A(\mac2.sum_lvl1_ff[85] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold163 (.A(\mac2.sum_lvl1_ff[39] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold164 (.A(\mac1.sum_lvl1_ff[12] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold165 (.A(\mac2.sum_lvl2_ff[46] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold166 (.A(\mac1.sum_lvl1_ff[45] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold167 (.A(\mac1.products_ff[140] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold168 (.A(\mac1.sum_lvl1_ff[51] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold169 (.A(\mac1.sum_lvl2_ff[45] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold170 (.A(\mac2.sum_lvl1_ff[38] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold171 (.A(\mac1.sum_lvl1_ff[41] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold172 (.A(\mac1.sum_lvl1_ff[36] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold173 (.A(\mac1.sum_lvl2_ff[51] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold174 (.A(\mac2.products_ff[72] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold175 (.A(\mac1.sum_lvl1_ff[73] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold176 (.A(\mac1.sum_lvl2_ff[44] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold177 (.A(\mac1.products_ff[69] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold178 (.A(\mac2.products_ff[69] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold179 (.A(\mac1.products_ff[1] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold180 (.A(\mac2.products_ff[1] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold181 (.A(\mac2.sum_lvl1_ff[7] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold182 (.A(\mac2.sum_lvl1_ff[3] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold183 (.A(\mac1.products_ff[150] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold184 (.A(\mac2.products_ff[79] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold185 (.A(\mac2.products_ff[12] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold186 (.A(\mac1.sum_lvl1_ff[11] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold187 (.A(\mac2.sum_lvl1_ff[5] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold188 (.A(\mac1.products_ff[145] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold189 (.A(\mac1.sum_lvl1_ff[86] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold190 (.A(\mac1.products_ff[80] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold191 (.A(\mac2.sum_lvl1_ff[41] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold192 (.A(\mac2.products_ff[148] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold193 (.A(\mac2.products_ff[150] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold194 (.A(\mac1.sum_lvl1_ff[2] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold195 (.A(\mac2.products_ff[8] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold196 (.A(\mac2.products_ff[146] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold197 (.A(\mac1.products_ff[73] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold198 (.A(\mac2.products_ff[71] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold199 (.A(\mac1.products_ff[68] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold200 (.A(\mac2.products_ff[83] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold201 (.A(\mac1.products_ff[77] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold202 (.A(\mac2.products_ff[13] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold203 (.A(\mac1.sum_lvl1_ff[80] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold204 (.A(\mac1.sum_lvl1_ff[79] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold205 (.A(\mac2.products_ff[78] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold206 (.A(\mac1.products_ff[10] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold207 (.A(\mac2.sum_lvl1_ff[8] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold208 (.A(\mac1.sum_lvl1_ff[84] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold209 (.A(\mac2.products_ff[5] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold210 (.A(\mac2.sum_lvl1_ff[13] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold211 (.A(\mac2.sum_lvl1_ff[12] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold212 (.A(\mac2.products_ff[77] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold213 (.A(\mac1.products_ff[81] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold214 (.A(\mac1.sum_lvl1_ff[76] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold215 (.A(\mac1.sum_lvl1_ff[40] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold216 (.A(\mac2.sum_lvl1_ff[11] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold217 (.A(\mac2.sum_lvl1_ff[10] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold218 (.A(\mac2.products_ff[149] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold219 (.A(\mac2.sum_lvl1_ff[9] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold220 (.A(\mac1.sum_lvl1_ff[43] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold221 (.A(\mac2.products_ff[6] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold222 (.A(\mac1.sum_lvl1_ff[46] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold223 (.A(\mac1.products_ff[148] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold224 (.A(\mac1.products_ff[151] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold225 (.A(\mac1.sum_lvl3_ff[0] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0016_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold227 (.A(\mac1.sum_lvl2_ff[0] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0000_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold229 (.A(\DP_4.matrix[76] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold230 (.A(\DP_4.matrix[75] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold231 (.A(\mac2.sum_lvl2_ff[0] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0032_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold233 (.A(\DP_3.matrix[80] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold234 (.A(\DP_2.matrix[44] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold235 (.A(\DP_3.matrix[72] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold236 (.A(\DP_3.matrix[79] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold237 (.A(\DP_3.matrix[77] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold238 (.A(\DP_4.matrix[80] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold239 (.A(\DP_3.matrix[78] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold240 (.A(\DP_1.matrix[7] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0179_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold242 (.A(\DP_1.matrix[5] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0177_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold244 (.A(\mac1.sum_lvl2_ff[15] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold245 (.A(_2157_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0006_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold247 (.A(\mac1.sum_lvl2_ff[19] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0007_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold249 (.A(\mac1.sum_lvl3_ff[15] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold250 (.A(_2214_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0022_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold252 (.A(\mac1.sum_lvl3_ff[20] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0023_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold254 (.A(\mac1.sum_lvl2_ff[5] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold255 (.A(_2117_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0011_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold257 (.A(\mac2.sum_lvl3_ff[14] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold258 (.A(_2325_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold259 (.A(_0053_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold260 (.A(\DP_2.matrix[43] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold261 (.A(\DP_3.matrix[75] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold262 (.A(\DP_3.matrix[8] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold263 (.A(\mac1.sum_lvl2_ff[14] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold264 (.A(_2155_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold265 (.A(_0005_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold266 (.A(\DP_2.matrix[38] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold267 (.A(\DP_3.matrix[74] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold268 (.A(\mac2.sum_lvl2_ff[19] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0039_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold270 (.A(\DP_3.matrix[73] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold271 (.A(\DP_2.matrix[77] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold272 (.A(\DP_1.matrix[39] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold273 (.A(\DP_1.matrix[40] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold274 (.A(\DP_1.matrix[75] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold275 (.A(\mac2.sum_lvl3_ff[9] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold276 (.A(_2302_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0063_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold278 (.A(\DP_4.matrix[77] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold279 (.A(\mac1.sum_lvl2_ff[12] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold280 (.A(_2144_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0003_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold282 (.A(\DP_2.matrix[0] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold283 (.A(\DP_1.matrix[41] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold284 (.A(\DP_4.matrix[79] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold285 (.A(\mac2.sum_lvl3_ff[0] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0048_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold287 (.A(\DP_4.matrix[8] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold288 (.A(\DP_1.matrix[36] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold289 (.A(\DP_4.matrix[38] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold290 (.A(\DP_4.matrix[40] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold291 (.A(\mac1.sum_lvl3_ff[14] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold292 (.A(_2212_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0021_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold294 (.A(\DP_4.matrix[43] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold295 (.A(\DP_4.matrix[42] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold296 (.A(\DP_1.matrix[0] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold297 (.A(\DP_3.matrix[40] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold298 (.A(\DP_3.matrix[37] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold299 (.A(\DP_3.matrix[38] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold300 (.A(\mac1.sum_lvl2_ff[4] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold301 (.A(_2114_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0010_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold303 (.A(\DP_4.matrix[36] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold304 (.A(\DP_4.matrix[44] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold305 (.A(\DP_3.matrix[6] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold306 (.A(\mac2.sum_lvl3_ff[10] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold307 (.A(_2306_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0049_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold309 (.A(\DP_3.matrix[36] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold310 (.A(\mac2.sum_lvl2_ff[2] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold311 (.A(_2221_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0040_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold313 (.A(\DP_3.matrix[76] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold314 (.A(\DP_3.matrix[44] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold315 (.A(\DP_3.matrix[0] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold316 (.A(\DP_3.matrix[41] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold317 (.A(\DP_4.matrix[6] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold318 (.A(_0250_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold319 (.A(\mac2.sum_lvl3_ff[5] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold320 (.A(_2286_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold321 (.A(_0059_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold322 (.A(\DP_1.matrix[44] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold323 (.A(\DP_2.matrix[36] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold324 (.A(\DP_4.matrix[41] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold325 (.A(\mac1.sum_lvl2_ff[29] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold326 (.A(_2134_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold327 (.A(_2141_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold328 (.A(_0002_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold329 (.A(\DP_1.matrix[42] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold330 (.A(\DP_4.matrix[74] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold331 (.A(\DP_4.matrix[4] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0248_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold333 (.A(\DP_4.matrix[37] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold334 (.A(\DP_4.matrix[0] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0244_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold336 (.A(\DP_4.matrix[72] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold337 (.A(\DP_2.matrix[7] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold338 (.A(_0203_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold339 (.A(\DP_4.matrix[2] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0246_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold341 (.A(\mac1.sum_lvl3_ff[2] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold342 (.A(_2164_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold343 (.A(_0024_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold344 (.A(\DP_4.matrix[3] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0247_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold346 (.A(\DP_2.matrix[80] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold347 (.A(\DP_3.matrix[3] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0223_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold349 (.A(\mac1.sum_lvl2_ff[2] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold350 (.A(_2108_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0008_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold352 (.A(\mac1.sum_lvl2_ff[8] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold353 (.A(_2127_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold354 (.A(_2128_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0014_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold356 (.A(\DP_1.matrix[4] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0176_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold358 (.A(\DP_4.matrix[39] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold359 (.A(\DP_1.matrix[43] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold360 (.A(\DP_2.matrix[41] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold361 (.A(\mac2.sum_lvl3_ff[30] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold362 (.A(_2311_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold363 (.A(_0050_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold364 (.A(\DP_2.matrix[76] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold365 (.A(\DP_4.matrix[7] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold366 (.A(\DP_2.matrix[3] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0199_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold368 (.A(\DP_1.matrix[6] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold369 (.A(_0178_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold370 (.A(\mac2.sum_lvl3_ff[13] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold371 (.A(_2319_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold372 (.A(_2320_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0052_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold374 (.A(\DP_2.matrix[4] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold375 (.A(\DP_2.matrix[42] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold376 (.A(\DP_2.matrix[6] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold377 (.A(_0202_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold378 (.A(\DP_1.matrix[80] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold379 (.A(\DP_4.matrix[78] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold380 (.A(\DP_3.matrix[4] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold381 (.A(_0224_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold382 (.A(\DP_3.matrix[1] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold383 (.A(_0221_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold384 (.A(\DP_1.matrix[72] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold385 (.A(\DP_1.matrix[2] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold386 (.A(\DP_2.matrix[78] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold387 (.A(\mac1.sum_lvl3_ff[13] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold388 (.A(_2206_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold389 (.A(_2207_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold390 (.A(_0020_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold391 (.A(\DP_2.matrix[39] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold392 (.A(\mac2.sum_lvl2_ff[3] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold393 (.A(_2224_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold394 (.A(_0041_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold395 (.A(\DP_3.matrix[2] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold396 (.A(_0222_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold397 (.A(\mac2.sum_lvl3_ff[35] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold398 (.A(_2327_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0054_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold400 (.A(\DP_2.matrix[2] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold401 (.A(\mac1.sum_lvl3_ff[3] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold402 (.A(_2167_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold403 (.A(_0025_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold404 (.A(\mac2.sum_lvl3_ff[4] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold405 (.A(_2283_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold406 (.A(_0058_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold407 (.A(\DP_3.matrix[5] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold408 (.A(\DP_1.matrix[37] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold409 (.A(_0617_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold410 (.A(\DP_4.matrix[5] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold411 (.A(\DP_3.matrix[7] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold412 (.A(\DP_2.matrix[40] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold413 (.A(\DP_1.matrix[3] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold414 (.A(\mac2.sum_lvl3_ff[27] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold415 (.A(_2292_),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold416 (.A(_2299_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold417 (.A(_0062_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold418 (.A(\mac1.sum_lvl2_ff[27] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold419 (.A(_0015_),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold420 (.A(\DP_2.matrix[5] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold421 (.A(\mac1.sum_lvl2_ff[6] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold422 (.A(_2119_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold423 (.A(_2122_),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold424 (.A(_0012_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold425 (.A(\mac1.sum_lvl2_ff[13] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold426 (.A(_2150_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold427 (.A(_2151_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold428 (.A(_0004_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold429 (.A(\mac2.sum_lvl2_ff[5] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold430 (.A(_2230_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold431 (.A(_0043_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold432 (.A(\DP_2.matrix[1] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold433 (.A(\DP_4.matrix[73] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold434 (.A(\DP_4.matrix[1] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold435 (.A(\mac1.sum_lvl2_ff[3] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold436 (.A(_2111_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold437 (.A(_0009_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold438 (.A(\mac1.sum_lvl2_ff[10] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold439 (.A(_0001_),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold440 (.A(\mac2.sum_lvl3_ff[20] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold441 (.A(_0055_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold442 (.A(\DP_2.matrix[74] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold443 (.A(\DP_3.matrix[39] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold444 (.A(\mac2.sum_lvl2_ff[15] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold445 (.A(_2270_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold446 (.A(_0038_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold447 (.A(\mac2.sum_lvl3_ff[26] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold448 (.A(_2288_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold449 (.A(_2291_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold450 (.A(_0060_),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold451 (.A(\DP_2.matrix[72] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold452 (.A(\DP_1.matrix[74] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold453 (.A(\DP_1.matrix[38] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold454 (.A(\mac1.sum_lvl3_ff[8] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold455 (.A(_2184_),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold456 (.A(_2185_),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold457 (.A(_0030_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold458 (.A(\mac2.sum_lvl3_ff[2] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold459 (.A(_2277_),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold460 (.A(_0056_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold461 (.A(\mac2.sum_lvl3_ff[3] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold462 (.A(_2280_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold463 (.A(_0057_),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold464 (.A(\DP_1.matrix[1] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold465 (.A(\DP_3.Q_range.out_data[4] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold466 (.A(_2473_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold467 (.A(_2475_),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold468 (.A(_0245_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold469 (.A(\mac1.sum_lvl3_ff[9] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold470 (.A(_2189_),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold471 (.A(_0031_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold472 (.A(\mac2.sum_lvl2_ff[4] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold473 (.A(_2227_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold474 (.A(_0042_),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold475 (.A(\DP_1.matrix[73] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold476 (.A(_2637_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold477 (.A(\mac2.sum_lvl2_ff[8] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold478 (.A(_2240_),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold479 (.A(_2241_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold480 (.A(_0046_),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold481 (.A(\mac1.sum_lvl3_ff[10] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold482 (.A(_2193_),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold483 (.A(\DP_2.matrix[79] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold484 (.A(\DP_2.matrix[37] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold485 (.A(\mac1.sum_lvl3_ff[30] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold486 (.A(_0018_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold487 (.A(\DP_2.matrix[8] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold488 (.A(\DP_1.matrix[76] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold489 (.A(\DP_3.matrix[43] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold490 (.A(\mac2.sum_lvl3_ff[12] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold491 (.A(_2313_),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold492 (.A(\mac1.sum_lvl3_ff[6] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold493 (.A(_2175_),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold494 (.A(_2178_),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold495 (.A(\mac1.sum_lvl2_ff[7] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold496 (.A(_2124_),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold497 (.A(_2125_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold498 (.A(_0013_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold499 (.A(\DP_3.matrix[42] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold500 (.A(\mac1.sum_lvl3_ff[12] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold501 (.A(_2200_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold502 (.A(\DP_1.matrix[77] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold503 (.A(\DP_2.matrix[73] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold504 (.A(\DP_1.matrix[78] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold505 (.A(\mac2.sum_lvl3_ff[7] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold506 (.A(\mac1.sum_lvl3_ff[5] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold507 (.A(_2173_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold508 (.A(\mac2.sum_lvl2_ff[24] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold509 (.A(_2235_),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold510 (.A(\DP_2.matrix[75] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold511 (.A(\mac1.sum_lvl3_ff[4] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold512 (.A(\mac2.sum_lvl2_ff[14] ),
    .X(net552));
 sg13g2_fill_2 FILLER_0_0 ();
 sg13g2_fill_1 FILLER_0_2 ();
 sg13g2_fill_2 FILLER_0_155 ();
 sg13g2_fill_1 FILLER_0_157 ();
 sg13g2_fill_1 FILLER_0_163 ();
 sg13g2_fill_1 FILLER_0_173 ();
 sg13g2_fill_1 FILLER_0_191 ();
 sg13g2_fill_2 FILLER_0_197 ();
 sg13g2_fill_1 FILLER_0_199 ();
 sg13g2_fill_1 FILLER_0_205 ();
 sg13g2_fill_1 FILLER_0_225 ();
 sg13g2_decap_8 FILLER_0_263 ();
 sg13g2_decap_8 FILLER_0_270 ();
 sg13g2_fill_2 FILLER_0_277 ();
 sg13g2_fill_1 FILLER_0_279 ();
 sg13g2_fill_1 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_369 ();
 sg13g2_fill_2 FILLER_0_403 ();
 sg13g2_fill_2 FILLER_0_445 ();
 sg13g2_decap_8 FILLER_0_452 ();
 sg13g2_decap_8 FILLER_0_459 ();
 sg13g2_decap_8 FILLER_0_466 ();
 sg13g2_fill_2 FILLER_0_473 ();
 sg13g2_fill_1 FILLER_0_488 ();
 sg13g2_fill_2 FILLER_0_569 ();
 sg13g2_fill_1 FILLER_0_612 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_fill_2 FILLER_0_714 ();
 sg13g2_fill_1 FILLER_0_716 ();
 sg13g2_decap_8 FILLER_0_722 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_decap_8 FILLER_0_875 ();
 sg13g2_decap_8 FILLER_0_882 ();
 sg13g2_decap_8 FILLER_0_889 ();
 sg13g2_decap_8 FILLER_0_896 ();
 sg13g2_decap_8 FILLER_0_903 ();
 sg13g2_decap_8 FILLER_0_910 ();
 sg13g2_decap_8 FILLER_0_917 ();
 sg13g2_decap_8 FILLER_0_924 ();
 sg13g2_decap_8 FILLER_0_931 ();
 sg13g2_decap_8 FILLER_0_938 ();
 sg13g2_decap_8 FILLER_0_945 ();
 sg13g2_decap_8 FILLER_0_952 ();
 sg13g2_decap_8 FILLER_0_959 ();
 sg13g2_decap_8 FILLER_0_966 ();
 sg13g2_decap_8 FILLER_0_973 ();
 sg13g2_decap_8 FILLER_0_980 ();
 sg13g2_decap_8 FILLER_0_987 ();
 sg13g2_decap_8 FILLER_0_994 ();
 sg13g2_decap_8 FILLER_0_1001 ();
 sg13g2_decap_8 FILLER_0_1008 ();
 sg13g2_decap_8 FILLER_0_1015 ();
 sg13g2_decap_8 FILLER_0_1022 ();
 sg13g2_fill_2 FILLER_1_27 ();
 sg13g2_fill_1 FILLER_1_29 ();
 sg13g2_fill_1 FILLER_1_179 ();
 sg13g2_fill_2 FILLER_1_220 ();
 sg13g2_fill_1 FILLER_1_222 ();
 sg13g2_decap_4 FILLER_1_231 ();
 sg13g2_decap_4 FILLER_1_250 ();
 sg13g2_fill_1 FILLER_1_270 ();
 sg13g2_fill_2 FILLER_1_361 ();
 sg13g2_fill_2 FILLER_1_520 ();
 sg13g2_fill_1 FILLER_1_522 ();
 sg13g2_fill_2 FILLER_1_550 ();
 sg13g2_fill_2 FILLER_1_678 ();
 sg13g2_fill_2 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_767 ();
 sg13g2_decap_8 FILLER_1_774 ();
 sg13g2_decap_8 FILLER_1_781 ();
 sg13g2_decap_8 FILLER_1_788 ();
 sg13g2_decap_8 FILLER_1_795 ();
 sg13g2_decap_8 FILLER_1_802 ();
 sg13g2_decap_8 FILLER_1_809 ();
 sg13g2_decap_8 FILLER_1_816 ();
 sg13g2_decap_8 FILLER_1_823 ();
 sg13g2_decap_8 FILLER_1_830 ();
 sg13g2_decap_8 FILLER_1_837 ();
 sg13g2_decap_8 FILLER_1_844 ();
 sg13g2_decap_8 FILLER_1_851 ();
 sg13g2_decap_8 FILLER_1_858 ();
 sg13g2_decap_8 FILLER_1_865 ();
 sg13g2_decap_8 FILLER_1_872 ();
 sg13g2_decap_8 FILLER_1_879 ();
 sg13g2_decap_8 FILLER_1_886 ();
 sg13g2_decap_8 FILLER_1_893 ();
 sg13g2_decap_8 FILLER_1_900 ();
 sg13g2_decap_8 FILLER_1_907 ();
 sg13g2_decap_8 FILLER_1_914 ();
 sg13g2_decap_8 FILLER_1_921 ();
 sg13g2_decap_8 FILLER_1_928 ();
 sg13g2_decap_8 FILLER_1_935 ();
 sg13g2_decap_8 FILLER_1_942 ();
 sg13g2_decap_8 FILLER_1_949 ();
 sg13g2_decap_8 FILLER_1_956 ();
 sg13g2_decap_8 FILLER_1_963 ();
 sg13g2_decap_8 FILLER_1_970 ();
 sg13g2_decap_8 FILLER_1_977 ();
 sg13g2_decap_8 FILLER_1_984 ();
 sg13g2_decap_8 FILLER_1_991 ();
 sg13g2_decap_8 FILLER_1_998 ();
 sg13g2_decap_8 FILLER_1_1005 ();
 sg13g2_decap_8 FILLER_1_1012 ();
 sg13g2_decap_8 FILLER_1_1019 ();
 sg13g2_fill_2 FILLER_1_1026 ();
 sg13g2_fill_1 FILLER_1_1028 ();
 sg13g2_fill_1 FILLER_2_0 ();
 sg13g2_fill_2 FILLER_2_68 ();
 sg13g2_fill_1 FILLER_2_151 ();
 sg13g2_fill_2 FILLER_2_167 ();
 sg13g2_fill_2 FILLER_2_214 ();
 sg13g2_fill_1 FILLER_2_216 ();
 sg13g2_fill_2 FILLER_2_270 ();
 sg13g2_fill_2 FILLER_2_299 ();
 sg13g2_fill_2 FILLER_2_318 ();
 sg13g2_fill_2 FILLER_2_395 ();
 sg13g2_fill_1 FILLER_2_513 ();
 sg13g2_fill_1 FILLER_2_567 ();
 sg13g2_fill_1 FILLER_2_609 ();
 sg13g2_fill_1 FILLER_2_637 ();
 sg13g2_fill_1 FILLER_2_671 ();
 sg13g2_fill_1 FILLER_2_752 ();
 sg13g2_decap_8 FILLER_2_780 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_decap_8 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_2_868 ();
 sg13g2_decap_8 FILLER_2_875 ();
 sg13g2_decap_8 FILLER_2_882 ();
 sg13g2_decap_8 FILLER_2_889 ();
 sg13g2_decap_8 FILLER_2_896 ();
 sg13g2_decap_8 FILLER_2_903 ();
 sg13g2_decap_8 FILLER_2_910 ();
 sg13g2_decap_8 FILLER_2_917 ();
 sg13g2_decap_8 FILLER_2_924 ();
 sg13g2_decap_8 FILLER_2_931 ();
 sg13g2_decap_8 FILLER_2_938 ();
 sg13g2_decap_8 FILLER_2_945 ();
 sg13g2_decap_8 FILLER_2_952 ();
 sg13g2_decap_8 FILLER_2_959 ();
 sg13g2_decap_8 FILLER_2_966 ();
 sg13g2_decap_8 FILLER_2_973 ();
 sg13g2_decap_8 FILLER_2_980 ();
 sg13g2_decap_8 FILLER_2_987 ();
 sg13g2_decap_8 FILLER_2_994 ();
 sg13g2_decap_8 FILLER_2_1001 ();
 sg13g2_decap_8 FILLER_2_1008 ();
 sg13g2_decap_8 FILLER_2_1015 ();
 sg13g2_decap_8 FILLER_2_1022 ();
 sg13g2_fill_1 FILLER_3_0 ();
 sg13g2_fill_2 FILLER_3_82 ();
 sg13g2_fill_1 FILLER_3_84 ();
 sg13g2_fill_2 FILLER_3_120 ();
 sg13g2_fill_1 FILLER_3_131 ();
 sg13g2_fill_2 FILLER_3_137 ();
 sg13g2_fill_1 FILLER_3_158 ();
 sg13g2_fill_2 FILLER_3_173 ();
 sg13g2_fill_1 FILLER_3_175 ();
 sg13g2_fill_2 FILLER_3_204 ();
 sg13g2_fill_1 FILLER_3_206 ();
 sg13g2_fill_2 FILLER_3_212 ();
 sg13g2_decap_8 FILLER_3_219 ();
 sg13g2_decap_4 FILLER_3_262 ();
 sg13g2_fill_2 FILLER_3_266 ();
 sg13g2_fill_1 FILLER_3_397 ();
 sg13g2_fill_1 FILLER_3_433 ();
 sg13g2_fill_2 FILLER_3_450 ();
 sg13g2_fill_1 FILLER_3_481 ();
 sg13g2_fill_2 FILLER_3_536 ();
 sg13g2_fill_1 FILLER_3_538 ();
 sg13g2_fill_2 FILLER_3_596 ();
 sg13g2_fill_1 FILLER_3_598 ();
 sg13g2_fill_2 FILLER_3_608 ();
 sg13g2_fill_2 FILLER_3_677 ();
 sg13g2_fill_2 FILLER_3_704 ();
 sg13g2_fill_1 FILLER_3_714 ();
 sg13g2_fill_2 FILLER_3_773 ();
 sg13g2_fill_1 FILLER_3_775 ();
 sg13g2_decap_8 FILLER_3_804 ();
 sg13g2_decap_8 FILLER_3_811 ();
 sg13g2_decap_8 FILLER_3_818 ();
 sg13g2_decap_8 FILLER_3_825 ();
 sg13g2_decap_8 FILLER_3_832 ();
 sg13g2_decap_8 FILLER_3_839 ();
 sg13g2_decap_8 FILLER_3_846 ();
 sg13g2_decap_8 FILLER_3_853 ();
 sg13g2_decap_8 FILLER_3_860 ();
 sg13g2_decap_8 FILLER_3_867 ();
 sg13g2_decap_8 FILLER_3_874 ();
 sg13g2_decap_8 FILLER_3_881 ();
 sg13g2_decap_8 FILLER_3_888 ();
 sg13g2_decap_8 FILLER_3_895 ();
 sg13g2_decap_8 FILLER_3_902 ();
 sg13g2_decap_8 FILLER_3_909 ();
 sg13g2_decap_8 FILLER_3_916 ();
 sg13g2_decap_8 FILLER_3_923 ();
 sg13g2_decap_8 FILLER_3_930 ();
 sg13g2_decap_8 FILLER_3_937 ();
 sg13g2_decap_8 FILLER_3_944 ();
 sg13g2_decap_8 FILLER_3_951 ();
 sg13g2_decap_8 FILLER_3_958 ();
 sg13g2_decap_8 FILLER_3_965 ();
 sg13g2_decap_8 FILLER_3_972 ();
 sg13g2_decap_8 FILLER_3_979 ();
 sg13g2_decap_8 FILLER_3_986 ();
 sg13g2_decap_8 FILLER_3_993 ();
 sg13g2_decap_8 FILLER_3_1000 ();
 sg13g2_decap_8 FILLER_3_1007 ();
 sg13g2_decap_8 FILLER_3_1014 ();
 sg13g2_decap_8 FILLER_3_1021 ();
 sg13g2_fill_1 FILLER_3_1028 ();
 sg13g2_fill_2 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_2 ();
 sg13g2_fill_1 FILLER_4_78 ();
 sg13g2_fill_2 FILLER_4_115 ();
 sg13g2_fill_1 FILLER_4_173 ();
 sg13g2_fill_2 FILLER_4_195 ();
 sg13g2_fill_1 FILLER_4_197 ();
 sg13g2_fill_2 FILLER_4_231 ();
 sg13g2_fill_2 FILLER_4_266 ();
 sg13g2_fill_2 FILLER_4_340 ();
 sg13g2_fill_1 FILLER_4_362 ();
 sg13g2_fill_1 FILLER_4_393 ();
 sg13g2_fill_1 FILLER_4_433 ();
 sg13g2_fill_2 FILLER_4_442 ();
 sg13g2_fill_1 FILLER_4_444 ();
 sg13g2_fill_2 FILLER_4_470 ();
 sg13g2_fill_2 FILLER_4_526 ();
 sg13g2_fill_1 FILLER_4_554 ();
 sg13g2_fill_2 FILLER_4_596 ();
 sg13g2_fill_2 FILLER_4_723 ();
 sg13g2_fill_2 FILLER_4_745 ();
 sg13g2_decap_8 FILLER_4_824 ();
 sg13g2_decap_8 FILLER_4_831 ();
 sg13g2_decap_8 FILLER_4_838 ();
 sg13g2_decap_8 FILLER_4_845 ();
 sg13g2_decap_8 FILLER_4_852 ();
 sg13g2_decap_8 FILLER_4_859 ();
 sg13g2_decap_8 FILLER_4_866 ();
 sg13g2_decap_8 FILLER_4_873 ();
 sg13g2_decap_8 FILLER_4_880 ();
 sg13g2_decap_8 FILLER_4_887 ();
 sg13g2_decap_8 FILLER_4_894 ();
 sg13g2_decap_8 FILLER_4_901 ();
 sg13g2_decap_8 FILLER_4_908 ();
 sg13g2_decap_8 FILLER_4_915 ();
 sg13g2_decap_8 FILLER_4_922 ();
 sg13g2_decap_8 FILLER_4_929 ();
 sg13g2_decap_8 FILLER_4_936 ();
 sg13g2_decap_8 FILLER_4_943 ();
 sg13g2_decap_8 FILLER_4_950 ();
 sg13g2_decap_8 FILLER_4_957 ();
 sg13g2_decap_8 FILLER_4_964 ();
 sg13g2_decap_8 FILLER_4_971 ();
 sg13g2_decap_8 FILLER_4_978 ();
 sg13g2_decap_8 FILLER_4_985 ();
 sg13g2_decap_8 FILLER_4_992 ();
 sg13g2_decap_8 FILLER_4_999 ();
 sg13g2_decap_8 FILLER_4_1006 ();
 sg13g2_decap_8 FILLER_4_1013 ();
 sg13g2_decap_8 FILLER_4_1020 ();
 sg13g2_fill_2 FILLER_4_1027 ();
 sg13g2_fill_1 FILLER_5_27 ();
 sg13g2_fill_2 FILLER_5_47 ();
 sg13g2_fill_1 FILLER_5_75 ();
 sg13g2_fill_2 FILLER_5_103 ();
 sg13g2_fill_1 FILLER_5_105 ();
 sg13g2_fill_2 FILLER_5_173 ();
 sg13g2_fill_1 FILLER_5_175 ();
 sg13g2_decap_4 FILLER_5_211 ();
 sg13g2_fill_2 FILLER_5_220 ();
 sg13g2_fill_1 FILLER_5_253 ();
 sg13g2_fill_1 FILLER_5_293 ();
 sg13g2_fill_1 FILLER_5_352 ();
 sg13g2_fill_2 FILLER_5_361 ();
 sg13g2_fill_2 FILLER_5_446 ();
 sg13g2_fill_1 FILLER_5_448 ();
 sg13g2_fill_2 FILLER_5_472 ();
 sg13g2_fill_1 FILLER_5_474 ();
 sg13g2_fill_2 FILLER_5_493 ();
 sg13g2_fill_1 FILLER_5_495 ();
 sg13g2_fill_2 FILLER_5_590 ();
 sg13g2_fill_1 FILLER_5_592 ();
 sg13g2_fill_1 FILLER_5_624 ();
 sg13g2_fill_2 FILLER_5_718 ();
 sg13g2_fill_2 FILLER_5_769 ();
 sg13g2_decap_8 FILLER_5_780 ();
 sg13g2_fill_1 FILLER_5_787 ();
 sg13g2_decap_4 FILLER_5_801 ();
 sg13g2_decap_8 FILLER_5_814 ();
 sg13g2_decap_8 FILLER_5_821 ();
 sg13g2_decap_8 FILLER_5_828 ();
 sg13g2_decap_8 FILLER_5_835 ();
 sg13g2_decap_8 FILLER_5_842 ();
 sg13g2_decap_8 FILLER_5_849 ();
 sg13g2_decap_8 FILLER_5_856 ();
 sg13g2_decap_8 FILLER_5_863 ();
 sg13g2_decap_8 FILLER_5_870 ();
 sg13g2_decap_8 FILLER_5_877 ();
 sg13g2_decap_8 FILLER_5_884 ();
 sg13g2_decap_8 FILLER_5_891 ();
 sg13g2_decap_8 FILLER_5_898 ();
 sg13g2_decap_8 FILLER_5_905 ();
 sg13g2_decap_8 FILLER_5_912 ();
 sg13g2_decap_8 FILLER_5_919 ();
 sg13g2_decap_8 FILLER_5_926 ();
 sg13g2_decap_8 FILLER_5_933 ();
 sg13g2_decap_8 FILLER_5_940 ();
 sg13g2_decap_8 FILLER_5_947 ();
 sg13g2_decap_8 FILLER_5_954 ();
 sg13g2_decap_8 FILLER_5_961 ();
 sg13g2_decap_8 FILLER_5_968 ();
 sg13g2_decap_8 FILLER_5_975 ();
 sg13g2_decap_8 FILLER_5_982 ();
 sg13g2_decap_8 FILLER_5_989 ();
 sg13g2_decap_8 FILLER_5_996 ();
 sg13g2_decap_8 FILLER_5_1003 ();
 sg13g2_decap_8 FILLER_5_1010 ();
 sg13g2_decap_8 FILLER_5_1017 ();
 sg13g2_decap_4 FILLER_5_1024 ();
 sg13g2_fill_1 FILLER_5_1028 ();
 sg13g2_fill_2 FILLER_6_76 ();
 sg13g2_fill_2 FILLER_6_87 ();
 sg13g2_fill_2 FILLER_6_131 ();
 sg13g2_fill_1 FILLER_6_133 ();
 sg13g2_fill_1 FILLER_6_162 ();
 sg13g2_fill_2 FILLER_6_176 ();
 sg13g2_fill_1 FILLER_6_178 ();
 sg13g2_decap_8 FILLER_6_213 ();
 sg13g2_fill_1 FILLER_6_220 ();
 sg13g2_fill_2 FILLER_6_256 ();
 sg13g2_fill_1 FILLER_6_258 ();
 sg13g2_fill_2 FILLER_6_276 ();
 sg13g2_fill_2 FILLER_6_314 ();
 sg13g2_fill_1 FILLER_6_316 ();
 sg13g2_fill_1 FILLER_6_339 ();
 sg13g2_fill_2 FILLER_6_363 ();
 sg13g2_fill_1 FILLER_6_365 ();
 sg13g2_fill_2 FILLER_6_472 ();
 sg13g2_fill_2 FILLER_6_486 ();
 sg13g2_fill_1 FILLER_6_488 ();
 sg13g2_fill_1 FILLER_6_552 ();
 sg13g2_fill_1 FILLER_6_624 ();
 sg13g2_fill_2 FILLER_6_676 ();
 sg13g2_fill_2 FILLER_6_726 ();
 sg13g2_fill_2 FILLER_6_756 ();
 sg13g2_fill_2 FILLER_6_776 ();
 sg13g2_decap_8 FILLER_6_832 ();
 sg13g2_decap_8 FILLER_6_839 ();
 sg13g2_decap_8 FILLER_6_846 ();
 sg13g2_decap_8 FILLER_6_853 ();
 sg13g2_decap_8 FILLER_6_860 ();
 sg13g2_decap_8 FILLER_6_867 ();
 sg13g2_decap_8 FILLER_6_874 ();
 sg13g2_decap_8 FILLER_6_881 ();
 sg13g2_decap_8 FILLER_6_888 ();
 sg13g2_decap_8 FILLER_6_895 ();
 sg13g2_decap_8 FILLER_6_902 ();
 sg13g2_decap_8 FILLER_6_909 ();
 sg13g2_decap_8 FILLER_6_916 ();
 sg13g2_decap_8 FILLER_6_923 ();
 sg13g2_decap_8 FILLER_6_930 ();
 sg13g2_decap_8 FILLER_6_937 ();
 sg13g2_decap_8 FILLER_6_944 ();
 sg13g2_decap_8 FILLER_6_951 ();
 sg13g2_decap_8 FILLER_6_958 ();
 sg13g2_decap_8 FILLER_6_965 ();
 sg13g2_decap_8 FILLER_6_972 ();
 sg13g2_decap_8 FILLER_6_979 ();
 sg13g2_decap_8 FILLER_6_986 ();
 sg13g2_decap_8 FILLER_6_993 ();
 sg13g2_decap_8 FILLER_6_1000 ();
 sg13g2_decap_8 FILLER_6_1007 ();
 sg13g2_decap_8 FILLER_6_1014 ();
 sg13g2_decap_8 FILLER_6_1021 ();
 sg13g2_fill_1 FILLER_6_1028 ();
 sg13g2_fill_1 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_130 ();
 sg13g2_fill_1 FILLER_7_140 ();
 sg13g2_decap_4 FILLER_7_215 ();
 sg13g2_fill_2 FILLER_7_231 ();
 sg13g2_fill_1 FILLER_7_233 ();
 sg13g2_fill_2 FILLER_7_239 ();
 sg13g2_fill_1 FILLER_7_241 ();
 sg13g2_fill_1 FILLER_7_247 ();
 sg13g2_fill_2 FILLER_7_257 ();
 sg13g2_fill_2 FILLER_7_304 ();
 sg13g2_fill_1 FILLER_7_306 ();
 sg13g2_fill_2 FILLER_7_320 ();
 sg13g2_fill_1 FILLER_7_322 ();
 sg13g2_fill_1 FILLER_7_360 ();
 sg13g2_fill_2 FILLER_7_367 ();
 sg13g2_fill_1 FILLER_7_369 ();
 sg13g2_fill_2 FILLER_7_379 ();
 sg13g2_fill_2 FILLER_7_409 ();
 sg13g2_fill_1 FILLER_7_411 ();
 sg13g2_fill_2 FILLER_7_442 ();
 sg13g2_fill_1 FILLER_7_444 ();
 sg13g2_fill_2 FILLER_7_485 ();
 sg13g2_fill_2 FILLER_7_514 ();
 sg13g2_fill_1 FILLER_7_555 ();
 sg13g2_fill_1 FILLER_7_640 ();
 sg13g2_fill_2 FILLER_7_691 ();
 sg13g2_fill_1 FILLER_7_693 ();
 sg13g2_fill_2 FILLER_7_723 ();
 sg13g2_fill_1 FILLER_7_725 ();
 sg13g2_decap_4 FILLER_7_802 ();
 sg13g2_fill_2 FILLER_7_806 ();
 sg13g2_decap_8 FILLER_7_835 ();
 sg13g2_decap_8 FILLER_7_842 ();
 sg13g2_decap_8 FILLER_7_849 ();
 sg13g2_decap_8 FILLER_7_856 ();
 sg13g2_decap_8 FILLER_7_863 ();
 sg13g2_decap_8 FILLER_7_870 ();
 sg13g2_decap_8 FILLER_7_877 ();
 sg13g2_decap_8 FILLER_7_884 ();
 sg13g2_decap_8 FILLER_7_891 ();
 sg13g2_decap_8 FILLER_7_898 ();
 sg13g2_decap_8 FILLER_7_905 ();
 sg13g2_decap_8 FILLER_7_912 ();
 sg13g2_decap_8 FILLER_7_919 ();
 sg13g2_decap_8 FILLER_7_926 ();
 sg13g2_decap_8 FILLER_7_933 ();
 sg13g2_decap_8 FILLER_7_940 ();
 sg13g2_decap_8 FILLER_7_947 ();
 sg13g2_decap_8 FILLER_7_954 ();
 sg13g2_decap_8 FILLER_7_961 ();
 sg13g2_decap_8 FILLER_7_968 ();
 sg13g2_decap_8 FILLER_7_975 ();
 sg13g2_decap_8 FILLER_7_982 ();
 sg13g2_decap_8 FILLER_7_989 ();
 sg13g2_decap_8 FILLER_7_996 ();
 sg13g2_decap_8 FILLER_7_1003 ();
 sg13g2_decap_8 FILLER_7_1010 ();
 sg13g2_decap_8 FILLER_7_1017 ();
 sg13g2_decap_4 FILLER_7_1024 ();
 sg13g2_fill_1 FILLER_7_1028 ();
 sg13g2_fill_2 FILLER_8_27 ();
 sg13g2_fill_2 FILLER_8_43 ();
 sg13g2_fill_1 FILLER_8_45 ();
 sg13g2_fill_2 FILLER_8_55 ();
 sg13g2_fill_1 FILLER_8_57 ();
 sg13g2_fill_2 FILLER_8_71 ();
 sg13g2_fill_1 FILLER_8_73 ();
 sg13g2_fill_2 FILLER_8_101 ();
 sg13g2_fill_2 FILLER_8_115 ();
 sg13g2_fill_1 FILLER_8_117 ();
 sg13g2_fill_2 FILLER_8_131 ();
 sg13g2_fill_2 FILLER_8_185 ();
 sg13g2_fill_1 FILLER_8_192 ();
 sg13g2_fill_2 FILLER_8_198 ();
 sg13g2_fill_2 FILLER_8_205 ();
 sg13g2_fill_1 FILLER_8_207 ();
 sg13g2_decap_4 FILLER_8_217 ();
 sg13g2_fill_2 FILLER_8_336 ();
 sg13g2_fill_1 FILLER_8_338 ();
 sg13g2_fill_2 FILLER_8_344 ();
 sg13g2_fill_1 FILLER_8_346 ();
 sg13g2_fill_2 FILLER_8_352 ();
 sg13g2_fill_2 FILLER_8_430 ();
 sg13g2_fill_2 FILLER_8_447 ();
 sg13g2_fill_1 FILLER_8_449 ();
 sg13g2_fill_2 FILLER_8_484 ();
 sg13g2_fill_1 FILLER_8_486 ();
 sg13g2_fill_2 FILLER_8_518 ();
 sg13g2_fill_1 FILLER_8_617 ();
 sg13g2_fill_2 FILLER_8_660 ();
 sg13g2_fill_1 FILLER_8_662 ();
 sg13g2_fill_2 FILLER_8_699 ();
 sg13g2_fill_1 FILLER_8_701 ();
 sg13g2_fill_2 FILLER_8_722 ();
 sg13g2_fill_2 FILLER_8_775 ();
 sg13g2_fill_1 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_807 ();
 sg13g2_decap_4 FILLER_8_814 ();
 sg13g2_fill_2 FILLER_8_818 ();
 sg13g2_decap_8 FILLER_8_857 ();
 sg13g2_decap_8 FILLER_8_864 ();
 sg13g2_decap_8 FILLER_8_871 ();
 sg13g2_decap_8 FILLER_8_878 ();
 sg13g2_decap_8 FILLER_8_885 ();
 sg13g2_decap_8 FILLER_8_892 ();
 sg13g2_decap_8 FILLER_8_899 ();
 sg13g2_decap_8 FILLER_8_906 ();
 sg13g2_decap_8 FILLER_8_913 ();
 sg13g2_decap_8 FILLER_8_920 ();
 sg13g2_decap_8 FILLER_8_927 ();
 sg13g2_decap_8 FILLER_8_934 ();
 sg13g2_decap_8 FILLER_8_941 ();
 sg13g2_decap_8 FILLER_8_948 ();
 sg13g2_decap_8 FILLER_8_955 ();
 sg13g2_decap_8 FILLER_8_962 ();
 sg13g2_decap_8 FILLER_8_969 ();
 sg13g2_decap_8 FILLER_8_976 ();
 sg13g2_decap_8 FILLER_8_983 ();
 sg13g2_decap_8 FILLER_8_990 ();
 sg13g2_decap_8 FILLER_8_997 ();
 sg13g2_decap_8 FILLER_8_1004 ();
 sg13g2_decap_8 FILLER_8_1011 ();
 sg13g2_decap_8 FILLER_8_1018 ();
 sg13g2_decap_4 FILLER_8_1025 ();
 sg13g2_fill_2 FILLER_9_92 ();
 sg13g2_fill_1 FILLER_9_140 ();
 sg13g2_fill_2 FILLER_9_169 ();
 sg13g2_fill_1 FILLER_9_171 ();
 sg13g2_fill_2 FILLER_9_188 ();
 sg13g2_decap_4 FILLER_9_194 ();
 sg13g2_fill_2 FILLER_9_198 ();
 sg13g2_decap_8 FILLER_9_204 ();
 sg13g2_decap_8 FILLER_9_211 ();
 sg13g2_fill_1 FILLER_9_218 ();
 sg13g2_fill_2 FILLER_9_231 ();
 sg13g2_fill_1 FILLER_9_233 ();
 sg13g2_fill_2 FILLER_9_239 ();
 sg13g2_fill_2 FILLER_9_251 ();
 sg13g2_fill_1 FILLER_9_268 ();
 sg13g2_fill_2 FILLER_9_277 ();
 sg13g2_fill_2 FILLER_9_326 ();
 sg13g2_fill_2 FILLER_9_347 ();
 sg13g2_fill_1 FILLER_9_349 ();
 sg13g2_fill_2 FILLER_9_381 ();
 sg13g2_fill_1 FILLER_9_411 ();
 sg13g2_fill_2 FILLER_9_421 ();
 sg13g2_fill_2 FILLER_9_460 ();
 sg13g2_fill_2 FILLER_9_467 ();
 sg13g2_fill_1 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_487 ();
 sg13g2_decap_8 FILLER_9_494 ();
 sg13g2_decap_8 FILLER_9_501 ();
 sg13g2_fill_2 FILLER_9_508 ();
 sg13g2_fill_1 FILLER_9_510 ();
 sg13g2_fill_2 FILLER_9_585 ();
 sg13g2_fill_2 FILLER_9_596 ();
 sg13g2_fill_1 FILLER_9_643 ();
 sg13g2_fill_2 FILLER_9_689 ();
 sg13g2_fill_1 FILLER_9_691 ();
 sg13g2_fill_1 FILLER_9_742 ();
 sg13g2_fill_2 FILLER_9_772 ();
 sg13g2_fill_1 FILLER_9_774 ();
 sg13g2_decap_8 FILLER_9_813 ();
 sg13g2_decap_8 FILLER_9_820 ();
 sg13g2_decap_8 FILLER_9_827 ();
 sg13g2_decap_8 FILLER_9_834 ();
 sg13g2_decap_4 FILLER_9_841 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_decap_8 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_9_868 ();
 sg13g2_decap_8 FILLER_9_875 ();
 sg13g2_decap_8 FILLER_9_882 ();
 sg13g2_decap_8 FILLER_9_889 ();
 sg13g2_decap_8 FILLER_9_896 ();
 sg13g2_decap_8 FILLER_9_903 ();
 sg13g2_decap_8 FILLER_9_910 ();
 sg13g2_decap_8 FILLER_9_917 ();
 sg13g2_decap_8 FILLER_9_924 ();
 sg13g2_decap_8 FILLER_9_931 ();
 sg13g2_decap_8 FILLER_9_938 ();
 sg13g2_decap_8 FILLER_9_945 ();
 sg13g2_decap_8 FILLER_9_952 ();
 sg13g2_decap_8 FILLER_9_959 ();
 sg13g2_decap_8 FILLER_9_966 ();
 sg13g2_decap_8 FILLER_9_973 ();
 sg13g2_decap_8 FILLER_9_980 ();
 sg13g2_decap_8 FILLER_9_987 ();
 sg13g2_decap_8 FILLER_9_994 ();
 sg13g2_decap_8 FILLER_9_1001 ();
 sg13g2_decap_8 FILLER_9_1008 ();
 sg13g2_decap_8 FILLER_9_1015 ();
 sg13g2_decap_8 FILLER_9_1022 ();
 sg13g2_fill_1 FILLER_10_117 ();
 sg13g2_fill_1 FILLER_10_144 ();
 sg13g2_fill_2 FILLER_10_204 ();
 sg13g2_fill_1 FILLER_10_223 ();
 sg13g2_fill_1 FILLER_10_237 ();
 sg13g2_fill_2 FILLER_10_263 ();
 sg13g2_fill_1 FILLER_10_265 ();
 sg13g2_fill_2 FILLER_10_296 ();
 sg13g2_fill_2 FILLER_10_308 ();
 sg13g2_fill_1 FILLER_10_337 ();
 sg13g2_fill_2 FILLER_10_373 ();
 sg13g2_fill_1 FILLER_10_423 ();
 sg13g2_fill_1 FILLER_10_433 ();
 sg13g2_fill_1 FILLER_10_444 ();
 sg13g2_fill_2 FILLER_10_450 ();
 sg13g2_fill_1 FILLER_10_452 ();
 sg13g2_decap_8 FILLER_10_506 ();
 sg13g2_fill_1 FILLER_10_612 ();
 sg13g2_decap_4 FILLER_10_739 ();
 sg13g2_fill_1 FILLER_10_743 ();
 sg13g2_decap_4 FILLER_10_765 ();
 sg13g2_fill_2 FILLER_10_769 ();
 sg13g2_decap_4 FILLER_10_775 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_decap_8 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_10_868 ();
 sg13g2_decap_8 FILLER_10_875 ();
 sg13g2_decap_8 FILLER_10_882 ();
 sg13g2_decap_8 FILLER_10_889 ();
 sg13g2_decap_8 FILLER_10_896 ();
 sg13g2_decap_8 FILLER_10_903 ();
 sg13g2_decap_8 FILLER_10_910 ();
 sg13g2_decap_8 FILLER_10_917 ();
 sg13g2_decap_8 FILLER_10_924 ();
 sg13g2_decap_8 FILLER_10_931 ();
 sg13g2_decap_8 FILLER_10_938 ();
 sg13g2_decap_8 FILLER_10_945 ();
 sg13g2_decap_8 FILLER_10_952 ();
 sg13g2_decap_8 FILLER_10_959 ();
 sg13g2_decap_8 FILLER_10_966 ();
 sg13g2_decap_8 FILLER_10_973 ();
 sg13g2_decap_8 FILLER_10_980 ();
 sg13g2_decap_8 FILLER_10_987 ();
 sg13g2_decap_8 FILLER_10_994 ();
 sg13g2_decap_8 FILLER_10_1001 ();
 sg13g2_decap_8 FILLER_10_1008 ();
 sg13g2_decap_8 FILLER_10_1015 ();
 sg13g2_decap_8 FILLER_10_1022 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_50 ();
 sg13g2_fill_2 FILLER_11_61 ();
 sg13g2_fill_1 FILLER_11_76 ();
 sg13g2_fill_2 FILLER_11_105 ();
 sg13g2_fill_2 FILLER_11_116 ();
 sg13g2_fill_2 FILLER_11_153 ();
 sg13g2_fill_1 FILLER_11_155 ();
 sg13g2_decap_4 FILLER_11_165 ();
 sg13g2_fill_1 FILLER_11_169 ();
 sg13g2_fill_2 FILLER_11_175 ();
 sg13g2_fill_1 FILLER_11_177 ();
 sg13g2_fill_2 FILLER_11_197 ();
 sg13g2_decap_4 FILLER_11_203 ();
 sg13g2_fill_1 FILLER_11_220 ();
 sg13g2_fill_1 FILLER_11_226 ();
 sg13g2_fill_2 FILLER_11_350 ();
 sg13g2_fill_1 FILLER_11_386 ();
 sg13g2_fill_2 FILLER_11_404 ();
 sg13g2_fill_1 FILLER_11_441 ();
 sg13g2_fill_1 FILLER_11_468 ();
 sg13g2_fill_1 FILLER_11_477 ();
 sg13g2_fill_2 FILLER_11_483 ();
 sg13g2_fill_1 FILLER_11_485 ();
 sg13g2_decap_4 FILLER_11_512 ();
 sg13g2_fill_2 FILLER_11_516 ();
 sg13g2_decap_4 FILLER_11_527 ();
 sg13g2_fill_1 FILLER_11_544 ();
 sg13g2_fill_2 FILLER_11_559 ();
 sg13g2_fill_1 FILLER_11_561 ();
 sg13g2_fill_2 FILLER_11_657 ();
 sg13g2_fill_1 FILLER_11_672 ();
 sg13g2_fill_1 FILLER_11_686 ();
 sg13g2_fill_2 FILLER_11_719 ();
 sg13g2_fill_1 FILLER_11_734 ();
 sg13g2_fill_2 FILLER_11_740 ();
 sg13g2_fill_1 FILLER_11_742 ();
 sg13g2_fill_2 FILLER_11_755 ();
 sg13g2_fill_1 FILLER_11_767 ();
 sg13g2_fill_2 FILLER_11_773 ();
 sg13g2_fill_2 FILLER_11_792 ();
 sg13g2_fill_1 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_decap_8 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_11_868 ();
 sg13g2_decap_8 FILLER_11_875 ();
 sg13g2_decap_8 FILLER_11_882 ();
 sg13g2_decap_8 FILLER_11_889 ();
 sg13g2_decap_8 FILLER_11_896 ();
 sg13g2_decap_8 FILLER_11_903 ();
 sg13g2_decap_8 FILLER_11_910 ();
 sg13g2_decap_8 FILLER_11_917 ();
 sg13g2_decap_8 FILLER_11_924 ();
 sg13g2_decap_8 FILLER_11_931 ();
 sg13g2_decap_8 FILLER_11_938 ();
 sg13g2_decap_8 FILLER_11_945 ();
 sg13g2_decap_8 FILLER_11_952 ();
 sg13g2_decap_8 FILLER_11_959 ();
 sg13g2_decap_8 FILLER_11_966 ();
 sg13g2_decap_8 FILLER_11_973 ();
 sg13g2_decap_8 FILLER_11_980 ();
 sg13g2_decap_8 FILLER_11_987 ();
 sg13g2_decap_8 FILLER_11_994 ();
 sg13g2_decap_8 FILLER_11_1001 ();
 sg13g2_decap_8 FILLER_11_1008 ();
 sg13g2_decap_8 FILLER_11_1015 ();
 sg13g2_decap_8 FILLER_11_1022 ();
 sg13g2_fill_2 FILLER_12_27 ();
 sg13g2_fill_2 FILLER_12_99 ();
 sg13g2_fill_1 FILLER_12_101 ();
 sg13g2_fill_2 FILLER_12_152 ();
 sg13g2_decap_8 FILLER_12_166 ();
 sg13g2_fill_1 FILLER_12_184 ();
 sg13g2_decap_8 FILLER_12_190 ();
 sg13g2_fill_2 FILLER_12_197 ();
 sg13g2_fill_2 FILLER_12_221 ();
 sg13g2_fill_1 FILLER_12_223 ();
 sg13g2_fill_1 FILLER_12_232 ();
 sg13g2_fill_2 FILLER_12_300 ();
 sg13g2_fill_1 FILLER_12_302 ();
 sg13g2_fill_2 FILLER_12_361 ();
 sg13g2_fill_1 FILLER_12_363 ();
 sg13g2_fill_2 FILLER_12_445 ();
 sg13g2_fill_1 FILLER_12_461 ();
 sg13g2_decap_4 FILLER_12_469 ();
 sg13g2_fill_1 FILLER_12_487 ();
 sg13g2_decap_8 FILLER_12_505 ();
 sg13g2_decap_8 FILLER_12_512 ();
 sg13g2_decap_4 FILLER_12_519 ();
 sg13g2_fill_1 FILLER_12_582 ();
 sg13g2_fill_2 FILLER_12_592 ();
 sg13g2_fill_1 FILLER_12_644 ();
 sg13g2_fill_1 FILLER_12_709 ();
 sg13g2_fill_1 FILLER_12_718 ();
 sg13g2_fill_2 FILLER_12_746 ();
 sg13g2_fill_1 FILLER_12_748 ();
 sg13g2_fill_2 FILLER_12_754 ();
 sg13g2_fill_1 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_799 ();
 sg13g2_decap_8 FILLER_12_806 ();
 sg13g2_decap_8 FILLER_12_813 ();
 sg13g2_decap_8 FILLER_12_820 ();
 sg13g2_decap_8 FILLER_12_843 ();
 sg13g2_decap_8 FILLER_12_850 ();
 sg13g2_decap_8 FILLER_12_857 ();
 sg13g2_decap_8 FILLER_12_864 ();
 sg13g2_decap_8 FILLER_12_871 ();
 sg13g2_decap_8 FILLER_12_878 ();
 sg13g2_decap_8 FILLER_12_885 ();
 sg13g2_decap_8 FILLER_12_892 ();
 sg13g2_decap_8 FILLER_12_899 ();
 sg13g2_decap_8 FILLER_12_906 ();
 sg13g2_decap_8 FILLER_12_913 ();
 sg13g2_decap_8 FILLER_12_920 ();
 sg13g2_decap_8 FILLER_12_927 ();
 sg13g2_decap_8 FILLER_12_934 ();
 sg13g2_decap_8 FILLER_12_941 ();
 sg13g2_decap_8 FILLER_12_948 ();
 sg13g2_decap_8 FILLER_12_955 ();
 sg13g2_decap_8 FILLER_12_962 ();
 sg13g2_decap_8 FILLER_12_969 ();
 sg13g2_decap_8 FILLER_12_976 ();
 sg13g2_decap_8 FILLER_12_983 ();
 sg13g2_decap_8 FILLER_12_990 ();
 sg13g2_decap_8 FILLER_12_997 ();
 sg13g2_decap_8 FILLER_12_1004 ();
 sg13g2_decap_8 FILLER_12_1011 ();
 sg13g2_decap_8 FILLER_12_1018 ();
 sg13g2_decap_4 FILLER_12_1025 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_10 ();
 sg13g2_fill_1 FILLER_13_12 ();
 sg13g2_fill_2 FILLER_13_40 ();
 sg13g2_fill_1 FILLER_13_42 ();
 sg13g2_fill_1 FILLER_13_132 ();
 sg13g2_fill_1 FILLER_13_194 ();
 sg13g2_fill_1 FILLER_13_232 ();
 sg13g2_fill_2 FILLER_13_246 ();
 sg13g2_fill_2 FILLER_13_275 ();
 sg13g2_fill_1 FILLER_13_401 ();
 sg13g2_fill_1 FILLER_13_428 ();
 sg13g2_fill_1 FILLER_13_458 ();
 sg13g2_decap_4 FILLER_13_464 ();
 sg13g2_fill_1 FILLER_13_468 ();
 sg13g2_decap_8 FILLER_13_474 ();
 sg13g2_decap_4 FILLER_13_493 ();
 sg13g2_fill_2 FILLER_13_545 ();
 sg13g2_fill_1 FILLER_13_547 ();
 sg13g2_fill_1 FILLER_13_584 ();
 sg13g2_decap_8 FILLER_13_709 ();
 sg13g2_fill_2 FILLER_13_771 ();
 sg13g2_fill_2 FILLER_13_780 ();
 sg13g2_fill_2 FILLER_13_827 ();
 sg13g2_decap_8 FILLER_13_856 ();
 sg13g2_decap_8 FILLER_13_863 ();
 sg13g2_decap_8 FILLER_13_870 ();
 sg13g2_decap_8 FILLER_13_877 ();
 sg13g2_decap_8 FILLER_13_884 ();
 sg13g2_decap_8 FILLER_13_891 ();
 sg13g2_decap_8 FILLER_13_898 ();
 sg13g2_decap_8 FILLER_13_905 ();
 sg13g2_decap_8 FILLER_13_912 ();
 sg13g2_decap_8 FILLER_13_919 ();
 sg13g2_decap_8 FILLER_13_926 ();
 sg13g2_decap_8 FILLER_13_933 ();
 sg13g2_decap_8 FILLER_13_940 ();
 sg13g2_decap_8 FILLER_13_947 ();
 sg13g2_decap_8 FILLER_13_954 ();
 sg13g2_decap_8 FILLER_13_961 ();
 sg13g2_decap_8 FILLER_13_968 ();
 sg13g2_decap_8 FILLER_13_975 ();
 sg13g2_decap_8 FILLER_13_982 ();
 sg13g2_decap_8 FILLER_13_989 ();
 sg13g2_decap_8 FILLER_13_996 ();
 sg13g2_decap_8 FILLER_13_1003 ();
 sg13g2_decap_8 FILLER_13_1010 ();
 sg13g2_decap_8 FILLER_13_1017 ();
 sg13g2_decap_4 FILLER_13_1024 ();
 sg13g2_fill_1 FILLER_13_1028 ();
 sg13g2_fill_1 FILLER_14_104 ();
 sg13g2_fill_2 FILLER_14_128 ();
 sg13g2_fill_2 FILLER_14_152 ();
 sg13g2_fill_2 FILLER_14_167 ();
 sg13g2_fill_1 FILLER_14_169 ();
 sg13g2_decap_8 FILLER_14_192 ();
 sg13g2_fill_1 FILLER_14_216 ();
 sg13g2_fill_2 FILLER_14_233 ();
 sg13g2_fill_2 FILLER_14_243 ();
 sg13g2_fill_2 FILLER_14_253 ();
 sg13g2_fill_1 FILLER_14_255 ();
 sg13g2_fill_2 FILLER_14_420 ();
 sg13g2_fill_1 FILLER_14_422 ();
 sg13g2_fill_2 FILLER_14_461 ();
 sg13g2_decap_4 FILLER_14_475 ();
 sg13g2_fill_2 FILLER_14_484 ();
 sg13g2_fill_1 FILLER_14_486 ();
 sg13g2_fill_1 FILLER_14_499 ();
 sg13g2_decap_4 FILLER_14_524 ();
 sg13g2_fill_1 FILLER_14_528 ();
 sg13g2_fill_1 FILLER_14_555 ();
 sg13g2_fill_1 FILLER_14_658 ();
 sg13g2_fill_2 FILLER_14_749 ();
 sg13g2_fill_1 FILLER_14_751 ();
 sg13g2_fill_1 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_4 FILLER_14_805 ();
 sg13g2_fill_1 FILLER_14_809 ();
 sg13g2_decap_8 FILLER_14_846 ();
 sg13g2_decap_8 FILLER_14_853 ();
 sg13g2_decap_8 FILLER_14_860 ();
 sg13g2_decap_8 FILLER_14_867 ();
 sg13g2_decap_8 FILLER_14_874 ();
 sg13g2_decap_8 FILLER_14_881 ();
 sg13g2_decap_8 FILLER_14_888 ();
 sg13g2_decap_8 FILLER_14_895 ();
 sg13g2_decap_8 FILLER_14_902 ();
 sg13g2_decap_8 FILLER_14_909 ();
 sg13g2_decap_8 FILLER_14_916 ();
 sg13g2_decap_8 FILLER_14_923 ();
 sg13g2_decap_8 FILLER_14_930 ();
 sg13g2_decap_8 FILLER_14_937 ();
 sg13g2_decap_8 FILLER_14_944 ();
 sg13g2_decap_8 FILLER_14_951 ();
 sg13g2_decap_8 FILLER_14_958 ();
 sg13g2_decap_8 FILLER_14_965 ();
 sg13g2_decap_8 FILLER_14_972 ();
 sg13g2_decap_8 FILLER_14_979 ();
 sg13g2_decap_8 FILLER_14_986 ();
 sg13g2_decap_8 FILLER_14_993 ();
 sg13g2_decap_8 FILLER_14_1000 ();
 sg13g2_decap_8 FILLER_14_1007 ();
 sg13g2_decap_8 FILLER_14_1014 ();
 sg13g2_decap_8 FILLER_14_1021 ();
 sg13g2_fill_1 FILLER_14_1028 ();
 sg13g2_fill_1 FILLER_15_36 ();
 sg13g2_fill_1 FILLER_15_94 ();
 sg13g2_fill_2 FILLER_15_137 ();
 sg13g2_fill_2 FILLER_15_169 ();
 sg13g2_decap_4 FILLER_15_192 ();
 sg13g2_fill_1 FILLER_15_196 ();
 sg13g2_fill_1 FILLER_15_220 ();
 sg13g2_fill_2 FILLER_15_226 ();
 sg13g2_fill_1 FILLER_15_228 ();
 sg13g2_fill_2 FILLER_15_244 ();
 sg13g2_fill_1 FILLER_15_316 ();
 sg13g2_fill_2 FILLER_15_332 ();
 sg13g2_fill_1 FILLER_15_334 ();
 sg13g2_fill_1 FILLER_15_383 ();
 sg13g2_fill_2 FILLER_15_431 ();
 sg13g2_fill_1 FILLER_15_433 ();
 sg13g2_fill_1 FILLER_15_448 ();
 sg13g2_decap_4 FILLER_15_459 ();
 sg13g2_fill_1 FILLER_15_492 ();
 sg13g2_fill_2 FILLER_15_512 ();
 sg13g2_decap_4 FILLER_15_523 ();
 sg13g2_fill_2 FILLER_15_527 ();
 sg13g2_fill_2 FILLER_15_583 ();
 sg13g2_fill_2 FILLER_15_637 ();
 sg13g2_fill_2 FILLER_15_656 ();
 sg13g2_fill_1 FILLER_15_658 ();
 sg13g2_fill_2 FILLER_15_681 ();
 sg13g2_fill_1 FILLER_15_683 ();
 sg13g2_fill_2 FILLER_15_752 ();
 sg13g2_fill_1 FILLER_15_754 ();
 sg13g2_fill_1 FILLER_15_776 ();
 sg13g2_fill_2 FILLER_15_785 ();
 sg13g2_decap_8 FILLER_15_796 ();
 sg13g2_decap_8 FILLER_15_803 ();
 sg13g2_fill_1 FILLER_15_810 ();
 sg13g2_decap_8 FILLER_15_824 ();
 sg13g2_decap_8 FILLER_15_831 ();
 sg13g2_decap_8 FILLER_15_838 ();
 sg13g2_fill_2 FILLER_15_845 ();
 sg13g2_fill_1 FILLER_15_847 ();
 sg13g2_decap_8 FILLER_15_876 ();
 sg13g2_decap_8 FILLER_15_883 ();
 sg13g2_decap_8 FILLER_15_890 ();
 sg13g2_decap_8 FILLER_15_897 ();
 sg13g2_decap_8 FILLER_15_904 ();
 sg13g2_decap_8 FILLER_15_911 ();
 sg13g2_decap_8 FILLER_15_918 ();
 sg13g2_decap_8 FILLER_15_925 ();
 sg13g2_decap_8 FILLER_15_932 ();
 sg13g2_decap_8 FILLER_15_939 ();
 sg13g2_decap_8 FILLER_15_946 ();
 sg13g2_decap_8 FILLER_15_953 ();
 sg13g2_decap_8 FILLER_15_960 ();
 sg13g2_decap_8 FILLER_15_967 ();
 sg13g2_decap_8 FILLER_15_974 ();
 sg13g2_decap_8 FILLER_15_981 ();
 sg13g2_decap_8 FILLER_15_988 ();
 sg13g2_decap_8 FILLER_15_995 ();
 sg13g2_decap_8 FILLER_15_1002 ();
 sg13g2_decap_8 FILLER_15_1009 ();
 sg13g2_decap_8 FILLER_15_1016 ();
 sg13g2_decap_4 FILLER_15_1023 ();
 sg13g2_fill_2 FILLER_15_1027 ();
 sg13g2_fill_2 FILLER_16_27 ();
 sg13g2_fill_1 FILLER_16_64 ();
 sg13g2_fill_1 FILLER_16_78 ();
 sg13g2_fill_2 FILLER_16_100 ();
 sg13g2_fill_1 FILLER_16_102 ();
 sg13g2_fill_2 FILLER_16_121 ();
 sg13g2_fill_1 FILLER_16_123 ();
 sg13g2_fill_2 FILLER_16_152 ();
 sg13g2_fill_2 FILLER_16_170 ();
 sg13g2_fill_2 FILLER_16_192 ();
 sg13g2_fill_1 FILLER_16_194 ();
 sg13g2_fill_2 FILLER_16_219 ();
 sg13g2_fill_1 FILLER_16_221 ();
 sg13g2_fill_2 FILLER_16_238 ();
 sg13g2_fill_1 FILLER_16_245 ();
 sg13g2_fill_2 FILLER_16_287 ();
 sg13g2_fill_2 FILLER_16_332 ();
 sg13g2_fill_1 FILLER_16_334 ();
 sg13g2_fill_2 FILLER_16_404 ();
 sg13g2_fill_1 FILLER_16_419 ();
 sg13g2_fill_2 FILLER_16_449 ();
 sg13g2_fill_1 FILLER_16_451 ();
 sg13g2_decap_8 FILLER_16_457 ();
 sg13g2_decap_4 FILLER_16_464 ();
 sg13g2_fill_1 FILLER_16_468 ();
 sg13g2_fill_2 FILLER_16_473 ();
 sg13g2_fill_2 FILLER_16_488 ();
 sg13g2_fill_1 FILLER_16_490 ();
 sg13g2_decap_8 FILLER_16_499 ();
 sg13g2_fill_2 FILLER_16_506 ();
 sg13g2_fill_1 FILLER_16_528 ();
 sg13g2_fill_1 FILLER_16_565 ();
 sg13g2_fill_1 FILLER_16_640 ();
 sg13g2_fill_2 FILLER_16_667 ();
 sg13g2_fill_2 FILLER_16_686 ();
 sg13g2_fill_1 FILLER_16_688 ();
 sg13g2_fill_2 FILLER_16_699 ();
 sg13g2_fill_1 FILLER_16_701 ();
 sg13g2_fill_2 FILLER_16_723 ();
 sg13g2_fill_2 FILLER_16_746 ();
 sg13g2_fill_1 FILLER_16_748 ();
 sg13g2_fill_1 FILLER_16_775 ();
 sg13g2_decap_8 FILLER_16_797 ();
 sg13g2_decap_8 FILLER_16_804 ();
 sg13g2_decap_8 FILLER_16_811 ();
 sg13g2_decap_8 FILLER_16_818 ();
 sg13g2_decap_8 FILLER_16_825 ();
 sg13g2_decap_8 FILLER_16_832 ();
 sg13g2_decap_8 FILLER_16_839 ();
 sg13g2_decap_4 FILLER_16_846 ();
 sg13g2_fill_2 FILLER_16_850 ();
 sg13g2_decap_8 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_16_868 ();
 sg13g2_decap_8 FILLER_16_875 ();
 sg13g2_decap_8 FILLER_16_882 ();
 sg13g2_decap_8 FILLER_16_889 ();
 sg13g2_decap_8 FILLER_16_896 ();
 sg13g2_decap_8 FILLER_16_903 ();
 sg13g2_decap_8 FILLER_16_910 ();
 sg13g2_decap_8 FILLER_16_917 ();
 sg13g2_decap_8 FILLER_16_924 ();
 sg13g2_decap_8 FILLER_16_931 ();
 sg13g2_decap_8 FILLER_16_938 ();
 sg13g2_decap_8 FILLER_16_945 ();
 sg13g2_decap_8 FILLER_16_952 ();
 sg13g2_decap_8 FILLER_16_959 ();
 sg13g2_decap_8 FILLER_16_966 ();
 sg13g2_decap_8 FILLER_16_973 ();
 sg13g2_decap_8 FILLER_16_980 ();
 sg13g2_decap_8 FILLER_16_987 ();
 sg13g2_decap_8 FILLER_16_994 ();
 sg13g2_decap_8 FILLER_16_1001 ();
 sg13g2_decap_8 FILLER_16_1008 ();
 sg13g2_decap_8 FILLER_16_1015 ();
 sg13g2_decap_8 FILLER_16_1022 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_2 ();
 sg13g2_fill_1 FILLER_17_43 ();
 sg13g2_fill_2 FILLER_17_92 ();
 sg13g2_fill_1 FILLER_17_107 ();
 sg13g2_fill_2 FILLER_17_126 ();
 sg13g2_fill_1 FILLER_17_136 ();
 sg13g2_fill_1 FILLER_17_145 ();
 sg13g2_fill_1 FILLER_17_168 ();
 sg13g2_fill_2 FILLER_17_190 ();
 sg13g2_fill_1 FILLER_17_192 ();
 sg13g2_fill_1 FILLER_17_213 ();
 sg13g2_fill_2 FILLER_17_233 ();
 sg13g2_fill_2 FILLER_17_269 ();
 sg13g2_fill_1 FILLER_17_339 ();
 sg13g2_fill_2 FILLER_17_354 ();
 sg13g2_fill_1 FILLER_17_356 ();
 sg13g2_fill_1 FILLER_17_366 ();
 sg13g2_fill_2 FILLER_17_404 ();
 sg13g2_fill_2 FILLER_17_414 ();
 sg13g2_fill_2 FILLER_17_439 ();
 sg13g2_decap_4 FILLER_17_474 ();
 sg13g2_fill_1 FILLER_17_478 ();
 sg13g2_fill_1 FILLER_17_484 ();
 sg13g2_decap_4 FILLER_17_499 ();
 sg13g2_fill_2 FILLER_17_522 ();
 sg13g2_fill_2 FILLER_17_583 ();
 sg13g2_fill_1 FILLER_17_585 ();
 sg13g2_fill_2 FILLER_17_643 ();
 sg13g2_fill_2 FILLER_17_658 ();
 sg13g2_fill_1 FILLER_17_668 ();
 sg13g2_decap_4 FILLER_17_694 ();
 sg13g2_fill_2 FILLER_17_715 ();
 sg13g2_fill_1 FILLER_17_717 ();
 sg13g2_fill_2 FILLER_17_767 ();
 sg13g2_fill_1 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_797 ();
 sg13g2_decap_8 FILLER_17_804 ();
 sg13g2_decap_8 FILLER_17_811 ();
 sg13g2_decap_8 FILLER_17_818 ();
 sg13g2_fill_2 FILLER_17_825 ();
 sg13g2_fill_1 FILLER_17_827 ();
 sg13g2_decap_8 FILLER_17_841 ();
 sg13g2_decap_8 FILLER_17_848 ();
 sg13g2_decap_8 FILLER_17_855 ();
 sg13g2_decap_8 FILLER_17_862 ();
 sg13g2_decap_8 FILLER_17_869 ();
 sg13g2_decap_8 FILLER_17_876 ();
 sg13g2_decap_8 FILLER_17_883 ();
 sg13g2_decap_8 FILLER_17_890 ();
 sg13g2_decap_8 FILLER_17_897 ();
 sg13g2_decap_8 FILLER_17_904 ();
 sg13g2_decap_8 FILLER_17_911 ();
 sg13g2_decap_8 FILLER_17_918 ();
 sg13g2_decap_8 FILLER_17_925 ();
 sg13g2_decap_8 FILLER_17_932 ();
 sg13g2_decap_8 FILLER_17_939 ();
 sg13g2_decap_8 FILLER_17_946 ();
 sg13g2_decap_8 FILLER_17_953 ();
 sg13g2_decap_8 FILLER_17_960 ();
 sg13g2_decap_8 FILLER_17_967 ();
 sg13g2_decap_8 FILLER_17_974 ();
 sg13g2_decap_8 FILLER_17_981 ();
 sg13g2_decap_8 FILLER_17_988 ();
 sg13g2_decap_8 FILLER_17_995 ();
 sg13g2_decap_8 FILLER_17_1002 ();
 sg13g2_decap_8 FILLER_17_1009 ();
 sg13g2_decap_8 FILLER_17_1016 ();
 sg13g2_decap_4 FILLER_17_1023 ();
 sg13g2_fill_2 FILLER_17_1027 ();
 sg13g2_fill_2 FILLER_18_4 ();
 sg13g2_fill_2 FILLER_18_91 ();
 sg13g2_fill_1 FILLER_18_93 ();
 sg13g2_fill_2 FILLER_18_125 ();
 sg13g2_fill_1 FILLER_18_127 ();
 sg13g2_fill_1 FILLER_18_133 ();
 sg13g2_fill_1 FILLER_18_139 ();
 sg13g2_fill_2 FILLER_18_163 ();
 sg13g2_fill_1 FILLER_18_165 ();
 sg13g2_fill_2 FILLER_18_179 ();
 sg13g2_fill_1 FILLER_18_181 ();
 sg13g2_decap_4 FILLER_18_194 ();
 sg13g2_fill_1 FILLER_18_198 ();
 sg13g2_fill_1 FILLER_18_220 ();
 sg13g2_fill_1 FILLER_18_261 ();
 sg13g2_fill_1 FILLER_18_288 ();
 sg13g2_fill_2 FILLER_18_329 ();
 sg13g2_fill_1 FILLER_18_331 ();
 sg13g2_fill_1 FILLER_18_380 ();
 sg13g2_fill_1 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_422 ();
 sg13g2_fill_1 FILLER_18_424 ();
 sg13g2_decap_8 FILLER_18_438 ();
 sg13g2_decap_8 FILLER_18_445 ();
 sg13g2_fill_1 FILLER_18_452 ();
 sg13g2_fill_2 FILLER_18_486 ();
 sg13g2_fill_1 FILLER_18_488 ();
 sg13g2_fill_1 FILLER_18_496 ();
 sg13g2_decap_4 FILLER_18_527 ();
 sg13g2_fill_2 FILLER_18_565 ();
 sg13g2_fill_2 FILLER_18_625 ();
 sg13g2_fill_1 FILLER_18_627 ();
 sg13g2_fill_2 FILLER_18_646 ();
 sg13g2_fill_1 FILLER_18_648 ();
 sg13g2_decap_4 FILLER_18_658 ();
 sg13g2_fill_1 FILLER_18_678 ();
 sg13g2_fill_1 FILLER_18_687 ();
 sg13g2_fill_1 FILLER_18_696 ();
 sg13g2_fill_1 FILLER_18_734 ();
 sg13g2_fill_1 FILLER_18_753 ();
 sg13g2_fill_2 FILLER_18_775 ();
 sg13g2_fill_1 FILLER_18_777 ();
 sg13g2_decap_8 FILLER_18_800 ();
 sg13g2_decap_8 FILLER_18_807 ();
 sg13g2_decap_8 FILLER_18_814 ();
 sg13g2_decap_4 FILLER_18_821 ();
 sg13g2_decap_8 FILLER_18_834 ();
 sg13g2_decap_8 FILLER_18_841 ();
 sg13g2_decap_4 FILLER_18_848 ();
 sg13g2_decap_8 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_18_868 ();
 sg13g2_decap_8 FILLER_18_875 ();
 sg13g2_decap_8 FILLER_18_882 ();
 sg13g2_decap_8 FILLER_18_889 ();
 sg13g2_decap_8 FILLER_18_896 ();
 sg13g2_decap_8 FILLER_18_903 ();
 sg13g2_decap_8 FILLER_18_910 ();
 sg13g2_decap_8 FILLER_18_917 ();
 sg13g2_decap_8 FILLER_18_924 ();
 sg13g2_decap_8 FILLER_18_931 ();
 sg13g2_decap_8 FILLER_18_938 ();
 sg13g2_decap_8 FILLER_18_945 ();
 sg13g2_decap_8 FILLER_18_952 ();
 sg13g2_decap_8 FILLER_18_959 ();
 sg13g2_decap_8 FILLER_18_966 ();
 sg13g2_decap_8 FILLER_18_973 ();
 sg13g2_decap_8 FILLER_18_980 ();
 sg13g2_decap_8 FILLER_18_987 ();
 sg13g2_decap_8 FILLER_18_994 ();
 sg13g2_decap_8 FILLER_18_1001 ();
 sg13g2_decap_8 FILLER_18_1008 ();
 sg13g2_decap_8 FILLER_18_1015 ();
 sg13g2_decap_8 FILLER_18_1022 ();
 sg13g2_fill_1 FILLER_19_32 ();
 sg13g2_fill_1 FILLER_19_45 ();
 sg13g2_decap_8 FILLER_19_106 ();
 sg13g2_decap_8 FILLER_19_134 ();
 sg13g2_decap_4 FILLER_19_141 ();
 sg13g2_decap_8 FILLER_19_158 ();
 sg13g2_fill_2 FILLER_19_165 ();
 sg13g2_fill_1 FILLER_19_167 ();
 sg13g2_decap_4 FILLER_19_194 ();
 sg13g2_decap_4 FILLER_19_215 ();
 sg13g2_fill_2 FILLER_19_219 ();
 sg13g2_fill_2 FILLER_19_228 ();
 sg13g2_fill_2 FILLER_19_257 ();
 sg13g2_fill_1 FILLER_19_345 ();
 sg13g2_fill_1 FILLER_19_386 ();
 sg13g2_fill_2 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_406 ();
 sg13g2_fill_2 FILLER_19_435 ();
 sg13g2_fill_2 FILLER_19_449 ();
 sg13g2_fill_1 FILLER_19_451 ();
 sg13g2_decap_8 FILLER_19_495 ();
 sg13g2_fill_1 FILLER_19_502 ();
 sg13g2_fill_1 FILLER_19_508 ();
 sg13g2_fill_2 FILLER_19_528 ();
 sg13g2_fill_2 FILLER_19_557 ();
 sg13g2_fill_1 FILLER_19_634 ();
 sg13g2_decap_4 FILLER_19_652 ();
 sg13g2_fill_2 FILLER_19_660 ();
 sg13g2_fill_1 FILLER_19_662 ();
 sg13g2_decap_8 FILLER_19_694 ();
 sg13g2_fill_1 FILLER_19_701 ();
 sg13g2_fill_1 FILLER_19_714 ();
 sg13g2_decap_4 FILLER_19_725 ();
 sg13g2_fill_1 FILLER_19_729 ();
 sg13g2_fill_2 FILLER_19_771 ();
 sg13g2_fill_1 FILLER_19_773 ();
 sg13g2_fill_2 FILLER_19_794 ();
 sg13g2_fill_1 FILLER_19_796 ();
 sg13g2_fill_1 FILLER_19_824 ();
 sg13g2_fill_2 FILLER_19_852 ();
 sg13g2_decap_8 FILLER_19_867 ();
 sg13g2_decap_8 FILLER_19_874 ();
 sg13g2_decap_8 FILLER_19_881 ();
 sg13g2_decap_8 FILLER_19_888 ();
 sg13g2_decap_8 FILLER_19_895 ();
 sg13g2_decap_8 FILLER_19_902 ();
 sg13g2_decap_8 FILLER_19_909 ();
 sg13g2_decap_8 FILLER_19_916 ();
 sg13g2_decap_8 FILLER_19_923 ();
 sg13g2_decap_8 FILLER_19_930 ();
 sg13g2_decap_8 FILLER_19_937 ();
 sg13g2_decap_8 FILLER_19_944 ();
 sg13g2_decap_8 FILLER_19_951 ();
 sg13g2_decap_8 FILLER_19_958 ();
 sg13g2_decap_8 FILLER_19_965 ();
 sg13g2_decap_8 FILLER_19_972 ();
 sg13g2_decap_8 FILLER_19_979 ();
 sg13g2_decap_8 FILLER_19_986 ();
 sg13g2_decap_8 FILLER_19_993 ();
 sg13g2_decap_8 FILLER_19_1000 ();
 sg13g2_decap_8 FILLER_19_1007 ();
 sg13g2_decap_8 FILLER_19_1014 ();
 sg13g2_decap_8 FILLER_19_1021 ();
 sg13g2_fill_1 FILLER_19_1028 ();
 sg13g2_fill_2 FILLER_20_16 ();
 sg13g2_fill_2 FILLER_20_63 ();
 sg13g2_fill_1 FILLER_20_70 ();
 sg13g2_fill_2 FILLER_20_102 ();
 sg13g2_fill_1 FILLER_20_104 ();
 sg13g2_fill_2 FILLER_20_126 ();
 sg13g2_decap_4 FILLER_20_136 ();
 sg13g2_decap_8 FILLER_20_165 ();
 sg13g2_decap_4 FILLER_20_172 ();
 sg13g2_fill_1 FILLER_20_176 ();
 sg13g2_fill_1 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_227 ();
 sg13g2_fill_2 FILLER_20_315 ();
 sg13g2_fill_1 FILLER_20_416 ();
 sg13g2_fill_2 FILLER_20_430 ();
 sg13g2_fill_2 FILLER_20_449 ();
 sg13g2_fill_1 FILLER_20_451 ();
 sg13g2_fill_1 FILLER_20_479 ();
 sg13g2_decap_8 FILLER_20_484 ();
 sg13g2_decap_4 FILLER_20_491 ();
 sg13g2_fill_1 FILLER_20_503 ();
 sg13g2_fill_2 FILLER_20_557 ();
 sg13g2_fill_1 FILLER_20_559 ();
 sg13g2_fill_1 FILLER_20_629 ();
 sg13g2_fill_1 FILLER_20_638 ();
 sg13g2_fill_2 FILLER_20_662 ();
 sg13g2_fill_1 FILLER_20_664 ();
 sg13g2_decap_8 FILLER_20_690 ();
 sg13g2_fill_1 FILLER_20_697 ();
 sg13g2_decap_8 FILLER_20_722 ();
 sg13g2_decap_4 FILLER_20_729 ();
 sg13g2_fill_2 FILLER_20_733 ();
 sg13g2_fill_2 FILLER_20_816 ();
 sg13g2_fill_1 FILLER_20_818 ();
 sg13g2_decap_4 FILLER_20_846 ();
 sg13g2_fill_1 FILLER_20_850 ();
 sg13g2_decap_8 FILLER_20_887 ();
 sg13g2_decap_8 FILLER_20_894 ();
 sg13g2_decap_8 FILLER_20_901 ();
 sg13g2_decap_8 FILLER_20_908 ();
 sg13g2_decap_8 FILLER_20_915 ();
 sg13g2_decap_8 FILLER_20_922 ();
 sg13g2_decap_8 FILLER_20_929 ();
 sg13g2_decap_8 FILLER_20_936 ();
 sg13g2_decap_8 FILLER_20_943 ();
 sg13g2_decap_8 FILLER_20_950 ();
 sg13g2_decap_8 FILLER_20_957 ();
 sg13g2_decap_8 FILLER_20_964 ();
 sg13g2_decap_8 FILLER_20_971 ();
 sg13g2_decap_8 FILLER_20_978 ();
 sg13g2_decap_8 FILLER_20_985 ();
 sg13g2_decap_8 FILLER_20_992 ();
 sg13g2_decap_8 FILLER_20_999 ();
 sg13g2_decap_8 FILLER_20_1006 ();
 sg13g2_decap_8 FILLER_20_1013 ();
 sg13g2_decap_8 FILLER_20_1020 ();
 sg13g2_fill_2 FILLER_20_1027 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_28 ();
 sg13g2_fill_1 FILLER_21_30 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_4 FILLER_21_105 ();
 sg13g2_fill_1 FILLER_21_109 ();
 sg13g2_decap_8 FILLER_21_127 ();
 sg13g2_decap_8 FILLER_21_134 ();
 sg13g2_fill_1 FILLER_21_141 ();
 sg13g2_fill_1 FILLER_21_152 ();
 sg13g2_decap_8 FILLER_21_177 ();
 sg13g2_decap_8 FILLER_21_184 ();
 sg13g2_decap_4 FILLER_21_191 ();
 sg13g2_fill_2 FILLER_21_195 ();
 sg13g2_decap_4 FILLER_21_201 ();
 sg13g2_fill_2 FILLER_21_237 ();
 sg13g2_fill_2 FILLER_21_279 ();
 sg13g2_fill_1 FILLER_21_343 ();
 sg13g2_fill_1 FILLER_21_379 ();
 sg13g2_fill_1 FILLER_21_449 ();
 sg13g2_fill_1 FILLER_21_458 ();
 sg13g2_fill_1 FILLER_21_475 ();
 sg13g2_fill_2 FILLER_21_484 ();
 sg13g2_fill_1 FILLER_21_486 ();
 sg13g2_fill_2 FILLER_21_565 ();
 sg13g2_fill_1 FILLER_21_615 ();
 sg13g2_fill_2 FILLER_21_629 ();
 sg13g2_decap_8 FILLER_21_649 ();
 sg13g2_fill_2 FILLER_21_656 ();
 sg13g2_fill_1 FILLER_21_658 ();
 sg13g2_fill_2 FILLER_21_667 ();
 sg13g2_fill_2 FILLER_21_693 ();
 sg13g2_fill_1 FILLER_21_695 ();
 sg13g2_fill_2 FILLER_21_726 ();
 sg13g2_decap_8 FILLER_21_741 ();
 sg13g2_decap_4 FILLER_21_748 ();
 sg13g2_fill_2 FILLER_21_752 ();
 sg13g2_decap_4 FILLER_21_780 ();
 sg13g2_fill_1 FILLER_21_784 ();
 sg13g2_fill_2 FILLER_21_871 ();
 sg13g2_decap_8 FILLER_21_901 ();
 sg13g2_decap_8 FILLER_21_908 ();
 sg13g2_decap_8 FILLER_21_915 ();
 sg13g2_decap_8 FILLER_21_922 ();
 sg13g2_decap_8 FILLER_21_929 ();
 sg13g2_decap_8 FILLER_21_936 ();
 sg13g2_decap_8 FILLER_21_943 ();
 sg13g2_decap_8 FILLER_21_950 ();
 sg13g2_decap_8 FILLER_21_957 ();
 sg13g2_decap_8 FILLER_21_964 ();
 sg13g2_decap_8 FILLER_21_971 ();
 sg13g2_decap_8 FILLER_21_978 ();
 sg13g2_decap_8 FILLER_21_985 ();
 sg13g2_decap_8 FILLER_21_992 ();
 sg13g2_decap_8 FILLER_21_999 ();
 sg13g2_decap_8 FILLER_21_1006 ();
 sg13g2_decap_8 FILLER_21_1013 ();
 sg13g2_decap_8 FILLER_21_1020 ();
 sg13g2_fill_2 FILLER_21_1027 ();
 sg13g2_fill_1 FILLER_22_27 ();
 sg13g2_decap_8 FILLER_22_102 ();
 sg13g2_decap_8 FILLER_22_109 ();
 sg13g2_decap_8 FILLER_22_116 ();
 sg13g2_decap_4 FILLER_22_123 ();
 sg13g2_fill_2 FILLER_22_127 ();
 sg13g2_decap_4 FILLER_22_174 ();
 sg13g2_fill_1 FILLER_22_178 ();
 sg13g2_decap_8 FILLER_22_206 ();
 sg13g2_decap_8 FILLER_22_213 ();
 sg13g2_decap_4 FILLER_22_220 ();
 sg13g2_fill_2 FILLER_22_224 ();
 sg13g2_fill_2 FILLER_22_306 ();
 sg13g2_fill_2 FILLER_22_362 ();
 sg13g2_fill_2 FILLER_22_434 ();
 sg13g2_fill_2 FILLER_22_446 ();
 sg13g2_fill_1 FILLER_22_470 ();
 sg13g2_decap_8 FILLER_22_476 ();
 sg13g2_decap_4 FILLER_22_483 ();
 sg13g2_fill_1 FILLER_22_491 ();
 sg13g2_fill_1 FILLER_22_589 ();
 sg13g2_decap_8 FILLER_22_638 ();
 sg13g2_decap_8 FILLER_22_645 ();
 sg13g2_decap_8 FILLER_22_652 ();
 sg13g2_decap_8 FILLER_22_659 ();
 sg13g2_fill_2 FILLER_22_675 ();
 sg13g2_fill_1 FILLER_22_677 ();
 sg13g2_decap_8 FILLER_22_683 ();
 sg13g2_fill_2 FILLER_22_690 ();
 sg13g2_fill_1 FILLER_22_692 ();
 sg13g2_decap_8 FILLER_22_725 ();
 sg13g2_decap_8 FILLER_22_737 ();
 sg13g2_decap_8 FILLER_22_744 ();
 sg13g2_fill_2 FILLER_22_751 ();
 sg13g2_fill_1 FILLER_22_753 ();
 sg13g2_fill_2 FILLER_22_758 ();
 sg13g2_fill_1 FILLER_22_760 ();
 sg13g2_fill_2 FILLER_22_778 ();
 sg13g2_fill_2 FILLER_22_820 ();
 sg13g2_fill_2 FILLER_22_880 ();
 sg13g2_fill_1 FILLER_22_882 ();
 sg13g2_decap_8 FILLER_22_896 ();
 sg13g2_decap_8 FILLER_22_903 ();
 sg13g2_decap_8 FILLER_22_910 ();
 sg13g2_decap_8 FILLER_22_917 ();
 sg13g2_decap_8 FILLER_22_924 ();
 sg13g2_decap_8 FILLER_22_931 ();
 sg13g2_decap_8 FILLER_22_938 ();
 sg13g2_decap_8 FILLER_22_945 ();
 sg13g2_decap_8 FILLER_22_952 ();
 sg13g2_decap_8 FILLER_22_959 ();
 sg13g2_decap_8 FILLER_22_966 ();
 sg13g2_decap_8 FILLER_22_973 ();
 sg13g2_decap_8 FILLER_22_980 ();
 sg13g2_decap_8 FILLER_22_987 ();
 sg13g2_decap_8 FILLER_22_994 ();
 sg13g2_decap_8 FILLER_22_1001 ();
 sg13g2_decap_8 FILLER_22_1008 ();
 sg13g2_decap_8 FILLER_22_1015 ();
 sg13g2_decap_8 FILLER_22_1022 ();
 sg13g2_fill_2 FILLER_23_34 ();
 sg13g2_fill_2 FILLER_23_41 ();
 sg13g2_fill_1 FILLER_23_70 ();
 sg13g2_fill_2 FILLER_23_110 ();
 sg13g2_fill_1 FILLER_23_112 ();
 sg13g2_fill_2 FILLER_23_120 ();
 sg13g2_fill_1 FILLER_23_122 ();
 sg13g2_fill_2 FILLER_23_155 ();
 sg13g2_fill_1 FILLER_23_157 ();
 sg13g2_fill_2 FILLER_23_239 ();
 sg13g2_fill_1 FILLER_23_241 ();
 sg13g2_fill_1 FILLER_23_300 ();
 sg13g2_fill_2 FILLER_23_344 ();
 sg13g2_fill_2 FILLER_23_377 ();
 sg13g2_fill_1 FILLER_23_379 ();
 sg13g2_fill_2 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_427 ();
 sg13g2_fill_1 FILLER_23_434 ();
 sg13g2_decap_8 FILLER_23_451 ();
 sg13g2_fill_2 FILLER_23_458 ();
 sg13g2_fill_1 FILLER_23_460 ();
 sg13g2_fill_2 FILLER_23_481 ();
 sg13g2_fill_2 FILLER_23_529 ();
 sg13g2_fill_1 FILLER_23_540 ();
 sg13g2_fill_2 FILLER_23_567 ();
 sg13g2_fill_1 FILLER_23_583 ();
 sg13g2_decap_8 FILLER_23_615 ();
 sg13g2_decap_4 FILLER_23_622 ();
 sg13g2_fill_1 FILLER_23_626 ();
 sg13g2_decap_4 FILLER_23_663 ();
 sg13g2_fill_2 FILLER_23_667 ();
 sg13g2_decap_8 FILLER_23_691 ();
 sg13g2_decap_4 FILLER_23_698 ();
 sg13g2_fill_1 FILLER_23_702 ();
 sg13g2_fill_2 FILLER_23_708 ();
 sg13g2_fill_1 FILLER_23_710 ();
 sg13g2_decap_4 FILLER_23_718 ();
 sg13g2_fill_2 FILLER_23_722 ();
 sg13g2_fill_2 FILLER_23_729 ();
 sg13g2_fill_2 FILLER_23_750 ();
 sg13g2_decap_8 FILLER_23_784 ();
 sg13g2_fill_2 FILLER_23_791 ();
 sg13g2_fill_1 FILLER_23_793 ();
 sg13g2_fill_1 FILLER_23_798 ();
 sg13g2_fill_1 FILLER_23_826 ();
 sg13g2_fill_1 FILLER_23_881 ();
 sg13g2_decap_8 FILLER_23_909 ();
 sg13g2_decap_8 FILLER_23_916 ();
 sg13g2_decap_8 FILLER_23_923 ();
 sg13g2_decap_8 FILLER_23_930 ();
 sg13g2_decap_8 FILLER_23_937 ();
 sg13g2_decap_8 FILLER_23_944 ();
 sg13g2_decap_8 FILLER_23_951 ();
 sg13g2_decap_8 FILLER_23_958 ();
 sg13g2_decap_8 FILLER_23_965 ();
 sg13g2_decap_8 FILLER_23_972 ();
 sg13g2_decap_8 FILLER_23_979 ();
 sg13g2_decap_8 FILLER_23_986 ();
 sg13g2_decap_8 FILLER_23_993 ();
 sg13g2_decap_8 FILLER_23_1000 ();
 sg13g2_decap_8 FILLER_23_1007 ();
 sg13g2_decap_8 FILLER_23_1014 ();
 sg13g2_decap_8 FILLER_23_1021 ();
 sg13g2_fill_1 FILLER_23_1028 ();
 sg13g2_fill_1 FILLER_24_4 ();
 sg13g2_fill_1 FILLER_24_75 ();
 sg13g2_fill_2 FILLER_24_105 ();
 sg13g2_fill_1 FILLER_24_139 ();
 sg13g2_decap_4 FILLER_24_148 ();
 sg13g2_fill_1 FILLER_24_173 ();
 sg13g2_fill_2 FILLER_24_187 ();
 sg13g2_fill_1 FILLER_24_189 ();
 sg13g2_fill_1 FILLER_24_199 ();
 sg13g2_fill_1 FILLER_24_258 ();
 sg13g2_fill_2 FILLER_24_300 ();
 sg13g2_fill_1 FILLER_24_337 ();
 sg13g2_fill_2 FILLER_24_367 ();
 sg13g2_fill_1 FILLER_24_369 ();
 sg13g2_fill_1 FILLER_24_388 ();
 sg13g2_fill_1 FILLER_24_397 ();
 sg13g2_fill_2 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_406 ();
 sg13g2_fill_2 FILLER_24_421 ();
 sg13g2_fill_1 FILLER_24_451 ();
 sg13g2_decap_4 FILLER_24_460 ();
 sg13g2_decap_8 FILLER_24_487 ();
 sg13g2_decap_8 FILLER_24_494 ();
 sg13g2_decap_4 FILLER_24_501 ();
 sg13g2_fill_1 FILLER_24_505 ();
 sg13g2_fill_1 FILLER_24_537 ();
 sg13g2_fill_2 FILLER_24_555 ();
 sg13g2_fill_1 FILLER_24_634 ();
 sg13g2_fill_2 FILLER_24_643 ();
 sg13g2_fill_1 FILLER_24_662 ();
 sg13g2_decap_8 FILLER_24_699 ();
 sg13g2_fill_2 FILLER_24_706 ();
 sg13g2_fill_2 FILLER_24_720 ();
 sg13g2_fill_1 FILLER_24_722 ();
 sg13g2_decap_8 FILLER_24_740 ();
 sg13g2_decap_4 FILLER_24_747 ();
 sg13g2_fill_2 FILLER_24_751 ();
 sg13g2_decap_8 FILLER_24_779 ();
 sg13g2_decap_4 FILLER_24_786 ();
 sg13g2_fill_1 FILLER_24_830 ();
 sg13g2_decap_8 FILLER_24_912 ();
 sg13g2_decap_8 FILLER_24_919 ();
 sg13g2_decap_8 FILLER_24_926 ();
 sg13g2_decap_8 FILLER_24_933 ();
 sg13g2_decap_8 FILLER_24_940 ();
 sg13g2_decap_8 FILLER_24_947 ();
 sg13g2_decap_8 FILLER_24_954 ();
 sg13g2_decap_8 FILLER_24_961 ();
 sg13g2_decap_8 FILLER_24_968 ();
 sg13g2_decap_8 FILLER_24_975 ();
 sg13g2_decap_8 FILLER_24_982 ();
 sg13g2_decap_8 FILLER_24_989 ();
 sg13g2_decap_8 FILLER_24_996 ();
 sg13g2_decap_8 FILLER_24_1003 ();
 sg13g2_decap_8 FILLER_24_1010 ();
 sg13g2_decap_8 FILLER_24_1017 ();
 sg13g2_decap_4 FILLER_24_1024 ();
 sg13g2_fill_1 FILLER_24_1028 ();
 sg13g2_fill_1 FILLER_25_8 ();
 sg13g2_fill_2 FILLER_25_30 ();
 sg13g2_fill_1 FILLER_25_32 ();
 sg13g2_fill_2 FILLER_25_73 ();
 sg13g2_fill_1 FILLER_25_160 ();
 sg13g2_fill_2 FILLER_25_168 ();
 sg13g2_fill_2 FILLER_25_226 ();
 sg13g2_fill_1 FILLER_25_331 ();
 sg13g2_fill_2 FILLER_25_345 ();
 sg13g2_fill_1 FILLER_25_347 ();
 sg13g2_fill_1 FILLER_25_361 ();
 sg13g2_fill_2 FILLER_25_375 ();
 sg13g2_fill_1 FILLER_25_377 ();
 sg13g2_fill_1 FILLER_25_389 ();
 sg13g2_fill_2 FILLER_25_403 ();
 sg13g2_fill_1 FILLER_25_405 ();
 sg13g2_fill_1 FILLER_25_414 ();
 sg13g2_decap_8 FILLER_25_425 ();
 sg13g2_decap_4 FILLER_25_432 ();
 sg13g2_fill_2 FILLER_25_436 ();
 sg13g2_fill_2 FILLER_25_458 ();
 sg13g2_fill_2 FILLER_25_508 ();
 sg13g2_fill_1 FILLER_25_575 ();
 sg13g2_decap_4 FILLER_25_603 ();
 sg13g2_decap_8 FILLER_25_654 ();
 sg13g2_decap_8 FILLER_25_661 ();
 sg13g2_fill_2 FILLER_25_668 ();
 sg13g2_fill_1 FILLER_25_670 ();
 sg13g2_fill_1 FILLER_25_698 ();
 sg13g2_fill_2 FILLER_25_711 ();
 sg13g2_fill_1 FILLER_25_713 ();
 sg13g2_decap_4 FILLER_25_730 ();
 sg13g2_decap_8 FILLER_25_738 ();
 sg13g2_decap_8 FILLER_25_745 ();
 sg13g2_decap_4 FILLER_25_752 ();
 sg13g2_decap_4 FILLER_25_778 ();
 sg13g2_decap_8 FILLER_25_816 ();
 sg13g2_fill_2 FILLER_25_823 ();
 sg13g2_fill_1 FILLER_25_825 ();
 sg13g2_decap_8 FILLER_25_844 ();
 sg13g2_fill_1 FILLER_25_851 ();
 sg13g2_decap_4 FILLER_25_898 ();
 sg13g2_fill_1 FILLER_25_902 ();
 sg13g2_decap_8 FILLER_25_912 ();
 sg13g2_decap_8 FILLER_25_919 ();
 sg13g2_decap_8 FILLER_25_926 ();
 sg13g2_decap_8 FILLER_25_933 ();
 sg13g2_decap_8 FILLER_25_940 ();
 sg13g2_decap_8 FILLER_25_947 ();
 sg13g2_decap_8 FILLER_25_954 ();
 sg13g2_decap_8 FILLER_25_961 ();
 sg13g2_decap_8 FILLER_25_968 ();
 sg13g2_decap_8 FILLER_25_975 ();
 sg13g2_decap_8 FILLER_25_982 ();
 sg13g2_decap_8 FILLER_25_989 ();
 sg13g2_decap_8 FILLER_25_996 ();
 sg13g2_decap_8 FILLER_25_1003 ();
 sg13g2_decap_8 FILLER_25_1010 ();
 sg13g2_decap_8 FILLER_25_1017 ();
 sg13g2_decap_4 FILLER_25_1024 ();
 sg13g2_fill_1 FILLER_25_1028 ();
 sg13g2_fill_1 FILLER_26_8 ();
 sg13g2_fill_2 FILLER_26_41 ();
 sg13g2_fill_1 FILLER_26_43 ();
 sg13g2_fill_1 FILLER_26_207 ();
 sg13g2_fill_1 FILLER_26_266 ();
 sg13g2_fill_2 FILLER_26_328 ();
 sg13g2_fill_1 FILLER_26_330 ();
 sg13g2_fill_2 FILLER_26_376 ();
 sg13g2_fill_2 FILLER_26_383 ();
 sg13g2_fill_1 FILLER_26_389 ();
 sg13g2_fill_2 FILLER_26_394 ();
 sg13g2_fill_1 FILLER_26_396 ();
 sg13g2_decap_8 FILLER_26_414 ();
 sg13g2_fill_2 FILLER_26_421 ();
 sg13g2_fill_1 FILLER_26_423 ();
 sg13g2_fill_1 FILLER_26_432 ();
 sg13g2_decap_4 FILLER_26_438 ();
 sg13g2_decap_8 FILLER_26_455 ();
 sg13g2_fill_2 FILLER_26_462 ();
 sg13g2_fill_1 FILLER_26_464 ();
 sg13g2_fill_2 FILLER_26_477 ();
 sg13g2_fill_1 FILLER_26_479 ();
 sg13g2_decap_4 FILLER_26_497 ();
 sg13g2_decap_4 FILLER_26_510 ();
 sg13g2_fill_2 FILLER_26_523 ();
 sg13g2_fill_1 FILLER_26_552 ();
 sg13g2_fill_1 FILLER_26_580 ();
 sg13g2_fill_1 FILLER_26_626 ();
 sg13g2_decap_4 FILLER_26_652 ();
 sg13g2_fill_1 FILLER_26_656 ();
 sg13g2_fill_1 FILLER_26_675 ();
 sg13g2_decap_4 FILLER_26_683 ();
 sg13g2_decap_8 FILLER_26_693 ();
 sg13g2_decap_4 FILLER_26_700 ();
 sg13g2_fill_2 FILLER_26_704 ();
 sg13g2_fill_2 FILLER_26_711 ();
 sg13g2_fill_2 FILLER_26_735 ();
 sg13g2_decap_8 FILLER_26_771 ();
 sg13g2_decap_4 FILLER_26_778 ();
 sg13g2_fill_1 FILLER_26_782 ();
 sg13g2_fill_1 FILLER_26_799 ();
 sg13g2_decap_4 FILLER_26_898 ();
 sg13g2_decap_8 FILLER_26_929 ();
 sg13g2_decap_8 FILLER_26_936 ();
 sg13g2_decap_8 FILLER_26_943 ();
 sg13g2_decap_8 FILLER_26_950 ();
 sg13g2_decap_8 FILLER_26_957 ();
 sg13g2_decap_8 FILLER_26_964 ();
 sg13g2_decap_8 FILLER_26_971 ();
 sg13g2_decap_8 FILLER_26_978 ();
 sg13g2_decap_8 FILLER_26_985 ();
 sg13g2_decap_8 FILLER_26_992 ();
 sg13g2_decap_8 FILLER_26_999 ();
 sg13g2_decap_8 FILLER_26_1006 ();
 sg13g2_decap_8 FILLER_26_1013 ();
 sg13g2_decap_8 FILLER_26_1020 ();
 sg13g2_fill_2 FILLER_26_1027 ();
 sg13g2_fill_2 FILLER_27_158 ();
 sg13g2_fill_1 FILLER_27_283 ();
 sg13g2_fill_2 FILLER_27_302 ();
 sg13g2_fill_2 FILLER_27_369 ();
 sg13g2_fill_1 FILLER_27_371 ();
 sg13g2_fill_2 FILLER_27_397 ();
 sg13g2_fill_1 FILLER_27_404 ();
 sg13g2_decap_4 FILLER_27_418 ();
 sg13g2_fill_1 FILLER_27_446 ();
 sg13g2_decap_8 FILLER_27_452 ();
 sg13g2_decap_8 FILLER_27_459 ();
 sg13g2_fill_2 FILLER_27_466 ();
 sg13g2_fill_1 FILLER_27_468 ();
 sg13g2_decap_4 FILLER_27_517 ();
 sg13g2_fill_1 FILLER_27_556 ();
 sg13g2_fill_2 FILLER_27_583 ();
 sg13g2_fill_1 FILLER_27_605 ();
 sg13g2_fill_2 FILLER_27_627 ();
 sg13g2_fill_1 FILLER_27_629 ();
 sg13g2_fill_2 FILLER_27_640 ();
 sg13g2_fill_1 FILLER_27_642 ();
 sg13g2_decap_8 FILLER_27_650 ();
 sg13g2_fill_2 FILLER_27_657 ();
 sg13g2_fill_1 FILLER_27_659 ();
 sg13g2_fill_1 FILLER_27_664 ();
 sg13g2_fill_2 FILLER_27_690 ();
 sg13g2_fill_1 FILLER_27_692 ();
 sg13g2_decap_4 FILLER_27_726 ();
 sg13g2_fill_2 FILLER_27_744 ();
 sg13g2_fill_1 FILLER_27_746 ();
 sg13g2_fill_1 FILLER_27_755 ();
 sg13g2_decap_4 FILLER_27_777 ();
 sg13g2_fill_2 FILLER_27_786 ();
 sg13g2_decap_8 FILLER_27_811 ();
 sg13g2_decap_4 FILLER_27_845 ();
 sg13g2_decap_4 FILLER_27_876 ();
 sg13g2_fill_2 FILLER_27_885 ();
 sg13g2_fill_1 FILLER_27_887 ();
 sg13g2_fill_1 FILLER_27_915 ();
 sg13g2_fill_2 FILLER_27_925 ();
 sg13g2_fill_1 FILLER_27_927 ();
 sg13g2_decap_8 FILLER_27_944 ();
 sg13g2_decap_8 FILLER_27_951 ();
 sg13g2_decap_8 FILLER_27_958 ();
 sg13g2_decap_8 FILLER_27_965 ();
 sg13g2_decap_8 FILLER_27_972 ();
 sg13g2_decap_8 FILLER_27_979 ();
 sg13g2_decap_8 FILLER_27_986 ();
 sg13g2_decap_8 FILLER_27_993 ();
 sg13g2_decap_8 FILLER_27_1000 ();
 sg13g2_decap_8 FILLER_27_1007 ();
 sg13g2_decap_8 FILLER_27_1014 ();
 sg13g2_decap_8 FILLER_27_1021 ();
 sg13g2_fill_1 FILLER_27_1028 ();
 sg13g2_fill_1 FILLER_28_4 ();
 sg13g2_fill_2 FILLER_28_18 ();
 sg13g2_fill_1 FILLER_28_20 ();
 sg13g2_fill_1 FILLER_28_75 ();
 sg13g2_fill_2 FILLER_28_129 ();
 sg13g2_fill_1 FILLER_28_131 ();
 sg13g2_fill_2 FILLER_28_196 ();
 sg13g2_fill_1 FILLER_28_198 ();
 sg13g2_fill_2 FILLER_28_265 ();
 sg13g2_fill_1 FILLER_28_284 ();
 sg13g2_fill_1 FILLER_28_312 ();
 sg13g2_fill_1 FILLER_28_338 ();
 sg13g2_fill_1 FILLER_28_353 ();
 sg13g2_fill_1 FILLER_28_367 ();
 sg13g2_fill_1 FILLER_28_376 ();
 sg13g2_fill_2 FILLER_28_384 ();
 sg13g2_fill_2 FILLER_28_394 ();
 sg13g2_fill_1 FILLER_28_396 ();
 sg13g2_decap_4 FILLER_28_415 ();
 sg13g2_fill_1 FILLER_28_419 ();
 sg13g2_decap_8 FILLER_28_442 ();
 sg13g2_decap_8 FILLER_28_449 ();
 sg13g2_decap_8 FILLER_28_456 ();
 sg13g2_decap_8 FILLER_28_463 ();
 sg13g2_fill_1 FILLER_28_470 ();
 sg13g2_decap_8 FILLER_28_507 ();
 sg13g2_fill_1 FILLER_28_514 ();
 sg13g2_decap_4 FILLER_28_528 ();
 sg13g2_fill_1 FILLER_28_532 ();
 sg13g2_fill_1 FILLER_28_555 ();
 sg13g2_fill_1 FILLER_28_586 ();
 sg13g2_fill_2 FILLER_28_593 ();
 sg13g2_fill_2 FILLER_28_621 ();
 sg13g2_decap_4 FILLER_28_631 ();
 sg13g2_fill_2 FILLER_28_635 ();
 sg13g2_decap_8 FILLER_28_651 ();
 sg13g2_decap_4 FILLER_28_658 ();
 sg13g2_fill_2 FILLER_28_662 ();
 sg13g2_decap_4 FILLER_28_695 ();
 sg13g2_decap_4 FILLER_28_735 ();
 sg13g2_decap_4 FILLER_28_744 ();
 sg13g2_fill_2 FILLER_28_748 ();
 sg13g2_fill_2 FILLER_28_758 ();
 sg13g2_fill_2 FILLER_28_777 ();
 sg13g2_fill_1 FILLER_28_779 ();
 sg13g2_fill_1 FILLER_28_796 ();
 sg13g2_decap_4 FILLER_28_810 ();
 sg13g2_fill_2 FILLER_28_814 ();
 sg13g2_decap_4 FILLER_28_821 ();
 sg13g2_decap_4 FILLER_28_838 ();
 sg13g2_fill_2 FILLER_28_842 ();
 sg13g2_fill_2 FILLER_28_923 ();
 sg13g2_decap_8 FILLER_28_953 ();
 sg13g2_decap_8 FILLER_28_960 ();
 sg13g2_decap_8 FILLER_28_967 ();
 sg13g2_decap_8 FILLER_28_974 ();
 sg13g2_decap_8 FILLER_28_981 ();
 sg13g2_decap_8 FILLER_28_988 ();
 sg13g2_decap_8 FILLER_28_995 ();
 sg13g2_decap_8 FILLER_28_1002 ();
 sg13g2_decap_8 FILLER_28_1009 ();
 sg13g2_decap_8 FILLER_28_1016 ();
 sg13g2_decap_4 FILLER_28_1023 ();
 sg13g2_fill_2 FILLER_28_1027 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_69 ();
 sg13g2_fill_1 FILLER_29_71 ();
 sg13g2_fill_2 FILLER_29_108 ();
 sg13g2_fill_2 FILLER_29_171 ();
 sg13g2_fill_1 FILLER_29_186 ();
 sg13g2_fill_1 FILLER_29_200 ();
 sg13g2_fill_2 FILLER_29_219 ();
 sg13g2_fill_1 FILLER_29_284 ();
 sg13g2_fill_2 FILLER_29_307 ();
 sg13g2_fill_1 FILLER_29_309 ();
 sg13g2_fill_2 FILLER_29_389 ();
 sg13g2_fill_1 FILLER_29_391 ();
 sg13g2_fill_1 FILLER_29_416 ();
 sg13g2_decap_4 FILLER_29_451 ();
 sg13g2_fill_1 FILLER_29_482 ();
 sg13g2_decap_4 FILLER_29_488 ();
 sg13g2_fill_2 FILLER_29_492 ();
 sg13g2_fill_2 FILLER_29_599 ();
 sg13g2_fill_1 FILLER_29_601 ();
 sg13g2_fill_2 FILLER_29_656 ();
 sg13g2_fill_2 FILLER_29_686 ();
 sg13g2_fill_1 FILLER_29_688 ();
 sg13g2_decap_8 FILLER_29_699 ();
 sg13g2_fill_1 FILLER_29_728 ();
 sg13g2_fill_2 FILLER_29_738 ();
 sg13g2_decap_8 FILLER_29_748 ();
 sg13g2_fill_2 FILLER_29_755 ();
 sg13g2_fill_1 FILLER_29_757 ();
 sg13g2_fill_1 FILLER_29_762 ();
 sg13g2_fill_1 FILLER_29_780 ();
 sg13g2_decap_8 FILLER_29_796 ();
 sg13g2_fill_2 FILLER_29_875 ();
 sg13g2_fill_1 FILLER_29_877 ();
 sg13g2_fill_2 FILLER_29_886 ();
 sg13g2_fill_1 FILLER_29_888 ();
 sg13g2_fill_1 FILLER_29_930 ();
 sg13g2_decap_8 FILLER_29_947 ();
 sg13g2_decap_8 FILLER_29_954 ();
 sg13g2_decap_8 FILLER_29_961 ();
 sg13g2_decap_8 FILLER_29_968 ();
 sg13g2_decap_8 FILLER_29_975 ();
 sg13g2_decap_8 FILLER_29_982 ();
 sg13g2_decap_8 FILLER_29_989 ();
 sg13g2_decap_8 FILLER_29_996 ();
 sg13g2_decap_8 FILLER_29_1003 ();
 sg13g2_decap_8 FILLER_29_1010 ();
 sg13g2_decap_8 FILLER_29_1017 ();
 sg13g2_decap_4 FILLER_29_1024 ();
 sg13g2_fill_1 FILLER_29_1028 ();
 sg13g2_fill_1 FILLER_30_4 ();
 sg13g2_fill_1 FILLER_30_90 ();
 sg13g2_fill_1 FILLER_30_100 ();
 sg13g2_fill_1 FILLER_30_183 ();
 sg13g2_fill_1 FILLER_30_229 ();
 sg13g2_fill_2 FILLER_30_265 ();
 sg13g2_fill_2 FILLER_30_303 ();
 sg13g2_fill_1 FILLER_30_305 ();
 sg13g2_fill_2 FILLER_30_342 ();
 sg13g2_decap_4 FILLER_30_413 ();
 sg13g2_fill_2 FILLER_30_417 ();
 sg13g2_fill_2 FILLER_30_436 ();
 sg13g2_fill_2 FILLER_30_456 ();
 sg13g2_fill_1 FILLER_30_458 ();
 sg13g2_fill_2 FILLER_30_622 ();
 sg13g2_fill_1 FILLER_30_624 ();
 sg13g2_fill_2 FILLER_30_636 ();
 sg13g2_fill_1 FILLER_30_638 ();
 sg13g2_fill_2 FILLER_30_688 ();
 sg13g2_fill_2 FILLER_30_694 ();
 sg13g2_fill_2 FILLER_30_708 ();
 sg13g2_fill_1 FILLER_30_710 ();
 sg13g2_fill_2 FILLER_30_761 ();
 sg13g2_fill_1 FILLER_30_771 ();
 sg13g2_decap_4 FILLER_30_790 ();
 sg13g2_fill_1 FILLER_30_794 ();
 sg13g2_fill_1 FILLER_30_816 ();
 sg13g2_decap_4 FILLER_30_834 ();
 sg13g2_fill_2 FILLER_30_838 ();
 sg13g2_fill_1 FILLER_30_857 ();
 sg13g2_fill_2 FILLER_30_878 ();
 sg13g2_fill_1 FILLER_30_880 ();
 sg13g2_fill_2 FILLER_30_899 ();
 sg13g2_fill_1 FILLER_30_901 ();
 sg13g2_decap_4 FILLER_30_932 ();
 sg13g2_fill_1 FILLER_30_936 ();
 sg13g2_decap_8 FILLER_30_964 ();
 sg13g2_decap_8 FILLER_30_971 ();
 sg13g2_decap_8 FILLER_30_978 ();
 sg13g2_decap_8 FILLER_30_985 ();
 sg13g2_decap_8 FILLER_30_992 ();
 sg13g2_decap_8 FILLER_30_999 ();
 sg13g2_decap_8 FILLER_30_1006 ();
 sg13g2_decap_8 FILLER_30_1013 ();
 sg13g2_decap_8 FILLER_30_1020 ();
 sg13g2_fill_2 FILLER_30_1027 ();
 sg13g2_fill_2 FILLER_31_4 ();
 sg13g2_fill_2 FILLER_31_73 ();
 sg13g2_fill_1 FILLER_31_75 ();
 sg13g2_fill_2 FILLER_31_150 ();
 sg13g2_fill_1 FILLER_31_152 ();
 sg13g2_fill_1 FILLER_31_213 ();
 sg13g2_fill_2 FILLER_31_263 ();
 sg13g2_fill_1 FILLER_31_320 ();
 sg13g2_fill_2 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_411 ();
 sg13g2_decap_8 FILLER_31_418 ();
 sg13g2_decap_4 FILLER_31_425 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_decap_8 FILLER_31_450 ();
 sg13g2_fill_1 FILLER_31_461 ();
 sg13g2_fill_1 FILLER_31_498 ();
 sg13g2_decap_8 FILLER_31_519 ();
 sg13g2_fill_2 FILLER_31_620 ();
 sg13g2_fill_2 FILLER_31_657 ();
 sg13g2_fill_2 FILLER_31_678 ();
 sg13g2_decap_4 FILLER_31_685 ();
 sg13g2_fill_2 FILLER_31_689 ();
 sg13g2_decap_4 FILLER_31_700 ();
 sg13g2_fill_2 FILLER_31_714 ();
 sg13g2_fill_1 FILLER_31_716 ();
 sg13g2_fill_2 FILLER_31_730 ();
 sg13g2_fill_1 FILLER_31_732 ();
 sg13g2_fill_1 FILLER_31_738 ();
 sg13g2_fill_1 FILLER_31_744 ();
 sg13g2_fill_1 FILLER_31_784 ();
 sg13g2_fill_2 FILLER_31_793 ();
 sg13g2_fill_1 FILLER_31_795 ();
 sg13g2_fill_2 FILLER_31_808 ();
 sg13g2_fill_2 FILLER_31_823 ();
 sg13g2_fill_1 FILLER_31_825 ();
 sg13g2_fill_2 FILLER_31_855 ();
 sg13g2_decap_8 FILLER_31_930 ();
 sg13g2_decap_8 FILLER_31_964 ();
 sg13g2_decap_8 FILLER_31_971 ();
 sg13g2_decap_8 FILLER_31_978 ();
 sg13g2_decap_8 FILLER_31_985 ();
 sg13g2_decap_8 FILLER_31_992 ();
 sg13g2_decap_8 FILLER_31_999 ();
 sg13g2_decap_8 FILLER_31_1006 ();
 sg13g2_decap_8 FILLER_31_1013 ();
 sg13g2_decap_8 FILLER_31_1020 ();
 sg13g2_fill_2 FILLER_31_1027 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_2 ();
 sg13g2_fill_1 FILLER_32_43 ();
 sg13g2_fill_1 FILLER_32_89 ();
 sg13g2_fill_1 FILLER_32_170 ();
 sg13g2_fill_1 FILLER_32_211 ();
 sg13g2_fill_1 FILLER_32_244 ();
 sg13g2_fill_1 FILLER_32_339 ();
 sg13g2_fill_2 FILLER_32_397 ();
 sg13g2_fill_1 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_427 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_4 FILLER_32_447 ();
 sg13g2_fill_1 FILLER_32_489 ();
 sg13g2_fill_2 FILLER_32_523 ();
 sg13g2_fill_2 FILLER_32_565 ();
 sg13g2_fill_1 FILLER_32_567 ();
 sg13g2_fill_1 FILLER_32_581 ();
 sg13g2_fill_1 FILLER_32_635 ();
 sg13g2_fill_1 FILLER_32_650 ();
 sg13g2_fill_2 FILLER_32_664 ();
 sg13g2_fill_1 FILLER_32_666 ();
 sg13g2_decap_4 FILLER_32_676 ();
 sg13g2_fill_2 FILLER_32_680 ();
 sg13g2_fill_2 FILLER_32_695 ();
 sg13g2_fill_1 FILLER_32_697 ();
 sg13g2_fill_2 FILLER_32_729 ();
 sg13g2_fill_2 FILLER_32_740 ();
 sg13g2_fill_2 FILLER_32_790 ();
 sg13g2_fill_1 FILLER_32_792 ();
 sg13g2_fill_2 FILLER_32_821 ();
 sg13g2_decap_4 FILLER_32_831 ();
 sg13g2_fill_1 FILLER_32_835 ();
 sg13g2_fill_1 FILLER_32_871 ();
 sg13g2_fill_2 FILLER_32_877 ();
 sg13g2_fill_2 FILLER_32_886 ();
 sg13g2_fill_2 FILLER_32_924 ();
 sg13g2_fill_1 FILLER_32_926 ();
 sg13g2_decap_8 FILLER_32_970 ();
 sg13g2_decap_8 FILLER_32_977 ();
 sg13g2_decap_8 FILLER_32_984 ();
 sg13g2_decap_8 FILLER_32_991 ();
 sg13g2_decap_8 FILLER_32_998 ();
 sg13g2_decap_8 FILLER_32_1005 ();
 sg13g2_decap_8 FILLER_32_1012 ();
 sg13g2_decap_8 FILLER_32_1019 ();
 sg13g2_fill_2 FILLER_32_1026 ();
 sg13g2_fill_1 FILLER_32_1028 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_23 ();
 sg13g2_fill_1 FILLER_33_25 ();
 sg13g2_fill_2 FILLER_33_107 ();
 sg13g2_fill_2 FILLER_33_123 ();
 sg13g2_fill_1 FILLER_33_125 ();
 sg13g2_fill_2 FILLER_33_135 ();
 sg13g2_fill_2 FILLER_33_150 ();
 sg13g2_fill_1 FILLER_33_152 ();
 sg13g2_fill_2 FILLER_33_197 ();
 sg13g2_fill_1 FILLER_33_349 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_1 FILLER_33_456 ();
 sg13g2_fill_2 FILLER_33_513 ();
 sg13g2_fill_1 FILLER_33_515 ();
 sg13g2_fill_2 FILLER_33_533 ();
 sg13g2_fill_1 FILLER_33_535 ();
 sg13g2_fill_2 FILLER_33_569 ();
 sg13g2_fill_2 FILLER_33_588 ();
 sg13g2_fill_1 FILLER_33_614 ();
 sg13g2_fill_2 FILLER_33_632 ();
 sg13g2_fill_2 FILLER_33_696 ();
 sg13g2_fill_2 FILLER_33_747 ();
 sg13g2_fill_2 FILLER_33_778 ();
 sg13g2_fill_2 FILLER_33_788 ();
 sg13g2_fill_2 FILLER_33_807 ();
 sg13g2_decap_4 FILLER_33_830 ();
 sg13g2_fill_2 FILLER_33_834 ();
 sg13g2_fill_2 FILLER_33_860 ();
 sg13g2_fill_2 FILLER_33_889 ();
 sg13g2_fill_2 FILLER_33_936 ();
 sg13g2_decap_8 FILLER_33_974 ();
 sg13g2_decap_8 FILLER_33_981 ();
 sg13g2_decap_8 FILLER_33_988 ();
 sg13g2_decap_8 FILLER_33_995 ();
 sg13g2_decap_8 FILLER_33_1002 ();
 sg13g2_decap_8 FILLER_33_1009 ();
 sg13g2_decap_8 FILLER_33_1016 ();
 sg13g2_decap_4 FILLER_33_1023 ();
 sg13g2_fill_2 FILLER_33_1027 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_29 ();
 sg13g2_fill_1 FILLER_34_66 ();
 sg13g2_fill_1 FILLER_34_94 ();
 sg13g2_fill_2 FILLER_34_122 ();
 sg13g2_fill_1 FILLER_34_124 ();
 sg13g2_fill_1 FILLER_34_186 ();
 sg13g2_fill_1 FILLER_34_203 ();
 sg13g2_fill_2 FILLER_34_244 ();
 sg13g2_fill_1 FILLER_34_246 ();
 sg13g2_fill_2 FILLER_34_274 ();
 sg13g2_fill_2 FILLER_34_343 ();
 sg13g2_fill_1 FILLER_34_376 ();
 sg13g2_fill_2 FILLER_34_440 ();
 sg13g2_fill_1 FILLER_34_442 ();
 sg13g2_fill_2 FILLER_34_540 ();
 sg13g2_fill_1 FILLER_34_542 ();
 sg13g2_fill_2 FILLER_34_642 ();
 sg13g2_fill_1 FILLER_34_644 ();
 sg13g2_fill_2 FILLER_34_658 ();
 sg13g2_fill_1 FILLER_34_660 ();
 sg13g2_fill_2 FILLER_34_744 ();
 sg13g2_fill_2 FILLER_34_752 ();
 sg13g2_fill_1 FILLER_34_754 ();
 sg13g2_fill_1 FILLER_34_809 ();
 sg13g2_fill_1 FILLER_34_831 ();
 sg13g2_fill_2 FILLER_34_850 ();
 sg13g2_decap_8 FILLER_34_865 ();
 sg13g2_fill_2 FILLER_34_872 ();
 sg13g2_decap_8 FILLER_34_976 ();
 sg13g2_decap_8 FILLER_34_983 ();
 sg13g2_decap_8 FILLER_34_990 ();
 sg13g2_decap_8 FILLER_34_997 ();
 sg13g2_decap_8 FILLER_34_1004 ();
 sg13g2_decap_8 FILLER_34_1011 ();
 sg13g2_decap_8 FILLER_34_1018 ();
 sg13g2_decap_4 FILLER_34_1025 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_162 ();
 sg13g2_fill_2 FILLER_35_181 ();
 sg13g2_fill_1 FILLER_35_183 ();
 sg13g2_fill_1 FILLER_35_202 ();
 sg13g2_fill_1 FILLER_35_302 ();
 sg13g2_fill_2 FILLER_35_503 ();
 sg13g2_fill_1 FILLER_35_522 ();
 sg13g2_fill_1 FILLER_35_630 ();
 sg13g2_fill_1 FILLER_35_694 ();
 sg13g2_fill_2 FILLER_35_699 ();
 sg13g2_fill_2 FILLER_35_738 ();
 sg13g2_fill_1 FILLER_35_762 ();
 sg13g2_fill_2 FILLER_35_781 ();
 sg13g2_fill_1 FILLER_35_783 ();
 sg13g2_fill_2 FILLER_35_805 ();
 sg13g2_fill_1 FILLER_35_807 ();
 sg13g2_decap_4 FILLER_35_832 ();
 sg13g2_fill_2 FILLER_35_836 ();
 sg13g2_fill_1 FILLER_35_842 ();
 sg13g2_decap_8 FILLER_35_855 ();
 sg13g2_fill_2 FILLER_35_911 ();
 sg13g2_decap_8 FILLER_35_985 ();
 sg13g2_decap_8 FILLER_35_992 ();
 sg13g2_decap_8 FILLER_35_999 ();
 sg13g2_decap_8 FILLER_35_1006 ();
 sg13g2_decap_8 FILLER_35_1013 ();
 sg13g2_decap_8 FILLER_35_1020 ();
 sg13g2_fill_2 FILLER_35_1027 ();
 sg13g2_fill_1 FILLER_36_81 ();
 sg13g2_fill_2 FILLER_36_122 ();
 sg13g2_fill_1 FILLER_36_124 ();
 sg13g2_fill_1 FILLER_36_179 ();
 sg13g2_fill_1 FILLER_36_213 ();
 sg13g2_fill_1 FILLER_36_232 ();
 sg13g2_fill_2 FILLER_36_260 ();
 sg13g2_fill_1 FILLER_36_262 ();
 sg13g2_fill_2 FILLER_36_297 ();
 sg13g2_fill_1 FILLER_36_299 ();
 sg13g2_fill_2 FILLER_36_332 ();
 sg13g2_fill_2 FILLER_36_475 ();
 sg13g2_fill_1 FILLER_36_548 ();
 sg13g2_fill_1 FILLER_36_585 ();
 sg13g2_fill_1 FILLER_36_715 ();
 sg13g2_fill_2 FILLER_36_765 ();
 sg13g2_fill_1 FILLER_36_767 ();
 sg13g2_fill_2 FILLER_36_810 ();
 sg13g2_fill_2 FILLER_36_819 ();
 sg13g2_fill_1 FILLER_36_821 ();
 sg13g2_fill_2 FILLER_36_838 ();
 sg13g2_fill_1 FILLER_36_840 ();
 sg13g2_fill_1 FILLER_36_876 ();
 sg13g2_decap_4 FILLER_36_930 ();
 sg13g2_fill_1 FILLER_36_934 ();
 sg13g2_decap_8 FILLER_36_980 ();
 sg13g2_decap_8 FILLER_36_987 ();
 sg13g2_decap_8 FILLER_36_994 ();
 sg13g2_decap_8 FILLER_36_1001 ();
 sg13g2_decap_8 FILLER_36_1008 ();
 sg13g2_decap_8 FILLER_36_1015 ();
 sg13g2_decap_8 FILLER_36_1022 ();
 sg13g2_fill_2 FILLER_37_52 ();
 sg13g2_fill_1 FILLER_37_67 ();
 sg13g2_fill_1 FILLER_37_225 ();
 sg13g2_fill_1 FILLER_37_240 ();
 sg13g2_fill_2 FILLER_37_321 ();
 sg13g2_fill_2 FILLER_37_385 ();
 sg13g2_fill_1 FILLER_37_387 ();
 sg13g2_fill_2 FILLER_37_401 ();
 sg13g2_fill_1 FILLER_37_403 ();
 sg13g2_fill_1 FILLER_37_426 ();
 sg13g2_decap_8 FILLER_37_503 ();
 sg13g2_fill_2 FILLER_37_518 ();
 sg13g2_fill_2 FILLER_37_547 ();
 sg13g2_fill_1 FILLER_37_561 ();
 sg13g2_fill_2 FILLER_37_577 ();
 sg13g2_fill_2 FILLER_37_632 ();
 sg13g2_fill_1 FILLER_37_634 ();
 sg13g2_fill_2 FILLER_37_670 ();
 sg13g2_fill_1 FILLER_37_672 ();
 sg13g2_fill_1 FILLER_37_726 ();
 sg13g2_fill_1 FILLER_37_767 ();
 sg13g2_fill_1 FILLER_37_789 ();
 sg13g2_fill_2 FILLER_37_805 ();
 sg13g2_fill_1 FILLER_37_816 ();
 sg13g2_fill_2 FILLER_37_835 ();
 sg13g2_fill_1 FILLER_37_837 ();
 sg13g2_decap_4 FILLER_37_850 ();
 sg13g2_fill_2 FILLER_37_854 ();
 sg13g2_fill_2 FILLER_37_905 ();
 sg13g2_decap_8 FILLER_37_974 ();
 sg13g2_decap_8 FILLER_37_981 ();
 sg13g2_decap_8 FILLER_37_988 ();
 sg13g2_decap_8 FILLER_37_995 ();
 sg13g2_decap_8 FILLER_37_1002 ();
 sg13g2_decap_8 FILLER_37_1009 ();
 sg13g2_decap_8 FILLER_37_1016 ();
 sg13g2_decap_4 FILLER_37_1023 ();
 sg13g2_fill_2 FILLER_37_1027 ();
 sg13g2_fill_2 FILLER_38_80 ();
 sg13g2_fill_2 FILLER_38_209 ();
 sg13g2_fill_1 FILLER_38_211 ();
 sg13g2_fill_2 FILLER_38_248 ();
 sg13g2_fill_1 FILLER_38_250 ();
 sg13g2_fill_2 FILLER_38_300 ();
 sg13g2_fill_1 FILLER_38_375 ();
 sg13g2_fill_1 FILLER_38_403 ();
 sg13g2_fill_1 FILLER_38_444 ();
 sg13g2_fill_2 FILLER_38_485 ();
 sg13g2_fill_2 FILLER_38_503 ();
 sg13g2_decap_4 FILLER_38_509 ();
 sg13g2_fill_2 FILLER_38_513 ();
 sg13g2_fill_2 FILLER_38_543 ();
 sg13g2_fill_1 FILLER_38_545 ();
 sg13g2_fill_2 FILLER_38_566 ();
 sg13g2_fill_1 FILLER_38_576 ();
 sg13g2_fill_1 FILLER_38_588 ();
 sg13g2_fill_2 FILLER_38_668 ();
 sg13g2_fill_1 FILLER_38_670 ();
 sg13g2_fill_2 FILLER_38_687 ();
 sg13g2_decap_4 FILLER_38_716 ();
 sg13g2_fill_1 FILLER_38_720 ();
 sg13g2_fill_1 FILLER_38_756 ();
 sg13g2_fill_2 FILLER_38_791 ();
 sg13g2_fill_1 FILLER_38_800 ();
 sg13g2_decap_8 FILLER_38_813 ();
 sg13g2_decap_4 FILLER_38_830 ();
 sg13g2_fill_1 FILLER_38_872 ();
 sg13g2_decap_4 FILLER_38_909 ();
 sg13g2_fill_2 FILLER_38_913 ();
 sg13g2_decap_8 FILLER_38_981 ();
 sg13g2_decap_8 FILLER_38_988 ();
 sg13g2_decap_8 FILLER_38_995 ();
 sg13g2_decap_8 FILLER_38_1002 ();
 sg13g2_decap_8 FILLER_38_1009 ();
 sg13g2_decap_8 FILLER_38_1016 ();
 sg13g2_decap_4 FILLER_38_1023 ();
 sg13g2_fill_2 FILLER_38_1027 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_159 ();
 sg13g2_fill_2 FILLER_39_187 ();
 sg13g2_fill_2 FILLER_39_243 ();
 sg13g2_fill_2 FILLER_39_317 ();
 sg13g2_fill_1 FILLER_39_319 ();
 sg13g2_fill_2 FILLER_39_369 ();
 sg13g2_fill_1 FILLER_39_473 ();
 sg13g2_fill_1 FILLER_39_486 ();
 sg13g2_fill_2 FILLER_39_509 ();
 sg13g2_decap_4 FILLER_39_516 ();
 sg13g2_fill_1 FILLER_39_520 ();
 sg13g2_fill_2 FILLER_39_540 ();
 sg13g2_fill_1 FILLER_39_542 ();
 sg13g2_fill_1 FILLER_39_575 ();
 sg13g2_fill_1 FILLER_39_605 ();
 sg13g2_fill_1 FILLER_39_611 ();
 sg13g2_fill_2 FILLER_39_637 ();
 sg13g2_fill_2 FILLER_39_669 ();
 sg13g2_fill_1 FILLER_39_671 ();
 sg13g2_decap_8 FILLER_39_717 ();
 sg13g2_fill_2 FILLER_39_724 ();
 sg13g2_fill_1 FILLER_39_738 ();
 sg13g2_fill_2 FILLER_39_781 ();
 sg13g2_fill_1 FILLER_39_783 ();
 sg13g2_decap_4 FILLER_39_809 ();
 sg13g2_fill_2 FILLER_39_839 ();
 sg13g2_decap_4 FILLER_39_922 ();
 sg13g2_fill_2 FILLER_39_926 ();
 sg13g2_decap_8 FILLER_39_972 ();
 sg13g2_decap_8 FILLER_39_979 ();
 sg13g2_decap_8 FILLER_39_986 ();
 sg13g2_decap_8 FILLER_39_993 ();
 sg13g2_decap_8 FILLER_39_1000 ();
 sg13g2_decap_8 FILLER_39_1007 ();
 sg13g2_decap_8 FILLER_39_1014 ();
 sg13g2_decap_8 FILLER_39_1021 ();
 sg13g2_fill_1 FILLER_39_1028 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_43 ();
 sg13g2_fill_1 FILLER_40_81 ();
 sg13g2_fill_2 FILLER_40_100 ();
 sg13g2_fill_1 FILLER_40_102 ();
 sg13g2_fill_2 FILLER_40_144 ();
 sg13g2_fill_1 FILLER_40_146 ();
 sg13g2_fill_1 FILLER_40_210 ();
 sg13g2_fill_2 FILLER_40_319 ();
 sg13g2_fill_1 FILLER_40_392 ();
 sg13g2_fill_2 FILLER_40_442 ();
 sg13g2_fill_1 FILLER_40_444 ();
 sg13g2_fill_1 FILLER_40_487 ();
 sg13g2_fill_2 FILLER_40_505 ();
 sg13g2_fill_1 FILLER_40_524 ();
 sg13g2_decap_8 FILLER_40_534 ();
 sg13g2_decap_4 FILLER_40_541 ();
 sg13g2_fill_1 FILLER_40_545 ();
 sg13g2_fill_2 FILLER_40_588 ();
 sg13g2_fill_1 FILLER_40_590 ();
 sg13g2_fill_1 FILLER_40_629 ();
 sg13g2_fill_2 FILLER_40_693 ();
 sg13g2_fill_1 FILLER_40_695 ();
 sg13g2_fill_2 FILLER_40_728 ();
 sg13g2_fill_1 FILLER_40_747 ();
 sg13g2_fill_1 FILLER_40_755 ();
 sg13g2_fill_2 FILLER_40_783 ();
 sg13g2_fill_1 FILLER_40_785 ();
 sg13g2_fill_2 FILLER_40_795 ();
 sg13g2_fill_2 FILLER_40_809 ();
 sg13g2_fill_1 FILLER_40_811 ();
 sg13g2_fill_1 FILLER_40_819 ();
 sg13g2_fill_1 FILLER_40_830 ();
 sg13g2_decap_8 FILLER_40_836 ();
 sg13g2_fill_2 FILLER_40_843 ();
 sg13g2_decap_8 FILLER_40_861 ();
 sg13g2_decap_8 FILLER_40_868 ();
 sg13g2_fill_1 FILLER_40_911 ();
 sg13g2_fill_1 FILLER_40_957 ();
 sg13g2_decap_8 FILLER_40_966 ();
 sg13g2_decap_8 FILLER_40_973 ();
 sg13g2_decap_8 FILLER_40_980 ();
 sg13g2_decap_8 FILLER_40_987 ();
 sg13g2_decap_8 FILLER_40_994 ();
 sg13g2_decap_8 FILLER_40_1001 ();
 sg13g2_decap_8 FILLER_40_1008 ();
 sg13g2_decap_8 FILLER_40_1015 ();
 sg13g2_decap_8 FILLER_40_1022 ();
 sg13g2_fill_1 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_35 ();
 sg13g2_fill_2 FILLER_41_67 ();
 sg13g2_fill_1 FILLER_41_69 ();
 sg13g2_fill_2 FILLER_41_99 ();
 sg13g2_fill_1 FILLER_41_101 ();
 sg13g2_fill_2 FILLER_41_147 ();
 sg13g2_fill_1 FILLER_41_149 ();
 sg13g2_fill_2 FILLER_41_155 ();
 sg13g2_fill_2 FILLER_41_211 ();
 sg13g2_fill_2 FILLER_41_233 ();
 sg13g2_fill_1 FILLER_41_235 ();
 sg13g2_fill_1 FILLER_41_329 ();
 sg13g2_fill_1 FILLER_41_420 ();
 sg13g2_fill_1 FILLER_41_439 ();
 sg13g2_fill_2 FILLER_41_461 ();
 sg13g2_fill_2 FILLER_41_481 ();
 sg13g2_fill_1 FILLER_41_483 ();
 sg13g2_fill_1 FILLER_41_489 ();
 sg13g2_fill_2 FILLER_41_495 ();
 sg13g2_fill_1 FILLER_41_538 ();
 sg13g2_fill_1 FILLER_41_556 ();
 sg13g2_fill_1 FILLER_41_625 ();
 sg13g2_fill_2 FILLER_41_651 ();
 sg13g2_fill_1 FILLER_41_653 ();
 sg13g2_fill_1 FILLER_41_690 ();
 sg13g2_fill_1 FILLER_41_703 ();
 sg13g2_fill_2 FILLER_41_716 ();
 sg13g2_decap_4 FILLER_41_730 ();
 sg13g2_fill_2 FILLER_41_744 ();
 sg13g2_fill_1 FILLER_41_746 ();
 sg13g2_fill_2 FILLER_41_777 ();
 sg13g2_fill_1 FILLER_41_779 ();
 sg13g2_fill_2 FILLER_41_801 ();
 sg13g2_fill_1 FILLER_41_803 ();
 sg13g2_decap_4 FILLER_41_829 ();
 sg13g2_fill_1 FILLER_41_833 ();
 sg13g2_fill_1 FILLER_41_838 ();
 sg13g2_decap_8 FILLER_41_860 ();
 sg13g2_decap_8 FILLER_41_867 ();
 sg13g2_fill_1 FILLER_41_874 ();
 sg13g2_fill_2 FILLER_41_883 ();
 sg13g2_fill_2 FILLER_41_912 ();
 sg13g2_decap_8 FILLER_41_972 ();
 sg13g2_decap_8 FILLER_41_979 ();
 sg13g2_decap_8 FILLER_41_986 ();
 sg13g2_decap_8 FILLER_41_993 ();
 sg13g2_decap_8 FILLER_41_1000 ();
 sg13g2_decap_8 FILLER_41_1007 ();
 sg13g2_decap_8 FILLER_41_1014 ();
 sg13g2_decap_8 FILLER_41_1021 ();
 sg13g2_fill_1 FILLER_41_1028 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_88 ();
 sg13g2_fill_1 FILLER_42_90 ();
 sg13g2_fill_2 FILLER_42_98 ();
 sg13g2_fill_1 FILLER_42_136 ();
 sg13g2_fill_1 FILLER_42_194 ();
 sg13g2_fill_2 FILLER_42_200 ();
 sg13g2_fill_1 FILLER_42_202 ();
 sg13g2_fill_1 FILLER_42_237 ();
 sg13g2_fill_2 FILLER_42_282 ();
 sg13g2_fill_1 FILLER_42_311 ();
 sg13g2_fill_1 FILLER_42_326 ();
 sg13g2_fill_2 FILLER_42_402 ();
 sg13g2_fill_1 FILLER_42_404 ();
 sg13g2_fill_2 FILLER_42_502 ();
 sg13g2_fill_1 FILLER_42_562 ();
 sg13g2_fill_2 FILLER_42_621 ();
 sg13g2_fill_2 FILLER_42_686 ();
 sg13g2_fill_1 FILLER_42_708 ();
 sg13g2_fill_1 FILLER_42_717 ();
 sg13g2_fill_2 FILLER_42_735 ();
 sg13g2_fill_1 FILLER_42_737 ();
 sg13g2_fill_2 FILLER_42_759 ();
 sg13g2_fill_1 FILLER_42_769 ();
 sg13g2_fill_1 FILLER_42_788 ();
 sg13g2_fill_1 FILLER_42_814 ();
 sg13g2_decap_4 FILLER_42_824 ();
 sg13g2_fill_1 FILLER_42_856 ();
 sg13g2_fill_1 FILLER_42_888 ();
 sg13g2_fill_2 FILLER_42_911 ();
 sg13g2_decap_8 FILLER_42_976 ();
 sg13g2_decap_8 FILLER_42_983 ();
 sg13g2_decap_8 FILLER_42_990 ();
 sg13g2_decap_8 FILLER_42_997 ();
 sg13g2_decap_8 FILLER_42_1004 ();
 sg13g2_decap_8 FILLER_42_1011 ();
 sg13g2_decap_8 FILLER_42_1018 ();
 sg13g2_decap_4 FILLER_42_1025 ();
 sg13g2_fill_1 FILLER_43_11 ();
 sg13g2_fill_2 FILLER_43_32 ();
 sg13g2_fill_1 FILLER_43_34 ();
 sg13g2_fill_2 FILLER_43_48 ();
 sg13g2_fill_1 FILLER_43_50 ();
 sg13g2_fill_2 FILLER_43_63 ();
 sg13g2_fill_2 FILLER_43_79 ();
 sg13g2_fill_1 FILLER_43_124 ();
 sg13g2_fill_2 FILLER_43_130 ();
 sg13g2_fill_2 FILLER_43_139 ();
 sg13g2_fill_1 FILLER_43_141 ();
 sg13g2_fill_2 FILLER_43_147 ();
 sg13g2_fill_1 FILLER_43_149 ();
 sg13g2_fill_2 FILLER_43_177 ();
 sg13g2_fill_1 FILLER_43_179 ();
 sg13g2_fill_1 FILLER_43_212 ();
 sg13g2_fill_2 FILLER_43_217 ();
 sg13g2_fill_1 FILLER_43_254 ();
 sg13g2_fill_2 FILLER_43_262 ();
 sg13g2_fill_2 FILLER_43_377 ();
 sg13g2_fill_2 FILLER_43_447 ();
 sg13g2_fill_1 FILLER_43_449 ();
 sg13g2_fill_1 FILLER_43_455 ();
 sg13g2_fill_2 FILLER_43_469 ();
 sg13g2_fill_1 FILLER_43_492 ();
 sg13g2_fill_1 FILLER_43_512 ();
 sg13g2_fill_1 FILLER_43_527 ();
 sg13g2_fill_1 FILLER_43_574 ();
 sg13g2_fill_2 FILLER_43_605 ();
 sg13g2_fill_1 FILLER_43_607 ();
 sg13g2_fill_1 FILLER_43_627 ();
 sg13g2_fill_2 FILLER_43_701 ();
 sg13g2_fill_1 FILLER_43_703 ();
 sg13g2_fill_2 FILLER_43_745 ();
 sg13g2_fill_2 FILLER_43_774 ();
 sg13g2_fill_2 FILLER_43_798 ();
 sg13g2_fill_2 FILLER_43_821 ();
 sg13g2_fill_1 FILLER_43_823 ();
 sg13g2_fill_2 FILLER_43_837 ();
 sg13g2_fill_2 FILLER_43_844 ();
 sg13g2_fill_1 FILLER_43_846 ();
 sg13g2_decap_4 FILLER_43_889 ();
 sg13g2_fill_1 FILLER_43_893 ();
 sg13g2_decap_4 FILLER_43_930 ();
 sg13g2_fill_2 FILLER_43_934 ();
 sg13g2_decap_8 FILLER_43_972 ();
 sg13g2_decap_8 FILLER_43_979 ();
 sg13g2_decap_8 FILLER_43_986 ();
 sg13g2_decap_8 FILLER_43_993 ();
 sg13g2_decap_8 FILLER_43_1000 ();
 sg13g2_decap_8 FILLER_43_1007 ();
 sg13g2_decap_8 FILLER_43_1014 ();
 sg13g2_decap_8 FILLER_43_1021 ();
 sg13g2_fill_1 FILLER_43_1028 ();
 sg13g2_fill_1 FILLER_44_12 ();
 sg13g2_fill_1 FILLER_44_21 ();
 sg13g2_fill_2 FILLER_44_37 ();
 sg13g2_fill_2 FILLER_44_66 ();
 sg13g2_fill_1 FILLER_44_104 ();
 sg13g2_fill_2 FILLER_44_122 ();
 sg13g2_fill_1 FILLER_44_151 ();
 sg13g2_fill_2 FILLER_44_199 ();
 sg13g2_fill_1 FILLER_44_234 ();
 sg13g2_fill_1 FILLER_44_269 ();
 sg13g2_fill_1 FILLER_44_301 ();
 sg13g2_fill_2 FILLER_44_314 ();
 sg13g2_fill_1 FILLER_44_316 ();
 sg13g2_fill_2 FILLER_44_395 ();
 sg13g2_fill_2 FILLER_44_414 ();
 sg13g2_fill_1 FILLER_44_416 ();
 sg13g2_fill_1 FILLER_44_458 ();
 sg13g2_fill_1 FILLER_44_486 ();
 sg13g2_fill_2 FILLER_44_496 ();
 sg13g2_fill_2 FILLER_44_562 ();
 sg13g2_fill_1 FILLER_44_585 ();
 sg13g2_fill_1 FILLER_44_600 ();
 sg13g2_fill_1 FILLER_44_609 ();
 sg13g2_fill_2 FILLER_44_637 ();
 sg13g2_fill_2 FILLER_44_679 ();
 sg13g2_fill_1 FILLER_44_681 ();
 sg13g2_fill_2 FILLER_44_799 ();
 sg13g2_decap_8 FILLER_44_825 ();
 sg13g2_decap_4 FILLER_44_832 ();
 sg13g2_fill_1 FILLER_44_836 ();
 sg13g2_fill_1 FILLER_44_850 ();
 sg13g2_fill_2 FILLER_44_860 ();
 sg13g2_fill_1 FILLER_44_862 ();
 sg13g2_fill_2 FILLER_44_868 ();
 sg13g2_decap_8 FILLER_44_964 ();
 sg13g2_decap_8 FILLER_44_971 ();
 sg13g2_decap_8 FILLER_44_978 ();
 sg13g2_decap_8 FILLER_44_985 ();
 sg13g2_decap_8 FILLER_44_992 ();
 sg13g2_decap_8 FILLER_44_999 ();
 sg13g2_decap_8 FILLER_44_1006 ();
 sg13g2_decap_8 FILLER_44_1013 ();
 sg13g2_decap_8 FILLER_44_1020 ();
 sg13g2_fill_2 FILLER_44_1027 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_2 ();
 sg13g2_fill_2 FILLER_45_13 ();
 sg13g2_fill_1 FILLER_45_32 ();
 sg13g2_fill_2 FILLER_45_43 ();
 sg13g2_fill_1 FILLER_45_45 ();
 sg13g2_fill_2 FILLER_45_80 ();
 sg13g2_fill_2 FILLER_45_98 ();
 sg13g2_fill_1 FILLER_45_129 ();
 sg13g2_fill_2 FILLER_45_166 ();
 sg13g2_fill_1 FILLER_45_168 ();
 sg13g2_fill_2 FILLER_45_202 ();
 sg13g2_fill_2 FILLER_45_220 ();
 sg13g2_fill_1 FILLER_45_222 ();
 sg13g2_fill_2 FILLER_45_252 ();
 sg13g2_fill_1 FILLER_45_272 ();
 sg13g2_fill_1 FILLER_45_301 ();
 sg13g2_fill_2 FILLER_45_315 ();
 sg13g2_fill_1 FILLER_45_333 ();
 sg13g2_fill_2 FILLER_45_367 ();
 sg13g2_fill_2 FILLER_45_390 ();
 sg13g2_fill_2 FILLER_45_446 ();
 sg13g2_fill_1 FILLER_45_448 ();
 sg13g2_fill_2 FILLER_45_472 ();
 sg13g2_fill_1 FILLER_45_500 ();
 sg13g2_fill_2 FILLER_45_540 ();
 sg13g2_fill_1 FILLER_45_542 ();
 sg13g2_fill_2 FILLER_45_566 ();
 sg13g2_fill_2 FILLER_45_606 ();
 sg13g2_fill_1 FILLER_45_608 ();
 sg13g2_fill_1 FILLER_45_627 ();
 sg13g2_fill_1 FILLER_45_669 ();
 sg13g2_fill_2 FILLER_45_692 ();
 sg13g2_fill_1 FILLER_45_694 ();
 sg13g2_fill_1 FILLER_45_732 ();
 sg13g2_fill_1 FILLER_45_737 ();
 sg13g2_fill_1 FILLER_45_742 ();
 sg13g2_fill_1 FILLER_45_749 ();
 sg13g2_fill_2 FILLER_45_755 ();
 sg13g2_fill_1 FILLER_45_774 ();
 sg13g2_fill_1 FILLER_45_783 ();
 sg13g2_fill_2 FILLER_45_792 ();
 sg13g2_fill_1 FILLER_45_794 ();
 sg13g2_fill_2 FILLER_45_800 ();
 sg13g2_fill_2 FILLER_45_810 ();
 sg13g2_fill_2 FILLER_45_833 ();
 sg13g2_fill_1 FILLER_45_843 ();
 sg13g2_decap_8 FILLER_45_865 ();
 sg13g2_fill_2 FILLER_45_884 ();
 sg13g2_decap_8 FILLER_45_894 ();
 sg13g2_fill_1 FILLER_45_901 ();
 sg13g2_decap_8 FILLER_45_929 ();
 sg13g2_fill_1 FILLER_45_936 ();
 sg13g2_decap_8 FILLER_45_965 ();
 sg13g2_decap_8 FILLER_45_972 ();
 sg13g2_decap_8 FILLER_45_979 ();
 sg13g2_decap_8 FILLER_45_986 ();
 sg13g2_decap_8 FILLER_45_993 ();
 sg13g2_decap_8 FILLER_45_1000 ();
 sg13g2_decap_8 FILLER_45_1007 ();
 sg13g2_decap_8 FILLER_45_1014 ();
 sg13g2_decap_8 FILLER_45_1021 ();
 sg13g2_fill_1 FILLER_45_1028 ();
 sg13g2_fill_1 FILLER_46_87 ();
 sg13g2_fill_2 FILLER_46_103 ();
 sg13g2_fill_2 FILLER_46_110 ();
 sg13g2_fill_2 FILLER_46_122 ();
 sg13g2_fill_2 FILLER_46_141 ();
 sg13g2_fill_1 FILLER_46_143 ();
 sg13g2_fill_1 FILLER_46_164 ();
 sg13g2_fill_2 FILLER_46_185 ();
 sg13g2_fill_1 FILLER_46_193 ();
 sg13g2_fill_1 FILLER_46_215 ();
 sg13g2_fill_1 FILLER_46_221 ();
 sg13g2_fill_1 FILLER_46_288 ();
 sg13g2_fill_1 FILLER_46_301 ();
 sg13g2_fill_1 FILLER_46_335 ();
 sg13g2_fill_2 FILLER_46_344 ();
 sg13g2_fill_2 FILLER_46_354 ();
 sg13g2_fill_1 FILLER_46_369 ();
 sg13g2_fill_1 FILLER_46_374 ();
 sg13g2_fill_2 FILLER_46_457 ();
 sg13g2_fill_1 FILLER_46_459 ();
 sg13g2_fill_1 FILLER_46_500 ();
 sg13g2_fill_2 FILLER_46_506 ();
 sg13g2_fill_1 FILLER_46_508 ();
 sg13g2_fill_1 FILLER_46_550 ();
 sg13g2_fill_1 FILLER_46_560 ();
 sg13g2_fill_1 FILLER_46_576 ();
 sg13g2_fill_2 FILLER_46_581 ();
 sg13g2_fill_1 FILLER_46_583 ();
 sg13g2_fill_1 FILLER_46_607 ();
 sg13g2_fill_1 FILLER_46_642 ();
 sg13g2_fill_2 FILLER_46_730 ();
 sg13g2_fill_1 FILLER_46_742 ();
 sg13g2_fill_2 FILLER_46_760 ();
 sg13g2_fill_2 FILLER_46_784 ();
 sg13g2_fill_1 FILLER_46_800 ();
 sg13g2_fill_2 FILLER_46_806 ();
 sg13g2_fill_2 FILLER_46_833 ();
 sg13g2_fill_1 FILLER_46_835 ();
 sg13g2_decap_4 FILLER_46_841 ();
 sg13g2_decap_8 FILLER_46_853 ();
 sg13g2_decap_4 FILLER_46_860 ();
 sg13g2_decap_8 FILLER_46_897 ();
 sg13g2_fill_2 FILLER_46_904 ();
 sg13g2_fill_1 FILLER_46_906 ();
 sg13g2_decap_8 FILLER_46_952 ();
 sg13g2_decap_8 FILLER_46_959 ();
 sg13g2_decap_8 FILLER_46_966 ();
 sg13g2_decap_8 FILLER_46_973 ();
 sg13g2_decap_8 FILLER_46_980 ();
 sg13g2_decap_8 FILLER_46_987 ();
 sg13g2_decap_8 FILLER_46_994 ();
 sg13g2_decap_8 FILLER_46_1001 ();
 sg13g2_decap_8 FILLER_46_1008 ();
 sg13g2_decap_8 FILLER_46_1015 ();
 sg13g2_decap_8 FILLER_46_1022 ();
 sg13g2_fill_2 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_44 ();
 sg13g2_fill_2 FILLER_47_83 ();
 sg13g2_fill_2 FILLER_47_105 ();
 sg13g2_fill_2 FILLER_47_112 ();
 sg13g2_fill_2 FILLER_47_139 ();
 sg13g2_fill_2 FILLER_47_225 ();
 sg13g2_fill_2 FILLER_47_275 ();
 sg13g2_fill_1 FILLER_47_277 ();
 sg13g2_fill_1 FILLER_47_293 ();
 sg13g2_fill_2 FILLER_47_335 ();
 sg13g2_fill_2 FILLER_47_423 ();
 sg13g2_fill_1 FILLER_47_425 ();
 sg13g2_fill_2 FILLER_47_485 ();
 sg13g2_fill_2 FILLER_47_506 ();
 sg13g2_fill_1 FILLER_47_508 ();
 sg13g2_fill_2 FILLER_47_598 ();
 sg13g2_fill_1 FILLER_47_709 ();
 sg13g2_fill_2 FILLER_47_731 ();
 sg13g2_fill_2 FILLER_47_739 ();
 sg13g2_fill_1 FILLER_47_747 ();
 sg13g2_fill_2 FILLER_47_753 ();
 sg13g2_fill_2 FILLER_47_760 ();
 sg13g2_fill_1 FILLER_47_762 ();
 sg13g2_fill_2 FILLER_47_771 ();
 sg13g2_fill_1 FILLER_47_814 ();
 sg13g2_fill_2 FILLER_47_822 ();
 sg13g2_fill_2 FILLER_47_837 ();
 sg13g2_fill_1 FILLER_47_839 ();
 sg13g2_fill_2 FILLER_47_858 ();
 sg13g2_fill_2 FILLER_47_922 ();
 sg13g2_fill_1 FILLER_47_924 ();
 sg13g2_decap_8 FILLER_47_938 ();
 sg13g2_decap_8 FILLER_47_945 ();
 sg13g2_decap_8 FILLER_47_952 ();
 sg13g2_decap_8 FILLER_47_959 ();
 sg13g2_decap_8 FILLER_47_966 ();
 sg13g2_decap_8 FILLER_47_973 ();
 sg13g2_decap_8 FILLER_47_980 ();
 sg13g2_decap_8 FILLER_47_987 ();
 sg13g2_decap_8 FILLER_47_994 ();
 sg13g2_decap_8 FILLER_47_1001 ();
 sg13g2_decap_8 FILLER_47_1008 ();
 sg13g2_decap_8 FILLER_47_1015 ();
 sg13g2_decap_8 FILLER_47_1022 ();
 sg13g2_fill_2 FILLER_48_8 ();
 sg13g2_fill_2 FILLER_48_64 ();
 sg13g2_fill_2 FILLER_48_92 ();
 sg13g2_fill_1 FILLER_48_94 ();
 sg13g2_fill_2 FILLER_48_111 ();
 sg13g2_fill_2 FILLER_48_139 ();
 sg13g2_fill_2 FILLER_48_164 ();
 sg13g2_fill_1 FILLER_48_174 ();
 sg13g2_fill_1 FILLER_48_192 ();
 sg13g2_fill_1 FILLER_48_327 ();
 sg13g2_fill_2 FILLER_48_346 ();
 sg13g2_fill_1 FILLER_48_348 ();
 sg13g2_fill_1 FILLER_48_386 ();
 sg13g2_fill_1 FILLER_48_503 ();
 sg13g2_fill_1 FILLER_48_537 ();
 sg13g2_fill_2 FILLER_48_742 ();
 sg13g2_fill_2 FILLER_48_772 ();
 sg13g2_fill_1 FILLER_48_774 ();
 sg13g2_fill_1 FILLER_48_780 ();
 sg13g2_fill_2 FILLER_48_810 ();
 sg13g2_fill_1 FILLER_48_812 ();
 sg13g2_fill_2 FILLER_48_821 ();
 sg13g2_fill_1 FILLER_48_823 ();
 sg13g2_fill_2 FILLER_48_840 ();
 sg13g2_decap_4 FILLER_48_847 ();
 sg13g2_fill_1 FILLER_48_859 ();
 sg13g2_fill_1 FILLER_48_876 ();
 sg13g2_decap_8 FILLER_48_898 ();
 sg13g2_decap_8 FILLER_48_905 ();
 sg13g2_decap_8 FILLER_48_912 ();
 sg13g2_decap_8 FILLER_48_928 ();
 sg13g2_decap_8 FILLER_48_935 ();
 sg13g2_decap_8 FILLER_48_942 ();
 sg13g2_decap_8 FILLER_48_949 ();
 sg13g2_decap_8 FILLER_48_956 ();
 sg13g2_decap_8 FILLER_48_963 ();
 sg13g2_decap_8 FILLER_48_970 ();
 sg13g2_decap_8 FILLER_48_977 ();
 sg13g2_decap_8 FILLER_48_984 ();
 sg13g2_decap_8 FILLER_48_991 ();
 sg13g2_decap_8 FILLER_48_998 ();
 sg13g2_decap_8 FILLER_48_1005 ();
 sg13g2_decap_8 FILLER_48_1012 ();
 sg13g2_decap_8 FILLER_48_1019 ();
 sg13g2_fill_2 FILLER_48_1026 ();
 sg13g2_fill_1 FILLER_48_1028 ();
 sg13g2_fill_1 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_23 ();
 sg13g2_fill_1 FILLER_49_25 ();
 sg13g2_fill_2 FILLER_49_31 ();
 sg13g2_fill_1 FILLER_49_33 ();
 sg13g2_fill_1 FILLER_49_44 ();
 sg13g2_fill_2 FILLER_49_50 ();
 sg13g2_fill_1 FILLER_49_57 ();
 sg13g2_fill_1 FILLER_49_76 ();
 sg13g2_fill_2 FILLER_49_87 ();
 sg13g2_fill_1 FILLER_49_89 ();
 sg13g2_fill_2 FILLER_49_111 ();
 sg13g2_fill_2 FILLER_49_132 ();
 sg13g2_fill_1 FILLER_49_134 ();
 sg13g2_fill_1 FILLER_49_156 ();
 sg13g2_fill_1 FILLER_49_163 ();
 sg13g2_fill_1 FILLER_49_185 ();
 sg13g2_fill_2 FILLER_49_211 ();
 sg13g2_fill_2 FILLER_49_221 ();
 sg13g2_fill_2 FILLER_49_245 ();
 sg13g2_fill_2 FILLER_49_267 ();
 sg13g2_fill_2 FILLER_49_276 ();
 sg13g2_fill_1 FILLER_49_278 ();
 sg13g2_fill_1 FILLER_49_298 ();
 sg13g2_fill_2 FILLER_49_333 ();
 sg13g2_fill_2 FILLER_49_344 ();
 sg13g2_fill_1 FILLER_49_363 ();
 sg13g2_fill_1 FILLER_49_413 ();
 sg13g2_fill_1 FILLER_49_455 ();
 sg13g2_fill_1 FILLER_49_484 ();
 sg13g2_fill_2 FILLER_49_550 ();
 sg13g2_fill_2 FILLER_49_562 ();
 sg13g2_fill_2 FILLER_49_622 ();
 sg13g2_fill_2 FILLER_49_665 ();
 sg13g2_fill_1 FILLER_49_667 ();
 sg13g2_fill_2 FILLER_49_690 ();
 sg13g2_fill_1 FILLER_49_692 ();
 sg13g2_fill_1 FILLER_49_711 ();
 sg13g2_fill_2 FILLER_49_745 ();
 sg13g2_fill_2 FILLER_49_784 ();
 sg13g2_fill_1 FILLER_49_786 ();
 sg13g2_fill_2 FILLER_49_799 ();
 sg13g2_fill_1 FILLER_49_801 ();
 sg13g2_fill_2 FILLER_49_807 ();
 sg13g2_fill_2 FILLER_49_820 ();
 sg13g2_decap_8 FILLER_49_843 ();
 sg13g2_fill_1 FILLER_49_850 ();
 sg13g2_decap_4 FILLER_49_856 ();
 sg13g2_fill_2 FILLER_49_864 ();
 sg13g2_decap_8 FILLER_49_871 ();
 sg13g2_fill_2 FILLER_49_878 ();
 sg13g2_decap_8 FILLER_49_889 ();
 sg13g2_decap_8 FILLER_49_896 ();
 sg13g2_decap_8 FILLER_49_903 ();
 sg13g2_decap_8 FILLER_49_910 ();
 sg13g2_decap_8 FILLER_49_917 ();
 sg13g2_decap_8 FILLER_49_924 ();
 sg13g2_decap_8 FILLER_49_931 ();
 sg13g2_decap_8 FILLER_49_938 ();
 sg13g2_decap_8 FILLER_49_945 ();
 sg13g2_decap_8 FILLER_49_952 ();
 sg13g2_decap_8 FILLER_49_959 ();
 sg13g2_decap_8 FILLER_49_966 ();
 sg13g2_decap_8 FILLER_49_973 ();
 sg13g2_decap_8 FILLER_49_980 ();
 sg13g2_decap_8 FILLER_49_987 ();
 sg13g2_decap_8 FILLER_49_994 ();
 sg13g2_decap_8 FILLER_49_1001 ();
 sg13g2_decap_8 FILLER_49_1008 ();
 sg13g2_decap_8 FILLER_49_1015 ();
 sg13g2_decap_8 FILLER_49_1022 ();
 assign uio_oe[0] = net33;
 assign uio_oe[1] = net34;
 assign uio_oe[2] = net35;
 assign uio_oe[3] = net36;
 assign uio_oe[4] = net37;
 assign uio_oe[5] = net38;
 assign uio_oe[6] = net39;
 assign uio_oe[7] = net40;
endmodule
