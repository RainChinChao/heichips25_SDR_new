* NGSPICE file created from heichips25_template.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_2 abstract view
.subckt sg13g2_and3_2 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_8 abstract view
.subckt sg13g2_inv_8 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

.subckt heichips25_template VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
XFILLER_39_222 VPWR VGND sg13g2_fill_2
XFILLER_39_244 VPWR VGND sg13g2_decap_8
X_3155_ net540 VGND VPWR net103 mac1.sum_lvl2_ff\[10\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_3086_ net526 VGND VPWR _0069_ mac1.products_ff\[73\] clknet_leaf_26_clk sg13g2_dfrbpq_1
X_2106_ _1390_ net450 net390 VPWR VGND sg13g2_nand2_1
XFILLER_39_288 VPWR VGND sg13g2_fill_1
X_2037_ _1328_ _1329_ _0019_ VPWR VGND sg13g2_and2_1
XFILLER_36_984 VPWR VGND sg13g2_decap_8
XFILLER_10_317 VPWR VGND sg13g2_decap_8
XFILLER_23_667 VPWR VGND sg13g2_decap_8
XFILLER_22_188 VPWR VGND sg13g2_decap_8
X_2939_ net485 net371 _0823_ VPWR VGND sg13g2_nor2_1
XFILLER_7_7 VPWR VGND sg13g2_decap_4
XFILLER_46_715 VPWR VGND sg13g2_fill_1
XFILLER_19_929 VPWR VGND sg13g2_decap_8
XFILLER_46_737 VPWR VGND sg13g2_decap_8
XFILLER_18_428 VPWR VGND sg13g2_decap_8
XFILLER_26_63 VPWR VGND sg13g2_decap_8
XFILLER_27_995 VPWR VGND sg13g2_decap_8
XFILLER_42_965 VPWR VGND sg13g2_decap_8
XFILLER_41_431 VPWR VGND sg13g2_decap_8
XFILLER_14_634 VPWR VGND sg13g2_decap_4
XFILLER_14_678 VPWR VGND sg13g2_fill_2
XFILLER_9_126 VPWR VGND sg13g2_decap_8
XFILLER_6_811 VPWR VGND sg13g2_decap_8
XFILLER_10_873 VPWR VGND sg13g2_decap_8
XFILLER_5_310 VPWR VGND sg13g2_decap_8
XFILLER_6_888 VPWR VGND sg13g2_decap_8
XFILLER_49_520 VPWR VGND sg13g2_decap_8
XFILLER_3_89 VPWR VGND sg13g2_decap_8
XFILLER_3_1018 VPWR VGND sg13g2_decap_8
XFILLER_37_759 VPWR VGND sg13g2_decap_8
XFILLER_18_951 VPWR VGND sg13g2_decap_8
XFILLER_45_781 VPWR VGND sg13g2_fill_1
XFILLER_33_910 VPWR VGND sg13g2_decap_8
XFILLER_33_987 VPWR VGND sg13g2_decap_8
XFILLER_20_626 VPWR VGND sg13g2_decap_4
XFILLER_32_497 VPWR VGND sg13g2_fill_2
XFILLER_20_659 VPWR VGND sg13g2_decap_8
X_2724_ _0620_ net479 net426 VPWR VGND sg13g2_nand2_1
XFILLER_8_170 VPWR VGND sg13g2_fill_1
X_2655_ _0518_ VPWR _0553_ VGND _0509_ _0519_ sg13g2_o21ai_1
X_1606_ _0936_ _0937_ _0927_ _0938_ VPWR VGND sg13g2_nand3_1
X_2586_ _0417_ VPWR _0486_ VGND _0482_ _0484_ sg13g2_o21ai_1
X_1537_ _0871_ net470 net410 VPWR VGND sg13g2_nand2_1
X_3207_ net530 VGND VPWR net110 mac1.sum_lvl1_ff\[86\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_3138_ net542 VGND VPWR net84 mac1.sum_lvl1_ff\[45\] clknet_leaf_24_clk sg13g2_dfrbpq_1
XFILLER_43_707 VPWR VGND sg13g2_decap_4
XFILLER_43_729 VPWR VGND sg13g2_decap_8
XFILLER_42_206 VPWR VGND sg13g2_decap_4
X_3069_ net548 VGND VPWR _0122_ DP_2.matrix\[40\] clknet_leaf_21_clk sg13g2_dfrbpq_1
XFILLER_23_420 VPWR VGND sg13g2_decap_8
XFILLER_24_943 VPWR VGND sg13g2_decap_8
XFILLER_3_836 VPWR VGND sg13g2_decap_8
Xhold170 DP_1.matrix\[40\] VPWR VGND net210 sg13g2_dlygate4sd3_1
Xhold192 _1330_ VPWR VGND net232 sg13g2_dlygate4sd3_1
Xhold181 DP_2.matrix\[1\] VPWR VGND net221 sg13g2_dlygate4sd3_1
XFILLER_15_921 VPWR VGND sg13g2_decap_8
XFILLER_42_740 VPWR VGND sg13g2_fill_2
XFILLER_14_420 VPWR VGND sg13g2_decap_8
XFILLER_15_998 VPWR VGND sg13g2_decap_8
XFILLER_30_913 VPWR VGND sg13g2_decap_8
XFILLER_14_475 VPWR VGND sg13g2_fill_1
XFILLER_6_685 VPWR VGND sg13g2_decap_8
X_2440_ _0345_ net492 net431 VPWR VGND sg13g2_nand2_1
X_2371_ VGND VPWR _0281_ _0280_ _0268_ sg13g2_or2_1
XFILLER_38_4 VPWR VGND sg13g2_decap_4
XFILLER_49_361 VPWR VGND sg13g2_decap_8
XFILLER_37_556 VPWR VGND sg13g2_decap_8
XFILLER_24_217 VPWR VGND sg13g2_decap_8
XFILLER_32_250 VPWR VGND sg13g2_fill_1
XFILLER_33_773 VPWR VGND sg13g2_decap_8
XFILLER_21_924 VPWR VGND sg13g2_decap_8
XFILLER_20_478 VPWR VGND sg13g2_decap_8
X_2707_ _0603_ _0591_ _0604_ VPWR VGND sg13g2_xor2_1
X_2638_ _0537_ _0535_ _0536_ VPWR VGND sg13g2_nand2_1
X_2569_ _0469_ net434 net479 net477 net438 VPWR VGND sg13g2_a22oi_1
XFILLER_0_839 VPWR VGND sg13g2_decap_8
XFILLER_28_523 VPWR VGND sg13g2_fill_1
XFILLER_16_707 VPWR VGND sg13g2_decap_8
XFILLER_43_504 VPWR VGND sg13g2_decap_8
XFILLER_16_718 VPWR VGND sg13g2_fill_1
XFILLER_24_762 VPWR VGND sg13g2_decap_8
XFILLER_24_795 VPWR VGND sg13g2_decap_8
XFILLER_8_928 VPWR VGND sg13g2_decap_8
XFILLER_11_434 VPWR VGND sg13g2_fill_2
XFILLER_12_968 VPWR VGND sg13g2_decap_8
XFILLER_23_64 VPWR VGND sg13g2_decap_4
XFILLER_11_467 VPWR VGND sg13g2_decap_8
XFILLER_23_75 VPWR VGND sg13g2_decap_8
XFILLER_3_633 VPWR VGND sg13g2_decap_8
XFILLER_2_143 VPWR VGND sg13g2_fill_1
XFILLER_2_176 VPWR VGND sg13g2_decap_8
Xfanout480 DP_1.matrix\[6\] net480 VPWR VGND sg13g2_buf_8
Xfanout491 DP_1.matrix\[1\] net491 VPWR VGND sg13g2_buf_8
XFILLER_47_843 VPWR VGND sg13g2_decap_8
XFILLER_46_342 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_19_567 VPWR VGND sg13g2_fill_1
XFILLER_34_548 VPWR VGND sg13g2_fill_2
XFILLER_9_11 VPWR VGND sg13g2_decap_4
X_1940_ _1248_ _1251_ net284 _1253_ VPWR VGND sg13g2_nand3_1
X_1871_ _0073_ _1194_ _1195_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_754 VPWR VGND sg13g2_decap_8
XFILLER_30_765 VPWR VGND sg13g2_fill_1
XFILLER_7_994 VPWR VGND sg13g2_decap_8
X_2423_ _0330_ _0320_ _0331_ VPWR VGND sg13g2_nor2b_1
X_2354_ _0250_ _0245_ _0252_ _0264_ VPWR VGND sg13g2_a21o_1
X_2285_ _0196_ _0197_ _0198_ VPWR VGND sg13g2_nor2b_1
XFILLER_38_854 VPWR VGND sg13g2_decap_8
XFILLER_40_507 VPWR VGND sg13g2_decap_8
XFILLER_21_710 VPWR VGND sg13g2_fill_2
XFILLER_21_798 VPWR VGND sg13g2_decap_8
XFILLER_5_909 VPWR VGND sg13g2_decap_8
XFILLER_0_636 VPWR VGND sg13g2_decap_8
XFILLER_47_117 VPWR VGND sg13g2_decap_8
XFILLER_29_854 VPWR VGND sg13g2_decap_4
XFILLER_44_824 VPWR VGND sg13g2_decap_8
XFILLER_18_86 VPWR VGND sg13g2_decap_8
XFILLER_12_721 VPWR VGND sg13g2_decap_8
XFILLER_31_529 VPWR VGND sg13g2_decap_8
XFILLER_11_231 VPWR VGND sg13g2_decap_4
XFILLER_8_725 VPWR VGND sg13g2_decap_8
XFILLER_4_931 VPWR VGND sg13g2_decap_8
XFILLER_3_441 VPWR VGND sg13g2_decap_8
XFILLER_38_106 VPWR VGND sg13g2_fill_2
XFILLER_47_640 VPWR VGND sg13g2_decap_8
X_2070_ _1354_ _1355_ _1356_ VPWR VGND sg13g2_nor2b_1
XFILLER_47_673 VPWR VGND sg13g2_decap_8
XFILLER_47_651 VPWR VGND sg13g2_fill_2
X_2972_ net496 _0083_ VPWR VGND sg13g2_buf_1
X_1923_ mac1.sum_lvl2_ff\[24\] net257 _1239_ VPWR VGND sg13g2_nor2_1
XFILLER_30_573 VPWR VGND sg13g2_fill_1
X_1854_ _1179_ net459 net402 VPWR VGND sg13g2_nand2_1
X_1785_ _1112_ _1111_ _1113_ VPWR VGND sg13g2_nor2b_1
XFILLER_7_791 VPWR VGND sg13g2_decap_8
X_2406_ _0051_ _0313_ _0314_ VPWR VGND sg13g2_xnor2_1
X_2337_ VGND VPWR _0248_ _0247_ _0204_ sg13g2_or2_1
X_2268_ _0135_ VPWR _0181_ VGND _1500_ _0136_ sg13g2_o21ai_1
XFILLER_37_150 VPWR VGND sg13g2_decap_8
X_2199_ _1469_ VPWR _1480_ VGND _1447_ _1470_ sg13g2_o21ai_1
XFILLER_25_301 VPWR VGND sg13g2_decap_8
XFILLER_37_161 VPWR VGND sg13g2_fill_2
XFILLER_37_172 VPWR VGND sg13g2_decap_8
XFILLER_41_805 VPWR VGND sg13g2_fill_1
XFILLER_26_868 VPWR VGND sg13g2_decap_4
XFILLER_5_706 VPWR VGND sg13g2_decap_8
XFILLER_20_32 VPWR VGND sg13g2_decap_8
XFILLER_1_912 VPWR VGND sg13g2_decap_8
XFILLER_20_98 VPWR VGND sg13g2_decap_8
XFILLER_49_916 VPWR VGND sg13g2_decap_8
XFILLER_0_433 VPWR VGND sg13g2_decap_8
XFILLER_1_989 VPWR VGND sg13g2_decap_8
Xhold30 mac1.sum_lvl1_ff\[73\] VPWR VGND net70 sg13g2_dlygate4sd3_1
Xhold41 mac1.products_ff\[76\] VPWR VGND net81 sg13g2_dlygate4sd3_1
Xhold74 mac1.sum_lvl2_ff\[42\] VPWR VGND net114 sg13g2_dlygate4sd3_1
Xhold52 mac1.sum_lvl2_ff\[48\] VPWR VGND net92 sg13g2_dlygate4sd3_1
Xhold63 mac1.sum_lvl1_ff\[10\] VPWR VGND net103 sg13g2_dlygate4sd3_1
Xhold85 mac1.products_ff\[142\] VPWR VGND net125 sg13g2_dlygate4sd3_1
Xhold96 mac1.sum_lvl2_ff\[46\] VPWR VGND net136 sg13g2_dlygate4sd3_1
XFILLER_21_1022 VPWR VGND sg13g2_decap_8
XFILLER_45_51 VPWR VGND sg13g2_decap_8
XFILLER_44_654 VPWR VGND sg13g2_decap_4
XFILLER_17_879 VPWR VGND sg13g2_decap_8
XFILLER_45_95 VPWR VGND sg13g2_decap_8
XFILLER_31_326 VPWR VGND sg13g2_decap_4
XFILLER_31_348 VPWR VGND sg13g2_fill_1
XFILLER_8_544 VPWR VGND sg13g2_decap_8
X_1570_ _0900_ _0901_ _0895_ _0903_ VPWR VGND sg13g2_nand3_1
XFILLER_3_293 VPWR VGND sg13g2_decap_8
X_3240_ net544 VGND VPWR net170 mac1.sum_lvl3_ff\[15\] clknet_leaf_19_clk sg13g2_dfrbpq_2
X_3171_ net540 VGND VPWR net102 mac1.sum_lvl2_ff\[29\] clknet_leaf_23_clk sg13g2_dfrbpq_1
XFILLER_20_4 VPWR VGND sg13g2_decap_8
X_2122_ _1403_ _1404_ _1379_ _1406_ VPWR VGND sg13g2_nand3_1
XFILLER_48_982 VPWR VGND sg13g2_decap_8
XFILLER_26_109 VPWR VGND sg13g2_fill_2
X_2053_ _1339_ _1340_ _0033_ VPWR VGND sg13g2_nor2_1
XFILLER_23_805 VPWR VGND sg13g2_decap_4
XFILLER_34_131 VPWR VGND sg13g2_decap_8
XFILLER_16_890 VPWR VGND sg13g2_decap_8
XFILLER_22_359 VPWR VGND sg13g2_fill_1
X_2955_ _0799_ _0797_ _0833_ VPWR VGND sg13g2_xor2_1
X_2886_ net371 net253 _0776_ VPWR VGND sg13g2_nor2b_1
X_1906_ _1226_ mac1.sum_lvl2_ff\[20\] mac1.sum_lvl2_ff\[1\] VPWR VGND sg13g2_nand2_1
X_1837_ _1161_ _1149_ _1163_ VPWR VGND sg13g2_xor2_1
X_1768_ _1096_ net460 net409 DP_1.matrix\[42\] net407 VPWR VGND sg13g2_a22oi_1
X_1699_ _0954_ _1026_ _1028_ _1029_ VPWR VGND sg13g2_or3_1
XFILLER_39_960 VPWR VGND sg13g2_decap_8
XFILLER_14_849 VPWR VGND sg13g2_decap_8
XFILLER_15_32 VPWR VGND sg13g2_decap_8
XFILLER_26_676 VPWR VGND sg13g2_decap_8
XFILLER_40_178 VPWR VGND sg13g2_decap_8
XFILLER_22_882 VPWR VGND sg13g2_decap_8
XFILLER_31_42 VPWR VGND sg13g2_fill_2
Xoutput31 net31 uo_out[6] VPWR VGND sg13g2_buf_1
Xoutput20 net20 uio_out[3] VPWR VGND sg13g2_buf_1
XFILLER_49_713 VPWR VGND sg13g2_decap_8
XFILLER_0_263 VPWR VGND sg13g2_decap_8
XFILLER_1_786 VPWR VGND sg13g2_decap_8
XFILLER_48_223 VPWR VGND sg13g2_decap_8
XFILLER_45_963 VPWR VGND sg13g2_decap_8
XFILLER_16_142 VPWR VGND sg13g2_fill_2
XFILLER_31_134 VPWR VGND sg13g2_decap_8
XFILLER_32_635 VPWR VGND sg13g2_fill_2
XFILLER_31_145 VPWR VGND sg13g2_fill_2
X_2740_ _0635_ _0628_ _0636_ VPWR VGND sg13g2_nor2b_1
X_2671_ _0569_ _0553_ _0567_ VPWR VGND sg13g2_xnor2_1
XFILLER_9_886 VPWR VGND sg13g2_decap_8
X_1622_ _0951_ _0952_ _0953_ VPWR VGND sg13g2_nor2b_1
X_1553_ _0885_ _0865_ _0046_ VPWR VGND sg13g2_xor2_1
XFILLER_28_1028 VPWR VGND sg13g2_fill_1
X_3223_ net530 VGND VPWR net75 mac1.sum_lvl3_ff\[34\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_3154_ net540 VGND VPWR net68 mac1.sum_lvl2_ff\[9\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_3085_ net525 VGND VPWR _0046_ mac1.products_ff\[72\] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_2105_ _1369_ VPWR _1389_ VGND _1367_ _1370_ sg13g2_o21ai_1
XFILLER_39_278 VPWR VGND sg13g2_fill_1
X_2036_ net292 _1325_ _1327_ _1329_ VPWR VGND sg13g2_or3_1
XFILLER_36_963 VPWR VGND sg13g2_decap_8
XFILLER_23_624 VPWR VGND sg13g2_fill_2
XFILLER_22_156 VPWR VGND sg13g2_fill_1
X_2938_ VGND VPWR net372 _0822_ _0089_ _0821_ sg13g2_a21oi_1
XFILLER_11_1010 VPWR VGND sg13g2_decap_8
X_2869_ net463 _0730_ _0759_ VPWR VGND sg13g2_nor2_1
XFILLER_18_407 VPWR VGND sg13g2_decap_8
XFILLER_19_908 VPWR VGND sg13g2_decap_8
XFILLER_45_215 VPWR VGND sg13g2_fill_2
XFILLER_39_790 VPWR VGND sg13g2_fill_2
XFILLER_26_42 VPWR VGND sg13g2_decap_8
XFILLER_27_974 VPWR VGND sg13g2_decap_8
Xclkbuf_3_6__f_clk clknet_0_clk clknet_3_6__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_42_944 VPWR VGND sg13g2_decap_8
XFILLER_41_410 VPWR VGND sg13g2_decap_8
XFILLER_13_101 VPWR VGND sg13g2_fill_2
XFILLER_41_476 VPWR VGND sg13g2_fill_1
XFILLER_41_454 VPWR VGND sg13g2_decap_8
XFILLER_9_105 VPWR VGND sg13g2_decap_8
XFILLER_10_852 VPWR VGND sg13g2_decap_8
XFILLER_6_867 VPWR VGND sg13g2_decap_8
XFILLER_5_399 VPWR VGND sg13g2_fill_2
XFILLER_3_46 VPWR VGND sg13g2_decap_8
XFILLER_1_583 VPWR VGND sg13g2_decap_8
XFILLER_18_930 VPWR VGND sg13g2_decap_8
XFILLER_36_204 VPWR VGND sg13g2_decap_8
XFILLER_37_738 VPWR VGND sg13g2_decap_8
XFILLER_36_248 VPWR VGND sg13g2_decap_8
XFILLER_36_259 VPWR VGND sg13g2_fill_1
XFILLER_33_966 VPWR VGND sg13g2_decap_8
XFILLER_34_1010 VPWR VGND sg13g2_decap_8
X_2723_ _0600_ _0593_ _0562_ _0619_ VPWR VGND sg13g2_a21o_2
XFILLER_13_690 VPWR VGND sg13g2_fill_1
X_2654_ _0552_ _0542_ _0550_ VPWR VGND sg13g2_xnor2_1
X_1605_ _0934_ _0933_ _0928_ _0937_ VPWR VGND sg13g2_a21o_1
X_2585_ _0417_ _0482_ _0484_ _0485_ VPWR VGND sg13g2_or3_1
X_1536_ VGND VPWR _0870_ _0858_ _0856_ sg13g2_or2_1
XFILLER_41_1025 VPWR VGND sg13g2_decap_4
X_3206_ net529 VGND VPWR net148 mac1.sum_lvl1_ff\[85\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_3137_ net543 VGND VPWR net81 mac1.sum_lvl1_ff\[44\] clknet_leaf_25_clk sg13g2_dfrbpq_1
XFILLER_27_204 VPWR VGND sg13g2_fill_2
XFILLER_27_226 VPWR VGND sg13g2_decap_8
XFILLER_28_738 VPWR VGND sg13g2_decap_8
XFILLER_24_922 VPWR VGND sg13g2_decap_8
X_3068_ net535 VGND VPWR _0121_ DP_2.matrix\[39\] clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_36_782 VPWR VGND sg13g2_fill_2
X_2019_ _0031_ _1311_ net182 VPWR VGND sg13g2_xnor2_1
XFILLER_24_999 VPWR VGND sg13g2_decap_8
XFILLER_12_55 VPWR VGND sg13g2_decap_4
XFILLER_3_815 VPWR VGND sg13g2_decap_8
Xhold160 mac1.sum_lvl3_ff\[23\] VPWR VGND net200 sg13g2_dlygate4sd3_1
Xhold171 DP_1.matrix\[42\] VPWR VGND net211 sg13g2_dlygate4sd3_1
Xhold193 _1331_ VPWR VGND net233 sg13g2_dlygate4sd3_1
Xhold182 _0111_ VPWR VGND net222 sg13g2_dlygate4sd3_1
XFILLER_46_579 VPWR VGND sg13g2_decap_8
XFILLER_15_900 VPWR VGND sg13g2_decap_8
XFILLER_42_774 VPWR VGND sg13g2_fill_1
XFILLER_14_454 VPWR VGND sg13g2_decap_4
XFILLER_15_977 VPWR VGND sg13g2_decap_8
XFILLER_30_969 VPWR VGND sg13g2_decap_8
XFILLER_6_664 VPWR VGND sg13g2_decap_8
X_2370_ _0278_ _0269_ _0280_ VPWR VGND sg13g2_xor2_1
XFILLER_2_881 VPWR VGND sg13g2_decap_8
XFILLER_49_340 VPWR VGND sg13g2_decap_8
XFILLER_49_384 VPWR VGND sg13g2_decap_8
XFILLER_37_513 VPWR VGND sg13g2_decap_8
XFILLER_18_771 VPWR VGND sg13g2_decap_8
XFILLER_37_568 VPWR VGND sg13g2_decap_8
XFILLER_21_903 VPWR VGND sg13g2_decap_8
XFILLER_33_752 VPWR VGND sg13g2_decap_8
XFILLER_20_446 VPWR VGND sg13g2_decap_8
XFILLER_32_295 VPWR VGND sg13g2_decap_4
X_2706_ _0601_ _0592_ _0603_ VPWR VGND sg13g2_xor2_1
X_2637_ _0488_ VPWR _0536_ VGND _0449_ _0489_ sg13g2_o21ai_1
X_2568_ net479 net477 net438 _0468_ VPWR VGND net434 sg13g2_nand4_1
XFILLER_0_818 VPWR VGND sg13g2_decap_8
X_1519_ _0846_ _0848_ _0854_ VPWR VGND sg13g2_nor2_1
X_2499_ _0398_ _0399_ _0393_ _0401_ VPWR VGND sg13g2_nand3_1
XFILLER_28_579 VPWR VGND sg13g2_decap_4
XFILLER_11_402 VPWR VGND sg13g2_decap_8
XFILLER_11_413 VPWR VGND sg13g2_fill_1
XFILLER_12_947 VPWR VGND sg13g2_decap_8
XFILLER_8_907 VPWR VGND sg13g2_decap_8
XFILLER_23_284 VPWR VGND sg13g2_decap_8
XFILLER_3_612 VPWR VGND sg13g2_decap_8
XFILLER_2_122 VPWR VGND sg13g2_decap_4
XFILLER_3_689 VPWR VGND sg13g2_decap_8
XFILLER_24_1020 VPWR VGND sg13g2_decap_8
XFILLER_47_822 VPWR VGND sg13g2_decap_8
Xfanout481 net483 net481 VPWR VGND sg13g2_buf_8
Xfanout470 net205 net470 VPWR VGND sg13g2_buf_8
Xfanout492 net194 net492 VPWR VGND sg13g2_buf_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_19_546 VPWR VGND sg13g2_decap_8
XFILLER_47_899 VPWR VGND sg13g2_decap_8
XFILLER_46_398 VPWR VGND sg13g2_decap_8
XFILLER_42_582 VPWR VGND sg13g2_decap_8
XFILLER_9_45 VPWR VGND sg13g2_fill_1
X_1870_ VGND VPWR _1171_ _1175_ _1195_ _1170_ sg13g2_a21oi_1
XFILLER_31_1013 VPWR VGND sg13g2_decap_8
XFILLER_7_973 VPWR VGND sg13g2_decap_8
X_2422_ _0330_ _0305_ _0329_ VPWR VGND sg13g2_xnor2_1
X_2353_ _0049_ _0262_ _0263_ VPWR VGND sg13g2_xnor2_1
X_2284_ _0197_ _0160_ _0195_ VPWR VGND sg13g2_nand2_1
XFILLER_21_744 VPWR VGND sg13g2_fill_2
XFILLER_21_777 VPWR VGND sg13g2_decap_8
X_1999_ mac1.sum_lvl3_ff\[6\] net261 _1298_ VPWR VGND sg13g2_and2_1
XFILLER_0_615 VPWR VGND sg13g2_decap_8
XFILLER_29_811 VPWR VGND sg13g2_fill_2
XFILLER_18_32 VPWR VGND sg13g2_decap_8
XFILLER_18_65 VPWR VGND sg13g2_fill_2
XFILLER_29_899 VPWR VGND sg13g2_decap_8
XFILLER_16_538 VPWR VGND sg13g2_decap_8
XFILLER_43_368 VPWR VGND sg13g2_fill_2
XFILLER_34_20 VPWR VGND sg13g2_decap_4
XFILLER_24_582 VPWR VGND sg13g2_decap_8
XFILLER_8_704 VPWR VGND sg13g2_decap_8
XFILLER_15_1019 VPWR VGND sg13g2_decap_8
XFILLER_24_593 VPWR VGND sg13g2_fill_1
XFILLER_12_777 VPWR VGND sg13g2_decap_8
XFILLER_7_247 VPWR VGND sg13g2_fill_2
XFILLER_7_236 VPWR VGND sg13g2_decap_8
XFILLER_4_910 VPWR VGND sg13g2_decap_8
XFILLER_4_987 VPWR VGND sg13g2_decap_8
XFILLER_19_310 VPWR VGND sg13g2_decap_8
XFILLER_34_357 VPWR VGND sg13g2_fill_1
XFILLER_43_880 VPWR VGND sg13g2_decap_8
X_2971_ net499 _0082_ VPWR VGND sg13g2_buf_1
XFILLER_42_390 VPWR VGND sg13g2_decap_8
X_1922_ VGND VPWR _1235_ _1237_ _1238_ _1236_ sg13g2_a21oi_1
X_1853_ _1178_ net465 net494 VPWR VGND sg13g2_nand2_1
XFILLER_7_770 VPWR VGND sg13g2_decap_8
X_1784_ VGND VPWR _1032_ _1075_ _1112_ _1074_ sg13g2_a21oi_1
X_2405_ VGND VPWR _0290_ _0293_ _0314_ _0289_ sg13g2_a21oi_1
XFILLER_29_118 VPWR VGND sg13g2_decap_8
X_2336_ _0247_ net446 net382 VPWR VGND sg13g2_nand2_2
X_2267_ _0180_ _0175_ _0179_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_630 VPWR VGND sg13g2_fill_1
X_2198_ _1478_ _1477_ _0055_ VPWR VGND sg13g2_xor2_1
XFILLER_38_1008 VPWR VGND sg13g2_decap_8
XFILLER_34_891 VPWR VGND sg13g2_decap_8
XFILLER_21_596 VPWR VGND sg13g2_fill_1
XFILLER_4_239 VPWR VGND sg13g2_decap_8
XFILLER_20_11 VPWR VGND sg13g2_decap_8
XFILLER_0_412 VPWR VGND sg13g2_decap_8
XFILLER_1_968 VPWR VGND sg13g2_decap_8
Xhold20 mac1.sum_lvl1_ff\[4\] VPWR VGND net60 sg13g2_dlygate4sd3_1
XFILLER_0_489 VPWR VGND sg13g2_decap_8
Xhold31 mac1.sum_lvl1_ff\[83\] VPWR VGND net71 sg13g2_dlygate4sd3_1
Xhold64 mac1.sum_lvl1_ff\[39\] VPWR VGND net104 sg13g2_dlygate4sd3_1
Xhold53 mac1.sum_lvl1_ff\[44\] VPWR VGND net93 sg13g2_dlygate4sd3_1
Xhold42 mac1.products_ff\[78\] VPWR VGND net82 sg13g2_dlygate4sd3_1
XFILLER_21_1001 VPWR VGND sg13g2_decap_8
XFILLER_29_64 VPWR VGND sg13g2_fill_2
XFILLER_29_86 VPWR VGND sg13g2_fill_2
Xhold86 mac1.sum_lvl1_ff\[75\] VPWR VGND net126 sg13g2_dlygate4sd3_1
Xhold75 mac1.sum_lvl2_ff\[40\] VPWR VGND net115 sg13g2_dlygate4sd3_1
Xhold97 mac1.products_ff\[68\] VPWR VGND net137 sg13g2_dlygate4sd3_1
XFILLER_44_611 VPWR VGND sg13g2_decap_8
XFILLER_28_173 VPWR VGND sg13g2_decap_4
XFILLER_45_74 VPWR VGND sg13g2_decap_8
XFILLER_43_176 VPWR VGND sg13g2_fill_1
XFILLER_40_883 VPWR VGND sg13g2_decap_8
XFILLER_8_534 VPWR VGND sg13g2_fill_1
XFILLER_12_585 VPWR VGND sg13g2_decap_4
XFILLER_4_784 VPWR VGND sg13g2_decap_8
XFILLER_6_1028 VPWR VGND sg13g2_fill_1
X_3170_ net542 VGND VPWR net77 mac1.sum_lvl2_ff\[28\] clknet_leaf_24_clk sg13g2_dfrbpq_1
X_2121_ _1403_ _1404_ _1405_ VPWR VGND sg13g2_and2_1
XFILLER_13_4 VPWR VGND sg13g2_decap_8
XFILLER_48_961 VPWR VGND sg13g2_decap_8
X_2052_ _1340_ net392 net457 net454 net397 VPWR VGND sg13g2_a22oi_1
XFILLER_47_493 VPWR VGND sg13g2_fill_1
XFILLER_22_305 VPWR VGND sg13g2_fill_1
XFILLER_15_390 VPWR VGND sg13g2_decap_8
X_2954_ _0832_ VPWR _0111_ VGND net374 _0831_ sg13g2_o21ai_1
X_2885_ _0775_ _0765_ net372 VPWR VGND sg13g2_nand2_1
X_1905_ _1225_ net235 net161 VPWR VGND sg13g2_nand2_1
XFILLER_31_894 VPWR VGND sg13g2_decap_8
X_1836_ VGND VPWR _1162_ _1161_ _1149_ sg13g2_or2_1
X_1767_ net408 net407 net463 net460 _1095_ VPWR VGND sg13g2_and4_1
X_1698_ VGND VPWR _1024_ _1025_ _1028_ _0990_ sg13g2_a21oi_1
X_2319_ _0231_ _0230_ _0229_ VPWR VGND sg13g2_nand2b_1
Xheichips25_template_33 VPWR VGND uio_oe[0] sg13g2_tiehi
XFILLER_26_600 VPWR VGND sg13g2_decap_8
XFILLER_26_655 VPWR VGND sg13g2_decap_8
XFILLER_14_817 VPWR VGND sg13g2_decap_4
XFILLER_15_11 VPWR VGND sg13g2_decap_4
XFILLER_26_688 VPWR VGND sg13g2_decap_8
XFILLER_40_102 VPWR VGND sg13g2_decap_8
XFILLER_13_349 VPWR VGND sg13g2_decap_8
XFILLER_15_77 VPWR VGND sg13g2_decap_8
XFILLER_21_393 VPWR VGND sg13g2_decap_8
Xoutput32 net32 uo_out[7] VPWR VGND sg13g2_buf_1
Xoutput21 net21 uio_out[4] VPWR VGND sg13g2_buf_1
XFILLER_1_765 VPWR VGND sg13g2_decap_8
XFILLER_48_202 VPWR VGND sg13g2_decap_8
XFILLER_49_769 VPWR VGND sg13g2_decap_8
XFILLER_36_408 VPWR VGND sg13g2_decap_8
XFILLER_48_279 VPWR VGND sg13g2_decap_8
XFILLER_45_942 VPWR VGND sg13g2_decap_8
XFILLER_16_154 VPWR VGND sg13g2_fill_1
XFILLER_31_113 VPWR VGND sg13g2_decap_8
XFILLER_40_680 VPWR VGND sg13g2_fill_2
XFILLER_13_883 VPWR VGND sg13g2_decap_8
X_2670_ _0568_ _0553_ _0567_ VPWR VGND sg13g2_nand2_1
XFILLER_9_865 VPWR VGND sg13g2_decap_8
XFILLER_8_386 VPWR VGND sg13g2_decap_8
X_1621_ net473 net403 net474 _0952_ VPWR VGND net402 sg13g2_nand4_1
X_1552_ _0865_ _0885_ _0886_ VPWR VGND sg13g2_nor2_1
XFILLER_28_1007 VPWR VGND sg13g2_decap_8
X_3222_ net523 VGND VPWR net142 mac1.sum_lvl3_ff\[33\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_3153_ net542 VGND VPWR net86 mac1.sum_lvl2_ff\[8\] clknet_leaf_24_clk sg13g2_dfrbpq_1
XFILLER_39_224 VPWR VGND sg13g2_fill_1
X_2104_ _1386_ _1383_ _1388_ VPWR VGND sg13g2_xor2_1
XFILLER_28_909 VPWR VGND sg13g2_decap_8
X_3084_ net525 VGND VPWR _0045_ mac1.products_ff\[71\] clknet_leaf_27_clk sg13g2_dfrbpq_1
XFILLER_47_290 VPWR VGND sg13g2_decap_8
X_2035_ net292 VPWR _1328_ VGND _1325_ _1327_ sg13g2_o21ai_1
XFILLER_36_942 VPWR VGND sg13g2_decap_8
XFILLER_22_102 VPWR VGND sg13g2_decap_8
XFILLER_22_113 VPWR VGND sg13g2_fill_1
XFILLER_22_135 VPWR VGND sg13g2_fill_2
X_2937_ _0750_ _0740_ _0822_ VPWR VGND sg13g2_xor2_1
X_2868_ _0758_ net443 _0732_ VPWR VGND sg13g2_nand2_1
X_2799_ _0692_ _0678_ _0693_ VPWR VGND sg13g2_xor2_1
X_1819_ _1132_ _1127_ _1134_ _1145_ VPWR VGND sg13g2_a21o_1
XFILLER_46_706 VPWR VGND sg13g2_decap_8
XFILLER_26_21 VPWR VGND sg13g2_decap_8
XFILLER_26_430 VPWR VGND sg13g2_fill_1
XFILLER_27_953 VPWR VGND sg13g2_decap_8
XFILLER_42_923 VPWR VGND sg13g2_decap_8
XFILLER_26_463 VPWR VGND sg13g2_decap_8
XFILLER_26_474 VPWR VGND sg13g2_fill_1
XFILLER_22_680 VPWR VGND sg13g2_decap_8
XFILLER_10_831 VPWR VGND sg13g2_decap_8
XFILLER_6_846 VPWR VGND sg13g2_decap_8
XFILLER_3_36 VPWR VGND sg13g2_fill_1
XFILLER_3_25 VPWR VGND sg13g2_decap_8
XFILLER_1_562 VPWR VGND sg13g2_decap_8
XFILLER_49_566 VPWR VGND sg13g2_decap_8
XFILLER_49_599 VPWR VGND sg13g2_decap_4
XFILLER_37_717 VPWR VGND sg13g2_decap_8
XFILLER_17_430 VPWR VGND sg13g2_fill_2
XFILLER_17_463 VPWR VGND sg13g2_decap_8
XFILLER_18_986 VPWR VGND sg13g2_decap_8
XFILLER_17_485 VPWR VGND sg13g2_fill_2
XFILLER_33_945 VPWR VGND sg13g2_decap_8
XFILLER_13_680 VPWR VGND sg13g2_decap_4
X_2722_ _0602_ VPWR _0618_ VGND _0591_ _0603_ sg13g2_o21ai_1
XFILLER_9_673 VPWR VGND sg13g2_decap_8
X_2653_ _0542_ _0550_ _0551_ VPWR VGND sg13g2_nor2_1
X_1604_ _0933_ _0934_ _0928_ _0936_ VPWR VGND sg13g2_nand3_1
X_2584_ VGND VPWR _0480_ _0481_ _0484_ _0450_ sg13g2_a21oi_1
X_1535_ _0866_ _0868_ _0869_ VPWR VGND sg13g2_nor2b_1
XFILLER_41_1004 VPWR VGND sg13g2_decap_8
X_3205_ net522 VGND VPWR net107 mac1.sum_lvl1_ff\[84\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_28_706 VPWR VGND sg13g2_decap_4
X_3136_ net536 VGND VPWR net43 mac1.sum_lvl1_ff\[43\] clknet_leaf_24_clk sg13g2_dfrbpq_1
XFILLER_28_717 VPWR VGND sg13g2_decap_8
X_3067_ net527 VGND VPWR _0120_ DP_2.matrix\[38\] clknet_leaf_22_clk sg13g2_dfrbpq_1
X_2018_ net182 VPWR _1314_ VGND _1307_ _1309_ sg13g2_o21ai_1
XFILLER_24_901 VPWR VGND sg13g2_decap_8
XFILLER_36_750 VPWR VGND sg13g2_decap_4
XFILLER_24_978 VPWR VGND sg13g2_decap_8
XFILLER_35_293 VPWR VGND sg13g2_decap_4
XFILLER_10_105 VPWR VGND sg13g2_fill_2
XFILLER_11_639 VPWR VGND sg13g2_decap_8
XFILLER_23_499 VPWR VGND sg13g2_decap_8
XFILLER_6_109 VPWR VGND sg13g2_decap_8
XFILLER_12_78 VPWR VGND sg13g2_decap_8
Xhold150 DP_2.matrix\[74\] VPWR VGND net190 sg13g2_dlygate4sd3_1
Xhold161 _1291_ VPWR VGND net201 sg13g2_dlygate4sd3_1
Xhold183 DP_2.matrix\[2\] VPWR VGND net223 sg13g2_dlygate4sd3_1
Xhold194 _0020_ VPWR VGND net234 sg13g2_dlygate4sd3_1
Xhold172 DP_1.matrix\[39\] VPWR VGND net212 sg13g2_dlygate4sd3_1
XFILLER_46_536 VPWR VGND sg13g2_decap_8
XFILLER_27_761 VPWR VGND sg13g2_fill_2
XFILLER_27_772 VPWR VGND sg13g2_decap_8
XFILLER_26_260 VPWR VGND sg13g2_fill_1
XFILLER_42_742 VPWR VGND sg13g2_fill_1
XFILLER_41_230 VPWR VGND sg13g2_decap_8
XFILLER_15_956 VPWR VGND sg13g2_decap_8
XFILLER_18_1028 VPWR VGND sg13g2_fill_1
XFILLER_41_274 VPWR VGND sg13g2_decap_8
XFILLER_14_488 VPWR VGND sg13g2_decap_8
XFILLER_30_948 VPWR VGND sg13g2_decap_8
XFILLER_10_661 VPWR VGND sg13g2_decap_4
XFILLER_6_610 VPWR VGND sg13g2_decap_8
XFILLER_10_683 VPWR VGND sg13g2_fill_1
XFILLER_6_643 VPWR VGND sg13g2_decap_8
XFILLER_5_197 VPWR VGND sg13g2_decap_8
XFILLER_2_860 VPWR VGND sg13g2_decap_8
XFILLER_32_241 VPWR VGND sg13g2_decap_8
XFILLER_33_742 VPWR VGND sg13g2_fill_2
XFILLER_21_959 VPWR VGND sg13g2_decap_8
X_2705_ _0602_ _0592_ _0601_ VPWR VGND sg13g2_nand2b_1
XFILLER_9_481 VPWR VGND sg13g2_decap_8
X_2636_ _0533_ _0534_ _0535_ VPWR VGND sg13g2_and2_1
X_2567_ net438 net480 net477 net434 _0467_ VPWR VGND sg13g2_and4_1
X_1518_ _0853_ net474 net408 VPWR VGND sg13g2_nand2_1
X_2498_ _0400_ _0393_ _0398_ _0399_ VPWR VGND sg13g2_and3_1
XFILLER_28_558 VPWR VGND sg13g2_decap_8
X_3119_ net536 VGND VPWR net87 mac1.sum_lvl1_ff\[6\] clknet_leaf_29_clk sg13g2_dfrbpq_1
XFILLER_43_539 VPWR VGND sg13g2_decap_8
XFILLER_24_731 VPWR VGND sg13g2_decap_8
XFILLER_36_580 VPWR VGND sg13g2_decap_8
XFILLER_24_742 VPWR VGND sg13g2_fill_2
XFILLER_12_926 VPWR VGND sg13g2_decap_8
XFILLER_23_11 VPWR VGND sg13g2_decap_8
XFILLER_11_436 VPWR VGND sg13g2_fill_1
XFILLER_7_429 VPWR VGND sg13g2_fill_1
XFILLER_20_981 VPWR VGND sg13g2_decap_8
XFILLER_3_668 VPWR VGND sg13g2_decap_8
XFILLER_2_156 VPWR VGND sg13g2_decap_8
XFILLER_48_63 VPWR VGND sg13g2_fill_1
Xfanout482 net483 net482 VPWR VGND sg13g2_buf_8
Xfanout471 DP_1.matrix\[38\] net471 VPWR VGND sg13g2_buf_8
Xfanout460 net461 net460 VPWR VGND sg13g2_buf_2
Xfanout493 DP_1.matrix\[0\] net493 VPWR VGND sg13g2_buf_1
XFILLER_46_311 VPWR VGND sg13g2_decap_8
XFILLER_19_525 VPWR VGND sg13g2_decap_8
XFILLER_47_878 VPWR VGND sg13g2_decap_8
XFILLER_34_517 VPWR VGND sg13g2_decap_8
XFILLER_30_778 VPWR VGND sg13g2_decap_8
XFILLER_7_952 VPWR VGND sg13g2_decap_8
XFILLER_6_473 VPWR VGND sg13g2_decap_8
X_2421_ _0327_ _0321_ _0329_ VPWR VGND sg13g2_xor2_1
XFILLER_9_1026 VPWR VGND sg13g2_fill_2
X_2352_ _0229_ _0234_ _0263_ VPWR VGND sg13g2_nor2_1
X_2283_ _0160_ _0195_ _0196_ VPWR VGND sg13g2_nor2_1
XFILLER_37_300 VPWR VGND sg13g2_decap_8
XFILLER_49_193 VPWR VGND sg13g2_decap_8
XFILLER_37_366 VPWR VGND sg13g2_decap_4
XFILLER_38_889 VPWR VGND sg13g2_decap_8
XFILLER_21_712 VPWR VGND sg13g2_fill_1
XFILLER_33_594 VPWR VGND sg13g2_decap_8
X_1998_ _0027_ _1295_ net179 VPWR VGND sg13g2_xnor2_1
X_2619_ _0515_ _0516_ _0510_ _0518_ VPWR VGND sg13g2_nand3_1
XFILLER_29_878 VPWR VGND sg13g2_decap_8
XFILLER_43_314 VPWR VGND sg13g2_fill_1
XFILLER_16_517 VPWR VGND sg13g2_fill_2
XFILLER_44_859 VPWR VGND sg13g2_decap_8
XFILLER_24_561 VPWR VGND sg13g2_decap_8
XFILLER_31_509 VPWR VGND sg13g2_fill_1
XFILLER_34_98 VPWR VGND sg13g2_fill_1
XFILLER_4_966 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_39_609 VPWR VGND sg13g2_decap_8
XFILLER_47_631 VPWR VGND sg13g2_decap_4
XFILLER_46_141 VPWR VGND sg13g2_fill_2
XFILLER_46_174 VPWR VGND sg13g2_fill_1
XFILLER_19_388 VPWR VGND sg13g2_fill_1
XFILLER_35_826 VPWR VGND sg13g2_decap_8
XFILLER_35_859 VPWR VGND sg13g2_decap_8
X_2970_ net156 _0080_ VPWR VGND sg13g2_buf_1
X_1921_ net266 _1235_ _0010_ VPWR VGND sg13g2_xor2_1
X_1852_ _1155_ VPWR _1177_ VGND _1152_ _1156_ sg13g2_o21ai_1
X_1783_ _1035_ _1077_ _1034_ _1111_ VPWR VGND sg13g2_nand3_1
X_2404_ _0311_ _0312_ _0313_ VPWR VGND sg13g2_and2_1
X_2335_ _0246_ DP_1.matrix\[75\] net502 VPWR VGND sg13g2_nand2_1
X_2266_ _0179_ _1494_ _0176_ VPWR VGND sg13g2_xnor2_1
X_2197_ _1479_ _1477_ _1478_ VPWR VGND sg13g2_nand2_1
XFILLER_26_804 VPWR VGND sg13g2_fill_1
XFILLER_25_336 VPWR VGND sg13g2_decap_8
XFILLER_26_859 VPWR VGND sg13g2_fill_2
XFILLER_41_829 VPWR VGND sg13g2_decap_8
XFILLER_34_870 VPWR VGND sg13g2_decap_8
XFILLER_20_89 VPWR VGND sg13g2_decap_4
XFILLER_1_947 VPWR VGND sg13g2_decap_8
Xhold10 mac1.sum_lvl2_ff\[38\] VPWR VGND net50 sg13g2_dlygate4sd3_1
XFILLER_0_468 VPWR VGND sg13g2_decap_8
Xhold21 mac1.products_ff\[5\] VPWR VGND net61 sg13g2_dlygate4sd3_1
Xhold32 mac1.sum_lvl1_ff\[11\] VPWR VGND net72 sg13g2_dlygate4sd3_1
Xhold65 mac1.sum_lvl1_ff\[38\] VPWR VGND net105 sg13g2_dlygate4sd3_1
Xhold54 mac1.sum_lvl1_ff\[36\] VPWR VGND net94 sg13g2_dlygate4sd3_1
Xhold43 mac1.sum_lvl1_ff\[85\] VPWR VGND net83 sg13g2_dlygate4sd3_1
Xhold87 mac1.products_ff\[15\] VPWR VGND net127 sg13g2_dlygate4sd3_1
Xhold98 mac1.sum_lvl2_ff\[44\] VPWR VGND net138 sg13g2_dlygate4sd3_1
Xhold76 mac1.sum_lvl1_ff\[3\] VPWR VGND net116 sg13g2_dlygate4sd3_1
XFILLER_29_653 VPWR VGND sg13g2_decap_4
XFILLER_45_20 VPWR VGND sg13g2_decap_4
XFILLER_16_303 VPWR VGND sg13g2_decap_8
XFILLER_29_697 VPWR VGND sg13g2_decap_8
XFILLER_44_667 VPWR VGND sg13g2_decap_8
XFILLER_28_196 VPWR VGND sg13g2_decap_4
XFILLER_43_155 VPWR VGND sg13g2_decap_8
XFILLER_16_369 VPWR VGND sg13g2_decap_8
XFILLER_25_892 VPWR VGND sg13g2_decap_8
XFILLER_40_862 VPWR VGND sg13g2_decap_8
XFILLER_12_531 VPWR VGND sg13g2_decap_4
XFILLER_6_36 VPWR VGND sg13g2_decap_8
XFILLER_4_763 VPWR VGND sg13g2_decap_8
XFILLER_39_417 VPWR VGND sg13g2_decap_8
XFILLER_6_1007 VPWR VGND sg13g2_decap_8
XFILLER_48_940 VPWR VGND sg13g2_decap_8
X_2120_ _1402_ _1401_ _1363_ _1404_ VPWR VGND sg13g2_a21o_1
X_2051_ _1339_ net454 net392 _0032_ VPWR VGND sg13g2_and3_2
XFILLER_47_472 VPWR VGND sg13g2_decap_4
XFILLER_23_818 VPWR VGND sg13g2_decap_8
XFILLER_34_166 VPWR VGND sg13g2_decap_4
XFILLER_34_188 VPWR VGND sg13g2_decap_4
X_2953_ _0832_ net433 net374 VPWR VGND sg13g2_nand2_1
X_1904_ net492 net437 _0037_ VPWR VGND sg13g2_and2_1
XFILLER_31_840 VPWR VGND sg13g2_fill_1
XFILLER_31_873 VPWR VGND sg13g2_decap_8
X_2884_ _0773_ net372 _0774_ VPWR VGND sg13g2_nor2b_1
XFILLER_30_372 VPWR VGND sg13g2_decap_8
X_1835_ _1159_ _1150_ _1161_ VPWR VGND sg13g2_xor2_1
X_1766_ _1094_ net406 net460 VPWR VGND sg13g2_nand2_1
X_1697_ _1024_ _1025_ _0990_ _1027_ VPWR VGND sg13g2_nand3_1
XFILLER_44_1013 VPWR VGND sg13g2_decap_8
X_2318_ _0194_ _0228_ _0192_ _0230_ VPWR VGND sg13g2_nand3_1
XFILLER_45_409 VPWR VGND sg13g2_decap_8
Xheichips25_template_34 VPWR VGND uio_oe[1] sg13g2_tiehi
XFILLER_39_995 VPWR VGND sg13g2_decap_8
X_2249_ _0145_ VPWR _0162_ VGND _1491_ _0146_ sg13g2_o21ai_1
XFILLER_26_612 VPWR VGND sg13g2_decap_8
XFILLER_26_623 VPWR VGND sg13g2_decap_4
XFILLER_15_23 VPWR VGND sg13g2_decap_4
XFILLER_41_626 VPWR VGND sg13g2_fill_2
XFILLER_40_147 VPWR VGND sg13g2_decap_8
XFILLER_21_372 VPWR VGND sg13g2_decap_8
XFILLER_31_44 VPWR VGND sg13g2_fill_1
XFILLER_5_538 VPWR VGND sg13g2_decap_8
XFILLER_31_99 VPWR VGND sg13g2_decap_8
Xoutput22 net22 uio_out[5] VPWR VGND sg13g2_buf_1
XFILLER_1_744 VPWR VGND sg13g2_decap_8
XFILLER_49_748 VPWR VGND sg13g2_decap_8
XFILLER_48_258 VPWR VGND sg13g2_decap_8
XFILLER_0_298 VPWR VGND sg13g2_decap_8
XFILLER_45_921 VPWR VGND sg13g2_decap_8
XFILLER_29_494 VPWR VGND sg13g2_decap_8
XFILLER_45_998 VPWR VGND sg13g2_decap_8
XFILLER_32_626 VPWR VGND sg13g2_decap_4
XFILLER_32_637 VPWR VGND sg13g2_fill_1
XFILLER_13_862 VPWR VGND sg13g2_decap_8
XFILLER_9_844 VPWR VGND sg13g2_decap_8
XFILLER_31_169 VPWR VGND sg13g2_fill_2
XFILLER_8_365 VPWR VGND sg13g2_decap_8
X_1620_ _0951_ net402 net475 net403 net473 VPWR VGND sg13g2_a22oi_1
X_1551_ VGND VPWR _0885_ _0884_ _0882_ sg13g2_or2_1
X_3221_ net523 VGND VPWR net90 mac1.sum_lvl3_ff\[32\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_3152_ net536 VGND VPWR net100 mac1.sum_lvl2_ff\[7\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_2103_ _1387_ _1386_ _1383_ VPWR VGND sg13g2_nand2b_1
XFILLER_39_258 VPWR VGND sg13g2_fill_1
X_3083_ net520 VGND VPWR _0044_ mac1.products_ff\[70\] clknet_leaf_33_clk sg13g2_dfrbpq_1
XFILLER_27_409 VPWR VGND sg13g2_decap_8
XFILLER_36_921 VPWR VGND sg13g2_decap_8
X_2034_ VGND VPWR _1312_ _1314_ _1327_ _1326_ sg13g2_a21oi_1
XFILLER_23_604 VPWR VGND sg13g2_fill_2
XFILLER_35_453 VPWR VGND sg13g2_decap_8
XFILLER_36_998 VPWR VGND sg13g2_decap_8
XFILLER_23_626 VPWR VGND sg13g2_fill_1
XFILLER_22_147 VPWR VGND sg13g2_decap_8
X_2936_ net486 net372 _0821_ VPWR VGND sg13g2_nor2_1
X_2867_ _0757_ _0738_ _0756_ VPWR VGND sg13g2_nand2b_1
X_1818_ _1144_ _1143_ _0071_ VPWR VGND sg13g2_xor2_1
X_2798_ _0690_ _0664_ _0692_ VPWR VGND sg13g2_xor2_1
X_1749_ _0079_ _1037_ _1076_ VPWR VGND sg13g2_xnor2_1
XFILLER_45_217 VPWR VGND sg13g2_fill_1
XFILLER_45_239 VPWR VGND sg13g2_decap_8
XFILLER_26_11 VPWR VGND sg13g2_decap_4
XFILLER_27_932 VPWR VGND sg13g2_decap_8
XFILLER_38_280 VPWR VGND sg13g2_fill_2
XFILLER_42_902 VPWR VGND sg13g2_decap_8
XFILLER_13_103 VPWR VGND sg13g2_fill_1
XFILLER_14_615 VPWR VGND sg13g2_decap_8
XFILLER_26_77 VPWR VGND sg13g2_fill_2
XFILLER_26_88 VPWR VGND sg13g2_fill_2
XFILLER_26_497 VPWR VGND sg13g2_decap_8
XFILLER_42_979 VPWR VGND sg13g2_decap_8
XFILLER_42_43 VPWR VGND sg13g2_decap_8
XFILLER_10_810 VPWR VGND sg13g2_decap_8
XFILLER_42_87 VPWR VGND sg13g2_decap_8
XFILLER_10_887 VPWR VGND sg13g2_decap_8
XFILLER_6_825 VPWR VGND sg13g2_decap_8
XFILLER_5_324 VPWR VGND sg13g2_fill_1
XFILLER_5_379 VPWR VGND sg13g2_decap_8
XFILLER_49_534 VPWR VGND sg13g2_decap_8
XFILLER_18_965 VPWR VGND sg13g2_decap_8
XFILLER_45_795 VPWR VGND sg13g2_decap_8
XFILLER_33_924 VPWR VGND sg13g2_decap_8
XFILLER_32_478 VPWR VGND sg13g2_decap_4
X_2721_ _0588_ _0582_ _0590_ _0617_ VPWR VGND sg13g2_a21o_1
XFILLER_41_990 VPWR VGND sg13g2_decap_8
XFILLER_9_663 VPWR VGND sg13g2_fill_1
X_2652_ _0550_ _0543_ _0549_ VPWR VGND sg13g2_xnor2_1
X_1603_ _0935_ _0928_ _0933_ _0934_ VPWR VGND sg13g2_and3_1
X_2583_ _0480_ _0481_ _0450_ _0483_ VPWR VGND sg13g2_nand3_1
X_1534_ VGND VPWR _0868_ _0867_ _0853_ sg13g2_or2_1
X_3204_ net522 VGND VPWR net146 mac1.sum_lvl1_ff\[83\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_3135_ net534 VGND VPWR net62 mac1.sum_lvl1_ff\[42\] clknet_leaf_26_clk sg13g2_dfrbpq_1
X_3066_ net528 VGND VPWR _0119_ DP_2.matrix\[37\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_2017_ net181 mac1.sum_lvl3_ff\[9\] _1313_ VPWR VGND sg13g2_xor2_1
XFILLER_35_272 VPWR VGND sg13g2_decap_8
XFILLER_24_957 VPWR VGND sg13g2_decap_8
XFILLER_11_618 VPWR VGND sg13g2_decap_8
XFILLER_23_478 VPWR VGND sg13g2_decap_8
X_2919_ _0805_ _0807_ _0808_ VPWR VGND sg13g2_nor2_1
XFILLER_32_990 VPWR VGND sg13g2_decap_8
XFILLER_12_35 VPWR VGND sg13g2_decap_4
Xhold151 DP_2.matrix\[42\] VPWR VGND net191 sg13g2_dlygate4sd3_1
Xhold140 _0027_ VPWR VGND net180 sg13g2_dlygate4sd3_1
Xhold162 _0025_ VPWR VGND net202 sg13g2_dlygate4sd3_1
XFILLER_2_338 VPWR VGND sg13g2_decap_4
Xhold184 _0112_ VPWR VGND net224 sg13g2_dlygate4sd3_1
Xhold195 mac1.sum_lvl2_ff\[19\] VPWR VGND net235 sg13g2_dlygate4sd3_1
Xhold173 mac1.sum_lvl3_ff\[30\] VPWR VGND net213 sg13g2_dlygate4sd3_1
XFILLER_19_707 VPWR VGND sg13g2_decap_8
XFILLER_19_729 VPWR VGND sg13g2_decap_8
XFILLER_2_1021 VPWR VGND sg13g2_decap_8
XFILLER_37_98 VPWR VGND sg13g2_decap_8
XFILLER_15_935 VPWR VGND sg13g2_decap_8
XFILLER_14_434 VPWR VGND sg13g2_fill_1
XFILLER_18_1007 VPWR VGND sg13g2_decap_8
XFILLER_30_927 VPWR VGND sg13g2_decap_8
XFILLER_6_699 VPWR VGND sg13g2_decap_8
XFILLER_45_8 VPWR VGND sg13g2_fill_2
XFILLER_49_375 VPWR VGND sg13g2_decap_4
XFILLER_18_740 VPWR VGND sg13g2_decap_8
XFILLER_21_938 VPWR VGND sg13g2_decap_8
XFILLER_33_787 VPWR VGND sg13g2_decap_8
X_2704_ _0601_ _0593_ _0600_ VPWR VGND sg13g2_xnor2_1
X_2635_ _0531_ _0530_ _0532_ _0534_ VPWR VGND sg13g2_a21o_1
X_2566_ _0466_ net482 net431 VPWR VGND sg13g2_nand2_1
X_1517_ _0044_ _0850_ _0851_ VPWR VGND sg13g2_xnor2_1
X_2497_ _0394_ VPWR _0399_ VGND _0395_ _0397_ sg13g2_o21ai_1
XFILLER_4_80 VPWR VGND sg13g2_decap_8
X_3118_ net535 VGND VPWR net61 mac1.sum_lvl1_ff\[5\] clknet_leaf_28_clk sg13g2_dfrbpq_1
XFILLER_43_518 VPWR VGND sg13g2_decap_8
XFILLER_15_209 VPWR VGND sg13g2_fill_2
X_3049_ net515 VGND VPWR _0102_ DP_1.matrix\[72\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_12_905 VPWR VGND sg13g2_decap_8
XFILLER_23_253 VPWR VGND sg13g2_decap_8
XFILLER_20_960 VPWR VGND sg13g2_decap_8
XFILLER_23_89 VPWR VGND sg13g2_decap_8
XFILLER_3_647 VPWR VGND sg13g2_decap_8
XFILLER_3_4 VPWR VGND sg13g2_decap_8
XFILLER_48_42 VPWR VGND sg13g2_decap_8
Xfanout450 net451 net450 VPWR VGND sg13g2_buf_8
Xfanout483 net225 net483 VPWR VGND sg13g2_buf_8
Xfanout472 net473 net472 VPWR VGND sg13g2_buf_8
Xfanout461 net274 net461 VPWR VGND sg13g2_buf_8
XFILLER_47_857 VPWR VGND sg13g2_decap_8
Xfanout494 DP_2.matrix\[44\] net494 VPWR VGND sg13g2_buf_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_15_743 VPWR VGND sg13g2_fill_2
XFILLER_42_551 VPWR VGND sg13g2_fill_2
XFILLER_14_242 VPWR VGND sg13g2_decap_4
XFILLER_14_264 VPWR VGND sg13g2_decap_8
XFILLER_9_69 VPWR VGND sg13g2_decap_8
XFILLER_9_58 VPWR VGND sg13g2_fill_2
XFILLER_30_724 VPWR VGND sg13g2_decap_8
XFILLER_7_931 VPWR VGND sg13g2_decap_8
XFILLER_11_982 VPWR VGND sg13g2_decap_8
XFILLER_6_430 VPWR VGND sg13g2_decap_8
XFILLER_6_496 VPWR VGND sg13g2_decap_4
X_2420_ _0328_ _0321_ _0327_ VPWR VGND sg13g2_nand2_1
XFILLER_9_1005 VPWR VGND sg13g2_decap_8
X_2351_ _0260_ _0261_ _0262_ VPWR VGND sg13g2_nor2_1
X_2282_ _0195_ _0161_ _0193_ VPWR VGND sg13g2_xnor2_1
XFILLER_49_172 VPWR VGND sg13g2_decap_8
XFILLER_38_868 VPWR VGND sg13g2_decap_8
XFILLER_37_378 VPWR VGND sg13g2_decap_4
XFILLER_46_890 VPWR VGND sg13g2_decap_8
XFILLER_18_592 VPWR VGND sg13g2_decap_8
XFILLER_33_573 VPWR VGND sg13g2_decap_8
XFILLER_20_223 VPWR VGND sg13g2_fill_2
XFILLER_21_724 VPWR VGND sg13g2_fill_2
X_1997_ mac1.sum_lvl3_ff\[25\] net178 _1297_ VPWR VGND sg13g2_xor2_1
XFILLER_21_768 VPWR VGND sg13g2_fill_1
XFILLER_9_290 VPWR VGND sg13g2_fill_2
XFILLER_47_1011 VPWR VGND sg13g2_decap_8
X_2618_ _0517_ _0510_ _0515_ _0516_ VPWR VGND sg13g2_and3_1
X_2549_ VGND VPWR _0412_ _0447_ _0449_ _0446_ sg13g2_a21oi_1
XFILLER_18_67 VPWR VGND sg13g2_fill_1
XFILLER_44_838 VPWR VGND sg13g2_decap_8
XFILLER_12_735 VPWR VGND sg13g2_decap_8
XFILLER_8_739 VPWR VGND sg13g2_decap_8
XFILLER_11_289 VPWR VGND sg13g2_fill_2
XFILLER_4_945 VPWR VGND sg13g2_decap_8
XFILLER_47_621 VPWR VGND sg13g2_decap_4
XFILLER_19_345 VPWR VGND sg13g2_fill_2
XFILLER_35_805 VPWR VGND sg13g2_decap_8
XFILLER_47_687 VPWR VGND sg13g2_decap_8
XFILLER_19_367 VPWR VGND sg13g2_decap_8
XFILLER_34_304 VPWR VGND sg13g2_decap_8
X_1920_ net265 mac1.sum_lvl2_ff\[23\] _1237_ VPWR VGND sg13g2_xor2_1
XFILLER_15_573 VPWR VGND sg13g2_decap_8
XFILLER_30_521 VPWR VGND sg13g2_decap_8
X_1851_ _1158_ _1151_ _1160_ _1176_ VPWR VGND sg13g2_a21o_1
X_1782_ _1110_ _1109_ _1108_ VPWR VGND sg13g2_nand2b_1
X_2403_ _0284_ _0286_ _0310_ _0312_ VPWR VGND sg13g2_or3_1
X_2334_ VGND VPWR _0245_ _0218_ _0216_ sg13g2_or2_1
XFILLER_27_0 VPWR VGND sg13g2_decap_8
X_2265_ _1494_ _0176_ _0178_ VPWR VGND sg13g2_and2_1
XFILLER_38_610 VPWR VGND sg13g2_fill_1
X_2196_ _1440_ _1439_ _1438_ _1478_ VPWR VGND sg13g2_a21o_2
XFILLER_38_643 VPWR VGND sg13g2_decap_4
XFILLER_1_92 VPWR VGND sg13g2_decap_4
XFILLER_25_315 VPWR VGND sg13g2_decap_8
XFILLER_38_698 VPWR VGND sg13g2_decap_8
XFILLER_33_370 VPWR VGND sg13g2_decap_4
XFILLER_14_1010 VPWR VGND sg13g2_decap_8
XFILLER_21_587 VPWR VGND sg13g2_decap_8
XFILLER_20_46 VPWR VGND sg13g2_decap_4
XFILLER_1_926 VPWR VGND sg13g2_decap_8
Xhold22 mac1.products_ff\[74\] VPWR VGND net62 sg13g2_dlygate4sd3_1
XFILLER_0_447 VPWR VGND sg13g2_decap_8
XFILLER_29_22 VPWR VGND sg13g2_fill_1
XFILLER_29_44 VPWR VGND sg13g2_decap_8
Xhold11 mac1.products_ff\[151\] VPWR VGND net51 sg13g2_dlygate4sd3_1
Xhold55 mac1.products_ff\[4\] VPWR VGND net95 sg13g2_dlygate4sd3_1
Xhold33 mac1.products_ff\[73\] VPWR VGND net73 sg13g2_dlygate4sd3_1
Xhold44 mac1.products_ff\[77\] VPWR VGND net84 sg13g2_dlygate4sd3_1
XFILLER_29_66 VPWR VGND sg13g2_fill_1
Xhold77 mac1.products_ff\[13\] VPWR VGND net117 sg13g2_dlygate4sd3_1
Xhold66 mac1.products_ff\[7\] VPWR VGND net106 sg13g2_dlygate4sd3_1
Xhold88 mac1.products_ff\[139\] VPWR VGND net128 sg13g2_dlygate4sd3_1
Xhold99 mac1.sum_lvl1_ff\[76\] VPWR VGND net139 sg13g2_dlygate4sd3_1
XFILLER_29_88 VPWR VGND sg13g2_fill_1
XFILLER_29_665 VPWR VGND sg13g2_fill_2
XFILLER_17_827 VPWR VGND sg13g2_decap_8
XFILLER_28_153 VPWR VGND sg13g2_fill_1
XFILLER_29_676 VPWR VGND sg13g2_decap_8
XFILLER_43_134 VPWR VGND sg13g2_decap_8
XFILLER_12_510 VPWR VGND sg13g2_decap_8
XFILLER_40_841 VPWR VGND sg13g2_decap_8
XFILLER_24_392 VPWR VGND sg13g2_decap_8
XFILLER_8_525 VPWR VGND sg13g2_decap_8
XFILLER_8_558 VPWR VGND sg13g2_decap_8
XFILLER_6_15 VPWR VGND sg13g2_decap_8
XFILLER_4_742 VPWR VGND sg13g2_decap_8
X_2050_ net153 mac1.sum_lvl3_ff\[0\] _0016_ VPWR VGND sg13g2_xor2_1
XFILLER_48_996 VPWR VGND sg13g2_decap_8
XFILLER_47_451 VPWR VGND sg13g2_fill_1
XFILLER_19_164 VPWR VGND sg13g2_decap_8
XFILLER_35_613 VPWR VGND sg13g2_decap_8
XFILLER_35_624 VPWR VGND sg13g2_fill_1
XFILLER_19_197 VPWR VGND sg13g2_decap_8
XFILLER_34_112 VPWR VGND sg13g2_fill_2
XFILLER_35_657 VPWR VGND sg13g2_decap_8
XFILLER_34_145 VPWR VGND sg13g2_decap_8
X_2952_ _0796_ _0792_ _0831_ VPWR VGND sg13g2_xor2_1
X_1903_ net457 net397 _0032_ VPWR VGND sg13g2_and2_1
X_2883_ _0734_ _0771_ _0772_ _0773_ VPWR VGND sg13g2_nor3_1
XFILLER_30_351 VPWR VGND sg13g2_decap_8
X_1834_ _1159_ _1150_ _1160_ VPWR VGND sg13g2_nor2b_1
X_1765_ _1093_ net465 DP_2.matrix\[41\] VPWR VGND sg13g2_nand2_1
X_1696_ _1026_ _0990_ _1024_ _1025_ VPWR VGND sg13g2_and3_1
X_2317_ VGND VPWR _0192_ _0194_ _0229_ _0228_ sg13g2_a21oi_1
Xheichips25_template_35 VPWR VGND uio_oe[2] sg13g2_tiehi
X_2248_ _1489_ VPWR _0161_ VGND _1444_ _1490_ sg13g2_o21ai_1
XFILLER_39_974 VPWR VGND sg13g2_decap_8
X_2179_ _1457_ _1458_ _1460_ _1461_ VPWR VGND sg13g2_or3_1
XFILLER_25_134 VPWR VGND sg13g2_decap_8
XFILLER_25_145 VPWR VGND sg13g2_fill_1
XFILLER_41_649 VPWR VGND sg13g2_decap_8
XFILLER_40_126 VPWR VGND sg13g2_decap_8
XFILLER_15_46 VPWR VGND sg13g2_decap_8
XFILLER_22_896 VPWR VGND sg13g2_decap_8
Xoutput23 net23 uio_out[6] VPWR VGND sg13g2_buf_1
XFILLER_0_211 VPWR VGND sg13g2_decap_8
XFILLER_1_723 VPWR VGND sg13g2_decap_8
XFILLER_49_727 VPWR VGND sg13g2_decap_8
XFILLER_0_277 VPWR VGND sg13g2_decap_8
XFILLER_48_237 VPWR VGND sg13g2_decap_8
XFILLER_45_900 VPWR VGND sg13g2_decap_8
XFILLER_17_602 VPWR VGND sg13g2_decap_8
XFILLER_29_473 VPWR VGND sg13g2_decap_8
XFILLER_17_624 VPWR VGND sg13g2_decap_8
XFILLER_45_977 VPWR VGND sg13g2_decap_8
XFILLER_44_465 VPWR VGND sg13g2_decap_8
XFILLER_17_657 VPWR VGND sg13g2_fill_2
XFILLER_17_679 VPWR VGND sg13g2_decap_4
XFILLER_16_167 VPWR VGND sg13g2_fill_2
XFILLER_16_178 VPWR VGND sg13g2_decap_4
XFILLER_13_841 VPWR VGND sg13g2_decap_8
XFILLER_9_823 VPWR VGND sg13g2_decap_8
X_1550_ _0881_ _0880_ _0884_ VPWR VGND sg13g2_nor2b_1
X_3220_ net522 VGND VPWR net65 mac1.sum_lvl3_ff\[31\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_3151_ net536 VGND VPWR net44 mac1.sum_lvl2_ff\[6\] clknet_leaf_25_clk sg13g2_dfrbpq_1
XFILLER_39_215 VPWR VGND sg13g2_decap_8
X_2102_ _1385_ _1362_ _1386_ VPWR VGND sg13g2_xor2_1
XFILLER_39_237 VPWR VGND sg13g2_decap_8
X_3082_ net520 VGND VPWR net269 mac1.products_ff\[69\] clknet_leaf_33_clk sg13g2_dfrbpq_1
XFILLER_36_900 VPWR VGND sg13g2_decap_8
XFILLER_48_793 VPWR VGND sg13g2_decap_8
X_2033_ _1320_ _1317_ _1326_ VPWR VGND _1319_ sg13g2_nand3b_1
XFILLER_36_977 VPWR VGND sg13g2_decap_8
XFILLER_22_137 VPWR VGND sg13g2_fill_1
X_2935_ VGND VPWR net373 _0820_ _0088_ net250 sg13g2_a21oi_1
X_2866_ _0756_ _0755_ _0751_ VPWR VGND sg13g2_nand2b_1
X_1817_ _1108_ _1114_ _1144_ VPWR VGND sg13g2_nor2_1
X_2797_ _0664_ _0690_ _0691_ VPWR VGND sg13g2_nor2_1
XFILLER_11_1024 VPWR VGND sg13g2_decap_4
X_1748_ VPWR _1077_ _1076_ VGND sg13g2_inv_1
X_1679_ _0967_ VPWR _1009_ VGND _0965_ _0968_ sg13g2_o21ai_1
XFILLER_27_911 VPWR VGND sg13g2_decap_8
XFILLER_26_421 VPWR VGND sg13g2_decap_8
XFILLER_26_56 VPWR VGND sg13g2_decap_8
XFILLER_27_988 VPWR VGND sg13g2_decap_8
XFILLER_41_424 VPWR VGND sg13g2_decap_8
XFILLER_42_958 VPWR VGND sg13g2_decap_8
XFILLER_42_22 VPWR VGND sg13g2_decap_8
XFILLER_9_119 VPWR VGND sg13g2_decap_8
XFILLER_10_866 VPWR VGND sg13g2_decap_8
XFILLER_6_804 VPWR VGND sg13g2_decap_8
XFILLER_5_303 VPWR VGND sg13g2_decap_8
XFILLER_49_513 VPWR VGND sg13g2_decap_8
XFILLER_1_597 VPWR VGND sg13g2_decap_8
XFILLER_18_944 VPWR VGND sg13g2_decap_8
XFILLER_36_218 VPWR VGND sg13g2_decap_8
XFILLER_33_903 VPWR VGND sg13g2_decap_8
XFILLER_44_273 VPWR VGND sg13g2_decap_8
XFILLER_17_487 VPWR VGND sg13g2_fill_1
XFILLER_32_402 VPWR VGND sg13g2_decap_4
XFILLER_32_424 VPWR VGND sg13g2_decap_8
XFILLER_32_435 VPWR VGND sg13g2_decap_4
XFILLER_32_446 VPWR VGND sg13g2_fill_2
XFILLER_20_619 VPWR VGND sg13g2_decap_8
XFILLER_34_1024 VPWR VGND sg13g2_decap_4
X_2720_ _0615_ _0616_ _0059_ VPWR VGND sg13g2_nor2b_1
X_2651_ _0549_ _0544_ _0547_ VPWR VGND sg13g2_xnor2_1
XFILLER_8_163 VPWR VGND sg13g2_decap_8
XFILLER_12_192 VPWR VGND sg13g2_fill_1
XFILLER_9_697 VPWR VGND sg13g2_decap_8
X_1602_ _0929_ VPWR _0934_ VGND _0930_ _0932_ sg13g2_o21ai_1
X_2582_ _0482_ _0450_ _0480_ _0481_ VPWR VGND sg13g2_and3_1
XFILLER_5_881 VPWR VGND sg13g2_decap_8
X_1533_ _0867_ net473 net406 VPWR VGND sg13g2_nand2_2
X_3203_ net511 VGND VPWR net66 mac1.sum_lvl1_ff\[82\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3134_ net534 VGND VPWR net73 mac1.sum_lvl1_ff\[41\] clknet_leaf_26_clk sg13g2_dfrbpq_1
X_3065_ net527 VGND VPWR _0118_ DP_2.matrix\[36\] clknet_leaf_30_clk sg13g2_dfrbpq_2
X_2016_ _1312_ mac1.sum_lvl3_ff\[9\] net181 VPWR VGND sg13g2_nand2_1
XFILLER_23_413 VPWR VGND sg13g2_decap_8
XFILLER_24_936 VPWR VGND sg13g2_decap_8
XFILLER_10_107 VPWR VGND sg13g2_fill_1
X_2918_ _0807_ _0784_ _0806_ _0783_ net383 VPWR VGND sg13g2_a22oi_1
XFILLER_12_14 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_30_clk clknet_3_4__leaf_clk clknet_leaf_30_clk VPWR VGND sg13g2_buf_8
X_2849_ net468 net486 net379 _0739_ VPWR VGND sg13g2_mux2_1
XFILLER_3_829 VPWR VGND sg13g2_decap_8
Xhold152 DP_2.matrix\[43\] VPWR VGND net192 sg13g2_dlygate4sd3_1
Xhold141 mac1.sum_lvl3_ff\[29\] VPWR VGND net181 sg13g2_dlygate4sd3_1
Xhold130 _0006_ VPWR VGND net170 sg13g2_dlygate4sd3_1
Xhold185 DP_1.matrix\[5\] VPWR VGND net225 sg13g2_dlygate4sd3_1
Xhold174 _0017_ VPWR VGND net214 sg13g2_dlygate4sd3_1
Xhold163 DP_2.matrix\[39\] VPWR VGND net203 sg13g2_dlygate4sd3_1
Xhold196 _0007_ VPWR VGND net236 sg13g2_dlygate4sd3_1
XFILLER_46_516 VPWR VGND sg13g2_decap_4
XFILLER_2_1000 VPWR VGND sg13g2_decap_8
XFILLER_27_763 VPWR VGND sg13g2_fill_1
XFILLER_15_914 VPWR VGND sg13g2_decap_8
XFILLER_26_251 VPWR VGND sg13g2_decap_8
XFILLER_42_733 VPWR VGND sg13g2_decap_8
XFILLER_30_906 VPWR VGND sg13g2_decap_8
XFILLER_41_298 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_21_clk clknet_3_6__leaf_clk clknet_leaf_21_clk VPWR VGND sg13g2_buf_8
XFILLER_6_678 VPWR VGND sg13g2_decap_8
XFILLER_38_8 VPWR VGND sg13g2_fill_1
XFILLER_2_895 VPWR VGND sg13g2_decap_8
XFILLER_49_354 VPWR VGND sg13g2_decap_8
XFILLER_18_785 VPWR VGND sg13g2_decap_8
XFILLER_21_917 VPWR VGND sg13g2_decap_8
XFILLER_33_766 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_12_clk clknet_3_3__leaf_clk clknet_leaf_12_clk VPWR VGND sg13g2_buf_8
X_2703_ _0598_ _0599_ _0600_ VPWR VGND sg13g2_nor2b_1
X_2634_ _0531_ _0532_ _0530_ _0533_ VPWR VGND sg13g2_nand3_1
X_2565_ _0430_ VPWR _0465_ VGND _0428_ _0431_ sg13g2_o21ai_1
X_1516_ _0850_ _0042_ _0845_ _0852_ VPWR VGND sg13g2_nand3_1
X_2496_ _0394_ _0395_ _0397_ _0398_ VPWR VGND sg13g2_or3_1
X_3117_ net534 VGND VPWR net95 mac1.sum_lvl1_ff\[4\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_3048_ net537 VGND VPWR _0101_ DP_1.matrix\[43\] clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_24_788 VPWR VGND sg13g2_decap_8
XFILLER_11_427 VPWR VGND sg13g2_decap_8
XFILLER_23_298 VPWR VGND sg13g2_decap_4
XFILLER_23_57 VPWR VGND sg13g2_decap_8
XFILLER_23_68 VPWR VGND sg13g2_fill_2
XFILLER_3_626 VPWR VGND sg13g2_decap_8
XFILLER_48_21 VPWR VGND sg13g2_decap_8
Xfanout440 net441 net440 VPWR VGND sg13g2_buf_2
Xfanout473 net276 net473 VPWR VGND sg13g2_buf_8
Xfanout462 net463 net462 VPWR VGND sg13g2_buf_8
Xfanout451 net220 net451 VPWR VGND sg13g2_buf_8
Xfanout484 net485 net484 VPWR VGND sg13g2_buf_8
XFILLER_47_836 VPWR VGND sg13g2_decap_8
Xfanout495 net227 net495 VPWR VGND sg13g2_buf_8
XFILLER_46_335 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_15_711 VPWR VGND sg13g2_decap_8
XFILLER_9_15 VPWR VGND sg13g2_fill_2
XFILLER_42_596 VPWR VGND sg13g2_fill_2
XFILLER_7_910 VPWR VGND sg13g2_decap_8
XFILLER_11_961 VPWR VGND sg13g2_decap_8
XFILLER_31_1027 VPWR VGND sg13g2_fill_2
XFILLER_10_482 VPWR VGND sg13g2_decap_8
XFILLER_7_987 VPWR VGND sg13g2_decap_8
XFILLER_9_1028 VPWR VGND sg13g2_fill_1
X_2350_ VGND VPWR _0225_ _0227_ _0261_ _0258_ sg13g2_a21oi_1
XFILLER_2_692 VPWR VGND sg13g2_decap_8
X_2281_ _0194_ _0161_ _0193_ VPWR VGND sg13g2_nand2b_1
Xclkbuf_leaf_1_clk clknet_3_0__leaf_clk clknet_leaf_1_clk VPWR VGND sg13g2_buf_8
XFILLER_29_4 VPWR VGND sg13g2_fill_2
XFILLER_38_803 VPWR VGND sg13g2_decap_4
XFILLER_49_151 VPWR VGND sg13g2_decap_8
XFILLER_21_703 VPWR VGND sg13g2_decap_8
XFILLER_33_541 VPWR VGND sg13g2_decap_4
XFILLER_20_202 VPWR VGND sg13g2_decap_8
X_1996_ net178 mac1.sum_lvl3_ff\[25\] _1296_ VPWR VGND sg13g2_nor2_1
XFILLER_9_280 VPWR VGND sg13g2_fill_1
X_2617_ _0511_ VPWR _0516_ VGND _0512_ _0514_ sg13g2_o21ai_1
XFILLER_0_629 VPWR VGND sg13g2_decap_8
X_2548_ _0448_ _0412_ _0065_ VPWR VGND sg13g2_xor2_1
X_2479_ _0361_ VPWR _0382_ VGND _0352_ _0362_ sg13g2_o21ai_1
XFILLER_29_847 VPWR VGND sg13g2_decap_8
XFILLER_44_806 VPWR VGND sg13g2_fill_2
XFILLER_29_858 VPWR VGND sg13g2_fill_1
XFILLER_44_817 VPWR VGND sg13g2_decap_8
XFILLER_18_79 VPWR VGND sg13g2_decap_8
XFILLER_11_202 VPWR VGND sg13g2_fill_2
XFILLER_12_714 VPWR VGND sg13g2_decap_8
XFILLER_8_718 VPWR VGND sg13g2_decap_8
XFILLER_11_224 VPWR VGND sg13g2_decap_8
XFILLER_7_206 VPWR VGND sg13g2_fill_2
Xclkload0 clkload0/Y clknet_3_6__leaf_clk VPWR VGND sg13g2_inv_2
XFILLER_4_924 VPWR VGND sg13g2_decap_8
XFILLER_3_412 VPWR VGND sg13g2_decap_8
XFILLER_3_434 VPWR VGND sg13g2_decap_8
XFILLER_47_666 VPWR VGND sg13g2_decap_8
XFILLER_19_324 VPWR VGND sg13g2_fill_1
XFILLER_43_894 VPWR VGND sg13g2_decap_8
XFILLER_30_500 VPWR VGND sg13g2_decap_8
X_1850_ _1175_ _1171_ _0072_ VPWR VGND sg13g2_xor2_1
X_1781_ _1072_ _1107_ _1070_ _1109_ VPWR VGND sg13g2_nand3_1
XFILLER_30_566 VPWR VGND sg13g2_decap_8
XFILLER_7_784 VPWR VGND sg13g2_decap_8
XFILLER_6_283 VPWR VGND sg13g2_fill_2
XFILLER_6_272 VPWR VGND sg13g2_fill_2
X_2402_ _0310_ VPWR _0311_ VGND _0284_ _0286_ sg13g2_o21ai_1
XFILLER_3_990 VPWR VGND sg13g2_decap_8
X_2333_ _0206_ VPWR _0244_ VGND _0203_ _0207_ sg13g2_o21ai_1
X_2264_ VGND VPWR _0177_ _0176_ _1494_ sg13g2_or2_1
X_2195_ _1476_ _1412_ _1477_ VPWR VGND sg13g2_xor2_1
XFILLER_37_143 VPWR VGND sg13g2_decap_8
XFILLER_38_677 VPWR VGND sg13g2_fill_2
XFILLER_19_880 VPWR VGND sg13g2_decap_8
X_1979_ _1283_ mac1.sum_lvl3_ff\[1\] mac1.sum_lvl3_ff\[21\] VPWR VGND sg13g2_nand2_1
XFILLER_20_25 VPWR VGND sg13g2_decap_8
XFILLER_1_905 VPWR VGND sg13g2_decap_8
XFILLER_0_426 VPWR VGND sg13g2_decap_8
XFILLER_49_909 VPWR VGND sg13g2_decap_8
Xhold12 mac1.sum_lvl1_ff\[48\] VPWR VGND net52 sg13g2_dlygate4sd3_1
XFILLER_29_34 VPWR VGND sg13g2_decap_4
Xhold23 mac1.products_ff\[82\] VPWR VGND net63 sg13g2_dlygate4sd3_1
Xhold34 mac1.products_ff\[70\] VPWR VGND net74 sg13g2_dlygate4sd3_1
Xhold56 mac1.products_ff\[8\] VPWR VGND net96 sg13g2_dlygate4sd3_1
Xhold45 mac1.products_ff\[83\] VPWR VGND net85 sg13g2_dlygate4sd3_1
Xhold78 mac1.sum_lvl1_ff\[0\] VPWR VGND net118 sg13g2_dlygate4sd3_1
Xhold89 mac1.sum_lvl1_ff\[43\] VPWR VGND net129 sg13g2_dlygate4sd3_1
XFILLER_21_1015 VPWR VGND sg13g2_decap_8
Xhold67 mac1.products_ff\[148\] VPWR VGND net107 sg13g2_dlygate4sd3_1
XFILLER_44_658 VPWR VGND sg13g2_fill_1
XFILLER_44_647 VPWR VGND sg13g2_decap_8
XFILLER_44_625 VPWR VGND sg13g2_decap_8
XFILLER_43_113 VPWR VGND sg13g2_decap_4
XFILLER_45_88 VPWR VGND sg13g2_decap_8
XFILLER_12_500 VPWR VGND sg13g2_decap_4
XFILLER_40_897 VPWR VGND sg13g2_decap_8
XFILLER_4_721 VPWR VGND sg13g2_decap_8
XFILLER_4_798 VPWR VGND sg13g2_decap_8
XFILLER_3_286 VPWR VGND sg13g2_decap_8
XFILLER_3_275 VPWR VGND sg13g2_fill_2
XFILLER_0_993 VPWR VGND sg13g2_decap_8
XFILLER_47_430 VPWR VGND sg13g2_decap_8
XFILLER_19_121 VPWR VGND sg13g2_decap_8
XFILLER_48_975 VPWR VGND sg13g2_decap_8
XFILLER_34_124 VPWR VGND sg13g2_decap_8
XFILLER_16_883 VPWR VGND sg13g2_decap_8
X_2951_ _0110_ net437 net374 VPWR VGND sg13g2_xnor2_1
XFILLER_37_1022 VPWR VGND sg13g2_decap_8
X_1902_ _0075_ _1217_ _1224_ VPWR VGND sg13g2_xnor2_1
X_2882_ net253 _0731_ _0772_ VPWR VGND sg13g2_nor2_1
X_1833_ _1159_ _1151_ _1158_ VPWR VGND sg13g2_xnor2_1
X_1764_ VGND VPWR net415 net459 _1092_ _1060_ sg13g2_a21oi_1
X_1695_ _1001_ VPWR _1025_ VGND _1021_ _1023_ sg13g2_o21ai_1
X_2316_ _0226_ _0199_ _0228_ VPWR VGND sg13g2_xor2_1
XFILLER_39_953 VPWR VGND sg13g2_decap_8
X_2247_ _0150_ VPWR _0160_ VGND _1446_ _0151_ sg13g2_o21ai_1
Xheichips25_template_36 VPWR VGND uio_oe[3] sg13g2_tiehi
XFILLER_25_102 VPWR VGND sg13g2_decap_8
X_2178_ _1460_ net395 net442 net440 net399 VPWR VGND sg13g2_a22oi_1
XFILLER_38_496 VPWR VGND sg13g2_decap_4
XFILLER_26_669 VPWR VGND sg13g2_decap_8
XFILLER_34_680 VPWR VGND sg13g2_decap_8
XFILLER_22_875 VPWR VGND sg13g2_decap_8
XFILLER_1_702 VPWR VGND sg13g2_decap_8
Xoutput24 net24 uio_out[7] VPWR VGND sg13g2_buf_1
XFILLER_49_706 VPWR VGND sg13g2_decap_8
XFILLER_48_216 VPWR VGND sg13g2_decap_8
XFILLER_0_256 VPWR VGND sg13g2_decap_8
XFILLER_1_779 VPWR VGND sg13g2_decap_8
XFILLER_45_956 VPWR VGND sg13g2_decap_8
XFILLER_16_135 VPWR VGND sg13g2_decap_8
XFILLER_9_802 VPWR VGND sg13g2_decap_8
XFILLER_12_330 VPWR VGND sg13g2_decap_8
XFILLER_25_691 VPWR VGND sg13g2_fill_2
XFILLER_31_127 VPWR VGND sg13g2_fill_2
XFILLER_8_312 VPWR VGND sg13g2_decap_8
XFILLER_8_323 VPWR VGND sg13g2_fill_1
XFILLER_12_385 VPWR VGND sg13g2_decap_4
XFILLER_13_897 VPWR VGND sg13g2_decap_8
XFILLER_9_879 VPWR VGND sg13g2_decap_8
Xclkbuf_3_1__f_clk clknet_0_clk clknet_3_1__leaf_clk VPWR VGND sg13g2_buf_8
X_3150_ net535 VGND VPWR net101 mac1.sum_lvl2_ff\[5\] clknet_leaf_28_clk sg13g2_dfrbpq_1
XFILLER_0_790 VPWR VGND sg13g2_decap_8
X_3081_ net521 VGND VPWR _0042_ mac1.products_ff\[68\] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_2101_ _1385_ net452 net388 VPWR VGND sg13g2_nand2_1
XFILLER_48_772 VPWR VGND sg13g2_decap_8
XFILLER_11_4 VPWR VGND sg13g2_decap_8
X_2032_ _1320_ VPWR _1325_ VGND _1316_ _1319_ sg13g2_o21ai_1
XFILLER_47_260 VPWR VGND sg13g2_decap_8
XFILLER_35_400 VPWR VGND sg13g2_decap_8
XFILLER_36_956 VPWR VGND sg13g2_decap_8
XFILLER_23_617 VPWR VGND sg13g2_decap_8
XFILLER_23_639 VPWR VGND sg13g2_fill_1
X_2934_ _0749_ _0747_ _0820_ VPWR VGND sg13g2_xor2_1
XFILLER_30_182 VPWR VGND sg13g2_decap_8
X_2865_ _0752_ VPWR _0755_ VGND _0753_ _0754_ sg13g2_o21ai_1
XFILLER_11_1003 VPWR VGND sg13g2_decap_8
X_1816_ _1143_ _1140_ _1142_ VPWR VGND sg13g2_nand2_1
X_2796_ _0690_ _0649_ _0688_ VPWR VGND sg13g2_xnor2_1
X_1747_ _1076_ _1038_ _1073_ VPWR VGND sg13g2_xnor2_1
X_1678_ _1008_ _1003_ _1007_ VPWR VGND sg13g2_xnor2_1
XFILLER_39_772 VPWR VGND sg13g2_decap_8
XFILLER_38_260 VPWR VGND sg13g2_fill_2
XFILLER_38_282 VPWR VGND sg13g2_fill_1
XFILLER_26_35 VPWR VGND sg13g2_decap_8
XFILLER_26_444 VPWR VGND sg13g2_fill_1
XFILLER_27_967 VPWR VGND sg13g2_decap_8
XFILLER_42_937 VPWR VGND sg13g2_decap_8
XFILLER_26_79 VPWR VGND sg13g2_fill_1
XFILLER_13_127 VPWR VGND sg13g2_decap_4
XFILLER_10_845 VPWR VGND sg13g2_decap_8
XFILLER_1_576 VPWR VGND sg13g2_decap_8
XFILLER_37_709 VPWR VGND sg13g2_decap_4
XFILLER_45_720 VPWR VGND sg13g2_fill_1
XFILLER_18_923 VPWR VGND sg13g2_decap_8
XFILLER_17_477 VPWR VGND sg13g2_fill_2
XFILLER_33_959 VPWR VGND sg13g2_decap_8
XFILLER_13_650 VPWR VGND sg13g2_decap_8
XFILLER_34_1003 VPWR VGND sg13g2_decap_8
XFILLER_12_160 VPWR VGND sg13g2_decap_4
X_2650_ _0548_ _0547_ _0544_ VPWR VGND sg13g2_nand2b_1
XFILLER_9_687 VPWR VGND sg13g2_fill_1
X_1601_ _0929_ _0930_ _0932_ _0933_ VPWR VGND sg13g2_or3_1
XFILLER_5_860 VPWR VGND sg13g2_decap_8
X_2581_ _0456_ VPWR _0481_ VGND _0477_ _0479_ sg13g2_o21ai_1
X_1532_ _0866_ net406 net474 net408 net472 VPWR VGND sg13g2_a22oi_1
X_3202_ net513 VGND VPWR net88 mac1.sum_lvl1_ff\[81\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_41_1018 VPWR VGND sg13g2_decap_8
X_3133_ net526 VGND VPWR net135 mac1.sum_lvl1_ff\[40\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_3064_ net539 VGND VPWR _0117_ DP_2.matrix\[7\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_27_219 VPWR VGND sg13g2_decap_8
X_2015_ _1307_ _1309_ _1311_ VPWR VGND sg13g2_nor2_1
XFILLER_24_915 VPWR VGND sg13g2_decap_8
X_2917_ net404 net424 _0781_ _0806_ VPWR VGND sg13g2_mux2_1
XFILLER_12_59 VPWR VGND sg13g2_fill_2
X_2848_ _0733_ VPWR _0738_ VGND _0736_ _0737_ sg13g2_o21ai_1
X_2779_ VGND VPWR _0609_ _0642_ _0674_ _0643_ sg13g2_a21oi_1
XFILLER_3_808 VPWR VGND sg13g2_decap_8
Xhold153 DP_1.matrix\[80\] VPWR VGND net193 sg13g2_dlygate4sd3_1
Xhold120 DP_1.matrix\[6\] VPWR VGND net160 sg13g2_dlygate4sd3_1
Xhold142 _1313_ VPWR VGND net182 sg13g2_dlygate4sd3_1
Xhold131 mac1.sum_lvl2_ff\[14\] VPWR VGND net171 sg13g2_dlygate4sd3_1
Xhold164 DP_1.matrix\[41\] VPWR VGND net204 sg13g2_dlygate4sd3_1
Xhold175 DP_1.matrix\[74\] VPWR VGND net215 sg13g2_dlygate4sd3_1
Xhold186 DP_1.matrix\[4\] VPWR VGND net226 sg13g2_dlygate4sd3_1
Xhold197 DP_2.matrix\[4\] VPWR VGND net237 sg13g2_dlygate4sd3_1
XFILLER_42_756 VPWR VGND sg13g2_decap_4
XFILLER_14_447 VPWR VGND sg13g2_decap_8
XFILLER_41_244 VPWR VGND sg13g2_fill_2
XFILLER_14_458 VPWR VGND sg13g2_fill_2
XFILLER_41_288 VPWR VGND sg13g2_fill_1
XFILLER_10_631 VPWR VGND sg13g2_decap_8
XFILLER_6_657 VPWR VGND sg13g2_decap_8
XFILLER_5_134 VPWR VGND sg13g2_decap_8
XFILLER_1_362 VPWR VGND sg13g2_decap_4
XFILLER_2_874 VPWR VGND sg13g2_decap_8
XFILLER_37_506 VPWR VGND sg13g2_decap_8
XFILLER_37_539 VPWR VGND sg13g2_decap_4
XFILLER_17_252 VPWR VGND sg13g2_decap_8
XFILLER_45_594 VPWR VGND sg13g2_fill_2
XFILLER_17_296 VPWR VGND sg13g2_fill_2
XFILLER_32_222 VPWR VGND sg13g2_decap_8
XFILLER_20_406 VPWR VGND sg13g2_fill_1
XFILLER_32_288 VPWR VGND sg13g2_decap_8
XFILLER_32_299 VPWR VGND sg13g2_fill_2
X_2702_ _0594_ VPWR _0599_ VGND _0596_ _0597_ sg13g2_o21ai_1
XFILLER_9_495 VPWR VGND sg13g2_decap_8
X_2633_ _0483_ VPWR _0532_ VGND _0417_ _0484_ sg13g2_o21ai_1
X_2564_ _0464_ _0458_ _0463_ VPWR VGND sg13g2_xnor2_1
X_1515_ _0851_ _0845_ _0042_ VPWR VGND sg13g2_nand2_1
X_2495_ _0397_ net436 net484 net481 net439 VPWR VGND sg13g2_a22oi_1
X_3116_ net525 VGND VPWR net133 mac1.sum_lvl1_ff\[3\] clknet_leaf_27_clk sg13g2_dfrbpq_1
XFILLER_28_539 VPWR VGND sg13g2_decap_4
X_3047_ net535 VGND VPWR _0100_ DP_1.matrix\[42\] clknet_leaf_22_clk sg13g2_dfrbpq_2
XFILLER_36_550 VPWR VGND sg13g2_decap_8
XFILLER_23_25 VPWR VGND sg13g2_decap_4
XFILLER_23_277 VPWR VGND sg13g2_decap_8
XFILLER_20_995 VPWR VGND sg13g2_decap_8
XFILLER_3_605 VPWR VGND sg13g2_decap_8
XFILLER_2_126 VPWR VGND sg13g2_fill_2
Xfanout430 DP_2.matrix\[3\] net430 VPWR VGND sg13g2_buf_1
Xfanout441 DP_1.matrix\[79\] net441 VPWR VGND sg13g2_buf_8
XFILLER_47_815 VPWR VGND sg13g2_decap_8
Xfanout474 net196 net474 VPWR VGND sg13g2_buf_8
Xfanout452 net453 net452 VPWR VGND sg13g2_buf_8
XFILLER_24_1013 VPWR VGND sg13g2_decap_8
Xfanout463 net211 net463 VPWR VGND sg13g2_buf_8
Xfanout496 net193 net496 VPWR VGND sg13g2_buf_8
XFILLER_19_539 VPWR VGND sg13g2_decap_8
Xfanout485 net226 net485 VPWR VGND sg13g2_buf_8
XFILLER_15_701 VPWR VGND sg13g2_decap_4
XFILLER_42_575 VPWR VGND sg13g2_decap_8
XFILLER_30_737 VPWR VGND sg13g2_fill_1
XFILLER_11_940 VPWR VGND sg13g2_decap_8
XFILLER_31_1006 VPWR VGND sg13g2_decap_8
XFILLER_7_966 VPWR VGND sg13g2_decap_8
XFILLER_2_671 VPWR VGND sg13g2_decap_8
X_2280_ _0193_ _0162_ _0191_ VPWR VGND sg13g2_xnor2_1
XFILLER_49_130 VPWR VGND sg13g2_decap_8
XFILLER_25_509 VPWR VGND sg13g2_fill_2
XFILLER_33_520 VPWR VGND sg13g2_fill_2
XFILLER_21_726 VPWR VGND sg13g2_fill_1
X_1995_ VGND VPWR _1292_ _1294_ _1295_ _1293_ sg13g2_a21oi_1
XFILLER_20_225 VPWR VGND sg13g2_fill_1
X_2616_ _0511_ _0512_ _0514_ _0515_ VPWR VGND sg13g2_or3_1
XFILLER_0_608 VPWR VGND sg13g2_decap_8
X_2547_ _0446_ _0447_ _0448_ VPWR VGND sg13g2_nor2b_1
X_2478_ _0381_ _0369_ _0380_ VPWR VGND sg13g2_xnor2_1
XFILLER_29_804 VPWR VGND sg13g2_decap_8
XFILLER_18_25 VPWR VGND sg13g2_decap_8
XFILLER_18_58 VPWR VGND sg13g2_decap_8
XFILLER_28_347 VPWR VGND sg13g2_fill_1
XFILLER_34_13 VPWR VGND sg13g2_decap_8
XFILLER_36_380 VPWR VGND sg13g2_decap_8
XFILLER_34_24 VPWR VGND sg13g2_fill_1
XFILLER_24_575 VPWR VGND sg13g2_decap_8
XFILLER_11_269 VPWR VGND sg13g2_fill_1
Xclkload1 clknet_3_7__leaf_clk clkload1/X VPWR VGND sg13g2_buf_8
XFILLER_4_903 VPWR VGND sg13g2_decap_8
XFILLER_3_479 VPWR VGND sg13g2_decap_4
XFILLER_19_303 VPWR VGND sg13g2_decap_8
XFILLER_28_881 VPWR VGND sg13g2_decap_8
XFILLER_43_873 VPWR VGND sg13g2_decap_8
XFILLER_42_350 VPWR VGND sg13g2_fill_2
XFILLER_42_383 VPWR VGND sg13g2_decap_8
X_1780_ VGND VPWR _1070_ _1072_ _1108_ _1107_ sg13g2_a21oi_1
XFILLER_11_781 VPWR VGND sg13g2_decap_4
XFILLER_7_763 VPWR VGND sg13g2_decap_8
XFILLER_6_295 VPWR VGND sg13g2_decap_8
XFILLER_41_4 VPWR VGND sg13g2_decap_8
X_2401_ _0308_ _0294_ _0310_ VPWR VGND sg13g2_xor2_1
X_2332_ _0243_ _0237_ _0242_ VPWR VGND sg13g2_xnor2_1
X_2263_ _0176_ net442 net389 VPWR VGND sg13g2_nand2_1
X_2194_ _1476_ _1473_ _1475_ VPWR VGND sg13g2_nand2_1
XFILLER_37_199 VPWR VGND sg13g2_decap_4
XFILLER_34_884 VPWR VGND sg13g2_decap_8
XFILLER_21_556 VPWR VGND sg13g2_decap_8
XFILLER_33_394 VPWR VGND sg13g2_decap_8
X_1978_ _1282_ net166 net153 VPWR VGND sg13g2_nand2_1
XFILLER_0_405 VPWR VGND sg13g2_decap_8
Xhold13 mac1.products_ff\[80\] VPWR VGND net53 sg13g2_dlygate4sd3_1
Xhold24 mac1.sum_lvl1_ff\[37\] VPWR VGND net64 sg13g2_dlygate4sd3_1
Xhold46 mac1.sum_lvl1_ff\[8\] VPWR VGND net86 sg13g2_dlygate4sd3_1
Xhold35 mac1.sum_lvl2_ff\[52\] VPWR VGND net75 sg13g2_dlygate4sd3_1
Xhold57 mac1.sum_lvl1_ff\[12\] VPWR VGND net97 sg13g2_dlygate4sd3_1
Xhold68 mac1.products_ff\[141\] VPWR VGND net108 sg13g2_dlygate4sd3_1
Xhold79 mac1.products_ff\[140\] VPWR VGND net119 sg13g2_dlygate4sd3_1
XFILLER_29_79 VPWR VGND sg13g2_decap_8
XFILLER_29_623 VPWR VGND sg13g2_fill_2
XFILLER_44_604 VPWR VGND sg13g2_decap_8
XFILLER_16_328 VPWR VGND sg13g2_decap_4
XFILLER_28_177 VPWR VGND sg13g2_fill_1
XFILLER_43_169 VPWR VGND sg13g2_decap_8
XFILLER_40_876 VPWR VGND sg13g2_decap_8
XFILLER_12_578 VPWR VGND sg13g2_decap_8
XFILLER_12_589 VPWR VGND sg13g2_fill_1
XFILLER_4_700 VPWR VGND sg13g2_decap_8
XFILLER_3_210 VPWR VGND sg13g2_decap_8
XFILLER_4_777 VPWR VGND sg13g2_decap_8
XFILLER_0_972 VPWR VGND sg13g2_decap_8
XFILLER_48_954 VPWR VGND sg13g2_decap_8
XFILLER_19_100 VPWR VGND sg13g2_decap_4
XFILLER_16_862 VPWR VGND sg13g2_decap_8
XFILLER_37_1001 VPWR VGND sg13g2_decap_8
X_2950_ _0829_ VPWR _0093_ VGND _0775_ _0830_ sg13g2_o21ai_1
XFILLER_43_692 VPWR VGND sg13g2_fill_2
XFILLER_15_383 VPWR VGND sg13g2_decap_8
XFILLER_30_320 VPWR VGND sg13g2_decap_8
X_2881_ net499 net379 _0771_ VPWR VGND sg13g2_nor2_1
X_1901_ _1224_ _1218_ _1223_ VPWR VGND sg13g2_xnor2_1
X_1832_ _1158_ _1152_ _1157_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_887 VPWR VGND sg13g2_decap_8
X_1763_ _1064_ VPWR _1091_ VGND _1058_ _1065_ sg13g2_o21ai_1
XFILLER_7_582 VPWR VGND sg13g2_decap_4
XFILLER_7_571 VPWR VGND sg13g2_fill_2
X_1694_ _1001_ _1021_ _1023_ _1024_ VPWR VGND sg13g2_or3_1
XFILLER_44_1027 VPWR VGND sg13g2_fill_2
X_2315_ _0227_ _0226_ _0199_ VPWR VGND sg13g2_nand2b_1
XFILLER_39_932 VPWR VGND sg13g2_decap_8
X_2246_ _0155_ VPWR _0159_ VGND _1479_ _0157_ sg13g2_o21ai_1
Xheichips25_template_37 VPWR VGND uio_oe[4] sg13g2_tiehi
XFILLER_38_453 VPWR VGND sg13g2_fill_2
XFILLER_26_648 VPWR VGND sg13g2_decap_8
X_2177_ net442 net440 net399 _1459_ VPWR VGND net395 sg13g2_nand4_1
XFILLER_15_15 VPWR VGND sg13g2_fill_2
XFILLER_25_169 VPWR VGND sg13g2_decap_4
XFILLER_21_320 VPWR VGND sg13g2_decap_8
XFILLER_21_386 VPWR VGND sg13g2_decap_8
Xoutput25 net25 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_1_758 VPWR VGND sg13g2_decap_8
XFILLER_5_1021 VPWR VGND sg13g2_decap_8
XFILLER_29_442 VPWR VGND sg13g2_decap_4
XFILLER_45_935 VPWR VGND sg13g2_decap_8
XFILLER_16_114 VPWR VGND sg13g2_fill_2
XFILLER_17_659 VPWR VGND sg13g2_fill_1
XFILLER_16_169 VPWR VGND sg13g2_fill_1
XFILLER_31_106 VPWR VGND sg13g2_decap_8
XFILLER_24_180 VPWR VGND sg13g2_fill_1
XFILLER_25_681 VPWR VGND sg13g2_decap_4
XFILLER_13_876 VPWR VGND sg13g2_decap_8
XFILLER_24_191 VPWR VGND sg13g2_decap_8
XFILLER_9_858 VPWR VGND sg13g2_decap_8
XFILLER_8_379 VPWR VGND sg13g2_decap_8
XFILLER_4_563 VPWR VGND sg13g2_decap_4
X_3080_ net538 VGND VPWR _0133_ DP_2.matrix\[79\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_2100_ _1384_ net452 net386 VPWR VGND sg13g2_nand2_1
XFILLER_48_751 VPWR VGND sg13g2_decap_8
X_2031_ net291 mac1.sum_lvl3_ff\[12\] _1324_ VPWR VGND sg13g2_xor2_1
XFILLER_36_935 VPWR VGND sg13g2_decap_8
XFILLER_35_467 VPWR VGND sg13g2_fill_2
XFILLER_35_489 VPWR VGND sg13g2_fill_2
X_2933_ net488 net373 _0819_ VPWR VGND sg13g2_nor2_1
X_2864_ net376 VPWR _0754_ VGND net485 _0731_ sg13g2_o21ai_1
X_2795_ _0649_ _0688_ _0689_ VPWR VGND sg13g2_nor2_1
X_1815_ VPWR _1142_ _1141_ VGND sg13g2_inv_1
X_1746_ _1075_ _1038_ _1073_ VPWR VGND sg13g2_nand2_1
X_1677_ _1007_ _0958_ _1005_ VPWR VGND sg13g2_xnor2_1
XFILLER_39_751 VPWR VGND sg13g2_decap_8
X_2229_ _1498_ VPWR _0143_ VGND _0139_ _0141_ sg13g2_o21ai_1
XFILLER_27_946 VPWR VGND sg13g2_decap_8
XFILLER_26_456 VPWR VGND sg13g2_decap_8
XFILLER_42_916 VPWR VGND sg13g2_decap_8
XFILLER_22_651 VPWR VGND sg13g2_decap_8
XFILLER_10_824 VPWR VGND sg13g2_decap_8
XFILLER_6_839 VPWR VGND sg13g2_decap_8
XFILLER_3_18 VPWR VGND sg13g2_decap_8
XFILLER_1_555 VPWR VGND sg13g2_decap_8
XFILLER_49_548 VPWR VGND sg13g2_decap_4
XFILLER_49_559 VPWR VGND sg13g2_decap_8
XFILLER_18_902 VPWR VGND sg13g2_decap_8
XFILLER_45_732 VPWR VGND sg13g2_decap_8
XFILLER_44_220 VPWR VGND sg13g2_fill_2
XFILLER_18_979 VPWR VGND sg13g2_decap_8
XFILLER_33_938 VPWR VGND sg13g2_decap_8
XFILLER_16_80 VPWR VGND sg13g2_decap_4
XFILLER_32_448 VPWR VGND sg13g2_fill_1
XFILLER_8_121 VPWR VGND sg13g2_decap_4
XFILLER_13_684 VPWR VGND sg13g2_fill_2
X_1600_ _0932_ net463 net419 net464 net414 VPWR VGND sg13g2_a22oi_1
XFILLER_8_198 VPWR VGND sg13g2_fill_2
X_2580_ _0456_ _0477_ _0479_ _0480_ VPWR VGND sg13g2_or3_1
X_1531_ _0045_ _0852_ _0864_ VPWR VGND sg13g2_xnor2_1
X_3201_ net512 VGND VPWR net46 mac1.sum_lvl1_ff\[80\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3132_ net525 VGND VPWR net69 mac1.sum_lvl1_ff\[39\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_3063_ net538 VGND VPWR _0116_ DP_2.matrix\[6\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_48_592 VPWR VGND sg13g2_decap_8
X_2014_ _1309_ net241 _0030_ VPWR VGND sg13g2_nor2b_1
XFILLER_36_743 VPWR VGND sg13g2_decap_8
XFILLER_36_754 VPWR VGND sg13g2_fill_1
XFILLER_35_286 VPWR VGND sg13g2_decap_8
XFILLER_35_297 VPWR VGND sg13g2_fill_2
X_2916_ VGND VPWR _0805_ _0804_ _0788_ sg13g2_or2_1
XFILLER_12_16 VPWR VGND sg13g2_fill_1
X_2847_ net376 VPWR _0737_ VGND net483 _0731_ sg13g2_o21ai_1
X_2778_ _0671_ _0670_ _0673_ VPWR VGND sg13g2_xor2_1
Xhold110 mac1.products_ff\[2\] VPWR VGND net150 sg13g2_dlygate4sd3_1
Xhold121 mac1.sum_lvl2_ff\[0\] VPWR VGND net161 sg13g2_dlygate4sd3_1
Xhold143 _0031_ VPWR VGND net183 sg13g2_dlygate4sd3_1
X_1729_ _1058_ _1053_ _1057_ VPWR VGND sg13g2_xnor2_1
Xhold132 _1279_ VPWR VGND net172 sg13g2_dlygate4sd3_1
Xhold176 DP_1.matrix\[7\] VPWR VGND net216 sg13g2_dlygate4sd3_1
Xhold165 DP_1.matrix\[38\] VPWR VGND net205 sg13g2_dlygate4sd3_1
Xhold154 DP_1.matrix\[0\] VPWR VGND net194 sg13g2_dlygate4sd3_1
Xhold187 DP_2.matrix\[8\] VPWR VGND net227 sg13g2_dlygate4sd3_1
Xhold198 DP_2.matrix\[40\] VPWR VGND net238 sg13g2_dlygate4sd3_1
XFILLER_39_592 VPWR VGND sg13g2_decap_4
XFILLER_27_754 VPWR VGND sg13g2_decap_8
XFILLER_15_949 VPWR VGND sg13g2_decap_8
XFILLER_41_267 VPWR VGND sg13g2_decap_8
XFILLER_23_982 VPWR VGND sg13g2_decap_8
XFILLER_10_654 VPWR VGND sg13g2_decap_8
XFILLER_6_603 VPWR VGND sg13g2_decap_8
XFILLER_10_676 VPWR VGND sg13g2_decap_8
XFILLER_10_665 VPWR VGND sg13g2_fill_2
XFILLER_6_636 VPWR VGND sg13g2_decap_8
XFILLER_5_168 VPWR VGND sg13g2_decap_4
XFILLER_2_853 VPWR VGND sg13g2_decap_8
XFILLER_49_312 VPWR VGND sg13g2_decap_8
XFILLER_33_735 VPWR VGND sg13g2_decap_8
XFILLER_32_234 VPWR VGND sg13g2_decap_8
XFILLER_14_982 VPWR VGND sg13g2_decap_8
X_2701_ _0594_ _0596_ _0597_ _0598_ VPWR VGND sg13g2_nor3_1
XFILLER_41_790 VPWR VGND sg13g2_fill_2
XFILLER_13_492 VPWR VGND sg13g2_decap_8
X_2632_ _0455_ VPWR _0531_ VGND _0527_ _0529_ sg13g2_o21ai_1
X_2563_ _0463_ _0422_ _0460_ VPWR VGND sg13g2_xnor2_1
X_1514_ net474 net417 _0042_ VPWR VGND sg13g2_and2_1
X_2494_ net484 net481 net439 _0396_ VPWR VGND net436 sg13g2_nand4_1
XFILLER_4_94 VPWR VGND sg13g2_decap_8
X_3115_ net525 VGND VPWR net150 mac1.sum_lvl1_ff\[2\] clknet_leaf_32_clk sg13g2_dfrbpq_1
XFILLER_28_507 VPWR VGND sg13g2_decap_8
X_3046_ net527 VGND VPWR _0099_ DP_1.matrix\[41\] clknet_leaf_22_clk sg13g2_dfrbpq_2
XFILLER_36_573 VPWR VGND sg13g2_decap_8
XFILLER_12_919 VPWR VGND sg13g2_decap_8
XFILLER_20_974 VPWR VGND sg13g2_decap_8
XFILLER_2_149 VPWR VGND sg13g2_decap_8
Xfanout431 net223 net431 VPWR VGND sg13g2_buf_8
Xfanout420 DP_2.matrix\[36\] net420 VPWR VGND sg13g2_buf_1
XFILLER_48_67 VPWR VGND sg13g2_decap_4
XFILLER_48_56 VPWR VGND sg13g2_decap_8
Xfanout475 DP_1.matrix\[36\] net475 VPWR VGND sg13g2_buf_1
Xfanout464 net204 net464 VPWR VGND sg13g2_buf_8
Xfanout453 net215 net453 VPWR VGND sg13g2_buf_8
Xfanout442 net443 net442 VPWR VGND sg13g2_buf_8
XFILLER_46_304 VPWR VGND sg13g2_decap_8
Xfanout497 DP_1.matrix\[80\] net497 VPWR VGND sg13g2_buf_1
Xfanout486 net260 net486 VPWR VGND sg13g2_buf_8
XFILLER_42_510 VPWR VGND sg13g2_decap_8
XFILLER_30_705 VPWR VGND sg13g2_decap_4
XFILLER_42_598 VPWR VGND sg13g2_fill_1
XFILLER_14_278 VPWR VGND sg13g2_decap_8
XFILLER_7_945 VPWR VGND sg13g2_decap_8
XFILLER_11_996 VPWR VGND sg13g2_decap_8
XFILLER_6_466 VPWR VGND sg13g2_decap_8
XFILLER_9_1019 VPWR VGND sg13g2_decap_8
XFILLER_2_650 VPWR VGND sg13g2_decap_8
XFILLER_29_6 VPWR VGND sg13g2_fill_1
XFILLER_49_186 VPWR VGND sg13g2_decap_8
XFILLER_33_587 VPWR VGND sg13g2_decap_8
X_1994_ net218 _1292_ _0026_ VPWR VGND sg13g2_xor2_1
XFILLER_9_260 VPWR VGND sg13g2_decap_4
X_2615_ _0514_ net434 net477 net500 net438 VPWR VGND sg13g2_a22oi_1
XFILLER_47_1025 VPWR VGND sg13g2_decap_4
X_2546_ _0413_ VPWR _0447_ VGND _0444_ _0445_ sg13g2_o21ai_1
X_2477_ _0380_ _0377_ _0379_ VPWR VGND sg13g2_nand2_1
X_3029_ net527 VGND VPWR _0082_ DP_1.matrix\[44\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_37_882 VPWR VGND sg13g2_decap_8
XFILLER_12_749 VPWR VGND sg13g2_decap_4
XFILLER_7_208 VPWR VGND sg13g2_fill_1
Xclkload2 clkload2/Y clknet_leaf_1_clk VPWR VGND sg13g2_inv_8
XFILLER_4_959 VPWR VGND sg13g2_decap_8
XFILLER_19_337 VPWR VGND sg13g2_fill_2
XFILLER_35_819 VPWR VGND sg13g2_decap_8
XFILLER_27_370 VPWR VGND sg13g2_decap_8
XFILLER_34_318 VPWR VGND sg13g2_decap_8
XFILLER_43_852 VPWR VGND sg13g2_decap_8
XFILLER_15_587 VPWR VGND sg13g2_fill_2
XFILLER_30_535 VPWR VGND sg13g2_decap_4
XFILLER_24_91 VPWR VGND sg13g2_decap_8
XFILLER_7_742 VPWR VGND sg13g2_decap_8
XFILLER_6_285 VPWR VGND sg13g2_fill_1
X_2400_ _0309_ _0294_ _0308_ VPWR VGND sg13g2_nand2_1
XFILLER_34_4 VPWR VGND sg13g2_decap_4
X_2331_ _0241_ _0238_ _0242_ VPWR VGND sg13g2_xor2_1
X_2262_ _0175_ net448 net384 VPWR VGND sg13g2_nand2_1
X_2193_ _1472_ _1471_ _1441_ _1475_ VPWR VGND sg13g2_a21o_1
XFILLER_37_112 VPWR VGND sg13g2_decap_8
XFILLER_25_329 VPWR VGND sg13g2_decap_8
XFILLER_37_167 VPWR VGND sg13g2_fill_1
XFILLER_34_863 VPWR VGND sg13g2_decap_8
XFILLER_21_524 VPWR VGND sg13g2_decap_8
XFILLER_14_1024 VPWR VGND sg13g2_decap_4
X_1977_ net161 mac1.sum_lvl2_ff\[19\] _0000_ VPWR VGND sg13g2_xor2_1
X_2529_ net481 net480 net439 _0430_ VPWR VGND net435 sg13g2_nand4_1
Xhold14 mac1.sum_lvl1_ff\[78\] VPWR VGND net54 sg13g2_dlygate4sd3_1
Xhold47 mac1.products_ff\[6\] VPWR VGND net87 sg13g2_dlygate4sd3_1
Xhold25 mac1.sum_lvl2_ff\[49\] VPWR VGND net65 sg13g2_dlygate4sd3_1
Xhold36 mac1.sum_lvl2_ff\[53\] VPWR VGND net76 sg13g2_dlygate4sd3_1
XFILLER_29_602 VPWR VGND sg13g2_decap_8
Xhold58 mac1.sum_lvl1_ff\[41\] VPWR VGND net98 sg13g2_dlygate4sd3_1
Xhold69 mac1.sum_lvl1_ff\[79\] VPWR VGND net109 sg13g2_dlygate4sd3_1
XFILLER_28_112 VPWR VGND sg13g2_decap_8
XFILLER_28_123 VPWR VGND sg13g2_fill_2
XFILLER_29_646 VPWR VGND sg13g2_decap_8
XFILLER_45_13 VPWR VGND sg13g2_decap_8
XFILLER_28_167 VPWR VGND sg13g2_fill_1
XFILLER_43_148 VPWR VGND sg13g2_decap_8
XFILLER_25_885 VPWR VGND sg13g2_decap_8
XFILLER_40_855 VPWR VGND sg13g2_decap_8
XFILLER_12_524 VPWR VGND sg13g2_decap_8
XFILLER_12_535 VPWR VGND sg13g2_fill_1
XFILLER_6_29 VPWR VGND sg13g2_decap_8
XFILLER_4_756 VPWR VGND sg13g2_decap_8
XFILLER_0_951 VPWR VGND sg13g2_decap_8
XFILLER_48_933 VPWR VGND sg13g2_decap_8
XFILLER_47_465 VPWR VGND sg13g2_decap_8
XFILLER_47_476 VPWR VGND sg13g2_fill_1
XFILLER_19_178 VPWR VGND sg13g2_decap_4
XFILLER_16_841 VPWR VGND sg13g2_decap_8
XFILLER_43_671 VPWR VGND sg13g2_fill_1
XFILLER_34_159 VPWR VGND sg13g2_decap_8
X_2880_ DP_1.Q_range.out_data\[3\] DP_1.Q_range.out_data\[5\] _0766_ _0769_ _0770_
+ VPWR VGND sg13g2_and4_1
X_1900_ _1223_ _1210_ _1222_ VPWR VGND sg13g2_xnor2_1
XFILLER_42_192 VPWR VGND sg13g2_fill_1
X_1831_ _1154_ _1156_ _1157_ VPWR VGND sg13g2_nor2_1
XFILLER_30_365 VPWR VGND sg13g2_decap_8
X_1762_ _1088_ _1080_ _1090_ VPWR VGND sg13g2_xor2_1
X_1693_ VGND VPWR _1019_ _1020_ _1023_ _1002_ sg13g2_a21oi_1
XFILLER_44_1006 VPWR VGND sg13g2_decap_8
XFILLER_39_911 VPWR VGND sg13g2_decap_8
X_2314_ _0224_ _0200_ _0226_ VPWR VGND sg13g2_xor2_1
X_2245_ _0157_ _1479_ _0056_ VPWR VGND sg13g2_xor2_1
XFILLER_39_988 VPWR VGND sg13g2_decap_8
Xheichips25_template_38 VPWR VGND uio_oe[5] sg13g2_tiehi
X_2176_ net399 net442 net440 net394 _1458_ VPWR VGND sg13g2_and4_1
XFILLER_25_126 VPWR VGND sg13g2_decap_4
XFILLER_41_619 VPWR VGND sg13g2_decap_8
XFILLER_21_365 VPWR VGND sg13g2_decap_8
Xoutput26 net26 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_0_225 VPWR VGND sg13g2_decap_8
XFILLER_1_737 VPWR VGND sg13g2_decap_8
XFILLER_5_1000 VPWR VGND sg13g2_decap_8
XFILLER_29_421 VPWR VGND sg13g2_decap_8
XFILLER_29_454 VPWR VGND sg13g2_fill_2
XFILLER_45_914 VPWR VGND sg13g2_decap_8
XFILLER_17_638 VPWR VGND sg13g2_decap_4
XFILLER_44_479 VPWR VGND sg13g2_decap_4
XFILLER_25_660 VPWR VGND sg13g2_fill_1
XFILLER_13_822 VPWR VGND sg13g2_fill_1
XFILLER_31_129 VPWR VGND sg13g2_fill_1
XFILLER_40_663 VPWR VGND sg13g2_decap_4
XFILLER_13_855 VPWR VGND sg13g2_decap_8
XFILLER_9_837 VPWR VGND sg13g2_decap_8
XFILLER_8_358 VPWR VGND sg13g2_decap_8
XFILLER_12_398 VPWR VGND sg13g2_decap_8
XFILLER_21_81 VPWR VGND sg13g2_decap_8
XFILLER_48_730 VPWR VGND sg13g2_decap_8
X_2030_ _1323_ mac1.sum_lvl3_ff\[12\] mac1.sum_lvl3_ff\[32\] VPWR VGND sg13g2_nand2_1
XFILLER_36_914 VPWR VGND sg13g2_decap_8
XFILLER_35_446 VPWR VGND sg13g2_decap_8
XFILLER_16_693 VPWR VGND sg13g2_decap_8
X_2932_ VGND VPWR net373 _0818_ _0087_ net247 sg13g2_a21oi_1
XFILLER_15_181 VPWR VGND sg13g2_decap_8
X_2863_ net466 net379 _0753_ VPWR VGND sg13g2_nor2_1
X_2794_ _0688_ _0679_ _0687_ VPWR VGND sg13g2_xnor2_1
X_1814_ VGND VPWR _1104_ _1106_ _1141_ _1139_ sg13g2_a21oi_1
XFILLER_7_50 VPWR VGND sg13g2_fill_1
X_1745_ _1038_ _1073_ _1074_ VPWR VGND sg13g2_nor2_1
X_1676_ VGND VPWR _1006_ _1004_ _0959_ sg13g2_or2_1
X_2228_ _1498_ _0139_ _0141_ _0142_ VPWR VGND sg13g2_or3_1
XFILLER_26_15 VPWR VGND sg13g2_fill_2
XFILLER_26_402 VPWR VGND sg13g2_fill_1
XFILLER_27_925 VPWR VGND sg13g2_decap_8
X_2159_ _1433_ VPWR _1441_ VGND _1413_ _1434_ sg13g2_o21ai_1
XFILLER_14_608 VPWR VGND sg13g2_decap_8
XFILLER_41_438 VPWR VGND sg13g2_fill_2
XFILLER_10_803 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_33_clk clknet_3_1__leaf_clk clknet_leaf_33_clk VPWR VGND sg13g2_buf_8
XFILLER_42_36 VPWR VGND sg13g2_decap_8
XFILLER_22_674 VPWR VGND sg13g2_fill_2
XFILLER_22_696 VPWR VGND sg13g2_decap_8
XFILLER_6_818 VPWR VGND sg13g2_decap_8
XFILLER_21_195 VPWR VGND sg13g2_fill_2
XFILLER_5_317 VPWR VGND sg13g2_decap_8
XFILLER_27_1023 VPWR VGND sg13g2_decap_4
XFILLER_49_527 VPWR VGND sg13g2_decap_8
XFILLER_17_402 VPWR VGND sg13g2_decap_4
XFILLER_17_446 VPWR VGND sg13g2_fill_1
XFILLER_18_958 VPWR VGND sg13g2_decap_8
XFILLER_45_777 VPWR VGND sg13g2_decap_4
XFILLER_33_917 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_24_clk clknet_3_5__leaf_clk clknet_leaf_24_clk VPWR VGND sg13g2_buf_8
XFILLER_41_983 VPWR VGND sg13g2_decap_8
XFILLER_40_460 VPWR VGND sg13g2_decap_8
XFILLER_8_100 VPWR VGND sg13g2_decap_4
XFILLER_9_656 VPWR VGND sg13g2_decap_8
X_1530_ _0865_ _0864_ VPWR VGND _0852_ sg13g2_nand2b_2
XFILLER_5_895 VPWR VGND sg13g2_decap_8
X_3200_ net512 VGND VPWR net113 mac1.sum_lvl1_ff\[79\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3131_ net520 VGND VPWR net74 mac1.sum_lvl1_ff\[38\] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_3062_ net539 VGND VPWR _0115_ DP_2.matrix\[5\] clknet_leaf_13_clk sg13g2_dfrbpq_2
X_2013_ _1305_ _1308_ net240 _1310_ VPWR VGND sg13g2_nand3_1
XFILLER_35_232 VPWR VGND sg13g2_decap_8
XFILLER_35_265 VPWR VGND sg13g2_decap_8
XFILLER_17_991 VPWR VGND sg13g2_decap_8
XFILLER_23_427 VPWR VGND sg13g2_decap_8
X_2915_ VGND VPWR _0804_ _0803_ _0801_ sg13g2_or2_1
XFILLER_32_983 VPWR VGND sg13g2_decap_8
X_2846_ net464 net379 _0736_ VPWR VGND sg13g2_nor2_1
XFILLER_12_28 VPWR VGND sg13g2_decap_8
X_2777_ _0670_ _0671_ _0672_ VPWR VGND sg13g2_nor2_1
Xhold100 mac1.products_ff\[0\] VPWR VGND net140 sg13g2_dlygate4sd3_1
Xhold144 DP_2.matrix\[78\] VPWR VGND net184 sg13g2_dlygate4sd3_1
Xhold122 _0000_ VPWR VGND net162 sg13g2_dlygate4sd3_1
XFILLER_2_309 VPWR VGND sg13g2_fill_2
X_1728_ _1057_ _1004_ _1054_ VPWR VGND sg13g2_xnor2_1
Xhold133 _0005_ VPWR VGND net173 sg13g2_dlygate4sd3_1
Xhold111 mac1.products_ff\[10\] VPWR VGND net151 sg13g2_dlygate4sd3_1
Xhold177 mac1.sum_lvl3_ff\[24\] VPWR VGND net217 sg13g2_dlygate4sd3_1
X_1659_ _0077_ _0948_ _0989_ VPWR VGND sg13g2_xnor2_1
Xhold166 mac1.sum_lvl3_ff\[10\] VPWR VGND net206 sg13g2_dlygate4sd3_1
Xhold155 _0086_ VPWR VGND net195 sg13g2_dlygate4sd3_1
Xhold188 _0084_ VPWR VGND net228 sg13g2_dlygate4sd3_1
Xhold199 mac1.sum_lvl3_ff\[27\] VPWR VGND net239 sg13g2_dlygate4sd3_1
XFILLER_39_560 VPWR VGND sg13g2_fill_1
XFILLER_2_1014 VPWR VGND sg13g2_decap_8
XFILLER_27_711 VPWR VGND sg13g2_decap_8
XFILLER_37_69 VPWR VGND sg13g2_fill_2
XFILLER_14_405 VPWR VGND sg13g2_fill_1
XFILLER_15_928 VPWR VGND sg13g2_decap_8
XFILLER_14_427 VPWR VGND sg13g2_decap_8
XFILLER_41_246 VPWR VGND sg13g2_fill_1
XFILLER_23_961 VPWR VGND sg13g2_decap_8
XFILLER_2_832 VPWR VGND sg13g2_decap_8
XFILLER_49_368 VPWR VGND sg13g2_decap_8
XFILLER_18_700 VPWR VGND sg13g2_decap_8
XFILLER_18_733 VPWR VGND sg13g2_decap_8
XFILLER_45_552 VPWR VGND sg13g2_fill_2
XFILLER_45_541 VPWR VGND sg13g2_decap_8
XFILLER_27_91 VPWR VGND sg13g2_decap_8
XFILLER_14_961 VPWR VGND sg13g2_decap_8
X_2700_ _0597_ net428 net479 net430 net476 VPWR VGND sg13g2_a22oi_1
X_2631_ _0455_ _0527_ _0529_ _0530_ VPWR VGND sg13g2_or3_1
X_2562_ _0422_ _0460_ _0462_ VPWR VGND sg13g2_and2_1
XFILLER_5_692 VPWR VGND sg13g2_decap_8
X_1513_ _0848_ _0849_ _0850_ VPWR VGND sg13g2_nor2b_1
X_2493_ net439 net485 net481 net436 _0395_ VPWR VGND sg13g2_and4_1
XFILLER_4_73 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_4_clk clknet_3_3__leaf_clk clknet_leaf_4_clk VPWR VGND sg13g2_buf_8
X_3114_ net520 VGND VPWR net123 mac1.sum_lvl1_ff\[1\] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_3045_ net543 VGND VPWR _0098_ DP_1.matrix\[40\] clknet_leaf_24_clk sg13g2_dfrbpq_2
XFILLER_48_390 VPWR VGND sg13g2_fill_1
XFILLER_23_202 VPWR VGND sg13g2_decap_8
XFILLER_24_714 VPWR VGND sg13g2_fill_2
XFILLER_24_769 VPWR VGND sg13g2_decap_8
XFILLER_20_953 VPWR VGND sg13g2_decap_8
X_2829_ _0710_ VPWR _0721_ VGND _0681_ _0708_ sg13g2_o21ai_1
Xfanout421 net423 net421 VPWR VGND sg13g2_buf_8
Xfanout432 DP_2.matrix\[2\] net432 VPWR VGND sg13g2_buf_1
Xfanout410 net197 net410 VPWR VGND sg13g2_buf_8
XFILLER_48_35 VPWR VGND sg13g2_decap_8
Xfanout443 DP_1.matrix\[78\] net443 VPWR VGND sg13g2_buf_8
Xfanout454 net456 net454 VPWR VGND sg13g2_buf_8
Xfanout465 DP_1.matrix\[41\] net465 VPWR VGND sg13g2_buf_8
Xfanout476 net478 net476 VPWR VGND sg13g2_buf_8
XFILLER_19_519 VPWR VGND sg13g2_fill_1
Xfanout498 net499 net498 VPWR VGND sg13g2_buf_8
Xfanout487 DP_1.matrix\[3\] net487 VPWR VGND sg13g2_buf_8
XFILLER_46_349 VPWR VGND sg13g2_fill_2
XFILLER_42_522 VPWR VGND sg13g2_fill_2
XFILLER_42_544 VPWR VGND sg13g2_decap_8
XFILLER_14_235 VPWR VGND sg13g2_decap_8
XFILLER_14_246 VPWR VGND sg13g2_fill_2
XFILLER_42_566 VPWR VGND sg13g2_fill_1
XFILLER_14_257 VPWR VGND sg13g2_decap_8
XFILLER_30_717 VPWR VGND sg13g2_decap_8
XFILLER_23_791 VPWR VGND sg13g2_decap_8
XFILLER_10_441 VPWR VGND sg13g2_decap_8
XFILLER_7_924 VPWR VGND sg13g2_decap_8
XFILLER_11_975 VPWR VGND sg13g2_decap_8
XFILLER_6_423 VPWR VGND sg13g2_decap_8
XFILLER_13_82 VPWR VGND sg13g2_fill_2
XFILLER_6_489 VPWR VGND sg13g2_decap_8
XFILLER_36_8 VPWR VGND sg13g2_decap_8
XFILLER_1_183 VPWR VGND sg13g2_fill_1
XFILLER_49_165 VPWR VGND sg13g2_decap_8
Xclkbuf_3_7__f_clk clknet_0_clk clknet_3_7__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_46_883 VPWR VGND sg13g2_decap_8
XFILLER_45_382 VPWR VGND sg13g2_decap_8
XFILLER_21_717 VPWR VGND sg13g2_decap_8
X_1993_ net217 mac1.sum_lvl3_ff\[4\] _1294_ VPWR VGND sg13g2_xor2_1
XFILLER_20_216 VPWR VGND sg13g2_decap_8
X_2614_ net477 net500 net438 _0513_ VPWR VGND net434 sg13g2_nand4_1
XFILLER_47_1004 VPWR VGND sg13g2_decap_8
X_2545_ _0413_ _0444_ _0445_ _0446_ VPWR VGND sg13g2_nor3_1
X_2476_ _0376_ _0375_ _0370_ _0379_ VPWR VGND sg13g2_a21o_1
XFILLER_37_861 VPWR VGND sg13g2_decap_8
X_3028_ net531 VGND VPWR _0081_ DP_1.matrix\[8\] clknet_leaf_12_clk sg13g2_dfrbpq_2
XFILLER_24_544 VPWR VGND sg13g2_decap_4
XFILLER_12_728 VPWR VGND sg13g2_decap_8
Xclkload3 clkload3/Y clknet_leaf_38_clk VPWR VGND sg13g2_inv_2
XFILLER_20_750 VPWR VGND sg13g2_decap_8
XFILLER_4_938 VPWR VGND sg13g2_decap_8
XFILLER_3_426 VPWR VGND sg13g2_decap_4
XFILLER_3_448 VPWR VGND sg13g2_fill_2
XFILLER_47_614 VPWR VGND sg13g2_decap_8
XFILLER_47_603 VPWR VGND sg13g2_decap_4
XFILLER_47_647 VPWR VGND sg13g2_decap_4
XFILLER_47_625 VPWR VGND sg13g2_fill_1
XFILLER_27_360 VPWR VGND sg13g2_fill_1
XFILLER_15_522 VPWR VGND sg13g2_decap_8
XFILLER_42_352 VPWR VGND sg13g2_fill_1
XFILLER_15_566 VPWR VGND sg13g2_fill_2
XFILLER_24_70 VPWR VGND sg13g2_decap_8
XFILLER_7_721 VPWR VGND sg13g2_decap_8
XFILLER_7_798 VPWR VGND sg13g2_decap_8
X_2330_ _0241_ _0215_ _0239_ VPWR VGND sg13g2_xnor2_1
XFILLER_2_481 VPWR VGND sg13g2_decap_4
X_2261_ _0140_ VPWR _0174_ VGND _1498_ _0141_ sg13g2_o21ai_1
XFILLER_38_603 VPWR VGND sg13g2_decap_8
X_2192_ VGND VPWR _1471_ _1472_ _1474_ _1441_ sg13g2_a21oi_1
XFILLER_38_636 VPWR VGND sg13g2_decap_8
XFILLER_38_647 VPWR VGND sg13g2_fill_1
XFILLER_37_157 VPWR VGND sg13g2_decap_4
XFILLER_19_894 VPWR VGND sg13g2_decap_8
XFILLER_25_308 VPWR VGND sg13g2_decap_8
XFILLER_37_179 VPWR VGND sg13g2_decap_8
XFILLER_45_190 VPWR VGND sg13g2_decap_8
XFILLER_33_363 VPWR VGND sg13g2_decap_8
XFILLER_14_1003 VPWR VGND sg13g2_decap_8
X_1976_ _0006_ _1280_ net169 VPWR VGND sg13g2_xnor2_1
XFILLER_20_39 VPWR VGND sg13g2_decap_8
XFILLER_1_919 VPWR VGND sg13g2_decap_8
X_2528_ net438 net481 net480 net435 _0429_ VPWR VGND sg13g2_and4_1
XFILLER_29_15 VPWR VGND sg13g2_decap_8
Xhold15 mac1.sum_lvl1_ff\[40\] VPWR VGND net55 sg13g2_dlygate4sd3_1
Xhold37 mac1.sum_lvl1_ff\[45\] VPWR VGND net77 sg13g2_dlygate4sd3_1
Xhold26 mac1.products_ff\[146\] VPWR VGND net66 sg13g2_dlygate4sd3_1
X_2459_ _0363_ _0352_ _0362_ VPWR VGND sg13g2_xnor2_1
Xhold59 mac1.sum_lvl1_ff\[13\] VPWR VGND net99 sg13g2_dlygate4sd3_1
Xhold48 mac1.products_ff\[145\] VPWR VGND net88 sg13g2_dlygate4sd3_1
XFILLER_28_146 VPWR VGND sg13g2_decap_8
XFILLER_45_58 VPWR VGND sg13g2_fill_2
XFILLER_8_518 VPWR VGND sg13g2_decap_8
XFILLER_12_558 VPWR VGND sg13g2_decap_8
XFILLER_4_735 VPWR VGND sg13g2_decap_8
XFILLER_3_245 VPWR VGND sg13g2_decap_4
XFILLER_10_72 VPWR VGND sg13g2_fill_1
XFILLER_0_930 VPWR VGND sg13g2_decap_8
XFILLER_48_912 VPWR VGND sg13g2_decap_8
XFILLER_48_989 VPWR VGND sg13g2_decap_8
XFILLER_47_444 VPWR VGND sg13g2_decap_8
XFILLER_19_81 VPWR VGND sg13g2_decap_8
XFILLER_19_157 VPWR VGND sg13g2_decap_8
XFILLER_35_606 VPWR VGND sg13g2_decap_8
XFILLER_34_138 VPWR VGND sg13g2_decap_8
XFILLER_27_190 VPWR VGND sg13g2_decap_8
XFILLER_43_694 VPWR VGND sg13g2_fill_1
XFILLER_16_897 VPWR VGND sg13g2_decap_8
XFILLER_31_823 VPWR VGND sg13g2_decap_4
X_1830_ _1156_ net401 net465 net403 net462 VPWR VGND sg13g2_a22oi_1
XFILLER_30_344 VPWR VGND sg13g2_decap_8
X_1761_ _1088_ _1080_ _1089_ VPWR VGND sg13g2_nor2b_1
X_1692_ _1019_ _1020_ _1002_ _1022_ VPWR VGND sg13g2_nand3_1
XFILLER_7_595 VPWR VGND sg13g2_fill_1
X_2313_ _0225_ _0200_ _0224_ VPWR VGND sg13g2_nand2_1
X_2244_ _1477_ _1478_ _0155_ _0156_ _0158_ VPWR VGND sg13g2_and4_1
XFILLER_39_967 VPWR VGND sg13g2_decap_8
Xheichips25_template_39 VPWR VGND uio_oe[6] sg13g2_tiehi
X_2175_ _1457_ net444 net391 VPWR VGND sg13g2_nand2_1
XFILLER_25_116 VPWR VGND sg13g2_decap_4
XFILLER_15_39 VPWR VGND sg13g2_decap_8
XFILLER_40_119 VPWR VGND sg13g2_decap_8
XFILLER_33_182 VPWR VGND sg13g2_decap_8
XFILLER_22_889 VPWR VGND sg13g2_decap_8
X_1959_ _1263_ VPWR _1268_ VGND _1259_ _1262_ sg13g2_o21ai_1
Xoutput27 net27 uo_out[2] VPWR VGND sg13g2_buf_1
XFILLER_1_716 VPWR VGND sg13g2_decap_8
XFILLER_0_204 VPWR VGND sg13g2_decap_8
XFILLER_29_400 VPWR VGND sg13g2_decap_8
XFILLER_17_617 VPWR VGND sg13g2_decap_8
XFILLER_29_466 VPWR VGND sg13g2_decap_8
XFILLER_40_620 VPWR VGND sg13g2_fill_2
XFILLER_13_834 VPWR VGND sg13g2_decap_8
XFILLER_40_642 VPWR VGND sg13g2_fill_1
XFILLER_9_816 VPWR VGND sg13g2_decap_8
XFILLER_12_344 VPWR VGND sg13g2_decap_8
XFILLER_21_60 VPWR VGND sg13g2_decap_8
XFILLER_47_230 VPWR VGND sg13g2_decap_8
XFILLER_48_786 VPWR VGND sg13g2_decap_8
XFILLER_47_241 VPWR VGND sg13g2_fill_1
XFILLER_35_414 VPWR VGND sg13g2_fill_2
XFILLER_35_425 VPWR VGND sg13g2_decap_8
XFILLER_16_661 VPWR VGND sg13g2_fill_2
XFILLER_35_469 VPWR VGND sg13g2_fill_1
XFILLER_44_992 VPWR VGND sg13g2_decap_8
XFILLER_15_160 VPWR VGND sg13g2_fill_1
X_2931_ _0746_ _0742_ _0818_ VPWR VGND sg13g2_xor2_1
XFILLER_43_491 VPWR VGND sg13g2_fill_2
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
XFILLER_31_642 VPWR VGND sg13g2_fill_1
XFILLER_31_653 VPWR VGND sg13g2_fill_2
XFILLER_31_675 VPWR VGND sg13g2_fill_2
X_2862_ _0752_ net449 _0732_ VPWR VGND sg13g2_nand2_1
X_2793_ _0687_ _0650_ _0685_ VPWR VGND sg13g2_xnor2_1
X_1813_ _1106_ _1139_ _1104_ _1140_ VPWR VGND sg13g2_nand3_1
XFILLER_30_196 VPWR VGND sg13g2_decap_4
XFILLER_11_1017 VPWR VGND sg13g2_decap_8
XFILLER_11_1028 VPWR VGND sg13g2_fill_1
X_1744_ _1073_ _1039_ _1071_ VPWR VGND sg13g2_xnor2_1
XFILLER_8_893 VPWR VGND sg13g2_decap_8
X_1675_ _1005_ net409 net465 VPWR VGND sg13g2_nand2_1
X_2227_ VGND VPWR _0137_ _0138_ _0141_ _1499_ sg13g2_a21oi_1
XFILLER_39_786 VPWR VGND sg13g2_decap_4
XFILLER_27_904 VPWR VGND sg13g2_decap_8
X_2158_ _1440_ _1439_ _0054_ VPWR VGND sg13g2_xor2_1
XFILLER_26_414 VPWR VGND sg13g2_decap_8
X_2089_ VGND VPWR _1371_ _1372_ _1374_ _1366_ sg13g2_a21oi_1
XFILLER_26_49 VPWR VGND sg13g2_decap_8
XFILLER_41_417 VPWR VGND sg13g2_decap_8
XFILLER_35_992 VPWR VGND sg13g2_decap_8
XFILLER_21_152 VPWR VGND sg13g2_decap_8
XFILLER_10_859 VPWR VGND sg13g2_decap_8
XFILLER_21_174 VPWR VGND sg13g2_decap_4
XFILLER_27_1002 VPWR VGND sg13g2_decap_8
XFILLER_49_506 VPWR VGND sg13g2_decap_8
XFILLER_18_937 VPWR VGND sg13g2_decap_8
XFILLER_29_241 VPWR VGND sg13g2_fill_2
XFILLER_32_406 VPWR VGND sg13g2_fill_1
XFILLER_32_417 VPWR VGND sg13g2_decap_8
XFILLER_32_439 VPWR VGND sg13g2_fill_2
XFILLER_41_962 VPWR VGND sg13g2_decap_8
XFILLER_13_620 VPWR VGND sg13g2_decap_8
XFILLER_34_1017 VPWR VGND sg13g2_decap_8
XFILLER_34_1028 VPWR VGND sg13g2_fill_1
XFILLER_8_156 VPWR VGND sg13g2_decap_8
XFILLER_5_874 VPWR VGND sg13g2_decap_8
XFILLER_4_373 VPWR VGND sg13g2_fill_1
XFILLER_4_362 VPWR VGND sg13g2_decap_8
X_3130_ net520 VGND VPWR net143 mac1.sum_lvl1_ff\[37\] clknet_leaf_33_clk sg13g2_dfrbpq_1
X_3061_ net538 VGND VPWR _0114_ DP_2.matrix\[4\] clknet_3_6__leaf_clk sg13g2_dfrbpq_1
X_2012_ VGND VPWR net240 _1305_ _1309_ _1308_ sg13g2_a21oi_1
XFILLER_35_211 VPWR VGND sg13g2_decap_8
XFILLER_24_929 VPWR VGND sg13g2_decap_8
XFILLER_17_970 VPWR VGND sg13g2_decap_8
XFILLER_23_406 VPWR VGND sg13g2_decap_8
X_2914_ _0803_ net377 _0802_ _0783_ net387 VPWR VGND sg13g2_a22oi_1
XFILLER_31_450 VPWR VGND sg13g2_decap_8
XFILLER_31_461 VPWR VGND sg13g2_fill_2
XFILLER_32_962 VPWR VGND sg13g2_decap_8
X_2845_ VPWR _0735_ _0734_ VGND sg13g2_inv_1
X_2776_ VGND VPWR _0618_ _0638_ _0671_ _0640_ sg13g2_a21oi_1
XFILLER_8_690 VPWR VGND sg13g2_decap_8
Xhold101 mac1.sum_lvl2_ff\[41\] VPWR VGND net141 sg13g2_dlygate4sd3_1
Xhold134 mac1.sum_lvl3_ff\[22\] VPWR VGND net174 sg13g2_dlygate4sd3_1
X_1727_ _1004_ _1054_ _1056_ VPWR VGND sg13g2_and2_1
Xhold123 mac1.sum_lvl3_ff\[35\] VPWR VGND net163 sg13g2_dlygate4sd3_1
Xhold112 mac1.products_ff\[9\] VPWR VGND net152 sg13g2_dlygate4sd3_1
Xhold145 DP_2.matrix\[79\] VPWR VGND net185 sg13g2_dlygate4sd3_1
X_1658_ _0986_ _0988_ _0989_ VPWR VGND sg13g2_nor2_1
Xhold167 _1316_ VPWR VGND net207 sg13g2_dlygate4sd3_1
Xhold156 DP_1.matrix\[36\] VPWR VGND net196 sg13g2_dlygate4sd3_1
Xhold189 DP_2.matrix\[3\] VPWR VGND net229 sg13g2_dlygate4sd3_1
Xhold178 _1294_ VPWR VGND net218 sg13g2_dlygate4sd3_1
X_1589_ _0903_ VPWR _0921_ VGND _0894_ _0904_ sg13g2_o21ai_1
XFILLER_46_509 VPWR VGND sg13g2_decap_8
X_3259_ net514 VGND VPWR net7 DP_1.Q_range.out_data\[4\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_27_701 VPWR VGND sg13g2_fill_2
XFILLER_26_211 VPWR VGND sg13g2_decap_4
XFILLER_15_907 VPWR VGND sg13g2_decap_8
XFILLER_26_244 VPWR VGND sg13g2_decap_8
XFILLER_42_726 VPWR VGND sg13g2_decap_8
XFILLER_23_940 VPWR VGND sg13g2_decap_8
XFILLER_2_811 VPWR VGND sg13g2_decap_8
XFILLER_2_888 VPWR VGND sg13g2_decap_8
XFILLER_49_347 VPWR VGND sg13g2_decap_8
XFILLER_45_564 VPWR VGND sg13g2_decap_8
XFILLER_17_222 VPWR VGND sg13g2_decap_4
XFILLER_18_778 VPWR VGND sg13g2_decap_8
XFILLER_45_575 VPWR VGND sg13g2_decap_8
XFILLER_17_266 VPWR VGND sg13g2_fill_2
XFILLER_32_203 VPWR VGND sg13g2_decap_4
XFILLER_14_940 VPWR VGND sg13g2_decap_8
XFILLER_33_759 VPWR VGND sg13g2_decap_8
X_2630_ VGND VPWR _0525_ _0526_ _0529_ _0491_ sg13g2_a21oi_1
X_2561_ VGND VPWR _0461_ _0459_ _0423_ sg13g2_or2_1
XFILLER_5_671 VPWR VGND sg13g2_decap_8
X_1512_ _0843_ VPWR _0849_ VGND _0846_ _0847_ sg13g2_o21ai_1
X_2492_ _0394_ net487 net431 VPWR VGND sg13g2_nand2_1
XFILLER_4_192 VPWR VGND sg13g2_fill_2
X_3113_ net521 VGND VPWR net140 mac1.sum_lvl1_ff\[0\] clknet_leaf_33_clk sg13g2_dfrbpq_1
XFILLER_49_881 VPWR VGND sg13g2_decap_8
X_3044_ net535 VGND VPWR _0097_ DP_1.matrix\[39\] clknet_leaf_22_clk sg13g2_dfrbpq_2
XFILLER_11_409 VPWR VGND sg13g2_decap_4
XFILLER_17_1012 VPWR VGND sg13g2_decap_8
XFILLER_20_932 VPWR VGND sg13g2_decap_8
XFILLER_23_39 VPWR VGND sg13g2_decap_8
X_2828_ VGND VPWR _0689_ _0713_ _0720_ _0715_ sg13g2_a21oi_1
X_2759_ _0654_ net484 net495 VPWR VGND sg13g2_nand2_1
XFILLER_3_619 VPWR VGND sg13g2_decap_8
Xfanout422 net423 net422 VPWR VGND sg13g2_buf_1
XFILLER_48_14 VPWR VGND sg13g2_decap_8
Xfanout411 DP_2.matrix\[38\] net411 VPWR VGND sg13g2_buf_1
Xfanout400 net290 net400 VPWR VGND sg13g2_buf_1
Xfanout466 DP_1.matrix\[40\] net466 VPWR VGND sg13g2_buf_8
Xfanout455 net456 net455 VPWR VGND sg13g2_buf_1
XFILLER_24_1027 VPWR VGND sg13g2_fill_2
Xfanout444 net445 net444 VPWR VGND sg13g2_buf_8
Xfanout433 net221 net433 VPWR VGND sg13g2_buf_8
XFILLER_47_829 VPWR VGND sg13g2_decap_8
Xfanout477 net478 net477 VPWR VGND sg13g2_buf_8
Xfanout499 net189 net499 VPWR VGND sg13g2_buf_8
Xfanout488 net249 net488 VPWR VGND sg13g2_buf_8
XFILLER_42_589 VPWR VGND sg13g2_decap_8
XFILLER_23_770 VPWR VGND sg13g2_decap_8
XFILLER_7_903 VPWR VGND sg13g2_decap_8
XFILLER_6_402 VPWR VGND sg13g2_decap_8
XFILLER_11_954 VPWR VGND sg13g2_decap_8
XFILLER_2_685 VPWR VGND sg13g2_decap_8
XFILLER_49_144 VPWR VGND sg13g2_decap_8
XFILLER_38_807 VPWR VGND sg13g2_fill_2
XFILLER_38_80 VPWR VGND sg13g2_decap_8
XFILLER_37_317 VPWR VGND sg13g2_fill_2
XFILLER_46_862 VPWR VGND sg13g2_decap_8
XFILLER_18_531 VPWR VGND sg13g2_decap_8
XFILLER_38_91 VPWR VGND sg13g2_fill_1
XFILLER_18_564 VPWR VGND sg13g2_decap_8
XFILLER_33_534 VPWR VGND sg13g2_decap_8
XFILLER_33_545 VPWR VGND sg13g2_fill_2
X_1992_ mac1.sum_lvl3_ff\[4\] net217 _1293_ VPWR VGND sg13g2_and2_1
XFILLER_14_781 VPWR VGND sg13g2_decap_4
Xclkload10 clknet_leaf_29_clk clkload10/Y VPWR VGND sg13g2_inv_4
X_2613_ net438 net477 net500 net434 _0512_ VPWR VGND sg13g2_and4_1
X_2544_ VGND VPWR _0442_ _0443_ _0445_ _0414_ sg13g2_a21oi_1
XFILLER_48_0 VPWR VGND sg13g2_decap_8
X_2475_ VGND VPWR _0375_ _0376_ _0378_ _0370_ sg13g2_a21oi_1
X_3027_ net538 VGND VPWR _0080_ DP_2.matrix\[80\] clknet_leaf_12_clk sg13g2_dfrbpq_2
XFILLER_36_394 VPWR VGND sg13g2_decap_4
XFILLER_34_38 VPWR VGND sg13g2_fill_2
XFILLER_11_217 VPWR VGND sg13g2_decap_8
XFILLER_24_589 VPWR VGND sg13g2_decap_4
Xclkload4 clkload4/Y clknet_leaf_2_clk VPWR VGND sg13g2_inv_8
XFILLER_4_917 VPWR VGND sg13g2_decap_8
XFILLER_3_405 VPWR VGND sg13g2_decap_8
XFILLER_19_317 VPWR VGND sg13g2_decap_8
XFILLER_19_339 VPWR VGND sg13g2_fill_1
XFILLER_28_895 VPWR VGND sg13g2_decap_8
XFILLER_43_887 VPWR VGND sg13g2_decap_8
XFILLER_15_589 VPWR VGND sg13g2_fill_1
XFILLER_7_700 VPWR VGND sg13g2_decap_8
XFILLER_6_210 VPWR VGND sg13g2_fill_2
XFILLER_7_777 VPWR VGND sg13g2_decap_8
XFILLER_6_221 VPWR VGND sg13g2_decap_8
XFILLER_3_983 VPWR VGND sg13g2_decap_8
X_2260_ _0173_ _0163_ _0171_ VPWR VGND sg13g2_xnor2_1
X_2191_ _1471_ _1472_ _1441_ _1473_ VPWR VGND sg13g2_nand3_1
XFILLER_38_626 VPWR VGND sg13g2_decap_4
XFILLER_19_873 VPWR VGND sg13g2_decap_8
XFILLER_46_692 VPWR VGND sg13g2_decap_8
XFILLER_21_504 VPWR VGND sg13g2_fill_2
XFILLER_34_898 VPWR VGND sg13g2_decap_8
X_1975_ _1281_ net168 mac1.sum_lvl2_ff\[15\] VPWR VGND sg13g2_xnor2_1
XFILLER_20_18 VPWR VGND sg13g2_decap_8
XFILLER_0_419 VPWR VGND sg13g2_decap_8
X_2527_ _0428_ net484 net431 VPWR VGND sg13g2_nand2_1
X_2458_ _0362_ _0353_ _0360_ VPWR VGND sg13g2_xnor2_1
Xhold16 mac1.sum_lvl1_ff\[72\] VPWR VGND net56 sg13g2_dlygate4sd3_1
Xhold38 mac1.sum_lvl1_ff\[81\] VPWR VGND net78 sg13g2_dlygate4sd3_1
Xhold27 mac1.products_ff\[79\] VPWR VGND net67 sg13g2_dlygate4sd3_1
XFILLER_29_27 VPWR VGND sg13g2_decap_8
XFILLER_29_38 VPWR VGND sg13g2_fill_2
X_2389_ _0298_ DP_1.matrix\[79\] net383 VPWR VGND sg13g2_nand2_1
Xhold49 mac1.sum_lvl2_ff\[39\] VPWR VGND net89 sg13g2_dlygate4sd3_1
XFILLER_21_1008 VPWR VGND sg13g2_decap_8
XFILLER_44_618 VPWR VGND sg13g2_decap_8
XFILLER_43_106 VPWR VGND sg13g2_decap_8
XFILLER_43_117 VPWR VGND sg13g2_fill_1
XFILLER_37_681 VPWR VGND sg13g2_decap_8
XFILLER_37_692 VPWR VGND sg13g2_fill_2
XFILLER_24_353 VPWR VGND sg13g2_fill_1
XFILLER_12_504 VPWR VGND sg13g2_fill_2
XFILLER_4_714 VPWR VGND sg13g2_decap_8
XFILLER_3_224 VPWR VGND sg13g2_decap_8
XFILLER_10_40 VPWR VGND sg13g2_decap_8
XFILLER_47_423 VPWR VGND sg13g2_decap_8
XFILLER_0_986 VPWR VGND sg13g2_decap_8
XFILLER_48_968 VPWR VGND sg13g2_decap_8
XFILLER_16_810 VPWR VGND sg13g2_decap_8
XFILLER_28_670 VPWR VGND sg13g2_decap_4
XFILLER_43_662 VPWR VGND sg13g2_decap_8
XFILLER_43_640 VPWR VGND sg13g2_decap_8
XFILLER_15_353 VPWR VGND sg13g2_fill_2
XFILLER_16_876 VPWR VGND sg13g2_decap_8
XFILLER_31_802 VPWR VGND sg13g2_decap_8
XFILLER_37_1015 VPWR VGND sg13g2_decap_8
XFILLER_42_161 VPWR VGND sg13g2_decap_8
XFILLER_15_397 VPWR VGND sg13g2_decap_8
X_1760_ _1088_ _1081_ _1087_ VPWR VGND sg13g2_xnor2_1
X_1691_ _1021_ _1002_ _1019_ _1020_ VPWR VGND sg13g2_and3_1
XFILLER_3_780 VPWR VGND sg13g2_decap_8
X_2312_ _0223_ _0211_ _0224_ VPWR VGND sg13g2_xor2_1
XFILLER_39_946 VPWR VGND sg13g2_decap_8
X_2243_ _0157_ _0155_ _0156_ VPWR VGND sg13g2_nand2_1
XFILLER_38_412 VPWR VGND sg13g2_fill_2
X_2174_ _1424_ VPWR _1456_ VGND _1422_ _1425_ sg13g2_o21ai_1
XFILLER_38_489 VPWR VGND sg13g2_decap_8
XFILLER_47_990 VPWR VGND sg13g2_decap_8
XFILLER_18_180 VPWR VGND sg13g2_decap_4
XFILLER_40_109 VPWR VGND sg13g2_fill_1
XFILLER_34_673 VPWR VGND sg13g2_decap_8
XFILLER_21_334 VPWR VGND sg13g2_decap_4
X_1958_ mac1.sum_lvl2_ff\[12\] mac1.sum_lvl2_ff\[31\] _1267_ VPWR VGND sg13g2_xor2_1
X_1889_ _1212_ _1202_ _1213_ VPWR VGND sg13g2_nor2b_1
Xoutput17 net17 uio_out[0] VPWR VGND sg13g2_buf_1
Xoutput28 net28 uo_out[3] VPWR VGND sg13g2_buf_1
XFILLER_0_249 VPWR VGND sg13g2_decap_8
XFILLER_48_209 VPWR VGND sg13g2_decap_8
XFILLER_29_456 VPWR VGND sg13g2_fill_1
XFILLER_45_949 VPWR VGND sg13g2_decap_8
XFILLER_16_128 VPWR VGND sg13g2_decap_8
XFILLER_12_323 VPWR VGND sg13g2_decap_8
XFILLER_8_305 VPWR VGND sg13g2_decap_8
XFILLER_12_378 VPWR VGND sg13g2_decap_8
XFILLER_0_783 VPWR VGND sg13g2_decap_8
XFILLER_47_220 VPWR VGND sg13g2_fill_1
XFILLER_48_765 VPWR VGND sg13g2_decap_8
XFILLER_47_253 VPWR VGND sg13g2_decap_8
XFILLER_47_297 VPWR VGND sg13g2_decap_4
XFILLER_29_990 VPWR VGND sg13g2_decap_8
XFILLER_36_949 VPWR VGND sg13g2_decap_8
XFILLER_44_971 VPWR VGND sg13g2_decap_8
XFILLER_22_109 VPWR VGND sg13g2_decap_4
X_2930_ net490 net373 _0817_ VPWR VGND sg13g2_nor2_1
XFILLER_30_142 VPWR VGND sg13g2_decap_8
X_2861_ _0751_ _0750_ _0740_ VPWR VGND sg13g2_nand2b_1
X_2792_ _0650_ _0685_ _0686_ VPWR VGND sg13g2_nor2b_1
XFILLER_7_30 VPWR VGND sg13g2_decap_4
X_1812_ _1137_ _1115_ _1139_ VPWR VGND sg13g2_xor2_1
XFILLER_30_175 VPWR VGND sg13g2_decap_8
XFILLER_31_698 VPWR VGND sg13g2_fill_1
XFILLER_8_872 VPWR VGND sg13g2_decap_8
X_1743_ _1072_ _1039_ _1071_ VPWR VGND sg13g2_nand2b_1
X_1674_ _1004_ net407 net465 VPWR VGND sg13g2_nand2_2
X_2226_ _0137_ _0138_ _1499_ _0140_ VPWR VGND sg13g2_nand3_1
XFILLER_38_220 VPWR VGND sg13g2_decap_8
XFILLER_39_765 VPWR VGND sg13g2_decap_8
XFILLER_38_242 VPWR VGND sg13g2_decap_8
X_2157_ _1406_ VPWR _1440_ VGND _1381_ _1407_ sg13g2_o21ai_1
XFILLER_26_28 VPWR VGND sg13g2_decap_8
X_2088_ _1371_ _1372_ _1366_ _1373_ VPWR VGND sg13g2_nand3_1
XFILLER_35_971 VPWR VGND sg13g2_decap_8
XFILLER_22_665 VPWR VGND sg13g2_fill_2
XFILLER_10_838 VPWR VGND sg13g2_decap_8
XFILLER_1_569 VPWR VGND sg13g2_decap_8
XFILLER_18_916 VPWR VGND sg13g2_decap_8
XFILLER_45_746 VPWR VGND sg13g2_decap_4
XFILLER_17_426 VPWR VGND sg13g2_decap_4
XFILLER_16_50 VPWR VGND sg13g2_decap_4
XFILLER_26_993 VPWR VGND sg13g2_decap_8
XFILLER_41_941 VPWR VGND sg13g2_decap_8
XFILLER_12_153 VPWR VGND sg13g2_decap_8
XFILLER_40_484 VPWR VGND sg13g2_decap_4
XFILLER_12_164 VPWR VGND sg13g2_fill_1
XFILLER_32_60 VPWR VGND sg13g2_decap_8
XFILLER_5_853 VPWR VGND sg13g2_decap_8
XFILLER_4_341 VPWR VGND sg13g2_decap_8
X_3060_ net538 VGND VPWR net230 DP_2.matrix\[3\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_0_580 VPWR VGND sg13g2_decap_8
X_2011_ _1308_ mac1.sum_lvl3_ff\[8\] mac1.sum_lvl3_ff\[28\] VPWR VGND sg13g2_xnor2_1
XFILLER_24_908 VPWR VGND sg13g2_decap_8
XFILLER_32_941 VPWR VGND sg13g2_decap_8
X_2913_ net406 net427 _0781_ _0802_ VPWR VGND sg13g2_mux2_1
X_2844_ _0734_ _0728_ _0729_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_495 VPWR VGND sg13g2_decap_8
X_2775_ _0668_ _0647_ _0670_ VPWR VGND sg13g2_xor2_1
Xhold113 mac1.sum_lvl3_ff\[20\] VPWR VGND net153 sg13g2_dlygate4sd3_1
Xhold135 _1288_ VPWR VGND net175 sg13g2_dlygate4sd3_1
Xhold102 mac1.sum_lvl2_ff\[51\] VPWR VGND net142 sg13g2_dlygate4sd3_1
X_1726_ VGND VPWR _1055_ _1054_ _1004_ sg13g2_or2_1
Xhold124 _1338_ VPWR VGND net164 sg13g2_dlygate4sd3_1
X_1657_ VGND VPWR _0984_ _0985_ _0988_ _0945_ sg13g2_a21oi_1
Xhold168 _1322_ VPWR VGND net208 sg13g2_dlygate4sd3_1
Xhold157 DP_2.matrix\[38\] VPWR VGND net197 sg13g2_dlygate4sd3_1
Xhold146 mac1.sum_lvl3_ff\[34\] VPWR VGND net186 sg13g2_dlygate4sd3_1
Xhold179 _0026_ VPWR VGND net219 sg13g2_dlygate4sd3_1
X_1588_ VPWR _0920_ _0919_ VGND sg13g2_inv_1
X_3258_ net514 VGND VPWR net6 DP_1.Q_range.out_data\[3\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_39_551 VPWR VGND sg13g2_decap_8
X_2209_ _1490_ _1481_ _1488_ VPWR VGND sg13g2_xnor2_1
X_3189_ net523 VGND VPWR net132 mac1.sum_lvl2_ff\[50\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_27_735 VPWR VGND sg13g2_decap_4
XFILLER_27_779 VPWR VGND sg13g2_decap_8
XFILLER_41_215 VPWR VGND sg13g2_decap_8
XFILLER_41_237 VPWR VGND sg13g2_decap_8
XFILLER_22_451 VPWR VGND sg13g2_fill_2
XFILLER_10_624 VPWR VGND sg13g2_decap_8
XFILLER_23_996 VPWR VGND sg13g2_decap_8
XFILLER_6_617 VPWR VGND sg13g2_fill_2
XFILLER_2_867 VPWR VGND sg13g2_decap_8
XFILLER_1_355 VPWR VGND sg13g2_decap_8
XFILLER_49_326 VPWR VGND sg13g2_fill_1
XFILLER_17_212 VPWR VGND sg13g2_fill_1
XFILLER_27_71 VPWR VGND sg13g2_fill_2
XFILLER_33_705 VPWR VGND sg13g2_fill_2
XFILLER_26_790 VPWR VGND sg13g2_decap_8
XFILLER_32_215 VPWR VGND sg13g2_decap_8
XFILLER_32_248 VPWR VGND sg13g2_fill_2
XFILLER_13_451 VPWR VGND sg13g2_decap_8
XFILLER_14_996 VPWR VGND sg13g2_decap_8
XFILLER_9_466 VPWR VGND sg13g2_fill_2
XFILLER_9_488 VPWR VGND sg13g2_decap_8
XFILLER_5_650 VPWR VGND sg13g2_decap_8
X_2560_ _0460_ net485 net429 VPWR VGND sg13g2_nand2_1
X_1511_ _0843_ _0846_ _0847_ _0848_ VPWR VGND sg13g2_nor3_1
X_2491_ _0373_ VPWR _0393_ VGND _0371_ _0374_ sg13g2_o21ai_1
XFILLER_49_860 VPWR VGND sg13g2_decap_8
X_3112_ net529 VGND VPWR _0053_ mac1.products_ff\[151\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_3043_ net527 VGND VPWR _0096_ DP_1.matrix\[38\] clknet_leaf_22_clk sg13g2_dfrbpq_2
XFILLER_36_543 VPWR VGND sg13g2_decap_8
XFILLER_36_565 VPWR VGND sg13g2_fill_2
XFILLER_24_738 VPWR VGND sg13g2_decap_4
XFILLER_23_18 VPWR VGND sg13g2_decap_8
XFILLER_20_911 VPWR VGND sg13g2_decap_8
XFILLER_23_29 VPWR VGND sg13g2_fill_1
XFILLER_31_281 VPWR VGND sg13g2_fill_1
X_2827_ _0718_ VPWR _0719_ VGND _0703_ _0716_ sg13g2_o21ai_1
XFILLER_20_988 VPWR VGND sg13g2_decap_8
X_2758_ _0622_ VPWR _0653_ VGND _0620_ _0623_ sg13g2_o21ai_1
X_1709_ _1027_ VPWR _1038_ VGND _0954_ _1028_ sg13g2_o21ai_1
X_2689_ VGND VPWR _0586_ _0584_ _0546_ sg13g2_or2_1
Xfanout423 net252 net423 VPWR VGND sg13g2_buf_2
Xfanout412 net416 net412 VPWR VGND sg13g2_buf_8
Xfanout401 net402 net401 VPWR VGND sg13g2_buf_8
Xfanout434 net435 net434 VPWR VGND sg13g2_buf_8
Xfanout456 net271 net456 VPWR VGND sg13g2_buf_8
XFILLER_24_1006 VPWR VGND sg13g2_decap_8
Xfanout445 net446 net445 VPWR VGND sg13g2_buf_2
XFILLER_47_808 VPWR VGND sg13g2_decap_8
Xfanout478 net216 net478 VPWR VGND sg13g2_buf_8
Xfanout467 net210 net467 VPWR VGND sg13g2_buf_8
Xfanout489 DP_1.matrix\[2\] net489 VPWR VGND sg13g2_buf_8
XFILLER_39_381 VPWR VGND sg13g2_decap_4
XFILLER_15_705 VPWR VGND sg13g2_fill_1
XFILLER_42_524 VPWR VGND sg13g2_fill_1
XFILLER_11_933 VPWR VGND sg13g2_decap_8
XFILLER_7_959 VPWR VGND sg13g2_decap_8
XFILLER_13_84 VPWR VGND sg13g2_fill_1
XFILLER_2_664 VPWR VGND sg13g2_decap_8
XFILLER_49_123 VPWR VGND sg13g2_decap_8
XFILLER_37_307 VPWR VGND sg13g2_fill_1
XFILLER_46_841 VPWR VGND sg13g2_decap_8
X_1991_ _1290_ VPWR _1292_ VGND _1289_ net201 sg13g2_o21ai_1
X_2612_ _0511_ net479 net432 VPWR VGND sg13g2_nand2_1
Xclkload11 VPWR clkload11/Y clknet_leaf_18_clk VGND sg13g2_inv_1
X_2543_ _0444_ _0414_ _0442_ _0443_ VPWR VGND sg13g2_and3_2
X_2474_ _0375_ _0376_ _0370_ _0377_ VPWR VGND sg13g2_nand3_1
XFILLER_24_502 VPWR VGND sg13g2_decap_8
X_3026_ net514 VGND VPWR net4 DP_1.I_range.out_data\[6\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_37_896 VPWR VGND sg13g2_decap_8
XFILLER_24_568 VPWR VGND sg13g2_decap_8
Xclkload5 VPWR clkload5/Y clknet_leaf_8_clk VGND sg13g2_inv_1
XFILLER_1_7 VPWR VGND sg13g2_decap_4
XFILLER_46_137 VPWR VGND sg13g2_decap_4
XFILLER_43_800 VPWR VGND sg13g2_decap_8
XFILLER_28_874 VPWR VGND sg13g2_decap_8
XFILLER_27_384 VPWR VGND sg13g2_decap_8
XFILLER_27_395 VPWR VGND sg13g2_decap_8
XFILLER_43_866 VPWR VGND sg13g2_decap_8
XFILLER_42_332 VPWR VGND sg13g2_decap_4
XFILLER_11_785 VPWR VGND sg13g2_fill_1
XFILLER_7_756 VPWR VGND sg13g2_decap_8
XFILLER_3_962 VPWR VGND sg13g2_decap_8
X_2190_ _1447_ VPWR _1472_ VGND _1468_ _1470_ sg13g2_o21ai_1
XFILLER_19_830 VPWR VGND sg13g2_decap_4
XFILLER_37_126 VPWR VGND sg13g2_decap_4
XFILLER_46_671 VPWR VGND sg13g2_decap_8
XFILLER_33_321 VPWR VGND sg13g2_decap_4
XFILLER_34_877 VPWR VGND sg13g2_decap_8
XFILLER_33_387 VPWR VGND sg13g2_decap_8
XFILLER_21_549 VPWR VGND sg13g2_decap_8
X_1974_ _1277_ VPWR _1280_ VGND _1276_ _1278_ sg13g2_o21ai_1
X_2526_ _0396_ VPWR _0427_ VGND _0394_ _0397_ sg13g2_o21ai_1
X_2457_ _0361_ _0353_ _0360_ VPWR VGND sg13g2_nand2_1
Xhold17 mac1.sum_lvl1_ff\[82\] VPWR VGND net57 sg13g2_dlygate4sd3_1
Xhold28 mac1.sum_lvl1_ff\[9\] VPWR VGND net68 sg13g2_dlygate4sd3_1
Xhold39 mac1.sum_lvl1_ff\[15\] VPWR VGND net79 sg13g2_dlygate4sd3_1
X_2388_ _0297_ DP_1.matrix\[79\] net381 VPWR VGND sg13g2_nand2_1
XFILLER_29_616 VPWR VGND sg13g2_decap_8
X_3009_ net525 VGND VPWR _0040_ mac1.products_ff\[3\] clknet_leaf_28_clk sg13g2_dfrbpq_1
XFILLER_24_332 VPWR VGND sg13g2_decap_8
XFILLER_40_825 VPWR VGND sg13g2_decap_8
XFILLER_25_899 VPWR VGND sg13g2_decap_8
XFILLER_40_869 VPWR VGND sg13g2_decap_8
XFILLER_20_593 VPWR VGND sg13g2_decap_8
XFILLER_3_203 VPWR VGND sg13g2_decap_8
XFILLER_0_965 VPWR VGND sg13g2_decap_8
XFILLER_48_947 VPWR VGND sg13g2_decap_8
XFILLER_16_800 VPWR VGND sg13g2_fill_1
XFILLER_15_310 VPWR VGND sg13g2_fill_2
XFILLER_16_855 VPWR VGND sg13g2_decap_8
XFILLER_43_685 VPWR VGND sg13g2_decap_8
XFILLER_42_140 VPWR VGND sg13g2_decap_8
XFILLER_30_313 VPWR VGND sg13g2_decap_8
XFILLER_30_379 VPWR VGND sg13g2_decap_4
X_1690_ _1008_ VPWR _1020_ VGND _1016_ _1018_ sg13g2_o21ai_1
X_2311_ _0221_ _0212_ _0223_ VPWR VGND sg13g2_xor2_1
XFILLER_39_925 VPWR VGND sg13g2_decap_8
X_2242_ _0153_ _0152_ _0154_ _0156_ VPWR VGND sg13g2_a21o_1
X_2173_ _1455_ _1449_ _1454_ VPWR VGND sg13g2_xnor2_1
XFILLER_19_693 VPWR VGND sg13g2_decap_8
XFILLER_46_490 VPWR VGND sg13g2_decap_4
XFILLER_34_652 VPWR VGND sg13g2_fill_1
XFILLER_21_313 VPWR VGND sg13g2_decap_8
XFILLER_21_379 VPWR VGND sg13g2_decap_8
X_1957_ _1266_ net278 mac1.sum_lvl2_ff\[12\] VPWR VGND sg13g2_nand2_1
X_1888_ _1212_ _1187_ _1211_ VPWR VGND sg13g2_xnor2_1
Xoutput29 net29 uo_out[4] VPWR VGND sg13g2_buf_1
Xoutput18 net18 uio_out[1] VPWR VGND sg13g2_buf_1
X_2509_ _0411_ _0383_ _0385_ VPWR VGND sg13g2_nand2_1
XFILLER_5_1014 VPWR VGND sg13g2_decap_8
XFILLER_29_435 VPWR VGND sg13g2_decap_8
XFILLER_45_928 VPWR VGND sg13g2_decap_8
XFILLER_44_416 VPWR VGND sg13g2_decap_8
XFILLER_16_107 VPWR VGND sg13g2_decap_8
XFILLER_38_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_36_clk clknet_3_0__leaf_clk clknet_leaf_36_clk VPWR VGND sg13g2_buf_8
XFILLER_24_162 VPWR VGND sg13g2_decap_8
XFILLER_25_674 VPWR VGND sg13g2_decap_8
XFILLER_25_685 VPWR VGND sg13g2_fill_2
XFILLER_13_869 VPWR VGND sg13g2_decap_8
XFILLER_4_567 VPWR VGND sg13g2_fill_2
XFILLER_4_556 VPWR VGND sg13g2_decap_8
XFILLER_21_95 VPWR VGND sg13g2_fill_2
XFILLER_43_1020 VPWR VGND sg13g2_decap_8
XFILLER_0_762 VPWR VGND sg13g2_decap_8
XFILLER_48_744 VPWR VGND sg13g2_decap_8
XFILLER_36_928 VPWR VGND sg13g2_decap_8
XFILLER_44_950 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_27_clk clknet_3_4__leaf_clk clknet_leaf_27_clk VPWR VGND sg13g2_buf_8
XFILLER_16_641 VPWR VGND sg13g2_fill_1
XFILLER_16_663 VPWR VGND sg13g2_fill_1
XFILLER_43_493 VPWR VGND sg13g2_fill_1
X_2860_ _0749_ _0747_ _0750_ VPWR VGND sg13g2_nor2b_1
X_1811_ _1137_ _1115_ _1138_ VPWR VGND sg13g2_nor2b_1
XFILLER_31_666 VPWR VGND sg13g2_decap_4
X_2791_ _0685_ _0680_ _0683_ VPWR VGND sg13g2_xnor2_1
XFILLER_12_891 VPWR VGND sg13g2_decap_8
XFILLER_8_851 VPWR VGND sg13g2_decap_8
XFILLER_7_64 VPWR VGND sg13g2_fill_2
X_1742_ _1071_ _1040_ _1069_ VPWR VGND sg13g2_xnor2_1
X_1673_ _1003_ net469 net405 VPWR VGND sg13g2_nand2_1
XFILLER_39_711 VPWR VGND sg13g2_fill_1
XFILLER_39_700 VPWR VGND sg13g2_decap_8
XFILLER_39_744 VPWR VGND sg13g2_decap_8
XFILLER_39_722 VPWR VGND sg13g2_fill_2
X_2225_ _0139_ _1499_ _0137_ _0138_ VPWR VGND sg13g2_and3_1
X_2156_ _1439_ _1409_ _1437_ VPWR VGND sg13g2_xnor2_1
XFILLER_27_939 VPWR VGND sg13g2_decap_8
XFILLER_42_909 VPWR VGND sg13g2_decap_8
X_2087_ _1367_ VPWR _1372_ VGND _1368_ _1370_ sg13g2_o21ai_1
XFILLER_26_449 VPWR VGND sg13g2_decap_8
XFILLER_35_950 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_18_clk clknet_3_6__leaf_clk clknet_leaf_18_clk VPWR VGND sg13g2_buf_8
XFILLER_22_644 VPWR VGND sg13g2_decap_8
XFILLER_34_493 VPWR VGND sg13g2_decap_4
XFILLER_10_817 VPWR VGND sg13g2_decap_8
X_2989_ net157 _0109_ VPWR VGND sg13g2_buf_1
XFILLER_45_703 VPWR VGND sg13g2_fill_2
XFILLER_45_725 VPWR VGND sg13g2_decap_8
XFILLER_44_202 VPWR VGND sg13g2_decap_8
XFILLER_44_235 VPWR VGND sg13g2_fill_2
XFILLER_26_972 VPWR VGND sg13g2_decap_8
XFILLER_41_920 VPWR VGND sg13g2_decap_8
XFILLER_16_73 VPWR VGND sg13g2_decap_8
XFILLER_16_84 VPWR VGND sg13g2_fill_1
XFILLER_40_430 VPWR VGND sg13g2_fill_1
XFILLER_12_132 VPWR VGND sg13g2_decap_8
XFILLER_41_997 VPWR VGND sg13g2_decap_8
XFILLER_40_474 VPWR VGND sg13g2_decap_4
XFILLER_8_125 VPWR VGND sg13g2_fill_2
XFILLER_8_114 VPWR VGND sg13g2_decap_8
XFILLER_32_83 VPWR VGND sg13g2_decap_4
XFILLER_5_832 VPWR VGND sg13g2_decap_8
XFILLER_48_541 VPWR VGND sg13g2_fill_2
X_2010_ mac1.sum_lvl3_ff\[8\] mac1.sum_lvl3_ff\[28\] _1307_ VPWR VGND sg13g2_and2_1
XFILLER_36_736 VPWR VGND sg13g2_decap_8
XFILLER_35_246 VPWR VGND sg13g2_decap_8
XFILLER_35_279 VPWR VGND sg13g2_fill_2
X_2912_ _0801_ _0800_ _0790_ VPWR VGND sg13g2_nand2b_1
XFILLER_32_920 VPWR VGND sg13g2_decap_8
XFILLER_32_997 VPWR VGND sg13g2_decap_8
X_2843_ _0733_ net446 _0732_ VPWR VGND sg13g2_nand2_1
X_2774_ _0668_ _0647_ _0669_ VPWR VGND sg13g2_nor2b_1
X_1725_ _1054_ net409 DP_1.matrix\[42\] VPWR VGND sg13g2_nand2_1
Xhold114 _0016_ VPWR VGND net154 sg13g2_dlygate4sd3_1
Xhold103 mac1.products_ff\[69\] VPWR VGND net143 sg13g2_dlygate4sd3_1
Xhold125 _0022_ VPWR VGND net165 sg13g2_dlygate4sd3_1
Xhold136 _0024_ VPWR VGND net176 sg13g2_dlygate4sd3_1
X_1656_ _0984_ _0985_ _0945_ _0987_ VPWR VGND sg13g2_nand3_1
Xhold147 _1336_ VPWR VGND net187 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_3_3__leaf_clk clknet_leaf_7_clk VPWR VGND sg13g2_buf_8
Xhold158 DP_2.matrix\[0\] VPWR VGND net198 sg13g2_dlygate4sd3_1
X_1587_ _0919_ _0916_ _0917_ VPWR VGND sg13g2_xnor2_1
Xhold169 _0018_ VPWR VGND net209 sg13g2_dlygate4sd3_1
X_3257_ net514 VGND VPWR net5 DP_1.Q_range.out_data\[2\] clknet_leaf_9_clk sg13g2_dfrbpq_2
XFILLER_39_596 VPWR VGND sg13g2_fill_2
XFILLER_2_1028 VPWR VGND sg13g2_fill_1
X_3188_ net522 VGND VPWR net71 mac1.sum_lvl2_ff\[49\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_2208_ _1489_ _1481_ _1488_ VPWR VGND sg13g2_nand2_1
X_2139_ _1422_ net447 net390 VPWR VGND sg13g2_nand2_1
XFILLER_35_791 VPWR VGND sg13g2_decap_8
XFILLER_22_430 VPWR VGND sg13g2_decap_8
XFILLER_23_975 VPWR VGND sg13g2_decap_8
XFILLER_10_647 VPWR VGND sg13g2_fill_2
XFILLER_6_629 VPWR VGND sg13g2_decap_8
XFILLER_5_106 VPWR VGND sg13g2_fill_1
XFILLER_2_846 VPWR VGND sg13g2_decap_8
XFILLER_49_305 VPWR VGND sg13g2_decap_8
XFILLER_40_1023 VPWR VGND sg13g2_decap_4
XFILLER_18_714 VPWR VGND sg13g2_decap_4
XFILLER_18_747 VPWR VGND sg13g2_decap_8
XFILLER_17_268 VPWR VGND sg13g2_fill_1
XFILLER_33_728 VPWR VGND sg13g2_decap_8
XFILLER_14_975 VPWR VGND sg13g2_decap_8
XFILLER_43_93 VPWR VGND sg13g2_fill_2
XFILLER_41_783 VPWR VGND sg13g2_decap_8
XFILLER_13_485 VPWR VGND sg13g2_decap_8
X_1510_ _0847_ net472 net412 net470 net417 VPWR VGND sg13g2_a22oi_1
X_2490_ _0392_ _0387_ _0390_ VPWR VGND sg13g2_xnor2_1
XFILLER_4_87 VPWR VGND sg13g2_decap_8
X_3111_ net529 VGND VPWR _0052_ mac1.products_ff\[150\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_3042_ net527 VGND VPWR _0095_ DP_1.matrix\[37\] clknet_leaf_30_clk sg13g2_dfrbpq_1
XFILLER_36_511 VPWR VGND sg13g2_decap_8
XFILLER_17_791 VPWR VGND sg13g2_fill_2
XFILLER_23_216 VPWR VGND sg13g2_fill_1
X_2826_ _0063_ _0702_ _0717_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_967 VPWR VGND sg13g2_decap_8
X_2757_ _0632_ VPWR _0652_ VGND _0630_ _0633_ sg13g2_o21ai_1
X_2688_ _0585_ net484 net424 VPWR VGND sg13g2_nand2_1
X_1708_ _1037_ _1032_ _1036_ VPWR VGND sg13g2_nand2_1
X_1639_ _0965_ VPWR _0970_ VGND _0966_ _0968_ sg13g2_o21ai_1
Xfanout402 net192 net402 VPWR VGND sg13g2_buf_8
Xfanout413 net416 net413 VPWR VGND sg13g2_buf_1
XFILLER_48_49 VPWR VGND sg13g2_decap_8
Xfanout424 net425 net424 VPWR VGND sg13g2_buf_8
Xfanout457 net458 net457 VPWR VGND sg13g2_buf_8
Xfanout446 net286 net446 VPWR VGND sg13g2_buf_2
Xfanout435 net436 net435 VPWR VGND sg13g2_buf_1
Xfanout479 net480 net479 VPWR VGND sg13g2_buf_8
Xfanout468 net212 net468 VPWR VGND sg13g2_buf_8
XFILLER_15_739 VPWR VGND sg13g2_decap_4
XFILLER_30_709 VPWR VGND sg13g2_fill_1
XFILLER_10_411 VPWR VGND sg13g2_decap_8
XFILLER_11_912 VPWR VGND sg13g2_decap_8
XFILLER_13_30 VPWR VGND sg13g2_decap_8
XFILLER_13_41 VPWR VGND sg13g2_fill_1
XFILLER_22_271 VPWR VGND sg13g2_fill_2
XFILLER_10_455 VPWR VGND sg13g2_decap_4
XFILLER_7_938 VPWR VGND sg13g2_decap_8
XFILLER_11_989 VPWR VGND sg13g2_decap_8
XFILLER_6_459 VPWR VGND sg13g2_decap_8
XFILLER_6_437 VPWR VGND sg13g2_decap_4
XFILLER_2_643 VPWR VGND sg13g2_decap_8
XFILLER_49_102 VPWR VGND sg13g2_decap_8
XFILLER_1_153 VPWR VGND sg13g2_fill_2
XFILLER_49_179 VPWR VGND sg13g2_decap_8
XFILLER_37_319 VPWR VGND sg13g2_fill_1
XFILLER_45_352 VPWR VGND sg13g2_decap_4
XFILLER_46_897 VPWR VGND sg13g2_decap_8
XFILLER_45_396 VPWR VGND sg13g2_fill_2
XFILLER_18_599 VPWR VGND sg13g2_fill_2
X_1990_ net201 _1289_ _0025_ VPWR VGND sg13g2_xor2_1
XFILLER_9_286 VPWR VGND sg13g2_decap_4
X_2611_ _0468_ VPWR _0510_ VGND _0466_ _0469_ sg13g2_o21ai_1
Xclkload12 clknet_leaf_21_clk clkload12/Y VPWR VGND sg13g2_inv_4
X_2542_ _0441_ _0439_ _0418_ _0443_ VPWR VGND sg13g2_a21o_1
XFILLER_47_1018 VPWR VGND sg13g2_decap_8
XFILLER_6_993 VPWR VGND sg13g2_decap_8
X_2473_ _0371_ VPWR _0376_ VGND _0372_ _0374_ sg13g2_o21ai_1
X_3025_ net514 VGND VPWR DP_1.I_range.data_plus_4\[6\] DP_1.I_range.out_data\[5\]
+ clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_36_330 VPWR VGND sg13g2_decap_8
XFILLER_37_875 VPWR VGND sg13g2_decap_8
XFILLER_20_731 VPWR VGND sg13g2_decap_4
XFILLER_20_775 VPWR VGND sg13g2_decap_8
Xclkload6 clknet_leaf_7_clk clkload6/Y VPWR VGND sg13g2_inv_4
X_2809_ _0699_ _0701_ _0702_ VPWR VGND sg13g2_nor2_1
XFILLER_30_1011 VPWR VGND sg13g2_decap_8
XFILLER_8_1012 VPWR VGND sg13g2_decap_8
XFILLER_15_503 VPWR VGND sg13g2_decap_8
XFILLER_43_845 VPWR VGND sg13g2_decap_8
XFILLER_42_311 VPWR VGND sg13g2_fill_2
XFILLER_15_536 VPWR VGND sg13g2_fill_2
XFILLER_42_366 VPWR VGND sg13g2_decap_4
XFILLER_30_528 VPWR VGND sg13g2_decap_8
XFILLER_24_84 VPWR VGND sg13g2_decap_8
XFILLER_30_539 VPWR VGND sg13g2_fill_2
XFILLER_11_753 VPWR VGND sg13g2_fill_1
XFILLER_10_285 VPWR VGND sg13g2_decap_4
XFILLER_7_735 VPWR VGND sg13g2_decap_8
XFILLER_40_72 VPWR VGND sg13g2_fill_2
XFILLER_3_941 VPWR VGND sg13g2_decap_8
XFILLER_34_8 VPWR VGND sg13g2_fill_1
XFILLER_27_7 VPWR VGND sg13g2_decap_8
XFILLER_37_105 VPWR VGND sg13g2_decap_8
XFILLER_19_820 VPWR VGND sg13g2_fill_1
XFILLER_34_856 VPWR VGND sg13g2_decap_8
XFILLER_21_506 VPWR VGND sg13g2_fill_1
X_1973_ _0005_ _1276_ net172 VPWR VGND sg13g2_xnor2_1
XFILLER_14_1017 VPWR VGND sg13g2_decap_8
XFILLER_14_1028 VPWR VGND sg13g2_fill_1
XFILLER_6_790 VPWR VGND sg13g2_decap_8
X_2525_ _0426_ _0421_ _0424_ VPWR VGND sg13g2_xnor2_1
X_2456_ _0358_ _0359_ _0360_ VPWR VGND sg13g2_nor2b_1
Xhold29 mac1.products_ff\[71\] VPWR VGND net69 sg13g2_dlygate4sd3_1
Xhold18 mac1.sum_lvl1_ff\[47\] VPWR VGND net58 sg13g2_dlygate4sd3_1
X_2387_ _0296_ net446 net502 VPWR VGND sg13g2_nand2_1
X_3008_ net523 VGND VPWR _0039_ mac1.products_ff\[2\] clknet_leaf_30_clk sg13g2_dfrbpq_1
XFILLER_24_311 VPWR VGND sg13g2_decap_8
XFILLER_36_182 VPWR VGND sg13g2_fill_2
XFILLER_12_517 VPWR VGND sg13g2_decap_8
XFILLER_40_848 VPWR VGND sg13g2_decap_8
XFILLER_24_399 VPWR VGND sg13g2_decap_4
XFILLER_20_572 VPWR VGND sg13g2_decap_8
XFILLER_4_749 VPWR VGND sg13g2_decap_8
XFILLER_0_944 VPWR VGND sg13g2_decap_8
XFILLER_48_926 VPWR VGND sg13g2_decap_8
XFILLER_35_61 VPWR VGND sg13g2_fill_1
XFILLER_30_358 VPWR VGND sg13g2_decap_8
X_2310_ _0222_ _0212_ _0221_ VPWR VGND sg13g2_nand2b_1
X_2241_ _0153_ _0154_ _0152_ _0155_ VPWR VGND sg13g2_nand3_1
XFILLER_39_904 VPWR VGND sg13g2_decap_8
XFILLER_25_4 VPWR VGND sg13g2_fill_2
X_2172_ _1454_ _1416_ _1451_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_436 VPWR VGND sg13g2_decap_4
XFILLER_34_631 VPWR VGND sg13g2_decap_8
XFILLER_21_303 VPWR VGND sg13g2_fill_1
XFILLER_33_152 VPWR VGND sg13g2_fill_1
XFILLER_33_196 VPWR VGND sg13g2_fill_2
X_1956_ _0002_ _1264_ _1265_ VPWR VGND sg13g2_xnor2_1
XFILLER_21_358 VPWR VGND sg13g2_decap_8
XFILLER_30_892 VPWR VGND sg13g2_decap_8
X_1887_ _1209_ _1203_ _1211_ VPWR VGND sg13g2_xor2_1
Xoutput19 net19 uio_out[2] VPWR VGND sg13g2_buf_1
XFILLER_0_218 VPWR VGND sg13g2_decap_8
X_2508_ _0408_ _0409_ _0410_ VPWR VGND sg13g2_and2_1
X_2439_ _0343_ _0344_ _0038_ VPWR VGND sg13g2_nor2_1
XFILLER_29_414 VPWR VGND sg13g2_decap_8
XFILLER_45_907 VPWR VGND sg13g2_decap_8
XFILLER_17_609 VPWR VGND sg13g2_decap_4
XFILLER_25_620 VPWR VGND sg13g2_decap_8
XFILLER_13_815 VPWR VGND sg13g2_decap_8
XFILLER_13_848 VPWR VGND sg13g2_decap_8
XFILLER_40_667 VPWR VGND sg13g2_fill_1
XFILLER_40_656 VPWR VGND sg13g2_decap_8
XFILLER_21_74 VPWR VGND sg13g2_decap_8
XFILLER_0_741 VPWR VGND sg13g2_decap_8
XFILLER_48_723 VPWR VGND sg13g2_decap_8
XFILLER_36_907 VPWR VGND sg13g2_decap_8
XFILLER_43_461 VPWR VGND sg13g2_decap_4
XFILLER_16_686 VPWR VGND sg13g2_decap_8
XFILLER_15_174 VPWR VGND sg13g2_decap_8
X_1810_ _1137_ _1116_ _1136_ VPWR VGND sg13g2_xnor2_1
X_2790_ _0684_ _0683_ _0680_ VPWR VGND sg13g2_nand2b_1
XFILLER_8_830 VPWR VGND sg13g2_decap_8
XFILLER_12_870 VPWR VGND sg13g2_decap_8
X_1741_ _1070_ _1040_ _1069_ VPWR VGND sg13g2_nand2_1
X_1672_ _0972_ VPWR _1002_ VGND _0963_ _0973_ sg13g2_o21ai_1
X_2224_ _1500_ VPWR _0138_ VGND _0134_ _0136_ sg13g2_o21ai_1
X_2155_ _1437_ _1409_ _1438_ VPWR VGND sg13g2_nor2b_1
XFILLER_27_918 VPWR VGND sg13g2_decap_8
XFILLER_38_233 VPWR VGND sg13g2_fill_1
XFILLER_26_428 VPWR VGND sg13g2_fill_2
XFILLER_38_288 VPWR VGND sg13g2_decap_4
X_2086_ _1367_ _1368_ _1370_ _1371_ VPWR VGND sg13g2_or3_1
XFILLER_22_612 VPWR VGND sg13g2_decap_8
XFILLER_22_623 VPWR VGND sg13g2_fill_1
XFILLER_34_472 VPWR VGND sg13g2_decap_8
XFILLER_42_29 VPWR VGND sg13g2_decap_8
XFILLER_22_667 VPWR VGND sg13g2_fill_1
X_2988_ net155 _0108_ VPWR VGND sg13g2_buf_1
X_1939_ VGND VPWR _1251_ _1252_ _1248_ net284 sg13g2_a21oi_2
XFILLER_27_1016 VPWR VGND sg13g2_decap_8
XFILLER_27_1027 VPWR VGND sg13g2_fill_2
XFILLER_26_951 VPWR VGND sg13g2_decap_8
XFILLER_12_111 VPWR VGND sg13g2_decap_4
XFILLER_13_634 VPWR VGND sg13g2_decap_8
XFILLER_41_976 VPWR VGND sg13g2_decap_8
XFILLER_40_453 VPWR VGND sg13g2_decap_8
XFILLER_8_104 VPWR VGND sg13g2_fill_1
XFILLER_5_811 VPWR VGND sg13g2_decap_8
XFILLER_10_1020 VPWR VGND sg13g2_decap_8
XFILLER_5_888 VPWR VGND sg13g2_decap_8
XFILLER_35_225 VPWR VGND sg13g2_decap_8
XFILLER_17_984 VPWR VGND sg13g2_decap_8
XFILLER_35_258 VPWR VGND sg13g2_fill_2
XFILLER_16_461 VPWR VGND sg13g2_decap_4
XFILLER_16_472 VPWR VGND sg13g2_fill_2
X_2911_ _0799_ _0797_ _0800_ VPWR VGND sg13g2_nor2b_1
XFILLER_32_976 VPWR VGND sg13g2_decap_8
XFILLER_31_475 VPWR VGND sg13g2_fill_1
X_2842_ _0728_ net379 _0732_ VPWR VGND sg13g2_and2_1
X_2773_ _0666_ _0665_ _0668_ VPWR VGND sg13g2_xor2_1
XFILLER_8_660 VPWR VGND sg13g2_fill_2
X_1724_ _1053_ net467 DP_2.matrix\[41\] VPWR VGND sg13g2_nand2_1
Xhold115 DP_1.matrix\[78\] VPWR VGND net155 sg13g2_dlygate4sd3_1
XFILLER_7_192 VPWR VGND sg13g2_decap_8
Xhold126 mac1.sum_lvl3_ff\[0\] VPWR VGND net166 sg13g2_dlygate4sd3_1
Xhold104 mac1.sum_lvl2_ff\[47\] VPWR VGND net144 sg13g2_dlygate4sd3_1
Xhold137 DP_2.matrix\[77\] VPWR VGND net177 sg13g2_dlygate4sd3_1
X_1655_ _0986_ _0945_ _0984_ _0985_ VPWR VGND sg13g2_and3_1
Xhold148 _0021_ VPWR VGND net188 sg13g2_dlygate4sd3_1
Xhold159 _0110_ VPWR VGND net199 sg13g2_dlygate4sd3_1
X_1586_ _0918_ _0916_ _0917_ VPWR VGND sg13g2_nand2b_1
X_3256_ net507 VGND VPWR net165 net24 clknet_leaf_6_clk sg13g2_dfrbpq_2
X_2207_ _1486_ _1482_ _1488_ VPWR VGND sg13g2_xor2_1
XFILLER_39_575 VPWR VGND sg13g2_decap_4
XFILLER_2_1007 VPWR VGND sg13g2_decap_8
X_3187_ net522 VGND VPWR net57 mac1.sum_lvl2_ff\[48\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2138_ _1392_ VPWR _1421_ VGND _1390_ _1393_ sg13g2_o21ai_1
X_2069_ _1350_ VPWR _1355_ VGND _1351_ _1353_ sg13g2_o21ai_1
XFILLER_26_258 VPWR VGND sg13g2_fill_2
XFILLER_35_770 VPWR VGND sg13g2_decap_8
XFILLER_22_453 VPWR VGND sg13g2_fill_1
XFILLER_23_954 VPWR VGND sg13g2_decap_8
XFILLER_6_619 VPWR VGND sg13g2_fill_1
XFILLER_2_825 VPWR VGND sg13g2_decap_8
XFILLER_1_302 VPWR VGND sg13g2_decap_8
XFILLER_40_1002 VPWR VGND sg13g2_decap_8
XFILLER_45_501 VPWR VGND sg13g2_decap_8
XFILLER_27_73 VPWR VGND sg13g2_fill_1
XFILLER_14_954 VPWR VGND sg13g2_decap_8
XFILLER_25_280 VPWR VGND sg13g2_decap_8
XFILLER_43_72 VPWR VGND sg13g2_decap_8
XFILLER_5_685 VPWR VGND sg13g2_decap_8
XFILLER_4_162 VPWR VGND sg13g2_fill_2
X_3110_ net529 VGND VPWR _0051_ mac1.products_ff\[149\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_1_891 VPWR VGND sg13g2_decap_8
XFILLER_49_895 VPWR VGND sg13g2_decap_8
X_3041_ net528 VGND VPWR _0094_ DP_1.matrix\[36\] clknet_leaf_30_clk sg13g2_dfrbpq_1
XFILLER_24_707 VPWR VGND sg13g2_decap_8
XFILLER_36_567 VPWR VGND sg13g2_fill_1
XFILLER_17_1026 VPWR VGND sg13g2_fill_2
X_2825_ _0717_ VPWR _0718_ VGND _0699_ _0701_ sg13g2_o21ai_1
XFILLER_20_946 VPWR VGND sg13g2_decap_8
Xclkbuf_3_2__f_clk clknet_0_clk clknet_3_2__leaf_clk VPWR VGND sg13g2_buf_8
X_2756_ _0651_ _0650_ _0648_ VPWR VGND sg13g2_nand2b_1
XFILLER_9_991 VPWR VGND sg13g2_decap_8
X_2687_ _0584_ net484 net421 VPWR VGND sg13g2_nand2_1
X_1707_ _1035_ _1034_ _0078_ VPWR VGND sg13g2_xor2_1
X_1638_ _0965_ _0966_ _0968_ _0969_ VPWR VGND sg13g2_or3_1
Xfanout414 net416 net414 VPWR VGND sg13g2_buf_8
Xfanout403 net404 net403 VPWR VGND sg13g2_buf_8
Xfanout425 net300 net425 VPWR VGND sg13g2_buf_8
XFILLER_48_28 VPWR VGND sg13g2_decap_8
X_1569_ _0902_ _0895_ _0900_ _0901_ VPWR VGND sg13g2_and3_1
Xfanout447 net448 net447 VPWR VGND sg13g2_buf_8
Xfanout436 DP_2.matrix\[1\] net436 VPWR VGND sg13g2_buf_1
Xfanout469 DP_1.matrix\[39\] net469 VPWR VGND sg13g2_buf_8
Xfanout458 net277 net458 VPWR VGND sg13g2_buf_8
X_3239_ net544 VGND VPWR net173 mac1.sum_lvl3_ff\[14\] clknet_leaf_19_clk sg13g2_dfrbpq_2
XFILLER_15_718 VPWR VGND sg13g2_decap_4
XFILLER_42_537 VPWR VGND sg13g2_decap_8
XFILLER_14_217 VPWR VGND sg13g2_fill_2
XFILLER_14_228 VPWR VGND sg13g2_decap_8
XFILLER_23_784 VPWR VGND sg13g2_decap_8
XFILLER_7_917 VPWR VGND sg13g2_decap_8
XFILLER_11_968 VPWR VGND sg13g2_decap_8
XFILLER_6_416 VPWR VGND sg13g2_decap_8
XFILLER_10_489 VPWR VGND sg13g2_decap_4
XFILLER_2_622 VPWR VGND sg13g2_decap_8
XFILLER_1_132 VPWR VGND sg13g2_fill_1
XFILLER_2_699 VPWR VGND sg13g2_decap_8
XFILLER_49_158 VPWR VGND sg13g2_decap_8
XFILLER_46_876 VPWR VGND sg13g2_decap_8
XFILLER_33_504 VPWR VGND sg13g2_fill_2
XFILLER_45_375 VPWR VGND sg13g2_decap_8
XFILLER_33_559 VPWR VGND sg13g2_fill_1
XFILLER_20_209 VPWR VGND sg13g2_decap_8
X_2610_ _0509_ _0504_ _0508_ VPWR VGND sg13g2_xnor2_1
Xclkload13 clknet_leaf_20_clk clkload13/Y VPWR VGND sg13g2_inv_4
XFILLER_6_972 VPWR VGND sg13g2_decap_8
X_2541_ _0439_ _0441_ _0418_ _0442_ VPWR VGND sg13g2_nand3_1
XFILLER_5_482 VPWR VGND sg13g2_fill_1
X_2472_ _0371_ _0372_ _0374_ _0375_ VPWR VGND sg13g2_or3_1
X_3024_ net514 VGND VPWR net3 DP_1.I_range.out_data\[4\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_37_854 VPWR VGND sg13g2_decap_8
XFILLER_20_743 VPWR VGND sg13g2_decap_8
Xclkload7 clkload7/Y clknet_leaf_12_clk VPWR VGND sg13g2_inv_2
X_2808_ _0701_ _0694_ _0700_ VPWR VGND sg13g2_nand2_1
X_2739_ _0635_ _0629_ _0634_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_419 VPWR VGND sg13g2_decap_8
XFILLER_47_607 VPWR VGND sg13g2_fill_2
XFILLER_28_810 VPWR VGND sg13g2_fill_2
XFILLER_27_331 VPWR VGND sg13g2_decap_8
XFILLER_27_342 VPWR VGND sg13g2_fill_1
XFILLER_24_30 VPWR VGND sg13g2_fill_2
XFILLER_30_507 VPWR VGND sg13g2_fill_2
XFILLER_24_63 VPWR VGND sg13g2_decap_8
XFILLER_7_714 VPWR VGND sg13g2_decap_8
XFILLER_6_235 VPWR VGND sg13g2_decap_8
XFILLER_40_40 VPWR VGND sg13g2_fill_1
XFILLER_3_920 VPWR VGND sg13g2_decap_8
XFILLER_3_997 VPWR VGND sg13g2_decap_8
XFILLER_2_474 VPWR VGND sg13g2_decap_8
XFILLER_49_60 VPWR VGND sg13g2_fill_1
XFILLER_2_485 VPWR VGND sg13g2_fill_2
XFILLER_19_843 VPWR VGND sg13g2_fill_1
XFILLER_46_651 VPWR VGND sg13g2_fill_1
XFILLER_19_887 VPWR VGND sg13g2_decap_8
XFILLER_45_183 VPWR VGND sg13g2_decap_8
XFILLER_33_334 VPWR VGND sg13g2_fill_1
X_1972_ net171 mac1.sum_lvl2_ff\[33\] _1279_ VPWR VGND sg13g2_xor2_1
XFILLER_46_0 VPWR VGND sg13g2_fill_2
X_2524_ _0425_ _0424_ _0421_ VPWR VGND sg13g2_nand2b_1
X_2455_ _0354_ VPWR _0359_ VGND _0355_ _0357_ sg13g2_o21ai_1
Xhold19 mac1.sum_lvl1_ff\[49\] VPWR VGND net59 sg13g2_dlygate4sd3_1
X_2386_ _0274_ VPWR _0295_ VGND _0271_ _0275_ sg13g2_o21ai_1
XFILLER_37_640 VPWR VGND sg13g2_decap_8
X_3007_ net524 VGND VPWR _0038_ mac1.products_ff\[1\] clknet_leaf_32_clk sg13g2_dfrbpq_1
XFILLER_24_301 VPWR VGND sg13g2_fill_1
XFILLER_36_172 VPWR VGND sg13g2_fill_2
XFILLER_20_551 VPWR VGND sg13g2_decap_8
XFILLER_4_728 VPWR VGND sg13g2_decap_8
XFILLER_10_54 VPWR VGND sg13g2_fill_2
XFILLER_10_65 VPWR VGND sg13g2_decap_8
XFILLER_0_923 VPWR VGND sg13g2_decap_8
XFILLER_48_905 VPWR VGND sg13g2_decap_8
XFILLER_47_437 VPWR VGND sg13g2_decap_8
XFILLER_19_63 VPWR VGND sg13g2_decap_8
XFILLER_19_74 VPWR VGND sg13g2_decap_8
XFILLER_19_128 VPWR VGND sg13g2_decap_8
XFILLER_16_824 VPWR VGND sg13g2_decap_4
XFILLER_27_161 VPWR VGND sg13g2_decap_8
XFILLER_28_662 VPWR VGND sg13g2_decap_4
XFILLER_43_654 VPWR VGND sg13g2_fill_2
XFILLER_15_312 VPWR VGND sg13g2_fill_1
XFILLER_27_183 VPWR VGND sg13g2_decap_8
XFILLER_28_695 VPWR VGND sg13g2_decap_4
XFILLER_31_816 VPWR VGND sg13g2_decap_8
XFILLER_42_197 VPWR VGND sg13g2_decap_4
XFILLER_30_337 VPWR VGND sg13g2_decap_8
XFILLER_7_500 VPWR VGND sg13g2_decap_8
XFILLER_3_794 VPWR VGND sg13g2_decap_8
X_2240_ _1473_ VPWR _0154_ VGND _1412_ _1474_ sg13g2_o21ai_1
XFILLER_18_4 VPWR VGND sg13g2_decap_4
X_2171_ _1416_ _1451_ _1453_ VPWR VGND sg13g2_and2_1
XFILLER_19_662 VPWR VGND sg13g2_decap_8
XFILLER_19_673 VPWR VGND sg13g2_decap_4
XFILLER_25_109 VPWR VGND sg13g2_decap_8
XFILLER_33_142 VPWR VGND sg13g2_fill_2
XFILLER_34_687 VPWR VGND sg13g2_fill_2
XFILLER_33_175 VPWR VGND sg13g2_decap_8
X_1955_ _1265_ _1259_ _1261_ VPWR VGND sg13g2_nand2_1
XFILLER_30_871 VPWR VGND sg13g2_decap_8
X_1886_ _1210_ _1203_ _1209_ VPWR VGND sg13g2_nand2_1
XFILLER_1_709 VPWR VGND sg13g2_decap_8
X_2507_ _0407_ _0405_ _0367_ _0409_ VPWR VGND sg13g2_a21o_1
X_2438_ _0344_ net433 net492 net490 net437 VPWR VGND sg13g2_a22oi_1
X_2369_ _0278_ _0269_ _0279_ VPWR VGND sg13g2_nor2b_1
XFILLER_37_492 VPWR VGND sg13g2_decap_8
XFILLER_40_635 VPWR VGND sg13g2_decap_8
XFILLER_40_613 VPWR VGND sg13g2_decap_8
XFILLER_9_809 VPWR VGND sg13g2_decap_8
XFILLER_13_827 VPWR VGND sg13g2_decap_8
XFILLER_24_186 VPWR VGND sg13g2_fill_2
XFILLER_8_319 VPWR VGND sg13g2_decap_4
XFILLER_12_337 VPWR VGND sg13g2_decap_8
XFILLER_21_882 VPWR VGND sg13g2_decap_8
XFILLER_20_392 VPWR VGND sg13g2_decap_8
XFILLER_21_20 VPWR VGND sg13g2_fill_2
XFILLER_21_42 VPWR VGND sg13g2_fill_2
XFILLER_21_53 VPWR VGND sg13g2_decap_8
XFILLER_0_720 VPWR VGND sg13g2_decap_8
XFILLER_48_713 VPWR VGND sg13g2_decap_4
XFILLER_0_797 VPWR VGND sg13g2_decap_8
XFILLER_48_779 VPWR VGND sg13g2_decap_8
XFILLER_47_267 VPWR VGND sg13g2_fill_1
XFILLER_35_407 VPWR VGND sg13g2_decap_8
XFILLER_46_94 VPWR VGND sg13g2_fill_2
XFILLER_28_481 VPWR VGND sg13g2_fill_2
XFILLER_44_985 VPWR VGND sg13g2_decap_8
XFILLER_16_654 VPWR VGND sg13g2_decap_8
XFILLER_43_484 VPWR VGND sg13g2_decap_8
XFILLER_31_624 VPWR VGND sg13g2_decap_4
XFILLER_7_11 VPWR VGND sg13g2_fill_1
XFILLER_7_341 VPWR VGND sg13g2_fill_2
XFILLER_11_381 VPWR VGND sg13g2_decap_4
X_1740_ _1068_ _1051_ _1069_ VPWR VGND sg13g2_xor2_1
XFILLER_30_189 VPWR VGND sg13g2_decap_8
XFILLER_8_886 VPWR VGND sg13g2_decap_8
XFILLER_7_66 VPWR VGND sg13g2_fill_1
X_1671_ _1001_ _0952_ _1000_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_591 VPWR VGND sg13g2_decap_8
X_2223_ _1500_ _0134_ _0136_ _0137_ VPWR VGND sg13g2_or3_1
XFILLER_38_201 VPWR VGND sg13g2_fill_1
XFILLER_39_779 VPWR VGND sg13g2_decap_8
X_2154_ _1437_ _1413_ _1436_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_407 VPWR VGND sg13g2_decap_8
XFILLER_38_256 VPWR VGND sg13g2_decap_4
X_2085_ _1370_ net393 net450 net447 net398 VPWR VGND sg13g2_a22oi_1
XFILLER_34_451 VPWR VGND sg13g2_decap_8
XFILLER_35_985 VPWR VGND sg13g2_decap_8
XFILLER_21_101 VPWR VGND sg13g2_decap_4
XFILLER_21_145 VPWR VGND sg13g2_decap_8
XFILLER_21_167 VPWR VGND sg13g2_decap_8
XFILLER_21_178 VPWR VGND sg13g2_fill_1
X_2987_ net445 _0107_ VPWR VGND sg13g2_buf_1
X_1938_ _1251_ mac1.sum_lvl2_ff\[27\] mac1.sum_lvl2_ff\[8\] VPWR VGND sg13g2_xnor2_1
XFILLER_30_690 VPWR VGND sg13g2_fill_2
X_1869_ _1192_ _1193_ _1194_ VPWR VGND sg13g2_and2_1
XFILLER_26_930 VPWR VGND sg13g2_decap_8
XFILLER_13_613 VPWR VGND sg13g2_decap_8
XFILLER_41_955 VPWR VGND sg13g2_decap_8
XFILLER_9_606 VPWR VGND sg13g2_decap_8
XFILLER_13_657 VPWR VGND sg13g2_fill_1
XFILLER_8_149 VPWR VGND sg13g2_decap_8
XFILLER_32_41 VPWR VGND sg13g2_fill_2
XFILLER_5_867 VPWR VGND sg13g2_decap_8
XFILLER_4_355 VPWR VGND sg13g2_decap_8
XFILLER_0_594 VPWR VGND sg13g2_decap_8
XFILLER_48_565 VPWR VGND sg13g2_decap_4
XFILLER_35_204 VPWR VGND sg13g2_decap_8
XFILLER_29_790 VPWR VGND sg13g2_decap_8
XFILLER_44_760 VPWR VGND sg13g2_decap_8
XFILLER_17_963 VPWR VGND sg13g2_decap_8
X_2910_ _0799_ net377 _0798_ _0783_ net391 VPWR VGND sg13g2_a22oi_1
XFILLER_31_432 VPWR VGND sg13g2_decap_4
XFILLER_32_955 VPWR VGND sg13g2_decap_8
X_2841_ DP_1.Q_range.out_data\[2\] DP_1.I_range.out_data\[2\] _0731_ VPWR VGND sg13g2_xor2_1
X_2772_ _0666_ _0665_ _0667_ VPWR VGND sg13g2_nor2b_1
X_1723_ _1017_ VPWR _1052_ VGND _1008_ _1018_ sg13g2_o21ai_1
Xhold116 DP_2.matrix\[80\] VPWR VGND net156 sg13g2_dlygate4sd3_1
Xhold105 mac1.sum_lvl1_ff\[1\] VPWR VGND net145 sg13g2_dlygate4sd3_1
Xhold138 mac1.sum_lvl3_ff\[5\] VPWR VGND net178 sg13g2_dlygate4sd3_1
Xhold127 _0023_ VPWR VGND net167 sg13g2_dlygate4sd3_1
X_1654_ _0918_ VPWR _0985_ VGND _0981_ _0983_ sg13g2_o21ai_1
Xhold149 DP_1.matrix\[44\] VPWR VGND net189 sg13g2_dlygate4sd3_1
X_1585_ _0917_ net475 net403 VPWR VGND sg13g2_nand2_1
X_3255_ net507 VGND VPWR net188 net23 clknet_leaf_5_clk sg13g2_dfrbpq_2
XFILLER_39_532 VPWR VGND sg13g2_decap_8
X_2206_ _1482_ _1486_ _1487_ VPWR VGND sg13g2_nor2_1
X_3186_ net511 VGND VPWR net78 mac1.sum_lvl2_ff\[47\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_26_204 VPWR VGND sg13g2_decap_8
X_2137_ _1420_ _1415_ _1418_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_215 VPWR VGND sg13g2_fill_2
XFILLER_42_719 VPWR VGND sg13g2_decap_8
X_2068_ _1350_ _1351_ _1353_ _1354_ VPWR VGND sg13g2_nor3_1
XFILLER_23_933 VPWR VGND sg13g2_decap_8
XFILLER_10_638 VPWR VGND sg13g2_decap_4
XFILLER_2_804 VPWR VGND sg13g2_decap_8
XFILLER_17_259 VPWR VGND sg13g2_decap_8
XFILLER_14_933 VPWR VGND sg13g2_decap_8
XFILLER_32_207 VPWR VGND sg13g2_fill_1
XFILLER_32_229 VPWR VGND sg13g2_fill_1
XFILLER_40_262 VPWR VGND sg13g2_fill_1
XFILLER_40_251 VPWR VGND sg13g2_fill_2
XFILLER_13_465 VPWR VGND sg13g2_decap_4
XFILLER_40_273 VPWR VGND sg13g2_decap_4
XFILLER_5_664 VPWR VGND sg13g2_decap_8
XFILLER_4_141 VPWR VGND sg13g2_decap_4
XFILLER_1_870 VPWR VGND sg13g2_decap_8
XFILLER_0_391 VPWR VGND sg13g2_decap_8
XFILLER_49_874 VPWR VGND sg13g2_decap_8
X_3040_ net539 VGND VPWR _0093_ DP_1.matrix\[7\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_17_1005 VPWR VGND sg13g2_decap_8
XFILLER_20_925 VPWR VGND sg13g2_decap_8
X_2824_ _0716_ _0703_ _0717_ VPWR VGND sg13g2_xor2_1
XFILLER_9_970 VPWR VGND sg13g2_decap_8
X_2755_ VGND VPWR _0650_ _0649_ _0595_ sg13g2_or2_1
X_2686_ _0583_ net489 net495 VPWR VGND sg13g2_nand2_1
X_1706_ _1036_ _1034_ _1035_ VPWR VGND sg13g2_nand2_1
X_1637_ _0968_ net461 net419 net462 net415 VPWR VGND sg13g2_a22oi_1
Xfanout404 net191 net404 VPWR VGND sg13g2_buf_8
X_1568_ _0896_ VPWR _0901_ VGND _0897_ _0899_ sg13g2_o21ai_1
Xfanout415 net416 net415 VPWR VGND sg13g2_buf_1
Xfanout437 net198 net437 VPWR VGND sg13g2_buf_8
Xfanout448 net449 net448 VPWR VGND sg13g2_buf_8
Xfanout426 net282 net426 VPWR VGND sg13g2_buf_8
Xfanout459 net461 net459 VPWR VGND sg13g2_buf_8
X_3238_ net527 VGND VPWR net281 mac1.sum_lvl3_ff\[13\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_27_502 VPWR VGND sg13g2_decap_4
X_3169_ net542 VGND VPWR net93 mac1.sum_lvl2_ff\[27\] clknet_leaf_25_clk sg13g2_dfrbpq_1
XFILLER_23_763 VPWR VGND sg13g2_decap_8
XFILLER_11_947 VPWR VGND sg13g2_decap_8
XFILLER_22_273 VPWR VGND sg13g2_fill_1
XFILLER_2_601 VPWR VGND sg13g2_decap_8
XFILLER_1_155 VPWR VGND sg13g2_fill_1
XFILLER_2_678 VPWR VGND sg13g2_decap_8
XFILLER_49_137 VPWR VGND sg13g2_decap_8
XFILLER_38_40 VPWR VGND sg13g2_decap_8
XFILLER_18_524 VPWR VGND sg13g2_decap_8
XFILLER_38_73 VPWR VGND sg13g2_decap_8
XFILLER_46_855 VPWR VGND sg13g2_decap_8
XFILLER_18_557 VPWR VGND sg13g2_decap_8
XFILLER_33_516 VPWR VGND sg13g2_decap_4
XFILLER_33_527 VPWR VGND sg13g2_decap_8
XFILLER_45_398 VPWR VGND sg13g2_fill_1
XFILLER_14_741 VPWR VGND sg13g2_decap_4
XFILLER_41_593 VPWR VGND sg13g2_fill_2
XFILLER_14_785 VPWR VGND sg13g2_fill_2
XFILLER_14_796 VPWR VGND sg13g2_decap_8
XFILLER_6_951 VPWR VGND sg13g2_decap_8
XFILLER_5_450 VPWR VGND sg13g2_decap_4
X_2540_ _0438_ _0437_ _0420_ _0441_ VPWR VGND sg13g2_a21o_1
X_2471_ _0374_ net436 net486 net485 net439 VPWR VGND sg13g2_a22oi_1
XFILLER_49_671 VPWR VGND sg13g2_fill_2
X_3023_ net514 VGND VPWR net2 DP_1.I_range.out_data\[3\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_48_181 VPWR VGND sg13g2_decap_8
XFILLER_36_387 VPWR VGND sg13g2_decap_8
Xclkload8 VPWR clkload8/Y clknet_leaf_22_clk VGND sg13g2_inv_1
X_2807_ _0700_ _0672_ _0695_ VPWR VGND sg13g2_nand2_1
X_2738_ _0633_ _0630_ _0634_ VPWR VGND sg13g2_xor2_1
X_2669_ _0566_ _0559_ _0567_ VPWR VGND sg13g2_xor2_1
XFILLER_39_192 VPWR VGND sg13g2_fill_2
XFILLER_28_888 VPWR VGND sg13g2_decap_8
XFILLER_23_593 VPWR VGND sg13g2_fill_1
XFILLER_10_298 VPWR VGND sg13g2_fill_2
XFILLER_2_420 VPWR VGND sg13g2_fill_1
XFILLER_3_976 VPWR VGND sg13g2_decap_8
XFILLER_2_464 VPWR VGND sg13g2_fill_1
XFILLER_38_619 VPWR VGND sg13g2_decap_8
XFILLER_19_866 VPWR VGND sg13g2_decap_8
XFILLER_46_685 VPWR VGND sg13g2_decap_8
XFILLER_18_387 VPWR VGND sg13g2_fill_2
X_1971_ mac1.sum_lvl2_ff\[33\] mac1.sum_lvl2_ff\[14\] _1278_ VPWR VGND sg13g2_nor2_1
X_2523_ _0423_ _0388_ _0424_ VPWR VGND sg13g2_xor2_1
X_2454_ _0354_ _0355_ _0357_ _0358_ VPWR VGND sg13g2_nor3_1
X_2385_ _0277_ _0270_ _0279_ _0294_ VPWR VGND sg13g2_a21o_1
Xinput1 ui_in[0] net1 VPWR VGND sg13g2_buf_1
XFILLER_28_129 VPWR VGND sg13g2_decap_4
X_3006_ net521 VGND VPWR _0037_ mac1.products_ff\[0\] clknet_leaf_33_clk sg13g2_dfrbpq_1
XFILLER_37_674 VPWR VGND sg13g2_decap_8
XFILLER_36_184 VPWR VGND sg13g2_fill_1
XFILLER_4_707 VPWR VGND sg13g2_decap_8
XFILLER_10_11 VPWR VGND sg13g2_decap_8
XFILLER_3_217 VPWR VGND sg13g2_decap_8
XFILLER_10_33 VPWR VGND sg13g2_decap_8
XFILLER_10_88 VPWR VGND sg13g2_decap_4
XFILLER_0_902 VPWR VGND sg13g2_decap_8
XFILLER_0_979 VPWR VGND sg13g2_decap_8
XFILLER_47_416 VPWR VGND sg13g2_decap_8
XFILLER_28_630 VPWR VGND sg13g2_fill_1
XFILLER_28_674 VPWR VGND sg13g2_fill_1
XFILLER_43_633 VPWR VGND sg13g2_decap_8
XFILLER_42_154 VPWR VGND sg13g2_decap_8
XFILLER_15_346 VPWR VGND sg13g2_decap_8
XFILLER_16_869 VPWR VGND sg13g2_decap_8
XFILLER_37_1008 VPWR VGND sg13g2_decap_8
XFILLER_24_880 VPWR VGND sg13g2_decap_8
XFILLER_3_773 VPWR VGND sg13g2_decap_8
XFILLER_39_939 VPWR VGND sg13g2_decap_8
X_2170_ VGND VPWR _1452_ _1450_ _1417_ sg13g2_or2_1
XFILLER_38_405 VPWR VGND sg13g2_decap_8
XFILLER_19_641 VPWR VGND sg13g2_decap_8
XFILLER_47_983 VPWR VGND sg13g2_decap_8
XFILLER_20_1023 VPWR VGND sg13g2_decap_4
XFILLER_46_482 VPWR VGND sg13g2_decap_4
XFILLER_18_173 VPWR VGND sg13g2_decap_8
XFILLER_18_184 VPWR VGND sg13g2_fill_2
XFILLER_34_611 VPWR VGND sg13g2_fill_1
XFILLER_34_666 VPWR VGND sg13g2_decap_8
XFILLER_21_327 VPWR VGND sg13g2_decap_8
XFILLER_21_338 VPWR VGND sg13g2_fill_2
X_1954_ _1264_ _1263_ _1262_ VPWR VGND sg13g2_nand2b_1
XFILLER_30_850 VPWR VGND sg13g2_decap_8
X_1885_ _1209_ _1204_ _1207_ VPWR VGND sg13g2_xnor2_1
X_2506_ _0405_ _0407_ _0367_ _0408_ VPWR VGND sg13g2_nand3_1
X_2437_ _0343_ net490 net433 _0037_ VPWR VGND sg13g2_and3_2
XFILLER_5_1028 VPWR VGND sg13g2_fill_1
X_2368_ _0278_ _0270_ _0277_ VPWR VGND sg13g2_xnor2_1
X_2299_ _0209_ _0201_ _0211_ VPWR VGND sg13g2_xor2_1
XFILLER_25_644 VPWR VGND sg13g2_fill_2
XFILLER_38_994 VPWR VGND sg13g2_decap_8
XFILLER_12_316 VPWR VGND sg13g2_decap_8
XFILLER_24_176 VPWR VGND sg13g2_decap_4
XFILLER_24_198 VPWR VGND sg13g2_decap_8
XFILLER_4_504 VPWR VGND sg13g2_fill_1
XFILLER_4_526 VPWR VGND sg13g2_fill_2
XFILLER_47_202 VPWR VGND sg13g2_decap_8
XFILLER_0_776 VPWR VGND sg13g2_decap_8
XFILLER_48_758 VPWR VGND sg13g2_decap_8
XFILLER_47_246 VPWR VGND sg13g2_decap_8
XFILLER_46_51 VPWR VGND sg13g2_decap_8
XFILLER_16_600 VPWR VGND sg13g2_decap_8
XFILLER_29_983 VPWR VGND sg13g2_decap_8
XFILLER_44_964 VPWR VGND sg13g2_decap_8
XFILLER_43_430 VPWR VGND sg13g2_decap_8
XFILLER_15_132 VPWR VGND sg13g2_decap_8
XFILLER_15_198 VPWR VGND sg13g2_decap_8
XFILLER_30_135 VPWR VGND sg13g2_decap_8
XFILLER_30_168 VPWR VGND sg13g2_decap_8
XFILLER_8_865 VPWR VGND sg13g2_decap_8
XFILLER_7_320 VPWR VGND sg13g2_decap_8
XFILLER_7_23 VPWR VGND sg13g2_decap_8
X_1670_ _1000_ _0991_ _0998_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_570 VPWR VGND sg13g2_decap_8
X_3271_ net517 VGND VPWR net12 DP_2.Q_range.out_data\[6\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_30_4 VPWR VGND sg13g2_decap_8
X_2222_ _0136_ net394 net440 net496 net400 VPWR VGND sg13g2_a22oi_1
XFILLER_39_758 VPWR VGND sg13g2_decap_8
X_2153_ _1436_ _1433_ _1435_ VPWR VGND sg13g2_nand2_1
X_2084_ net450 net447 net397 _1369_ VPWR VGND net392 sg13g2_nand4_1
XFILLER_46_290 VPWR VGND sg13g2_decap_8
XFILLER_35_964 VPWR VGND sg13g2_decap_8
XFILLER_21_124 VPWR VGND sg13g2_decap_4
XFILLER_22_658 VPWR VGND sg13g2_decap_8
X_2986_ net448 _0106_ VPWR VGND sg13g2_buf_1
X_1937_ mac1.sum_lvl2_ff\[27\] mac1.sum_lvl2_ff\[8\] _1250_ VPWR VGND sg13g2_and2_1
X_1868_ _1165_ _1167_ _1191_ _1193_ VPWR VGND sg13g2_or3_1
X_1799_ _1085_ VPWR _1126_ VGND _1082_ _1086_ sg13g2_o21ai_1
XFILLER_18_909 VPWR VGND sg13g2_decap_8
XFILLER_17_419 VPWR VGND sg13g2_decap_8
XFILLER_45_739 VPWR VGND sg13g2_decap_8
XFILLER_44_216 VPWR VGND sg13g2_decap_4
XFILLER_41_934 VPWR VGND sg13g2_decap_8
XFILLER_16_54 VPWR VGND sg13g2_fill_2
XFILLER_26_986 VPWR VGND sg13g2_decap_8
XFILLER_12_146 VPWR VGND sg13g2_decap_8
XFILLER_40_488 VPWR VGND sg13g2_fill_2
XFILLER_32_53 VPWR VGND sg13g2_decap_8
XFILLER_5_846 VPWR VGND sg13g2_decap_8
XFILLER_4_334 VPWR VGND sg13g2_decap_8
XFILLER_0_573 VPWR VGND sg13g2_decap_8
XFILLER_36_706 VPWR VGND sg13g2_fill_2
XFILLER_44_750 VPWR VGND sg13g2_fill_1
XFILLER_17_942 VPWR VGND sg13g2_decap_8
XFILLER_16_474 VPWR VGND sg13g2_fill_1
XFILLER_31_400 VPWR VGND sg13g2_fill_1
XFILLER_32_934 VPWR VGND sg13g2_decap_8
X_2840_ _0730_ DP_1.I_range.out_data\[2\] DP_1.Q_range.out_data\[2\] VPWR VGND sg13g2_xnor2_1
X_2771_ VGND VPWR _0626_ _0637_ _0666_ _0625_ sg13g2_a21oi_1
XFILLER_8_640 VPWR VGND sg13g2_fill_1
XFILLER_31_488 VPWR VGND sg13g2_decap_8
XFILLER_8_662 VPWR VGND sg13g2_fill_1
X_1722_ _1051_ _1041_ _1049_ VPWR VGND sg13g2_xnor2_1
Xhold117 DP_1.matrix\[79\] VPWR VGND net157 sg13g2_dlygate4sd3_1
X_1653_ _0918_ _0981_ _0983_ _0984_ VPWR VGND sg13g2_or3_1
Xhold106 mac1.products_ff\[147\] VPWR VGND net146 sg13g2_dlygate4sd3_1
Xhold139 _1297_ VPWR VGND net179 sg13g2_dlygate4sd3_1
Xhold128 mac1.sum_lvl2_ff\[34\] VPWR VGND net168 sg13g2_dlygate4sd3_1
X_1584_ _0891_ VPWR _0916_ VGND _0888_ _0892_ sg13g2_o21ai_1
XFILLER_39_511 VPWR VGND sg13g2_decap_8
X_3254_ net507 VGND VPWR net234 net22 clknet_leaf_5_clk sg13g2_dfrbpq_2
X_2205_ VGND VPWR _1486_ _1485_ _1484_ sg13g2_or2_1
X_3185_ net511 VGND VPWR net112 mac1.sum_lvl2_ff\[46\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2136_ _1419_ _1418_ _1415_ VPWR VGND sg13g2_nand2b_1
X_2067_ _1353_ net392 net452 net450 net397 VPWR VGND sg13g2_a22oi_1
XFILLER_41_208 VPWR VGND sg13g2_decap_8
XFILLER_23_912 VPWR VGND sg13g2_decap_8
XFILLER_22_444 VPWR VGND sg13g2_decap_8
XFILLER_23_989 VPWR VGND sg13g2_decap_8
X_2969_ _0841_ net423 net375 _0117_ VPWR VGND sg13g2_mux2_1
XFILLER_33_1022 VPWR VGND sg13g2_decap_8
XFILLER_49_319 VPWR VGND sg13g2_decap_8
XFILLER_17_205 VPWR VGND sg13g2_decap_8
XFILLER_27_53 VPWR VGND sg13g2_decap_4
XFILLER_27_64 VPWR VGND sg13g2_decap_8
XFILLER_14_912 VPWR VGND sg13g2_decap_8
XFILLER_25_260 VPWR VGND sg13g2_decap_4
XFILLER_26_783 VPWR VGND sg13g2_decap_8
XFILLER_41_731 VPWR VGND sg13g2_decap_8
XFILLER_13_433 VPWR VGND sg13g2_fill_2
XFILLER_13_444 VPWR VGND sg13g2_decap_8
XFILLER_14_989 VPWR VGND sg13g2_decap_8
XFILLER_40_296 VPWR VGND sg13g2_decap_8
XFILLER_9_459 VPWR VGND sg13g2_decap_8
XFILLER_5_643 VPWR VGND sg13g2_decap_8
XFILLER_4_131 VPWR VGND sg13g2_fill_1
XFILLER_4_164 VPWR VGND sg13g2_fill_1
XFILLER_49_853 VPWR VGND sg13g2_decap_8
XFILLER_36_525 VPWR VGND sg13g2_decap_4
XFILLER_36_536 VPWR VGND sg13g2_decap_8
XFILLER_16_271 VPWR VGND sg13g2_fill_2
XFILLER_16_282 VPWR VGND sg13g2_decap_8
XFILLER_32_720 VPWR VGND sg13g2_fill_2
XFILLER_32_731 VPWR VGND sg13g2_decap_8
XFILLER_17_1028 VPWR VGND sg13g2_fill_1
XFILLER_20_904 VPWR VGND sg13g2_decap_8
XFILLER_31_252 VPWR VGND sg13g2_fill_1
X_2823_ _0714_ _0704_ _0716_ VPWR VGND sg13g2_xor2_1
X_2754_ _0649_ net500 DP_2.matrix\[5\] VPWR VGND sg13g2_nand2_2
X_1705_ _0987_ VPWR _1035_ VGND _0948_ _0988_ sg13g2_o21ai_1
X_2685_ _0556_ VPWR _0582_ VGND _0554_ _0557_ sg13g2_o21ai_1
X_1636_ net415 net462 net419 _0967_ VPWR VGND net461 sg13g2_nand4_1
X_1567_ _0896_ _0897_ _0899_ _0900_ VPWR VGND sg13g2_or3_1
Xfanout405 DP_2.matrix\[41\] net405 VPWR VGND sg13g2_buf_8
Xfanout427 net237 net427 VPWR VGND sg13g2_buf_8
Xfanout438 net439 net438 VPWR VGND sg13g2_buf_2
Xfanout416 net268 net416 VPWR VGND sg13g2_buf_8
Xfanout449 net272 net449 VPWR VGND sg13g2_buf_2
X_3237_ net527 VGND VPWR _0003_ mac1.sum_lvl3_ff\[12\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_3168_ net537 VGND VPWR net129 mac1.sum_lvl2_ff\[26\] clknet_leaf_25_clk sg13g2_dfrbpq_1
XFILLER_39_363 VPWR VGND sg13g2_decap_4
XFILLER_39_385 VPWR VGND sg13g2_fill_2
XFILLER_39_396 VPWR VGND sg13g2_decap_8
X_2119_ _1401_ _1402_ _1363_ _1403_ VPWR VGND sg13g2_nand3_1
XFILLER_27_547 VPWR VGND sg13g2_decap_8
X_3099_ net508 VGND VPWR _0034_ mac1.products_ff\[138\] clknet_leaf_38_clk sg13g2_dfrbpq_1
XFILLER_23_742 VPWR VGND sg13g2_decap_4
XFILLER_35_580 VPWR VGND sg13g2_decap_8
XFILLER_10_425 VPWR VGND sg13g2_decap_8
XFILLER_11_926 VPWR VGND sg13g2_decap_8
XFILLER_13_11 VPWR VGND sg13g2_decap_8
XFILLER_1_123 VPWR VGND sg13g2_fill_1
XFILLER_2_657 VPWR VGND sg13g2_decap_8
XFILLER_49_116 VPWR VGND sg13g2_decap_8
XFILLER_46_834 VPWR VGND sg13g2_decap_8
XFILLER_41_572 VPWR VGND sg13g2_decap_8
XFILLER_9_212 VPWR VGND sg13g2_decap_8
XFILLER_6_930 VPWR VGND sg13g2_decap_8
XFILLER_10_992 VPWR VGND sg13g2_decap_8
X_2470_ net486 net485 net439 _0373_ VPWR VGND net436 sg13g2_nand4_1
XFILLER_49_650 VPWR VGND sg13g2_decap_8
XFILLER_23_1010 VPWR VGND sg13g2_decap_8
X_3022_ net514 VGND VPWR net1 DP_1.I_range.out_data\[2\] clknet_leaf_10_clk sg13g2_dfrbpq_2
XFILLER_37_889 VPWR VGND sg13g2_decap_8
XFILLER_32_572 VPWR VGND sg13g2_fill_1
Xclkload9 VPWR clkload9/Y clknet_leaf_25_clk VGND sg13g2_inv_1
X_2806_ VPWR VGND _0644_ _0698_ _0676_ _0612_ _0699_ _0675_ sg13g2_a221oi_1
XFILLER_30_1025 VPWR VGND sg13g2_decap_4
X_2737_ _0633_ _0584_ _0631_ VPWR VGND sg13g2_xnor2_1
X_2668_ _0566_ _0560_ _0564_ VPWR VGND sg13g2_xnor2_1
X_1619_ _0926_ VPWR _0950_ VGND _0889_ _0924_ sg13g2_o21ai_1
X_2599_ _0493_ _0497_ _0498_ VPWR VGND sg13g2_nor2_1
XFILLER_8_1026 VPWR VGND sg13g2_fill_2
XFILLER_27_377 VPWR VGND sg13g2_decap_8
XFILLER_43_859 VPWR VGND sg13g2_decap_8
XFILLER_42_336 VPWR VGND sg13g2_fill_1
XFILLER_42_325 VPWR VGND sg13g2_decap_8
XFILLER_24_32 VPWR VGND sg13g2_fill_1
XFILLER_23_572 VPWR VGND sg13g2_decap_8
XFILLER_10_222 VPWR VGND sg13g2_decap_4
XFILLER_24_98 VPWR VGND sg13g2_decap_8
XFILLER_10_255 VPWR VGND sg13g2_fill_2
XFILLER_7_749 VPWR VGND sg13g2_decap_8
XFILLER_3_955 VPWR VGND sg13g2_decap_8
XFILLER_49_95 VPWR VGND sg13g2_decap_8
XFILLER_37_119 VPWR VGND sg13g2_decap_8
XFILLER_46_642 VPWR VGND sg13g2_decap_8
XFILLER_18_322 VPWR VGND sg13g2_fill_1
XFILLER_46_664 VPWR VGND sg13g2_decap_8
XFILLER_34_815 VPWR VGND sg13g2_fill_2
XFILLER_34_826 VPWR VGND sg13g2_decap_4
X_1970_ _1277_ mac1.sum_lvl2_ff\[33\] mac1.sum_lvl2_ff\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_42_881 VPWR VGND sg13g2_decap_8
XFILLER_14_572 VPWR VGND sg13g2_decap_8
XFILLER_14_583 VPWR VGND sg13g2_fill_1
XFILLER_41_391 VPWR VGND sg13g2_fill_2
XFILLER_41_380 VPWR VGND sg13g2_decap_8
X_2522_ _0423_ net487 net429 VPWR VGND sg13g2_nand2_1
XFILLER_46_2 VPWR VGND sg13g2_fill_1
X_2453_ _0357_ DP_2.matrix\[1\] net488 net486 DP_2.matrix\[0\] VPWR VGND sg13g2_a22oi_1
X_2384_ _0293_ _0290_ _0050_ VPWR VGND sg13g2_xor2_1
XFILLER_29_609 VPWR VGND sg13g2_decap_8
XFILLER_28_119 VPWR VGND sg13g2_decap_4
Xinput2 ui_in[1] net2 VPWR VGND sg13g2_buf_1
X_3005_ net381 _0133_ VPWR VGND sg13g2_buf_1
XFILLER_24_325 VPWR VGND sg13g2_decap_8
XFILLER_36_196 VPWR VGND sg13g2_fill_2
XFILLER_20_586 VPWR VGND sg13g2_decap_8
XFILLER_0_958 VPWR VGND sg13g2_decap_8
XFILLER_43_601 VPWR VGND sg13g2_fill_2
XFILLER_16_848 VPWR VGND sg13g2_decap_8
XFILLER_35_42 VPWR VGND sg13g2_fill_1
XFILLER_43_656 VPWR VGND sg13g2_fill_1
XFILLER_42_133 VPWR VGND sg13g2_decap_8
XFILLER_35_75 VPWR VGND sg13g2_fill_1
XFILLER_42_188 VPWR VGND sg13g2_decap_4
XFILLER_30_306 VPWR VGND sg13g2_decap_8
XFILLER_11_597 VPWR VGND sg13g2_decap_4
XFILLER_3_752 VPWR VGND sg13g2_decap_8
XFILLER_2_251 VPWR VGND sg13g2_decap_8
XFILLER_32_8 VPWR VGND sg13g2_decap_4
XFILLER_39_918 VPWR VGND sg13g2_decap_8
XFILLER_20_1002 VPWR VGND sg13g2_decap_8
XFILLER_47_962 VPWR VGND sg13g2_decap_8
XFILLER_46_494 VPWR VGND sg13g2_fill_2
XFILLER_19_686 VPWR VGND sg13g2_decap_8
XFILLER_33_111 VPWR VGND sg13g2_decap_8
XFILLER_34_645 VPWR VGND sg13g2_decap_8
XFILLER_34_689 VPWR VGND sg13g2_fill_1
X_1953_ _1263_ mac1.sum_lvl2_ff\[30\] mac1.sum_lvl2_ff\[11\] VPWR VGND sg13g2_nand2_1
X_1884_ _1208_ _1207_ _1204_ VPWR VGND sg13g2_nand2b_1
X_2505_ _0404_ _0403_ _0386_ _0407_ VPWR VGND sg13g2_a21o_1
X_2436_ _0053_ _0335_ _0342_ VPWR VGND sg13g2_xnor2_1
XFILLER_5_1007 VPWR VGND sg13g2_decap_8
XFILLER_29_428 VPWR VGND sg13g2_decap_8
X_2367_ _0277_ _0271_ _0276_ VPWR VGND sg13g2_xnor2_1
X_2298_ _0209_ _0201_ _0210_ VPWR VGND sg13g2_nor2b_1
XFILLER_44_409 VPWR VGND sg13g2_decap_8
XFILLER_38_973 VPWR VGND sg13g2_decap_8
XFILLER_25_656 VPWR VGND sg13g2_decap_4
XFILLER_24_155 VPWR VGND sg13g2_decap_8
XFILLER_21_840 VPWR VGND sg13g2_decap_8
XFILLER_21_44 VPWR VGND sg13g2_fill_1
XFILLER_21_88 VPWR VGND sg13g2_decap_8
XFILLER_43_1013 VPWR VGND sg13g2_decap_8
XFILLER_0_755 VPWR VGND sg13g2_decap_8
XFILLER_48_737 VPWR VGND sg13g2_decap_8
XFILLER_46_30 VPWR VGND sg13g2_decap_8
XFILLER_29_962 VPWR VGND sg13g2_decap_8
XFILLER_44_943 VPWR VGND sg13g2_decap_8
XFILLER_16_634 VPWR VGND sg13g2_decap_8
XFILLER_46_96 VPWR VGND sg13g2_fill_1
XFILLER_15_111 VPWR VGND sg13g2_decap_8
XFILLER_15_188 VPWR VGND sg13g2_fill_1
XFILLER_31_648 VPWR VGND sg13g2_fill_1
XFILLER_31_659 VPWR VGND sg13g2_decap_8
XFILLER_8_844 VPWR VGND sg13g2_decap_8
XFILLER_7_46 VPWR VGND sg13g2_decap_4
XFILLER_12_884 VPWR VGND sg13g2_decap_8
XFILLER_7_343 VPWR VGND sg13g2_fill_1
X_3270_ net517 VGND VPWR DP_2.Q_range.data_plus_4\[6\] DP_2.Q_range.out_data\[5\]
+ clknet_leaf_11_clk sg13g2_dfrbpq_1
X_2221_ net440 net496 net399 _0135_ VPWR VGND net394 sg13g2_nand4_1
XFILLER_23_4 VPWR VGND sg13g2_decap_8
XFILLER_39_737 VPWR VGND sg13g2_decap_8
X_2152_ _1432_ _1431_ _1414_ _1435_ VPWR VGND sg13g2_a21o_1
X_2083_ net397 net450 net447 net393 _1368_ VPWR VGND sg13g2_and4_1
XFILLER_35_943 VPWR VGND sg13g2_decap_8
XFILLER_34_486 VPWR VGND sg13g2_decap_8
XFILLER_22_637 VPWR VGND sg13g2_decap_8
XFILLER_34_497 VPWR VGND sg13g2_fill_1
X_2985_ net451 _0105_ VPWR VGND sg13g2_buf_1
X_1936_ _1248_ _1249_ _0013_ VPWR VGND sg13g2_and2_1
XFILLER_30_681 VPWR VGND sg13g2_decap_4
XFILLER_30_692 VPWR VGND sg13g2_fill_1
X_1867_ _1191_ VPWR _1192_ VGND _1165_ _1167_ sg13g2_o21ai_1
X_1798_ _1125_ _1117_ _1122_ VPWR VGND sg13g2_xnor2_1
X_2419_ _0327_ _0322_ _0325_ VPWR VGND sg13g2_xnor2_1
XFILLER_45_718 VPWR VGND sg13g2_fill_2
XFILLER_16_11 VPWR VGND sg13g2_decap_8
XFILLER_16_22 VPWR VGND sg13g2_decap_8
XFILLER_26_965 VPWR VGND sg13g2_decap_8
XFILLER_37_280 VPWR VGND sg13g2_decap_8
XFILLER_41_913 VPWR VGND sg13g2_decap_8
XFILLER_12_125 VPWR VGND sg13g2_decap_8
XFILLER_40_478 VPWR VGND sg13g2_fill_2
XFILLER_40_467 VPWR VGND sg13g2_decap_8
XFILLER_32_43 VPWR VGND sg13g2_fill_1
XFILLER_32_76 VPWR VGND sg13g2_decap_8
XFILLER_32_87 VPWR VGND sg13g2_fill_2
XFILLER_5_825 VPWR VGND sg13g2_decap_8
XFILLER_0_552 VPWR VGND sg13g2_decap_8
XFILLER_48_556 VPWR VGND sg13g2_fill_1
XFILLER_17_921 VPWR VGND sg13g2_decap_8
XFILLER_36_729 VPWR VGND sg13g2_decap_8
XFILLER_35_239 VPWR VGND sg13g2_decap_8
XFILLER_17_998 VPWR VGND sg13g2_decap_8
XFILLER_32_913 VPWR VGND sg13g2_decap_8
XFILLER_43_294 VPWR VGND sg13g2_decap_8
X_2770_ _0663_ _0651_ _0665_ VPWR VGND sg13g2_xor2_1
XFILLER_12_681 VPWR VGND sg13g2_decap_8
XFILLER_11_191 VPWR VGND sg13g2_fill_2
XFILLER_12_692 VPWR VGND sg13g2_fill_2
X_1721_ _1041_ _1049_ _1050_ VPWR VGND sg13g2_nor2_1
Xhold107 mac1.sum_lvl1_ff\[74\] VPWR VGND net147 sg13g2_dlygate4sd3_1
X_1652_ VGND VPWR _0979_ _0980_ _0983_ _0949_ sg13g2_a21oi_1
Xhold118 DP_2.matrix\[41\] VPWR VGND net158 sg13g2_dlygate4sd3_1
Xhold129 _1281_ VPWR VGND net169 sg13g2_dlygate4sd3_1
X_1583_ _0908_ VPWR _0915_ VGND _0868_ _0909_ sg13g2_o21ai_1
X_3253_ net507 VGND VPWR net293 net21 clknet_leaf_30_clk sg13g2_dfrbpq_2
X_3184_ net511 VGND VPWR net109 mac1.sum_lvl2_ff\[45\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2204_ _1485_ net380 net456 net382 net453 VPWR VGND sg13g2_a22oi_1
X_2135_ _1417_ _1384_ _1418_ VPWR VGND sg13g2_xor2_1
XFILLER_27_718 VPWR VGND sg13g2_fill_2
X_2066_ net452 net450 net398 _1352_ VPWR VGND net392 sg13g2_nand4_1
XFILLER_35_784 VPWR VGND sg13g2_decap_8
XFILLER_23_968 VPWR VGND sg13g2_decap_8
XFILLER_33_1001 VPWR VGND sg13g2_decap_8
X_2968_ _0841_ _0786_ _0808_ VPWR VGND sg13g2_xnor2_1
X_1919_ mac1.sum_lvl2_ff\[23\] mac1.sum_lvl2_ff\[4\] _1236_ VPWR VGND sg13g2_and2_1
X_2899_ _0788_ net377 _0787_ _0783_ net385 VPWR VGND sg13g2_a22oi_1
XFILLER_1_316 VPWR VGND sg13g2_fill_2
XFILLER_2_839 VPWR VGND sg13g2_decap_8
XFILLER_40_1027 VPWR VGND sg13g2_fill_2
XFILLER_40_1016 VPWR VGND sg13g2_decap_8
XFILLER_18_707 VPWR VGND sg13g2_decap_8
XFILLER_18_718 VPWR VGND sg13g2_fill_2
XFILLER_45_515 VPWR VGND sg13g2_fill_2
XFILLER_45_548 VPWR VGND sg13g2_decap_4
XFILLER_17_239 VPWR VGND sg13g2_decap_4
XFILLER_27_98 VPWR VGND sg13g2_decap_4
XFILLER_25_294 VPWR VGND sg13g2_decap_8
XFILLER_41_776 VPWR VGND sg13g2_decap_8
XFILLER_40_253 VPWR VGND sg13g2_fill_1
XFILLER_14_968 VPWR VGND sg13g2_decap_8
XFILLER_43_86 VPWR VGND sg13g2_decap_8
XFILLER_13_478 VPWR VGND sg13g2_decap_8
XFILLER_5_699 VPWR VGND sg13g2_decap_8
XFILLER_49_832 VPWR VGND sg13g2_decap_8
XFILLER_36_504 VPWR VGND sg13g2_decap_8
XFILLER_1_1010 VPWR VGND sg13g2_decap_8
XFILLER_17_751 VPWR VGND sg13g2_decap_8
XFILLER_17_762 VPWR VGND sg13g2_fill_2
XFILLER_23_209 VPWR VGND sg13g2_decap_8
XFILLER_44_570 VPWR VGND sg13g2_decap_8
X_2822_ _0714_ _0704_ _0715_ VPWR VGND sg13g2_nor2b_1
X_2753_ _0648_ DP_2.matrix\[5\] net476 net428 net500 VPWR VGND sg13g2_a22oi_1
X_1704_ _1032_ _1033_ _1034_ VPWR VGND sg13g2_and2_1
X_2684_ _0548_ VPWR _0581_ VGND _0494_ _0546_ sg13g2_o21ai_1
X_1635_ net420 net414 net463 net461 _0966_ VPWR VGND sg13g2_and4_1
X_1566_ _0899_ net464 net419 net466 net413 VPWR VGND sg13g2_a22oi_1
Xfanout428 DP_2.matrix\[4\] net428 VPWR VGND sg13g2_buf_1
Xfanout417 net418 net417 VPWR VGND sg13g2_buf_8
Xfanout406 DP_2.matrix\[40\] net406 VPWR VGND sg13g2_buf_8
Xfanout439 DP_2.matrix\[0\] net439 VPWR VGND sg13g2_buf_2
X_3236_ net522 VGND VPWR _0002_ mac1.sum_lvl3_ff\[11\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_39_342 VPWR VGND sg13g2_decap_8
X_3167_ net536 VGND VPWR net122 mac1.sum_lvl2_ff\[25\] clknet_leaf_26_clk sg13g2_dfrbpq_1
X_3098_ net503 VGND VPWR _0033_ mac1.products_ff\[137\] clknet_leaf_38_clk sg13g2_dfrbpq_1
X_2118_ _1400_ _1399_ _1382_ _1402_ VPWR VGND sg13g2_a21o_1
X_2049_ _0022_ _1337_ net164 VPWR VGND sg13g2_xnor2_1
XFILLER_11_905 VPWR VGND sg13g2_decap_8
XFILLER_10_404 VPWR VGND sg13g2_decap_8
XFILLER_23_798 VPWR VGND sg13g2_decap_8
XFILLER_10_459 VPWR VGND sg13g2_fill_2
XFILLER_10_448 VPWR VGND sg13g2_decap_8
XFILLER_13_67 VPWR VGND sg13g2_fill_2
XFILLER_2_636 VPWR VGND sg13g2_decap_8
XFILLER_18_504 VPWR VGND sg13g2_decap_4
XFILLER_45_345 VPWR VGND sg13g2_decap_8
XFILLER_45_356 VPWR VGND sg13g2_fill_1
XFILLER_45_389 VPWR VGND sg13g2_decap_8
XFILLER_14_710 VPWR VGND sg13g2_decap_8
XFILLER_13_275 VPWR VGND sg13g2_fill_2
XFILLER_10_971 VPWR VGND sg13g2_decap_8
XFILLER_6_986 VPWR VGND sg13g2_decap_8
XFILLER_5_496 VPWR VGND sg13g2_decap_4
XFILLER_0_190 VPWR VGND sg13g2_decap_8
XFILLER_49_673 VPWR VGND sg13g2_fill_1
X_3021_ net547 VGND VPWR _0064_ mac1.products_ff\[15\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_36_323 VPWR VGND sg13g2_decap_8
XFILLER_37_868 VPWR VGND sg13g2_decap_8
XFILLER_17_570 VPWR VGND sg13g2_fill_2
XFILLER_32_540 VPWR VGND sg13g2_decap_8
XFILLER_20_724 VPWR VGND sg13g2_decap_8
X_2805_ _0698_ _0673_ _0696_ VPWR VGND sg13g2_nand2_1
XFILLER_20_757 VPWR VGND sg13g2_fill_1
XFILLER_20_768 VPWR VGND sg13g2_decap_8
XFILLER_30_1004 VPWR VGND sg13g2_decap_8
X_2736_ VGND VPWR _0632_ _0631_ _0584_ sg13g2_or2_1
X_2667_ _0565_ _0560_ _0564_ VPWR VGND sg13g2_nand2_1
X_1618_ _0941_ VPWR _0949_ VGND _0920_ _0942_ sg13g2_o21ai_1
XFILLER_8_1005 VPWR VGND sg13g2_decap_8
X_2598_ VGND VPWR _0497_ _0496_ _0495_ sg13g2_or2_1
X_1549_ _0883_ _0881_ _0880_ VPWR VGND sg13g2_nand2b_1
X_3219_ net522 VGND VPWR net92 mac1.sum_lvl3_ff\[30\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_27_301 VPWR VGND sg13g2_fill_1
XFILLER_43_838 VPWR VGND sg13g2_decap_8
XFILLER_42_304 VPWR VGND sg13g2_decap_8
XFILLER_15_529 VPWR VGND sg13g2_decap_8
XFILLER_23_540 VPWR VGND sg13g2_fill_2
XFILLER_11_724 VPWR VGND sg13g2_fill_2
XFILLER_24_77 VPWR VGND sg13g2_decap_8
XFILLER_7_728 VPWR VGND sg13g2_decap_8
XFILLER_3_934 VPWR VGND sg13g2_decap_8
XFILLER_2_400 VPWR VGND sg13g2_fill_2
XFILLER_2_411 VPWR VGND sg13g2_decap_8
XFILLER_18_312 VPWR VGND sg13g2_fill_1
XFILLER_18_389 VPWR VGND sg13g2_fill_1
XFILLER_27_890 VPWR VGND sg13g2_decap_8
XFILLER_45_197 VPWR VGND sg13g2_decap_4
XFILLER_42_860 VPWR VGND sg13g2_decap_8
X_2521_ _0422_ net487 net427 VPWR VGND sg13g2_nand2_1
XFILLER_6_783 VPWR VGND sg13g2_decap_8
X_2452_ net488 net486 net437 _0356_ VPWR VGND net433 sg13g2_nand4_1
X_2383_ VGND VPWR _0292_ _0293_ _0291_ _0233_ sg13g2_a21oi_2
XFILLER_37_610 VPWR VGND sg13g2_fill_2
X_3004_ net383 _0132_ VPWR VGND sg13g2_buf_1
Xinput3 ui_in[2] net3 VPWR VGND sg13g2_buf_1
XFILLER_37_621 VPWR VGND sg13g2_fill_2
XFILLER_37_654 VPWR VGND sg13g2_fill_1
XFILLER_33_882 VPWR VGND sg13g2_decap_8
XFILLER_20_565 VPWR VGND sg13g2_decap_8
X_2719_ _0612_ _0614_ _0611_ _0616_ VPWR VGND sg13g2_nand3_1
XFILLER_0_937 VPWR VGND sg13g2_decap_8
XFILLER_48_919 VPWR VGND sg13g2_decap_8
XFILLER_19_11 VPWR VGND sg13g2_fill_1
XFILLER_28_621 VPWR VGND sg13g2_decap_8
XFILLER_43_624 VPWR VGND sg13g2_fill_2
XFILLER_42_112 VPWR VGND sg13g2_fill_1
XFILLER_42_101 VPWR VGND sg13g2_decap_8
XFILLER_27_197 VPWR VGND sg13g2_decap_8
XFILLER_35_54 VPWR VGND sg13g2_decap_8
XFILLER_23_392 VPWR VGND sg13g2_decap_8
XFILLER_11_587 VPWR VGND sg13g2_fill_1
XFILLER_3_731 VPWR VGND sg13g2_decap_8
XFILLER_47_941 VPWR VGND sg13g2_decap_8
XFILLER_34_602 VPWR VGND sg13g2_decap_8
XFILLER_15_893 VPWR VGND sg13g2_decap_8
X_1952_ mac1.sum_lvl2_ff\[30\] mac1.sum_lvl2_ff\[11\] _1262_ VPWR VGND sg13g2_nor2_1
XFILLER_33_189 VPWR VGND sg13g2_decap_8
X_1883_ _1206_ _1179_ _1207_ VPWR VGND sg13g2_xor2_1
XFILLER_30_885 VPWR VGND sg13g2_decap_8
X_2504_ VGND VPWR _0403_ _0404_ _0406_ _0386_ sg13g2_a21oi_1
X_2435_ _0342_ _0336_ _0341_ VPWR VGND sg13g2_xnor2_1
XFILLER_29_407 VPWR VGND sg13g2_decap_8
X_2366_ _0273_ _0275_ _0276_ VPWR VGND sg13g2_nor2_1
X_2297_ _0209_ _0202_ _0208_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_952 VPWR VGND sg13g2_decap_8
XFILLER_25_602 VPWR VGND sg13g2_fill_2
XFILLER_37_462 VPWR VGND sg13g2_fill_2
XFILLER_24_112 VPWR VGND sg13g2_decap_4
XFILLER_25_646 VPWR VGND sg13g2_fill_1
XFILLER_24_145 VPWR VGND sg13g2_fill_1
XFILLER_21_896 VPWR VGND sg13g2_decap_8
XFILLER_4_528 VPWR VGND sg13g2_fill_1
XFILLER_21_67 VPWR VGND sg13g2_decap_8
XFILLER_0_734 VPWR VGND sg13g2_decap_8
XFILLER_47_237 VPWR VGND sg13g2_decap_4
XFILLER_29_941 VPWR VGND sg13g2_decap_8
XFILLER_44_922 VPWR VGND sg13g2_decap_8
XFILLER_44_999 VPWR VGND sg13g2_decap_8
XFILLER_30_115 VPWR VGND sg13g2_fill_1
XFILLER_31_638 VPWR VGND sg13g2_decap_4
XFILLER_8_823 VPWR VGND sg13g2_decap_8
XFILLER_12_863 VPWR VGND sg13g2_decap_8
XFILLER_11_395 VPWR VGND sg13g2_decap_8
X_2220_ net400 net440 net496 net394 _0134_ VPWR VGND sg13g2_and4_1
XFILLER_16_4 VPWR VGND sg13g2_decap_8
X_2151_ VGND VPWR _1431_ _1432_ _1434_ _1414_ sg13g2_a21oi_1
X_2082_ _1367_ net452 net390 VPWR VGND sg13g2_nand2_1
XFILLER_35_922 VPWR VGND sg13g2_decap_8
XFILLER_34_465 VPWR VGND sg13g2_decap_8
XFILLER_35_999 VPWR VGND sg13g2_decap_8
X_2984_ net453 _0104_ VPWR VGND sg13g2_buf_1
X_1935_ _1241_ _1244_ net305 _1249_ VPWR VGND sg13g2_or3_1
X_1866_ _1190_ _1176_ _1191_ VPWR VGND sg13g2_xor2_1
X_1797_ VGND VPWR _1124_ _1122_ _1117_ sg13g2_or2_1
XFILLER_27_1009 VPWR VGND sg13g2_decap_8
X_2418_ _0326_ _0325_ _0322_ VPWR VGND sg13g2_nand2b_1
X_2349_ VPWR _0260_ _0259_ VGND sg13g2_inv_1
XFILLER_29_226 VPWR VGND sg13g2_decap_8
XFILLER_26_944 VPWR VGND sg13g2_decap_8
XFILLER_12_104 VPWR VGND sg13g2_decap_8
XFILLER_12_115 VPWR VGND sg13g2_fill_2
XFILLER_13_627 VPWR VGND sg13g2_decap_8
XFILLER_41_969 VPWR VGND sg13g2_decap_8
XFILLER_21_660 VPWR VGND sg13g2_decap_4
XFILLER_5_804 VPWR VGND sg13g2_decap_8
XFILLER_20_181 VPWR VGND sg13g2_decap_8
XFILLER_10_1013 VPWR VGND sg13g2_decap_8
XFILLER_4_369 VPWR VGND sg13g2_decap_4
XFILLER_0_531 VPWR VGND sg13g2_decap_8
XFILLER_36_708 VPWR VGND sg13g2_fill_1
XFILLER_17_900 VPWR VGND sg13g2_decap_8
XFILLER_35_218 VPWR VGND sg13g2_decap_8
XFILLER_16_432 VPWR VGND sg13g2_decap_8
XFILLER_44_774 VPWR VGND sg13g2_decap_4
XFILLER_16_454 VPWR VGND sg13g2_decap_8
XFILLER_16_465 VPWR VGND sg13g2_fill_1
XFILLER_17_977 VPWR VGND sg13g2_decap_8
XFILLER_31_457 VPWR VGND sg13g2_decap_4
XFILLER_31_468 VPWR VGND sg13g2_decap_8
XFILLER_32_969 VPWR VGND sg13g2_decap_8
XFILLER_8_653 VPWR VGND sg13g2_decap_8
XFILLER_11_170 VPWR VGND sg13g2_decap_8
X_1720_ _1049_ _1042_ _1048_ VPWR VGND sg13g2_xnor2_1
XFILLER_8_697 VPWR VGND sg13g2_decap_8
X_1651_ _0979_ _0980_ _0949_ _0982_ VPWR VGND sg13g2_nand3_1
Xhold108 mac1.products_ff\[149\] VPWR VGND net148 sg13g2_dlygate4sd3_1
Xhold119 DP_2.matrix\[44\] VPWR VGND net159 sg13g2_dlygate4sd3_1
X_1582_ _0069_ _0886_ _0913_ VPWR VGND sg13g2_xnor2_1
X_3252_ net507 VGND VPWR net209 net20 clknet_leaf_30_clk sg13g2_dfrbpq_2
X_3183_ net512 VGND VPWR net54 mac1.sum_lvl2_ff\[44\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_2203_ net456 net453 net382 net380 _1484_ VPWR VGND sg13g2_and4_1
XFILLER_39_546 VPWR VGND sg13g2_fill_1
X_2134_ _1417_ net451 net388 VPWR VGND sg13g2_nand2_1
XFILLER_39_579 VPWR VGND sg13g2_fill_1
X_2065_ net397 net452 net450 net392 _1351_ VPWR VGND sg13g2_and4_1
XFILLER_19_270 VPWR VGND sg13g2_decap_8
XFILLER_22_402 VPWR VGND sg13g2_fill_1
XFILLER_23_947 VPWR VGND sg13g2_decap_8
X_2967_ _0840_ net424 net375 _0116_ VPWR VGND sg13g2_mux2_1
X_2898_ net405 net426 net378 _0787_ VPWR VGND sg13g2_mux2_1
X_1918_ _1233_ VPWR _1235_ VGND _1232_ _1234_ sg13g2_o21ai_1
X_1849_ _1175_ _1174_ _1142_ _1173_ _1111_ VPWR VGND sg13g2_a22oi_1
XFILLER_2_818 VPWR VGND sg13g2_decap_8
XFILLER_26_741 VPWR VGND sg13g2_fill_1
XFILLER_14_947 VPWR VGND sg13g2_decap_8
XFILLER_43_65 VPWR VGND sg13g2_decap_8
XFILLER_13_435 VPWR VGND sg13g2_fill_1
XFILLER_40_287 VPWR VGND sg13g2_decap_4
XFILLER_22_980 VPWR VGND sg13g2_decap_8
XFILLER_21_490 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_20_clk clknet_3_7__leaf_clk clknet_leaf_20_clk VPWR VGND sg13g2_buf_8
XFILLER_5_612 VPWR VGND sg13g2_decap_4
XFILLER_5_678 VPWR VGND sg13g2_decap_8
XFILLER_4_155 VPWR VGND sg13g2_decap_8
XFILLER_49_811 VPWR VGND sg13g2_decap_8
XFILLER_1_884 VPWR VGND sg13g2_decap_8
XFILLER_49_888 VPWR VGND sg13g2_decap_8
XFILLER_17_730 VPWR VGND sg13g2_decap_8
XFILLER_32_722 VPWR VGND sg13g2_fill_1
XFILLER_17_1019 VPWR VGND sg13g2_decap_8
X_2821_ _0714_ _0689_ _0713_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_939 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_11_clk clknet_3_2__leaf_clk clknet_leaf_11_clk VPWR VGND sg13g2_buf_8
X_2752_ _0634_ _0629_ _0636_ _0647_ VPWR VGND sg13g2_a21o_1
XFILLER_9_984 VPWR VGND sg13g2_decap_8
X_1703_ _1030_ _1029_ _1031_ _1033_ VPWR VGND sg13g2_a21o_1
X_2683_ _0568_ VPWR _0580_ VGND _0552_ _0569_ sg13g2_o21ai_1
X_1634_ _0965_ net411 net465 VPWR VGND sg13g2_nand2_1
X_1565_ net414 net466 net419 _0898_ VPWR VGND net464 sg13g2_nand4_1
Xfanout429 net229 net429 VPWR VGND sg13g2_buf_8
Xfanout418 net270 net418 VPWR VGND sg13g2_buf_8
Xfanout407 net238 net407 VPWR VGND sg13g2_buf_1
X_3235_ net523 VGND VPWR net303 mac1.sum_lvl3_ff\[10\] clknet_leaf_31_clk sg13g2_dfrbpq_1
XFILLER_39_321 VPWR VGND sg13g2_decap_8
X_3166_ net534 VGND VPWR net98 mac1.sum_lvl2_ff\[24\] clknet_leaf_26_clk sg13g2_dfrbpq_1
X_3097_ net507 VGND VPWR _0032_ mac1.products_ff\[136\] clknet_leaf_38_clk sg13g2_dfrbpq_1
X_2117_ _1399_ _1400_ _1382_ _1401_ VPWR VGND sg13g2_nand3_1
X_2048_ _1338_ mac1.sum_lvl3_ff\[15\] net163 VPWR VGND sg13g2_xnor2_1
XFILLER_22_232 VPWR VGND sg13g2_decap_8
XFILLER_22_243 VPWR VGND sg13g2_fill_1
XFILLER_13_24 VPWR VGND sg13g2_fill_2
XFILLER_23_777 VPWR VGND sg13g2_decap_8
XFILLER_6_409 VPWR VGND sg13g2_decap_8
XFILLER_2_615 VPWR VGND sg13g2_decap_8
XFILLER_38_54 VPWR VGND sg13g2_decap_4
XFILLER_38_87 VPWR VGND sg13g2_decap_4
XFILLER_46_869 VPWR VGND sg13g2_decap_8
XFILLER_45_368 VPWR VGND sg13g2_decap_8
XFILLER_41_552 VPWR VGND sg13g2_fill_2
XFILLER_41_541 VPWR VGND sg13g2_decap_8
XFILLER_10_950 VPWR VGND sg13g2_decap_8
XFILLER_6_965 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_1_681 VPWR VGND sg13g2_decap_8
X_3020_ net547 VGND VPWR _0063_ mac1.products_ff\[14\] clknet_leaf_16_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_0_clk clknet_3_0__leaf_clk clknet_leaf_0_clk VPWR VGND sg13g2_buf_8
XFILLER_48_195 VPWR VGND sg13g2_decap_8
XFILLER_37_847 VPWR VGND sg13g2_decap_8
X_2804_ _0062_ _0696_ _0697_ VPWR VGND sg13g2_xnor2_1
XFILLER_9_781 VPWR VGND sg13g2_decap_8
X_2735_ _0631_ net481 net424 VPWR VGND sg13g2_nand2_1
XFILLER_8_291 VPWR VGND sg13g2_decap_8
X_2666_ _0562_ _0563_ _0564_ VPWR VGND sg13g2_nor2_1
X_1617_ _0946_ VPWR _0948_ VGND _0912_ _0914_ sg13g2_o21ai_1
X_2597_ _0496_ net421 net491 net425 net489 VPWR VGND sg13g2_a22oi_1
XFILLER_8_1028 VPWR VGND sg13g2_fill_1
X_1548_ _0880_ _0881_ _0882_ VPWR VGND sg13g2_nor2b_1
X_3218_ net522 VGND VPWR net144 mac1.sum_lvl3_ff\[29\] clknet_leaf_31_clk sg13g2_dfrbpq_1
XFILLER_39_140 VPWR VGND sg13g2_decap_4
X_3149_ net534 VGND VPWR net60 mac1.sum_lvl2_ff\[4\] clknet_leaf_28_clk sg13g2_dfrbpq_1
XFILLER_27_324 VPWR VGND sg13g2_decap_8
XFILLER_24_23 VPWR VGND sg13g2_decap_8
XFILLER_24_45 VPWR VGND sg13g2_fill_2
XFILLER_24_56 VPWR VGND sg13g2_decap_8
XFILLER_7_707 VPWR VGND sg13g2_decap_8
XFILLER_10_257 VPWR VGND sg13g2_fill_1
XFILLER_6_206 VPWR VGND sg13g2_decap_4
XFILLER_6_228 VPWR VGND sg13g2_decap_8
XFILLER_3_913 VPWR VGND sg13g2_decap_8
XFILLER_46_1023 VPWR VGND sg13g2_decap_4
XFILLER_2_445 VPWR VGND sg13g2_decap_4
XFILLER_49_42 VPWR VGND sg13g2_decap_8
XFILLER_46_600 VPWR VGND sg13g2_fill_1
XFILLER_46_622 VPWR VGND sg13g2_decap_8
XFILLER_46_699 VPWR VGND sg13g2_decap_8
XFILLER_45_176 VPWR VGND sg13g2_decap_8
XFILLER_33_305 VPWR VGND sg13g2_decap_8
XFILLER_14_530 VPWR VGND sg13g2_decap_8
XFILLER_6_762 VPWR VGND sg13g2_decap_8
X_2520_ _0421_ net491 DP_2.matrix\[5\] VPWR VGND sg13g2_nand2_1
X_2451_ net437 net488 net486 net433 _0355_ VPWR VGND sg13g2_and4_1
X_2382_ VGND VPWR _0230_ _0259_ _0292_ _0261_ sg13g2_a21oi_1
XFILLER_49_493 VPWR VGND sg13g2_decap_4
X_3003_ net385 _0131_ VPWR VGND sg13g2_buf_1
Xinput4 ui_in[3] net4 VPWR VGND sg13g2_buf_1
XFILLER_36_165 VPWR VGND sg13g2_decap_8
XFILLER_37_688 VPWR VGND sg13g2_decap_4
XFILLER_24_349 VPWR VGND sg13g2_decap_4
XFILLER_36_198 VPWR VGND sg13g2_fill_1
XFILLER_20_533 VPWR VGND sg13g2_fill_1
XFILLER_32_371 VPWR VGND sg13g2_decap_8
X_2718_ VGND VPWR _0612_ _0614_ _0615_ _0611_ sg13g2_a21oi_1
X_2649_ _0546_ _0494_ _0547_ VPWR VGND sg13g2_xor2_1
XFILLER_10_47 VPWR VGND sg13g2_decap_8
XFILLER_0_916 VPWR VGND sg13g2_decap_8
XFILLER_16_817 VPWR VGND sg13g2_decap_8
XFILLER_28_655 VPWR VGND sg13g2_decap_8
XFILLER_43_603 VPWR VGND sg13g2_fill_1
XFILLER_16_828 VPWR VGND sg13g2_fill_1
XFILLER_27_154 VPWR VGND sg13g2_decap_8
XFILLER_27_176 VPWR VGND sg13g2_decap_8
XFILLER_28_688 VPWR VGND sg13g2_decap_8
XFILLER_28_699 VPWR VGND sg13g2_fill_2
XFILLER_43_669 VPWR VGND sg13g2_fill_2
XFILLER_43_647 VPWR VGND sg13g2_decap_8
XFILLER_31_809 VPWR VGND sg13g2_decap_8
XFILLER_42_168 VPWR VGND sg13g2_decap_8
XFILLER_11_511 VPWR VGND sg13g2_decap_8
XFILLER_24_894 VPWR VGND sg13g2_decap_8
XFILLER_3_710 VPWR VGND sg13g2_decap_8
XFILLER_3_787 VPWR VGND sg13g2_decap_8
XFILLER_47_920 VPWR VGND sg13g2_decap_8
XFILLER_19_611 VPWR VGND sg13g2_fill_1
XFILLER_46_441 VPWR VGND sg13g2_decap_8
XFILLER_18_121 VPWR VGND sg13g2_decap_8
XFILLER_19_655 VPWR VGND sg13g2_decap_8
XFILLER_47_997 VPWR VGND sg13g2_decap_8
XFILLER_19_677 VPWR VGND sg13g2_fill_1
XFILLER_33_135 VPWR VGND sg13g2_decap_8
XFILLER_15_872 VPWR VGND sg13g2_decap_8
XFILLER_33_168 VPWR VGND sg13g2_decap_8
X_1951_ net302 _1258_ _0001_ VPWR VGND sg13g2_xor2_1
XFILLER_30_864 VPWR VGND sg13g2_decap_8
X_1882_ _1206_ net404 net498 VPWR VGND sg13g2_nand2_1
X_2503_ _0403_ _0404_ _0386_ _0405_ VPWR VGND sg13g2_nand3_1
X_2434_ _0341_ _0328_ _0340_ VPWR VGND sg13g2_xnor2_1
XFILLER_37_0 VPWR VGND sg13g2_decap_8
X_2365_ _0275_ net381 net446 net383 net443 VPWR VGND sg13g2_a22oi_1
X_2296_ _0207_ _0203_ _0208_ VPWR VGND sg13g2_xor2_1
XFILLER_38_931 VPWR VGND sg13g2_decap_8
XFILLER_2_81 VPWR VGND sg13g2_decap_4
XFILLER_37_441 VPWR VGND sg13g2_decap_8
XFILLER_37_474 VPWR VGND sg13g2_decap_4
XFILLER_21_875 VPWR VGND sg13g2_decap_8
XFILLER_21_13 VPWR VGND sg13g2_decap_8
XFILLER_21_35 VPWR VGND sg13g2_decap_8
XFILLER_0_713 VPWR VGND sg13g2_decap_8
XFILLER_48_717 VPWR VGND sg13g2_fill_1
XFILLER_48_706 VPWR VGND sg13g2_decap_8
XFILLER_47_216 VPWR VGND sg13g2_decap_4
XFILLER_29_920 VPWR VGND sg13g2_decap_8
XFILLER_44_901 VPWR VGND sg13g2_decap_8
XFILLER_16_614 VPWR VGND sg13g2_decap_8
XFILLER_28_452 VPWR VGND sg13g2_fill_2
XFILLER_28_474 VPWR VGND sg13g2_decap_8
XFILLER_29_997 VPWR VGND sg13g2_decap_8
XFILLER_46_87 VPWR VGND sg13g2_decap_8
XFILLER_43_444 VPWR VGND sg13g2_decap_4
XFILLER_16_647 VPWR VGND sg13g2_decap_8
XFILLER_44_978 VPWR VGND sg13g2_decap_8
XFILLER_31_617 VPWR VGND sg13g2_decap_8
XFILLER_8_802 VPWR VGND sg13g2_decap_8
XFILLER_12_842 VPWR VGND sg13g2_decap_8
XFILLER_30_149 VPWR VGND sg13g2_decap_4
XFILLER_11_363 VPWR VGND sg13g2_decap_4
XFILLER_8_879 VPWR VGND sg13g2_decap_8
XFILLER_7_334 VPWR VGND sg13g2_decap_8
XFILLER_11_385 VPWR VGND sg13g2_fill_2
XFILLER_3_584 VPWR VGND sg13g2_decap_8
X_2150_ _1431_ _1432_ _1414_ _1433_ VPWR VGND sg13g2_nand3_1
XFILLER_38_227 VPWR VGND sg13g2_fill_2
X_2081_ _1352_ VPWR _1366_ VGND _1350_ _1353_ sg13g2_o21ai_1
XFILLER_38_249 VPWR VGND sg13g2_decap_8
XFILLER_35_901 VPWR VGND sg13g2_decap_8
XFILLER_47_794 VPWR VGND sg13g2_decap_4
XFILLER_34_444 VPWR VGND sg13g2_decap_8
XFILLER_35_978 VPWR VGND sg13g2_decap_8
X_2983_ net454 _0103_ VPWR VGND sg13g2_buf_1
XFILLER_21_105 VPWR VGND sg13g2_fill_2
X_1934_ _1247_ VPWR _1248_ VGND _1241_ _1244_ sg13g2_o21ai_1
X_1865_ _1188_ _1162_ _1190_ VPWR VGND sg13g2_xor2_1
X_1796_ _1117_ _1122_ _1123_ VPWR VGND sg13g2_and2_1
X_2417_ _0324_ _0297_ _0325_ VPWR VGND sg13g2_xor2_1
X_2348_ _0227_ _0258_ _0225_ _0259_ VPWR VGND sg13g2_nand3_1
X_2279_ _0192_ _0162_ _0191_ VPWR VGND sg13g2_nand2_1
XFILLER_26_923 VPWR VGND sg13g2_decap_8
XFILLER_25_433 VPWR VGND sg13g2_fill_2
XFILLER_37_271 VPWR VGND sg13g2_decap_4
XFILLER_41_948 VPWR VGND sg13g2_decap_8
XFILLER_32_12 VPWR VGND sg13g2_fill_1
XFILLER_4_315 VPWR VGND sg13g2_decap_4
XFILLER_4_348 VPWR VGND sg13g2_decap_8
XFILLER_0_510 VPWR VGND sg13g2_decap_8
XFILLER_0_587 VPWR VGND sg13g2_decap_8
XFILLER_48_569 VPWR VGND sg13g2_fill_2
XFILLER_29_783 VPWR VGND sg13g2_decap_8
XFILLER_16_411 VPWR VGND sg13g2_decap_8
XFILLER_16_422 VPWR VGND sg13g2_fill_2
XFILLER_17_956 VPWR VGND sg13g2_decap_8
XFILLER_43_252 VPWR VGND sg13g2_decap_8
XFILLER_43_285 VPWR VGND sg13g2_decap_4
XFILLER_31_425 VPWR VGND sg13g2_decap_8
XFILLER_32_948 VPWR VGND sg13g2_decap_8
XFILLER_31_436 VPWR VGND sg13g2_fill_2
XFILLER_40_981 VPWR VGND sg13g2_decap_8
XFILLER_11_160 VPWR VGND sg13g2_fill_1
X_1650_ _0981_ _0949_ _0979_ _0980_ VPWR VGND sg13g2_and3_1
X_1581_ _0865_ _0882_ _0884_ _0911_ _0914_ VPWR VGND sg13g2_nor4_1
Xhold109 mac1.sum_lvl1_ff\[51\] VPWR VGND net149 sg13g2_dlygate4sd3_1
XFILLER_4_882 VPWR VGND sg13g2_decap_8
X_3251_ net507 VGND VPWR net214 net19 clknet_leaf_31_clk sg13g2_dfrbpq_2
XFILLER_26_1021 VPWR VGND sg13g2_decap_8
XFILLER_39_525 VPWR VGND sg13g2_decap_8
X_3182_ net509 VGND VPWR net134 mac1.sum_lvl2_ff\[43\] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_2202_ _1483_ net453 net380 VPWR VGND sg13g2_nand2_1
XFILLER_39_569 VPWR VGND sg13g2_fill_1
XFILLER_39_558 VPWR VGND sg13g2_fill_2
X_2133_ _1416_ net450 net386 VPWR VGND sg13g2_nand2_1
X_2064_ _1350_ net454 net390 VPWR VGND sg13g2_nand2_1
XFILLER_35_742 VPWR VGND sg13g2_fill_1
XFILLER_23_926 VPWR VGND sg13g2_decap_8
XFILLER_34_296 VPWR VGND sg13g2_decap_4
X_2966_ _0807_ _0805_ _0840_ VPWR VGND sg13g2_xor2_1
X_2897_ _0786_ net377 _0785_ _0783_ net381 VPWR VGND sg13g2_a22oi_1
X_1917_ net244 _1232_ _0009_ VPWR VGND sg13g2_xor2_1
XFILLER_31_992 VPWR VGND sg13g2_decap_8
X_1848_ _1174_ _1109_ _1140_ VPWR VGND sg13g2_nand2_1
X_1779_ _1105_ _1078_ _1107_ VPWR VGND sg13g2_xor2_1
XFILLER_1_318 VPWR VGND sg13g2_fill_1
XFILLER_26_720 VPWR VGND sg13g2_fill_1
XFILLER_38_591 VPWR VGND sg13g2_decap_8
XFILLER_14_926 VPWR VGND sg13g2_decap_8
XFILLER_26_797 VPWR VGND sg13g2_decap_8
XFILLER_40_244 VPWR VGND sg13g2_decap_8
XFILLER_40_222 VPWR VGND sg13g2_decap_8
XFILLER_13_458 VPWR VGND sg13g2_decap_8
XFILLER_43_99 VPWR VGND sg13g2_decap_8
XFILLER_40_266 VPWR VGND sg13g2_decap_8
XFILLER_13_469 VPWR VGND sg13g2_fill_1
XFILLER_5_657 VPWR VGND sg13g2_decap_8
XFILLER_4_101 VPWR VGND sg13g2_decap_4
XFILLER_49_1021 VPWR VGND sg13g2_decap_8
XFILLER_4_145 VPWR VGND sg13g2_fill_1
XFILLER_1_863 VPWR VGND sg13g2_decap_8
XFILLER_49_867 VPWR VGND sg13g2_decap_8
XFILLER_0_384 VPWR VGND sg13g2_decap_8
XFILLER_48_388 VPWR VGND sg13g2_fill_2
XFILLER_16_296 VPWR VGND sg13g2_decap_8
XFILLER_31_222 VPWR VGND sg13g2_decap_8
X_2820_ _0711_ _0705_ _0713_ VPWR VGND sg13g2_xor2_1
XFILLER_13_981 VPWR VGND sg13g2_decap_8
XFILLER_20_918 VPWR VGND sg13g2_decap_8
XFILLER_9_963 VPWR VGND sg13g2_decap_8
XFILLER_8_440 VPWR VGND sg13g2_decap_8
X_2751_ _0646_ _0645_ _0060_ VPWR VGND sg13g2_xor2_1
X_2682_ VGND VPWR _0543_ _0549_ _0579_ _0551_ sg13g2_a21oi_1
X_1702_ _1030_ _1031_ _1029_ _1032_ VPWR VGND sg13g2_nand3_1
X_1633_ _0931_ VPWR _0964_ VGND _0929_ _0932_ sg13g2_o21ai_1
X_1564_ net419 net413 net466 net464 _0897_ VPWR VGND sg13g2_and4_1
Xfanout419 DP_2.matrix\[36\] net419 VPWR VGND sg13g2_buf_8
Xfanout408 net203 net408 VPWR VGND sg13g2_buf_8
X_3234_ net521 VGND VPWR _0015_ mac1.sum_lvl3_ff\[9\] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_3165_ net534 VGND VPWR net55 mac1.sum_lvl2_ff\[23\] clknet_leaf_26_clk sg13g2_dfrbpq_1
XFILLER_27_506 VPWR VGND sg13g2_fill_2
XFILLER_27_517 VPWR VGND sg13g2_fill_2
X_2116_ _1388_ VPWR _1400_ VGND _1396_ _1398_ sg13g2_o21ai_1
X_3096_ net546 VGND VPWR _0075_ mac1.products_ff\[83\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_2047_ _1334_ VPWR _1337_ VGND _1333_ _1335_ sg13g2_o21ai_1
XFILLER_23_701 VPWR VGND sg13g2_decap_8
XFILLER_23_712 VPWR VGND sg13g2_fill_2
XFILLER_35_561 VPWR VGND sg13g2_fill_2
XFILLER_23_756 VPWR VGND sg13g2_decap_8
X_2949_ _0762_ _0764_ _0830_ VPWR VGND sg13g2_nor2b_1
XFILLER_13_47 VPWR VGND sg13g2_fill_1
XFILLER_13_69 VPWR VGND sg13g2_fill_1
XFILLER_38_22 VPWR VGND sg13g2_decap_8
XFILLER_46_848 VPWR VGND sg13g2_decap_8
XFILLER_14_734 VPWR VGND sg13g2_decap_8
XFILLER_14_745 VPWR VGND sg13g2_fill_1
XFILLER_41_586 VPWR VGND sg13g2_decap_8
XFILLER_9_226 VPWR VGND sg13g2_decap_8
XFILLER_6_944 VPWR VGND sg13g2_decap_8
XFILLER_5_421 VPWR VGND sg13g2_fill_2
XFILLER_5_410 VPWR VGND sg13g2_decap_8
XFILLER_5_454 VPWR VGND sg13g2_fill_1
XFILLER_1_660 VPWR VGND sg13g2_decap_8
XFILLER_49_664 VPWR VGND sg13g2_decap_8
XFILLER_23_1024 VPWR VGND sg13g2_decap_4
XFILLER_49_686 VPWR VGND sg13g2_decap_8
XFILLER_48_174 VPWR VGND sg13g2_decap_8
XFILLER_24_509 VPWR VGND sg13g2_decap_8
X_2803_ VGND VPWR _0673_ _0677_ _0697_ _0672_ sg13g2_a21oi_1
XFILLER_9_760 VPWR VGND sg13g2_decap_8
X_2734_ _0630_ net487 net495 VPWR VGND sg13g2_nand2_1
X_2665_ _0563_ net432 net476 net434 net501 VPWR VGND sg13g2_a22oi_1
X_1616_ _0076_ _0914_ _0947_ VPWR VGND sg13g2_xnor2_1
X_2596_ net491 net489 net425 net421 _0495_ VPWR VGND sg13g2_and4_1
XFILLER_5_70 VPWR VGND sg13g2_fill_2
X_1547_ _0881_ _0861_ _0863_ VPWR VGND sg13g2_nand2_1
X_3217_ net511 VGND VPWR net136 mac1.sum_lvl3_ff\[28\] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_3148_ net526 VGND VPWR net116 mac1.sum_lvl2_ff\[3\] clknet_leaf_27_clk sg13g2_dfrbpq_1
XFILLER_39_185 VPWR VGND sg13g2_decap_8
XFILLER_43_807 VPWR VGND sg13g2_fill_2
X_3079_ net538 VGND VPWR _0132_ DP_2.matrix\[78\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_23_586 VPWR VGND sg13g2_decap_8
XFILLER_49_21 VPWR VGND sg13g2_decap_8
XFILLER_46_1002 VPWR VGND sg13g2_decap_8
XFILLER_6_4 VPWR VGND sg13g2_fill_2
XFILLER_3_969 VPWR VGND sg13g2_decap_8
XFILLER_2_457 VPWR VGND sg13g2_decap_8
XFILLER_19_804 VPWR VGND sg13g2_decap_4
XFILLER_46_678 VPWR VGND sg13g2_decap_8
XFILLER_41_350 VPWR VGND sg13g2_decap_8
XFILLER_42_895 VPWR VGND sg13g2_decap_8
XFILLER_6_741 VPWR VGND sg13g2_decap_8
X_2450_ _0354_ net490 net431 VPWR VGND sg13g2_nand2_1
X_2381_ VGND VPWR _0229_ _0259_ _0291_ _0261_ sg13g2_a21oi_1
XFILLER_39_4 VPWR VGND sg13g2_fill_2
XFILLER_49_472 VPWR VGND sg13g2_decap_8
Xinput5 ui_in[4] net5 VPWR VGND sg13g2_buf_1
X_3002_ net386 _0130_ VPWR VGND sg13g2_buf_1
XFILLER_37_612 VPWR VGND sg13g2_fill_1
XFILLER_37_623 VPWR VGND sg13g2_fill_1
XFILLER_36_111 VPWR VGND sg13g2_fill_2
XFILLER_37_667 VPWR VGND sg13g2_decap_8
XFILLER_18_881 VPWR VGND sg13g2_decap_8
XFILLER_24_339 VPWR VGND sg13g2_fill_1
X_2717_ VPWR _0614_ _0613_ VGND sg13g2_inv_1
X_2648_ _0546_ net487 net424 VPWR VGND sg13g2_nand2_1
X_2579_ VGND VPWR _0475_ _0476_ _0479_ _0457_ sg13g2_a21oi_1
XFILLER_47_409 VPWR VGND sg13g2_decap_8
XFILLER_27_133 VPWR VGND sg13g2_fill_2
XFILLER_15_339 VPWR VGND sg13g2_decap_8
XFILLER_42_147 VPWR VGND sg13g2_decap_8
XFILLER_24_851 VPWR VGND sg13g2_decap_8
XFILLER_13_1023 VPWR VGND sg13g2_decap_4
XFILLER_3_766 VPWR VGND sg13g2_decap_8
XFILLER_18_100 VPWR VGND sg13g2_fill_2
XFILLER_19_623 VPWR VGND sg13g2_fill_2
XFILLER_47_976 VPWR VGND sg13g2_decap_8
XFILLER_20_1016 VPWR VGND sg13g2_decap_8
XFILLER_20_1027 VPWR VGND sg13g2_fill_2
XFILLER_15_851 VPWR VGND sg13g2_decap_8
XFILLER_42_692 VPWR VGND sg13g2_decap_8
XFILLER_14_361 VPWR VGND sg13g2_decap_8
X_1950_ _1261_ _1258_ _1260_ VPWR VGND sg13g2_nand2_1
XFILLER_30_843 VPWR VGND sg13g2_decap_8
X_1881_ _1205_ net402 net499 VPWR VGND sg13g2_nand2_1
X_2502_ _0402_ _0401_ _0392_ _0404_ VPWR VGND sg13g2_a21o_1
X_2433_ _0340_ _0337_ _0339_ VPWR VGND sg13g2_xnor2_1
X_2364_ VGND VPWR _0274_ _0272_ _0247_ sg13g2_or2_1
X_2295_ _0207_ _0166_ _0205_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_910 VPWR VGND sg13g2_decap_8
XFILLER_49_291 VPWR VGND sg13g2_decap_8
XFILLER_38_987 VPWR VGND sg13g2_decap_8
XFILLER_24_169 VPWR VGND sg13g2_decap_8
XFILLER_36_1012 VPWR VGND sg13g2_decap_8
XFILLER_33_670 VPWR VGND sg13g2_decap_4
XFILLER_21_854 VPWR VGND sg13g2_fill_1
XFILLER_20_353 VPWR VGND sg13g2_fill_2
XFILLER_4_519 VPWR VGND sg13g2_decap_8
XFILLER_43_1027 VPWR VGND sg13g2_fill_2
XFILLER_0_769 VPWR VGND sg13g2_decap_8
XFILLER_46_44 VPWR VGND sg13g2_decap_8
XFILLER_29_976 VPWR VGND sg13g2_decap_8
XFILLER_44_957 VPWR VGND sg13g2_decap_8
XFILLER_43_423 VPWR VGND sg13g2_decap_8
XFILLER_15_125 VPWR VGND sg13g2_decap_8
XFILLER_15_147 VPWR VGND sg13g2_fill_1
XFILLER_12_821 VPWR VGND sg13g2_decap_8
XFILLER_30_128 VPWR VGND sg13g2_decap_8
XFILLER_11_320 VPWR VGND sg13g2_decap_8
XFILLER_7_313 VPWR VGND sg13g2_decap_8
XFILLER_7_16 VPWR VGND sg13g2_decap_8
XFILLER_12_898 VPWR VGND sg13g2_decap_8
XFILLER_8_858 VPWR VGND sg13g2_decap_8
XFILLER_3_563 VPWR VGND sg13g2_decap_8
XFILLER_39_707 VPWR VGND sg13g2_decap_4
XFILLER_38_206 VPWR VGND sg13g2_decap_8
X_2080_ VPWR _1365_ _1364_ VGND sg13g2_inv_1
XFILLER_19_442 VPWR VGND sg13g2_decap_8
XFILLER_46_283 VPWR VGND sg13g2_decap_8
XFILLER_35_957 VPWR VGND sg13g2_decap_8
X_2982_ net457 _0102_ VPWR VGND sg13g2_buf_1
X_1933_ net304 mac1.sum_lvl2_ff\[26\] _1247_ VPWR VGND sg13g2_xor2_1
XFILLER_21_128 VPWR VGND sg13g2_fill_2
XFILLER_30_662 VPWR VGND sg13g2_fill_2
X_1864_ _1162_ _1188_ _1189_ VPWR VGND sg13g2_nor2_1
X_1795_ _1121_ _1118_ _1122_ VPWR VGND sg13g2_xor2_1
X_2416_ _0324_ net497 net383 VPWR VGND sg13g2_nand2_1
X_2347_ _0256_ _0235_ _0258_ VPWR VGND sg13g2_xor2_1
X_2278_ _0190_ _0173_ _0191_ VPWR VGND sg13g2_xor2_1
XFILLER_44_209 VPWR VGND sg13g2_decap_8
XFILLER_26_902 VPWR VGND sg13g2_decap_8
XFILLER_37_250 VPWR VGND sg13g2_decap_8
XFILLER_37_294 VPWR VGND sg13g2_fill_1
XFILLER_26_979 VPWR VGND sg13g2_decap_8
XFILLER_41_927 VPWR VGND sg13g2_decap_8
XFILLER_12_139 VPWR VGND sg13g2_decap_8
XFILLER_5_839 VPWR VGND sg13g2_decap_8
XFILLER_48_515 VPWR VGND sg13g2_fill_2
XFILLER_0_566 VPWR VGND sg13g2_decap_8
XFILLER_17_935 VPWR VGND sg13g2_decap_8
XFILLER_28_272 VPWR VGND sg13g2_decap_8
XFILLER_43_231 VPWR VGND sg13g2_fill_2
XFILLER_43_220 VPWR VGND sg13g2_fill_1
XFILLER_25_990 VPWR VGND sg13g2_decap_8
XFILLER_32_927 VPWR VGND sg13g2_decap_8
XFILLER_40_960 VPWR VGND sg13g2_decap_8
X_1580_ _0913_ _0883_ _0911_ VPWR VGND sg13g2_xnor2_1
XFILLER_4_861 VPWR VGND sg13g2_decap_8
X_3250_ net504 VGND VPWR net183 net18 clknet_leaf_31_clk sg13g2_dfrbpq_2
XFILLER_26_1000 VPWR VGND sg13g2_decap_8
XFILLER_39_504 VPWR VGND sg13g2_decap_8
X_3181_ net509 VGND VPWR net139 mac1.sum_lvl2_ff\[42\] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_2201_ _1482_ net458 net502 VPWR VGND sg13g2_nand2_1
X_2132_ _1415_ net455 net384 VPWR VGND sg13g2_nand2_1
X_2063_ VGND VPWR _1349_ _1344_ _1342_ sg13g2_or2_1
XFILLER_23_905 VPWR VGND sg13g2_decap_8
XFILLER_34_253 VPWR VGND sg13g2_decap_4
XFILLER_34_264 VPWR VGND sg13g2_decap_4
XFILLER_35_798 VPWR VGND sg13g2_decap_8
XFILLER_22_437 VPWR VGND sg13g2_decap_8
X_2965_ _0839_ net426 net375 _0115_ VPWR VGND sg13g2_mux2_1
XFILLER_31_971 VPWR VGND sg13g2_decap_8
XFILLER_33_1015 VPWR VGND sg13g2_decap_8
X_2896_ net402 net423 net378 _0785_ VPWR VGND sg13g2_mux2_1
X_1916_ _1234_ mac1.sum_lvl2_ff\[22\] net243 VPWR VGND sg13g2_xnor2_1
XFILLER_8_70 VPWR VGND sg13g2_fill_2
X_1847_ _1112_ _1172_ _1173_ VPWR VGND sg13g2_nor2b_1
X_1778_ _1106_ _1105_ _1078_ VPWR VGND sg13g2_nand2b_1
XFILLER_27_46 VPWR VGND sg13g2_decap_8
XFILLER_27_57 VPWR VGND sg13g2_fill_1
XFILLER_38_570 VPWR VGND sg13g2_decap_8
XFILLER_14_905 VPWR VGND sg13g2_decap_8
XFILLER_25_231 VPWR VGND sg13g2_decap_8
XFILLER_25_242 VPWR VGND sg13g2_fill_2
XFILLER_26_765 VPWR VGND sg13g2_decap_4
XFILLER_41_724 VPWR VGND sg13g2_decap_8
XFILLER_41_713 VPWR VGND sg13g2_fill_2
XFILLER_25_253 VPWR VGND sg13g2_decap_8
XFILLER_25_264 VPWR VGND sg13g2_fill_2
XFILLER_13_426 VPWR VGND sg13g2_decap_8
XFILLER_21_470 VPWR VGND sg13g2_fill_2
XFILLER_49_1000 VPWR VGND sg13g2_decap_8
XFILLER_1_842 VPWR VGND sg13g2_decap_8
XFILLER_49_846 VPWR VGND sg13g2_decap_8
XFILLER_36_518 VPWR VGND sg13g2_decap_8
XFILLER_1_1024 VPWR VGND sg13g2_decap_4
XFILLER_17_710 VPWR VGND sg13g2_decap_8
XFILLER_17_721 VPWR VGND sg13g2_fill_1
XFILLER_36_529 VPWR VGND sg13g2_fill_2
XFILLER_44_540 VPWR VGND sg13g2_decap_8
XFILLER_16_242 VPWR VGND sg13g2_fill_2
XFILLER_44_584 VPWR VGND sg13g2_decap_4
XFILLER_13_960 VPWR VGND sg13g2_decap_8
XFILLER_31_245 VPWR VGND sg13g2_decap_8
X_2750_ _0609_ _0615_ _0646_ VPWR VGND sg13g2_nor2_1
XFILLER_9_942 VPWR VGND sg13g2_decap_8
X_1701_ _0982_ VPWR _1031_ VGND _0918_ _0983_ sg13g2_o21ai_1
X_2681_ _0068_ _0538_ _0577_ VPWR VGND sg13g2_xnor2_1
X_1632_ _0963_ _0957_ _0962_ VPWR VGND sg13g2_xnor2_1
X_1563_ _0896_ net410 net468 VPWR VGND sg13g2_nand2_1
Xfanout409 DP_2.matrix\[39\] net409 VPWR VGND sg13g2_buf_1
X_3233_ net521 VGND VPWR net285 mac1.sum_lvl3_ff\[8\] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_3164_ net526 VGND VPWR net104 mac1.sum_lvl2_ff\[22\] clknet_leaf_27_clk sg13g2_dfrbpq_1
XFILLER_39_356 VPWR VGND sg13g2_decap_8
X_2115_ _1388_ _1396_ _1398_ _1399_ VPWR VGND sg13g2_or3_1
X_3095_ net546 VGND VPWR _0074_ mac1.products_ff\[82\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_2046_ _0021_ _1333_ net187 VPWR VGND sg13g2_xnor2_1
XFILLER_23_735 VPWR VGND sg13g2_decap_8
XFILLER_23_746 VPWR VGND sg13g2_fill_2
XFILLER_11_919 VPWR VGND sg13g2_decap_8
X_2948_ _0829_ net478 net371 VPWR VGND sg13g2_nand2b_1
XFILLER_10_418 VPWR VGND sg13g2_decap_8
XFILLER_13_37 VPWR VGND sg13g2_decap_4
X_2879_ DP_1.I_range.out_data\[2\] DP_1.I_range.out_data\[4\] DP_1.Q_range.out_data\[2\]
+ _0768_ _0769_ VPWR VGND sg13g2_nor4_1
XFILLER_49_109 VPWR VGND sg13g2_decap_8
XFILLER_46_827 VPWR VGND sg13g2_decap_8
XFILLER_39_890 VPWR VGND sg13g2_decap_8
XFILLER_14_724 VPWR VGND sg13g2_fill_2
XFILLER_26_551 VPWR VGND sg13g2_fill_1
XFILLER_13_201 VPWR VGND sg13g2_decap_4
XFILLER_41_565 VPWR VGND sg13g2_decap_8
XFILLER_9_205 VPWR VGND sg13g2_decap_8
XFILLER_10_985 VPWR VGND sg13g2_decap_8
XFILLER_6_923 VPWR VGND sg13g2_decap_8
XFILLER_49_643 VPWR VGND sg13g2_decap_8
XFILLER_23_1003 VPWR VGND sg13g2_decap_8
XFILLER_17_540 VPWR VGND sg13g2_fill_2
XFILLER_36_337 VPWR VGND sg13g2_fill_2
XFILLER_45_893 VPWR VGND sg13g2_decap_8
XFILLER_17_595 VPWR VGND sg13g2_decap_8
XFILLER_32_565 VPWR VGND sg13g2_decap_8
X_2802_ _0694_ _0695_ _0696_ VPWR VGND sg13g2_and2_1
X_2733_ VGND VPWR _0629_ _0598_ _0596_ sg13g2_or2_1
XFILLER_30_1018 VPWR VGND sg13g2_decap_8
X_2664_ net476 net501 net435 net432 _0562_ VPWR VGND sg13g2_and4_1
X_2595_ _0494_ net489 net421 VPWR VGND sg13g2_nand2_1
X_1615_ _0947_ _0912_ _0946_ VPWR VGND sg13g2_xnor2_1
X_1546_ _0879_ _0869_ _0880_ VPWR VGND sg13g2_xor2_1
XFILLER_8_1019 VPWR VGND sg13g2_decap_8
X_3216_ net511 VGND VPWR net124 mac1.sum_lvl3_ff\[27\] clknet_leaf_31_clk sg13g2_dfrbpq_1
XFILLER_39_131 VPWR VGND sg13g2_decap_4
X_3147_ net525 VGND VPWR net49 mac1.sum_lvl2_ff\[2\] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_3078_ net538 VGND VPWR _0131_ DP_2.matrix\[77\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_42_318 VPWR VGND sg13g2_decap_8
X_2029_ _0018_ _1321_ net208 VPWR VGND sg13g2_xnor2_1
XFILLER_23_521 VPWR VGND sg13g2_fill_2
XFILLER_36_893 VPWR VGND sg13g2_decap_8
XFILLER_24_47 VPWR VGND sg13g2_fill_1
XFILLER_10_248 VPWR VGND sg13g2_decap_8
XFILLER_40_68 VPWR VGND sg13g2_decap_4
Xhold260 DP_2.matrix\[6\] VPWR VGND net300 sg13g2_dlygate4sd3_1
XFILLER_3_948 VPWR VGND sg13g2_decap_8
XFILLER_49_88 VPWR VGND sg13g2_decap_8
XFILLER_46_635 VPWR VGND sg13g2_decap_8
XFILLER_46_657 VPWR VGND sg13g2_decap_8
XFILLER_45_123 VPWR VGND sg13g2_decap_4
XFILLER_34_808 VPWR VGND sg13g2_decap_8
XFILLER_45_156 VPWR VGND sg13g2_decap_4
XFILLER_42_874 VPWR VGND sg13g2_decap_8
XFILLER_14_565 VPWR VGND sg13g2_decap_8
XFILLER_14_80 VPWR VGND sg13g2_decap_8
XFILLER_6_720 VPWR VGND sg13g2_decap_8
XFILLER_10_782 VPWR VGND sg13g2_decap_8
XFILLER_6_797 VPWR VGND sg13g2_decap_8
XFILLER_5_296 VPWR VGND sg13g2_decap_8
X_2380_ _0288_ _0287_ _0290_ VPWR VGND sg13g2_xor2_1
XFILLER_49_451 VPWR VGND sg13g2_decap_8
Xinput6 ui_in[5] net6 VPWR VGND sg13g2_buf_1
X_3001_ net388 _0129_ VPWR VGND sg13g2_buf_1
XFILLER_37_602 VPWR VGND sg13g2_fill_2
XFILLER_24_318 VPWR VGND sg13g2_decap_8
XFILLER_17_381 VPWR VGND sg13g2_decap_8
XFILLER_20_502 VPWR VGND sg13g2_decap_8
XFILLER_33_896 VPWR VGND sg13g2_decap_8
XFILLER_32_395 VPWR VGND sg13g2_decap_8
XFILLER_20_579 VPWR VGND sg13g2_decap_8
X_2716_ VGND VPWR _0533_ _0576_ _0613_ _0575_ sg13g2_a21oi_1
X_2647_ _0545_ net487 net421 VPWR VGND sg13g2_nand2_1
XFILLER_10_27 VPWR VGND sg13g2_fill_1
X_2578_ _0475_ _0476_ _0457_ _0478_ VPWR VGND sg13g2_nand3_1
X_1529_ _0864_ _0853_ _0862_ VPWR VGND sg13g2_xnor2_1
XFILLER_27_112 VPWR VGND sg13g2_decap_8
XFILLER_42_126 VPWR VGND sg13g2_decap_8
XFILLER_24_830 VPWR VGND sg13g2_decap_8
Xclkbuf_3_3__f_clk clknet_0_clk clknet_3_3__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_13_1002 VPWR VGND sg13g2_decap_8
XFILLER_3_745 VPWR VGND sg13g2_decap_8
XFILLER_2_211 VPWR VGND sg13g2_decap_8
XFILLER_2_266 VPWR VGND sg13g2_decap_4
XFILLER_47_955 VPWR VGND sg13g2_decap_8
XFILLER_18_156 VPWR VGND sg13g2_decap_4
XFILLER_33_104 VPWR VGND sg13g2_decap_8
XFILLER_34_638 VPWR VGND sg13g2_decap_8
XFILLER_33_148 VPWR VGND sg13g2_decap_4
XFILLER_30_822 VPWR VGND sg13g2_decap_8
X_1880_ _1204_ net462 net494 VPWR VGND sg13g2_nand2_1
XFILLER_30_899 VPWR VGND sg13g2_decap_8
X_2501_ _0401_ _0402_ _0392_ _0403_ VPWR VGND sg13g2_nand3_1
XFILLER_6_583 VPWR VGND sg13g2_fill_1
X_2432_ _0339_ _0323_ _0338_ VPWR VGND sg13g2_xnor2_1
X_2363_ _0247_ _0272_ _0273_ VPWR VGND sg13g2_nor2_1
XFILLER_2_61 VPWR VGND sg13g2_decap_4
X_2294_ VGND VPWR _0206_ _0204_ _0167_ sg13g2_or2_1
XFILLER_49_270 VPWR VGND sg13g2_decap_8
XFILLER_38_966 VPWR VGND sg13g2_decap_8
XFILLER_25_627 VPWR VGND sg13g2_fill_1
XFILLER_21_833 VPWR VGND sg13g2_decap_8
XFILLER_43_1006 VPWR VGND sg13g2_decap_8
XFILLER_0_748 VPWR VGND sg13g2_decap_8
XFILLER_29_955 VPWR VGND sg13g2_decap_8
XFILLER_44_936 VPWR VGND sg13g2_decap_8
XFILLER_15_104 VPWR VGND sg13g2_decap_8
XFILLER_12_800 VPWR VGND sg13g2_decap_8
XFILLER_8_837 VPWR VGND sg13g2_decap_8
XFILLER_11_343 VPWR VGND sg13g2_decap_8
XFILLER_12_877 VPWR VGND sg13g2_decap_8
XFILLER_3_553 VPWR VGND sg13g2_fill_1
XFILLER_3_542 VPWR VGND sg13g2_decap_8
XFILLER_47_730 VPWR VGND sg13g2_decap_8
XFILLER_4_1022 VPWR VGND sg13g2_decap_8
XFILLER_19_454 VPWR VGND sg13g2_decap_8
XFILLER_35_936 VPWR VGND sg13g2_decap_8
XFILLER_22_619 VPWR VGND sg13g2_decap_4
X_2981_ net459 _0101_ VPWR VGND sg13g2_buf_1
XFILLER_34_479 VPWR VGND sg13g2_decap_8
X_1932_ _1246_ net283 mac1.sum_lvl2_ff\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_30_641 VPWR VGND sg13g2_decap_8
X_1863_ _1188_ _1147_ _1186_ VPWR VGND sg13g2_xnor2_1
X_1794_ _1121_ _1094_ _1119_ VPWR VGND sg13g2_xnor2_1
X_2415_ _0323_ net497 net381 VPWR VGND sg13g2_nand2_1
X_2346_ _0256_ _0235_ _0257_ VPWR VGND sg13g2_nor2b_1
X_2277_ _0190_ _0174_ _0188_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_958 VPWR VGND sg13g2_decap_8
XFILLER_41_906 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_32_clk clknet_3_1__leaf_clk clknet_leaf_32_clk VPWR VGND sg13g2_buf_8
XFILLER_33_490 VPWR VGND sg13g2_decap_8
XFILLER_21_685 VPWR VGND sg13g2_decap_4
XFILLER_5_818 VPWR VGND sg13g2_decap_8
XFILLER_20_195 VPWR VGND sg13g2_decap_8
XFILLER_10_1027 VPWR VGND sg13g2_fill_2
XFILLER_0_545 VPWR VGND sg13g2_decap_8
XFILLER_17_914 VPWR VGND sg13g2_decap_8
XFILLER_29_741 VPWR VGND sg13g2_decap_8
XFILLER_28_251 VPWR VGND sg13g2_decap_8
XFILLER_16_446 VPWR VGND sg13g2_fill_2
XFILLER_32_906 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_23_clk clknet_3_5__leaf_clk clknet_leaf_23_clk VPWR VGND sg13g2_buf_8
XFILLER_7_166 VPWR VGND sg13g2_decap_4
XFILLER_11_184 VPWR VGND sg13g2_decap_8
XFILLER_7_199 VPWR VGND sg13g2_decap_8
XFILLER_4_840 VPWR VGND sg13g2_decap_8
XFILLER_3_383 VPWR VGND sg13g2_decap_4
X_2200_ _1452_ VPWR _1481_ VGND _1449_ _1453_ sg13g2_o21ai_1
X_3180_ net506 VGND VPWR net126 mac1.sum_lvl2_ff\[41\] clknet_leaf_36_clk sg13g2_dfrbpq_1
XFILLER_14_4 VPWR VGND sg13g2_decap_4
X_2131_ _1397_ VPWR _1414_ VGND _1388_ _1398_ sg13g2_o21ai_1
X_2062_ _1348_ net457 net388 VPWR VGND sg13g2_nand2_1
XFILLER_47_582 VPWR VGND sg13g2_decap_8
XFILLER_35_711 VPWR VGND sg13g2_fill_1
XFILLER_34_232 VPWR VGND sg13g2_decap_8
XFILLER_34_276 VPWR VGND sg13g2_decap_4
XFILLER_35_777 VPWR VGND sg13g2_decap_8
X_2964_ _0804_ _0788_ _0839_ VPWR VGND sg13g2_xor2_1
X_1915_ _1233_ mac1.sum_lvl2_ff\[22\] net243 VPWR VGND sg13g2_nand2_1
XFILLER_31_950 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_14_clk clknet_3_6__leaf_clk clknet_leaf_14_clk VPWR VGND sg13g2_buf_8
X_2895_ _0784_ _0780_ _0782_ VPWR VGND sg13g2_xnor2_1
XFILLER_8_93 VPWR VGND sg13g2_decap_8
X_1846_ VGND VPWR _1108_ _1140_ _1172_ _1141_ sg13g2_a21oi_1
XFILLER_30_493 VPWR VGND sg13g2_decap_8
X_1777_ _1103_ _1079_ _1105_ VPWR VGND sg13g2_xor2_1
XFILLER_1_309 VPWR VGND sg13g2_decap_8
XFILLER_40_1009 VPWR VGND sg13g2_decap_8
X_2329_ VGND VPWR _0240_ _0239_ _0215_ sg13g2_or2_1
XFILLER_45_508 VPWR VGND sg13g2_decap_8
XFILLER_27_25 VPWR VGND sg13g2_decap_4
XFILLER_38_560 VPWR VGND sg13g2_fill_1
XFILLER_25_210 VPWR VGND sg13g2_decap_8
XFILLER_25_287 VPWR VGND sg13g2_decap_8
XFILLER_43_79 VPWR VGND sg13g2_decap_8
XFILLER_41_769 VPWR VGND sg13g2_decap_8
XFILLER_22_994 VPWR VGND sg13g2_decap_8
XFILLER_1_821 VPWR VGND sg13g2_decap_8
XFILLER_49_825 VPWR VGND sg13g2_decap_8
XFILLER_0_342 VPWR VGND sg13g2_decap_8
XFILLER_1_898 VPWR VGND sg13g2_decap_8
XFILLER_1_1003 VPWR VGND sg13g2_decap_8
XFILLER_29_560 VPWR VGND sg13g2_decap_8
XFILLER_17_744 VPWR VGND sg13g2_decap_8
XFILLER_44_563 VPWR VGND sg13g2_decap_8
XFILLER_17_91 VPWR VGND sg13g2_decap_8
XFILLER_44_596 VPWR VGND sg13g2_fill_2
XFILLER_9_921 VPWR VGND sg13g2_decap_8
XFILLER_31_257 VPWR VGND sg13g2_fill_2
XFILLER_31_279 VPWR VGND sg13g2_fill_2
XFILLER_12_493 VPWR VGND sg13g2_decap_8
X_1700_ _0954_ VPWR _1030_ VGND _1026_ _1028_ sg13g2_o21ai_1
XFILLER_33_90 VPWR VGND sg13g2_decap_8
X_2680_ VPWR _0578_ _0577_ VGND sg13g2_inv_1
XFILLER_9_998 VPWR VGND sg13g2_decap_8
X_1631_ _0962_ _0923_ _0959_ VPWR VGND sg13g2_xnor2_1
X_1562_ _0873_ VPWR _0895_ VGND _0871_ _0874_ sg13g2_o21ai_1
X_3232_ net521 VGND VPWR _0013_ mac1.sum_lvl3_ff\[7\] clknet_leaf_32_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_3_clk clknet_3_3__leaf_clk clknet_leaf_3_clk VPWR VGND sg13g2_buf_8
X_3163_ net525 VGND VPWR net105 mac1.sum_lvl2_ff\[21\] clknet_leaf_27_clk sg13g2_dfrbpq_1
XFILLER_39_335 VPWR VGND sg13g2_decap_8
X_2114_ VGND VPWR _1394_ _1395_ _1398_ _1389_ sg13g2_a21oi_1
XFILLER_48_891 VPWR VGND sg13g2_decap_8
XFILLER_27_519 VPWR VGND sg13g2_fill_1
X_3094_ net541 VGND VPWR _0073_ mac1.products_ff\[81\] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_2045_ net186 mac1.sum_lvl3_ff\[14\] _1336_ VPWR VGND sg13g2_xor2_1
XFILLER_35_563 VPWR VGND sg13g2_fill_1
XFILLER_22_202 VPWR VGND sg13g2_decap_8
X_2947_ VGND VPWR net371 _0827_ _0092_ _0828_ sg13g2_a21oi_1
X_2878_ _0768_ DP_1.I_range.out_data\[5\] _0767_ VPWR VGND sg13g2_nand2_1
X_1829_ VGND VPWR _1155_ _1153_ _1129_ sg13g2_or2_1
XFILLER_2_629 VPWR VGND sg13g2_decap_8
XFILLER_45_338 VPWR VGND sg13g2_decap_8
XFILLER_14_703 VPWR VGND sg13g2_decap_8
XFILLER_26_563 VPWR VGND sg13g2_fill_1
XFILLER_10_964 VPWR VGND sg13g2_decap_8
XFILLER_6_902 VPWR VGND sg13g2_decap_8
XFILLER_6_979 VPWR VGND sg13g2_decap_8
XFILLER_49_633 VPWR VGND sg13g2_fill_2
XFILLER_1_695 VPWR VGND sg13g2_decap_8
XFILLER_0_183 VPWR VGND sg13g2_decap_8
XFILLER_36_316 VPWR VGND sg13g2_decap_8
XFILLER_36_349 VPWR VGND sg13g2_fill_1
XFILLER_45_872 VPWR VGND sg13g2_decap_8
XFILLER_17_563 VPWR VGND sg13g2_decap_8
X_2801_ _0667_ _0669_ _0693_ _0695_ VPWR VGND sg13g2_or3_1
X_2732_ _0586_ VPWR _0628_ VGND _0583_ _0587_ sg13g2_o21ai_1
XFILLER_9_795 VPWR VGND sg13g2_decap_8
X_2663_ _0561_ net501 net432 VPWR VGND sg13g2_nand2_1
X_1614_ _0946_ _0915_ _0944_ VPWR VGND sg13g2_xnor2_1
X_2594_ _0493_ net493 net495 VPWR VGND sg13g2_nand2_1
X_1545_ _0879_ _0878_ _0877_ VPWR VGND sg13g2_nand2b_1
X_3215_ net510 VGND VPWR net138 mac1.sum_lvl3_ff\[26\] clknet_leaf_35_clk sg13g2_dfrbpq_1
XFILLER_39_110 VPWR VGND sg13g2_decap_8
XFILLER_28_806 VPWR VGND sg13g2_decap_4
X_3146_ net520 VGND VPWR net145 mac1.sum_lvl2_ff\[1\] clknet_leaf_33_clk sg13g2_dfrbpq_1
XFILLER_43_809 VPWR VGND sg13g2_fill_1
XFILLER_27_338 VPWR VGND sg13g2_decap_4
X_3077_ net519 VGND VPWR _0130_ DP_2.matrix\[76\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2028_ _1322_ net207 _1318_ VPWR VGND sg13g2_nand2_1
XFILLER_36_872 VPWR VGND sg13g2_decap_8
XFILLER_35_371 VPWR VGND sg13g2_decap_4
XFILLER_23_566 VPWR VGND sg13g2_fill_2
XFILLER_35_393 VPWR VGND sg13g2_decap_8
XFILLER_11_717 VPWR VGND sg13g2_decap_8
XFILLER_3_927 VPWR VGND sg13g2_decap_8
Xhold261 mac1.sum_lvl2_ff\[29\] VPWR VGND net301 sg13g2_dlygate4sd3_1
Xhold250 DP_2.matrix\[72\] VPWR VGND net290 sg13g2_dlygate4sd3_1
XFILLER_49_56 VPWR VGND sg13g2_decap_4
XFILLER_45_102 VPWR VGND sg13g2_decap_8
XFILLER_18_305 VPWR VGND sg13g2_decap_8
XFILLER_27_883 VPWR VGND sg13g2_decap_8
XFILLER_42_853 VPWR VGND sg13g2_decap_8
XFILLER_14_544 VPWR VGND sg13g2_fill_2
XFILLER_10_761 VPWR VGND sg13g2_decap_8
XFILLER_6_776 VPWR VGND sg13g2_decap_8
XFILLER_2_993 VPWR VGND sg13g2_decap_8
X_3000_ net391 _0128_ VPWR VGND sg13g2_buf_1
Xinput7 ui_in[6] net7 VPWR VGND sg13g2_buf_1
XFILLER_36_113 VPWR VGND sg13g2_fill_1
XFILLER_36_135 VPWR VGND sg13g2_decap_4
XFILLER_37_647 VPWR VGND sg13g2_decap_8
XFILLER_17_360 VPWR VGND sg13g2_decap_8
XFILLER_33_875 VPWR VGND sg13g2_decap_8
XFILLER_20_558 VPWR VGND sg13g2_decap_8
XFILLER_9_592 VPWR VGND sg13g2_decap_8
X_2715_ _0536_ _0578_ _0535_ _0612_ VPWR VGND sg13g2_nand3_1
X_2646_ _0544_ net491 net495 VPWR VGND sg13g2_nand2_1
X_2577_ _0477_ _0457_ _0475_ _0476_ VPWR VGND sg13g2_and3_1
X_1528_ _0863_ _0862_ _0853_ VPWR VGND sg13g2_nand2b_1
XFILLER_28_614 VPWR VGND sg13g2_decap_8
XFILLER_27_102 VPWR VGND sg13g2_fill_2
XFILLER_43_617 VPWR VGND sg13g2_decap_8
X_3129_ net521 VGND VPWR net137 mac1.sum_lvl1_ff\[36\] clknet_leaf_34_clk sg13g2_dfrbpq_1
XFILLER_35_47 VPWR VGND sg13g2_decap_8
XFILLER_11_525 VPWR VGND sg13g2_fill_2
XFILLER_23_385 VPWR VGND sg13g2_decap_8
XFILLER_7_507 VPWR VGND sg13g2_fill_1
XFILLER_3_724 VPWR VGND sg13g2_decap_8
XFILLER_47_934 VPWR VGND sg13g2_decap_8
XFILLER_19_636 VPWR VGND sg13g2_fill_1
XFILLER_46_455 VPWR VGND sg13g2_fill_1
XFILLER_18_135 VPWR VGND sg13g2_fill_2
XFILLER_26_190 VPWR VGND sg13g2_decap_8
XFILLER_15_886 VPWR VGND sg13g2_decap_8
XFILLER_30_812 VPWR VGND sg13g2_fill_1
XFILLER_30_878 VPWR VGND sg13g2_decap_8
X_2500_ _0399_ _0398_ _0393_ _0402_ VPWR VGND sg13g2_a21o_1
X_2431_ _0338_ net441 net502 VPWR VGND sg13g2_nand2_1
X_2362_ _0272_ net443 net380 VPWR VGND sg13g2_nand2_2
XFILLER_2_790 VPWR VGND sg13g2_decap_8
X_2293_ _0205_ net448 net382 VPWR VGND sg13g2_nand2_1
XFILLER_38_945 VPWR VGND sg13g2_decap_8
XFILLER_37_455 VPWR VGND sg13g2_decap_8
XFILLER_18_680 VPWR VGND sg13g2_decap_8
XFILLER_24_105 VPWR VGND sg13g2_decap_8
XFILLER_24_116 VPWR VGND sg13g2_fill_2
XFILLER_37_499 VPWR VGND sg13g2_decap_8
XFILLER_24_138 VPWR VGND sg13g2_decap_8
XFILLER_21_812 VPWR VGND sg13g2_fill_1
XFILLER_32_182 VPWR VGND sg13g2_decap_8
XFILLER_21_889 VPWR VGND sg13g2_decap_8
XFILLER_20_399 VPWR VGND sg13g2_decap_8
X_2629_ _0525_ _0526_ _0491_ _0528_ VPWR VGND sg13g2_nand3_1
XFILLER_0_727 VPWR VGND sg13g2_decap_8
XFILLER_28_400 VPWR VGND sg13g2_decap_8
XFILLER_28_411 VPWR VGND sg13g2_fill_1
XFILLER_29_934 VPWR VGND sg13g2_decap_8
XFILLER_44_915 VPWR VGND sg13g2_decap_8
XFILLER_43_469 VPWR VGND sg13g2_decap_8
XFILLER_24_650 VPWR VGND sg13g2_decap_4
XFILLER_30_108 VPWR VGND sg13g2_decap_8
XFILLER_12_856 VPWR VGND sg13g2_decap_8
XFILLER_23_160 VPWR VGND sg13g2_fill_1
XFILLER_8_816 VPWR VGND sg13g2_decap_8
XFILLER_3_521 VPWR VGND sg13g2_decap_8
XFILLER_3_598 VPWR VGND sg13g2_decap_8
XFILLER_4_1001 VPWR VGND sg13g2_decap_8
Xfanout390 net391 net390 VPWR VGND sg13g2_buf_8
XFILLER_35_915 VPWR VGND sg13g2_decap_8
XFILLER_34_436 VPWR VGND sg13g2_fill_2
XFILLER_34_458 VPWR VGND sg13g2_decap_8
XFILLER_36_90 VPWR VGND sg13g2_decap_8
X_2980_ net463 _0100_ VPWR VGND sg13g2_buf_1
XFILLER_43_992 VPWR VGND sg13g2_decap_8
X_1931_ _1244_ net298 _0012_ VPWR VGND sg13g2_nor2b_2
XFILLER_15_694 VPWR VGND sg13g2_decap_8
XFILLER_30_664 VPWR VGND sg13g2_fill_1
X_1862_ _1147_ _1186_ _1187_ VPWR VGND sg13g2_nor2_1
Xinput10 uio_in[1] net10 VPWR VGND sg13g2_buf_1
X_1793_ VGND VPWR _1120_ _1119_ _1094_ sg13g2_or2_1
XFILLER_7_882 VPWR VGND sg13g2_decap_8
X_2414_ _0322_ net443 DP_2.matrix\[80\] VPWR VGND sg13g2_nand2_1
XFILLER_35_0 VPWR VGND sg13g2_fill_2
X_2345_ _0256_ _0236_ _0255_ VPWR VGND sg13g2_xnor2_1
X_2276_ _0189_ _0174_ _0188_ VPWR VGND sg13g2_nand2_1
XFILLER_29_219 VPWR VGND sg13g2_decap_8
XFILLER_26_937 VPWR VGND sg13g2_decap_8
XFILLER_21_653 VPWR VGND sg13g2_decap_8
XFILLER_21_664 VPWR VGND sg13g2_fill_1
XFILLER_20_163 VPWR VGND sg13g2_decap_4
XFILLER_10_1006 VPWR VGND sg13g2_decap_8
XFILLER_0_524 VPWR VGND sg13g2_decap_8
XFILLER_28_230 VPWR VGND sg13g2_decap_8
XFILLER_29_797 VPWR VGND sg13g2_decap_8
XFILLER_44_767 VPWR VGND sg13g2_decap_8
XFILLER_43_233 VPWR VGND sg13g2_fill_1
XFILLER_44_778 VPWR VGND sg13g2_fill_1
XFILLER_19_1020 VPWR VGND sg13g2_decap_8
XFILLER_8_602 VPWR VGND sg13g2_decap_8
XFILLER_40_995 VPWR VGND sg13g2_decap_8
XFILLER_8_646 VPWR VGND sg13g2_decap_8
XFILLER_22_70 VPWR VGND sg13g2_fill_1
XFILLER_4_896 VPWR VGND sg13g2_decap_8
XFILLER_3_362 VPWR VGND sg13g2_decap_8
XFILLER_3_351 VPWR VGND sg13g2_fill_2
XFILLER_39_539 VPWR VGND sg13g2_decap_8
X_2130_ _1411_ _1410_ _1413_ VPWR VGND sg13g2_xor2_1
X_2061_ _1346_ _1339_ _0034_ VPWR VGND sg13g2_xor2_1
XFILLER_47_561 VPWR VGND sg13g2_decap_8
XFILLER_19_263 VPWR VGND sg13g2_decap_8
XFILLER_19_296 VPWR VGND sg13g2_decap_8
XFILLER_34_222 VPWR VGND sg13g2_decap_4
X_2963_ _0838_ VPWR _0114_ VGND net375 _0837_ sg13g2_o21ai_1
XFILLER_16_981 VPWR VGND sg13g2_decap_8
XFILLER_34_288 VPWR VGND sg13g2_decap_4
X_1914_ VGND VPWR _1229_ _1231_ _1232_ _1230_ sg13g2_a21oi_1
X_2894_ net378 _0782_ _0783_ VPWR VGND sg13g2_and2_1
X_1845_ _1169_ _1168_ _1171_ VPWR VGND sg13g2_xor2_1
X_1776_ _1104_ _1079_ _1103_ VPWR VGND sg13g2_nand2_1
X_2328_ _0239_ net497 net389 VPWR VGND sg13g2_nand2_1
X_2259_ _0163_ _0171_ _0172_ VPWR VGND sg13g2_nor2_1
XFILLER_26_734 VPWR VGND sg13g2_decap_8
XFILLER_41_715 VPWR VGND sg13g2_fill_1
XFILLER_43_58 VPWR VGND sg13g2_decap_8
XFILLER_22_973 VPWR VGND sg13g2_decap_8
XFILLER_5_605 VPWR VGND sg13g2_decap_8
XFILLER_21_483 VPWR VGND sg13g2_decap_8
XFILLER_1_800 VPWR VGND sg13g2_decap_8
XFILLER_49_804 VPWR VGND sg13g2_decap_8
XFILLER_1_877 VPWR VGND sg13g2_decap_8
XFILLER_0_398 VPWR VGND sg13g2_decap_8
XFILLER_16_211 VPWR VGND sg13g2_decap_4
XFILLER_9_900 VPWR VGND sg13g2_decap_8
XFILLER_13_995 VPWR VGND sg13g2_decap_8
XFILLER_9_977 VPWR VGND sg13g2_decap_8
XFILLER_8_454 VPWR VGND sg13g2_fill_2
XFILLER_8_465 VPWR VGND sg13g2_decap_4
X_1630_ _0923_ _0959_ _0961_ VPWR VGND sg13g2_and2_1
X_1561_ _0894_ _0888_ _0893_ VPWR VGND sg13g2_xnor2_1
XFILLER_4_693 VPWR VGND sg13g2_decap_8
X_3231_ net510 VGND VPWR net299 mac1.sum_lvl3_ff\[6\] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_3162_ net520 VGND VPWR net64 mac1.sum_lvl2_ff\[20\] clknet_leaf_33_clk sg13g2_dfrbpq_1
XFILLER_39_314 VPWR VGND sg13g2_decap_8
X_2113_ _1394_ _1395_ _1389_ _1397_ VPWR VGND sg13g2_nand3_1
XFILLER_48_870 VPWR VGND sg13g2_decap_8
X_3093_ net541 VGND VPWR _0072_ mac1.products_ff\[80\] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_2044_ mac1.sum_lvl3_ff\[14\] mac1.sum_lvl3_ff\[34\] _1335_ VPWR VGND sg13g2_nor2_1
X_2946_ net160 net371 _0828_ VPWR VGND sg13g2_nor2_1
XFILLER_31_781 VPWR VGND sg13g2_decap_8
X_2877_ DP_1.I_range.out_data\[6\] DP_1.I_range.out_data\[3\] _0767_ VPWR VGND sg13g2_nor2_1
X_1828_ net465 net462 net403 net401 _1154_ VPWR VGND sg13g2_and4_1
XFILLER_2_608 VPWR VGND sg13g2_decap_8
X_1759_ _1086_ _1082_ _1087_ VPWR VGND sg13g2_xor2_1
XFILLER_38_47 VPWR VGND sg13g2_decap_8
XFILLER_38_58 VPWR VGND sg13g2_fill_2
XFILLER_26_542 VPWR VGND sg13g2_decap_8
XFILLER_41_534 VPWR VGND sg13g2_decap_8
XFILLER_41_512 VPWR VGND sg13g2_fill_2
XFILLER_14_726 VPWR VGND sg13g2_fill_1
XFILLER_26_575 VPWR VGND sg13g2_fill_2
XFILLER_13_247 VPWR VGND sg13g2_fill_1
XFILLER_16_1023 VPWR VGND sg13g2_decap_4
XFILLER_10_943 VPWR VGND sg13g2_decap_8
XFILLER_6_958 VPWR VGND sg13g2_decap_8
XFILLER_49_612 VPWR VGND sg13g2_decap_8
XFILLER_0_162 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_4
XFILLER_1_674 VPWR VGND sg13g2_decap_8
XFILLER_37_829 VPWR VGND sg13g2_fill_1
XFILLER_48_188 VPWR VGND sg13g2_decap_8
XFILLER_28_80 VPWR VGND sg13g2_decap_8
XFILLER_36_339 VPWR VGND sg13g2_fill_1
XFILLER_45_851 VPWR VGND sg13g2_decap_8
X_2800_ _0693_ VPWR _0694_ VGND _0667_ _0669_ sg13g2_o21ai_1
X_2731_ _0627_ _0619_ _0624_ VPWR VGND sg13g2_xnor2_1
XFILLER_9_774 VPWR VGND sg13g2_decap_8
X_2662_ _0513_ VPWR _0560_ VGND _0511_ _0514_ sg13g2_o21ai_1
X_1613_ _0944_ _0915_ _0945_ VPWR VGND sg13g2_nor2b_1
X_2593_ _0461_ VPWR _0492_ VGND _0458_ _0462_ sg13g2_o21ai_1
X_1544_ _0876_ _0875_ _0870_ _0878_ VPWR VGND sg13g2_a21o_1
X_3214_ net509 VGND VPWR net111 mac1.sum_lvl3_ff\[25\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_3145_ net520 VGND VPWR net118 mac1.sum_lvl2_ff\[0\] clknet_leaf_33_clk sg13g2_dfrbpq_1
XFILLER_39_144 VPWR VGND sg13g2_fill_1
X_3076_ net519 VGND VPWR _0129_ DP_2.matrix\[75\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_2027_ _1321_ _1320_ _1319_ VPWR VGND sg13g2_nand2b_1
XFILLER_39_1023 VPWR VGND sg13g2_decap_4
X_2929_ net373 net492 _0086_ VPWR VGND sg13g2_xor2_1
XFILLER_3_906 VPWR VGND sg13g2_decap_8
XFILLER_2_438 VPWR VGND sg13g2_decap_8
Xhold262 _1260_ VPWR VGND net302 sg13g2_dlygate4sd3_1
Xhold251 mac1.sum_lvl3_ff\[32\] VPWR VGND net291 sg13g2_dlygate4sd3_1
Xhold240 _1275_ VPWR VGND net280 sg13g2_dlygate4sd3_1
XFILLER_49_35 VPWR VGND sg13g2_decap_8
XFILLER_46_1027 VPWR VGND sg13g2_fill_2
XFILLER_46_1016 VPWR VGND sg13g2_decap_8
XFILLER_19_818 VPWR VGND sg13g2_fill_2
XFILLER_45_169 VPWR VGND sg13g2_decap_8
XFILLER_27_862 VPWR VGND sg13g2_decap_8
XFILLER_14_523 VPWR VGND sg13g2_decap_8
XFILLER_41_331 VPWR VGND sg13g2_fill_2
XFILLER_41_364 VPWR VGND sg13g2_decap_4
XFILLER_14_60 VPWR VGND sg13g2_fill_2
XFILLER_10_740 VPWR VGND sg13g2_decap_8
XFILLER_6_755 VPWR VGND sg13g2_decap_8
XFILLER_2_972 VPWR VGND sg13g2_decap_8
Xinput8 ui_in[7] net8 VPWR VGND sg13g2_buf_1
XFILLER_37_604 VPWR VGND sg13g2_fill_1
XFILLER_39_90 VPWR VGND sg13g2_decap_8
XFILLER_49_497 VPWR VGND sg13g2_fill_1
XFILLER_49_486 VPWR VGND sg13g2_decap_8
XFILLER_36_158 VPWR VGND sg13g2_decap_8
XFILLER_18_895 VPWR VGND sg13g2_decap_8
XFILLER_32_364 VPWR VGND sg13g2_decap_8
X_2714_ _0611_ _0610_ _0609_ VPWR VGND sg13g2_nand2b_1
X_2645_ _0507_ VPWR _0543_ VGND _0504_ _0508_ sg13g2_o21ai_1
XFILLER_0_909 VPWR VGND sg13g2_decap_8
X_2576_ _0464_ VPWR _0476_ VGND _0472_ _0474_ sg13g2_o21ai_1
X_1527_ _0862_ _0854_ _0860_ VPWR VGND sg13g2_xnor2_1
X_3128_ net547 VGND VPWR net127 mac1.sum_lvl1_ff\[15\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_28_648 VPWR VGND sg13g2_decap_8
XFILLER_27_147 VPWR VGND sg13g2_decap_8
X_3059_ net531 VGND VPWR net224 DP_2.matrix\[2\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_23_331 VPWR VGND sg13g2_decap_8
XFILLER_36_692 VPWR VGND sg13g2_decap_8
XFILLER_11_504 VPWR VGND sg13g2_decap_8
XFILLER_24_887 VPWR VGND sg13g2_decap_8
XFILLER_11_537 VPWR VGND sg13g2_decap_4
XFILLER_3_703 VPWR VGND sg13g2_decap_8
XFILLER_2_279 VPWR VGND sg13g2_fill_2
XFILLER_47_913 VPWR VGND sg13g2_decap_8
XFILLER_19_604 VPWR VGND sg13g2_decap_8
XFILLER_46_412 VPWR VGND sg13g2_fill_1
XFILLER_18_114 VPWR VGND sg13g2_fill_2
XFILLER_19_648 VPWR VGND sg13g2_decap_8
XFILLER_14_320 VPWR VGND sg13g2_decap_8
XFILLER_42_673 VPWR VGND sg13g2_decap_4
XFILLER_15_865 VPWR VGND sg13g2_decap_8
XFILLER_14_375 VPWR VGND sg13g2_decap_4
XFILLER_30_857 VPWR VGND sg13g2_decap_8
XFILLER_41_91 VPWR VGND sg13g2_decap_8
XFILLER_6_563 VPWR VGND sg13g2_decap_4
X_2430_ _0326_ VPWR _0337_ VGND _0297_ _0324_ sg13g2_o21ai_1
XFILLER_6_596 VPWR VGND sg13g2_decap_8
XFILLER_29_1011 VPWR VGND sg13g2_decap_8
X_2361_ _0271_ net449 net502 VPWR VGND sg13g2_nand2_1
X_2292_ _0204_ net449 net380 VPWR VGND sg13g2_nand2_1
XFILLER_38_924 VPWR VGND sg13g2_decap_8
XFILLER_2_74 VPWR VGND sg13g2_decap_8
XFILLER_2_85 VPWR VGND sg13g2_fill_1
XFILLER_37_434 VPWR VGND sg13g2_decap_8
XFILLER_37_478 VPWR VGND sg13g2_fill_2
XFILLER_17_191 VPWR VGND sg13g2_decap_8
XFILLER_33_640 VPWR VGND sg13g2_decap_8
XFILLER_36_1026 VPWR VGND sg13g2_fill_2
XFILLER_20_334 VPWR VGND sg13g2_fill_2
XFILLER_21_868 VPWR VGND sg13g2_decap_8
X_2628_ _0527_ _0491_ _0525_ _0526_ VPWR VGND sg13g2_and3_1
XFILLER_0_706 VPWR VGND sg13g2_decap_8
X_2559_ _0459_ net484 net427 VPWR VGND sg13g2_nand2_1
XFILLER_47_209 VPWR VGND sg13g2_decap_8
XFILLER_29_913 VPWR VGND sg13g2_decap_8
XFILLER_46_58 VPWR VGND sg13g2_fill_2
XFILLER_16_607 VPWR VGND sg13g2_decap_8
XFILLER_28_445 VPWR VGND sg13g2_decap_8
XFILLER_28_467 VPWR VGND sg13g2_decap_8
XFILLER_43_437 VPWR VGND sg13g2_decap_8
XFILLER_15_139 VPWR VGND sg13g2_decap_4
XFILLER_12_835 VPWR VGND sg13g2_decap_8
XFILLER_23_172 VPWR VGND sg13g2_decap_8
XFILLER_7_327 VPWR VGND sg13g2_decap_8
XFILLER_11_367 VPWR VGND sg13g2_fill_1
XFILLER_20_890 VPWR VGND sg13g2_decap_8
XFILLER_11_72 VPWR VGND sg13g2_decap_8
XFILLER_3_577 VPWR VGND sg13g2_decap_8
Xfanout391 net190 net391 VPWR VGND sg13g2_buf_8
Xfanout380 net381 net380 VPWR VGND sg13g2_buf_8
XFILLER_46_220 VPWR VGND sg13g2_fill_1
XFILLER_47_798 VPWR VGND sg13g2_fill_1
XFILLER_47_787 VPWR VGND sg13g2_decap_8
XFILLER_46_297 VPWR VGND sg13g2_decap_8
XFILLER_43_971 VPWR VGND sg13g2_decap_8
XFILLER_15_662 VPWR VGND sg13g2_decap_8
X_1930_ net297 VPWR _1245_ VGND _1239_ _1243_ sg13g2_o21ai_1
XFILLER_14_150 VPWR VGND sg13g2_decap_8
X_1861_ _1186_ _1177_ _1185_ VPWR VGND sg13g2_xnor2_1
Xinput11 uio_in[2] net11 VPWR VGND sg13g2_buf_1
XFILLER_30_698 VPWR VGND sg13g2_decap_8
XFILLER_7_861 VPWR VGND sg13g2_decap_8
X_1792_ _1119_ net408 net499 VPWR VGND sg13g2_nand2_1
X_2413_ _0300_ VPWR _0321_ VGND _0272_ _0298_ sg13g2_o21ai_1
X_2344_ _0253_ _0243_ _0255_ VPWR VGND sg13g2_xor2_1
X_2275_ _0187_ _0180_ _0188_ VPWR VGND sg13g2_xor2_1
XFILLER_26_916 VPWR VGND sg13g2_decap_8
XFILLER_37_264 VPWR VGND sg13g2_decap_8
XFILLER_37_275 VPWR VGND sg13g2_fill_1
XFILLER_25_448 VPWR VGND sg13g2_fill_1
XFILLER_33_470 VPWR VGND sg13g2_fill_1
XFILLER_34_982 VPWR VGND sg13g2_decap_8
XFILLER_21_632 VPWR VGND sg13g2_decap_8
XFILLER_20_142 VPWR VGND sg13g2_decap_8
XFILLER_4_319 VPWR VGND sg13g2_fill_2
XFILLER_4_308 VPWR VGND sg13g2_decap_8
XFILLER_0_503 VPWR VGND sg13g2_decap_8
XFILLER_29_732 VPWR VGND sg13g2_fill_1
XFILLER_44_702 VPWR VGND sg13g2_decap_8
XFILLER_16_448 VPWR VGND sg13g2_fill_1
XFILLER_17_949 VPWR VGND sg13g2_decap_8
XFILLER_28_286 VPWR VGND sg13g2_decap_8
XFILLER_43_245 VPWR VGND sg13g2_decap_8
XFILLER_11_120 VPWR VGND sg13g2_decap_8
XFILLER_40_974 VPWR VGND sg13g2_decap_8
XFILLER_8_625 VPWR VGND sg13g2_decap_4
XFILLER_4_875 VPWR VGND sg13g2_decap_8
XFILLER_26_1014 VPWR VGND sg13g2_decap_8
XFILLER_39_518 VPWR VGND sg13g2_decap_8
X_2060_ _1347_ _1339_ _1346_ VPWR VGND sg13g2_nand2_1
XFILLER_35_735 VPWR VGND sg13g2_decap_8
XFILLER_16_960 VPWR VGND sg13g2_decap_8
XFILLER_23_919 VPWR VGND sg13g2_decap_8
X_2962_ _0838_ net427 net375 VPWR VGND sg13g2_nand2_1
X_1913_ net255 _1229_ _0008_ VPWR VGND sg13g2_xor2_1
X_2893_ _0782_ DP_2.I_range.out_data\[3\] DP_2.Q_range.out_data\[3\] VPWR VGND sg13g2_xnor2_1
XFILLER_30_451 VPWR VGND sg13g2_decap_8
XFILLER_31_985 VPWR VGND sg13g2_decap_8
XFILLER_8_84 VPWR VGND sg13g2_fill_1
X_1844_ _1168_ _1169_ _1170_ VPWR VGND sg13g2_nor2_1
X_1775_ _1102_ _1090_ _1103_ VPWR VGND sg13g2_xor2_1
X_2327_ _0238_ net443 net384 VPWR VGND sg13g2_nand2_1
X_2258_ _0171_ _0164_ _0170_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_702 VPWR VGND sg13g2_decap_8
XFILLER_38_551 VPWR VGND sg13g2_fill_2
X_2189_ _1447_ _1468_ _1470_ _1471_ VPWR VGND sg13g2_or3_1
XFILLER_38_584 VPWR VGND sg13g2_decap_8
XFILLER_14_919 VPWR VGND sg13g2_decap_8
XFILLER_40_215 VPWR VGND sg13g2_decap_8
XFILLER_40_237 VPWR VGND sg13g2_decap_8
XFILLER_22_952 VPWR VGND sg13g2_decap_8
XFILLER_34_790 VPWR VGND sg13g2_decap_4
XFILLER_4_105 VPWR VGND sg13g2_fill_2
XFILLER_49_1014 VPWR VGND sg13g2_decap_8
XFILLER_1_856 VPWR VGND sg13g2_decap_8
XFILLER_44_521 VPWR VGND sg13g2_fill_2
XFILLER_29_595 VPWR VGND sg13g2_decap_8
XFILLER_44_554 VPWR VGND sg13g2_decap_4
XFILLER_17_60 VPWR VGND sg13g2_fill_2
XFILLER_32_705 VPWR VGND sg13g2_decap_4
XFILLER_44_598 VPWR VGND sg13g2_fill_1
XFILLER_16_289 VPWR VGND sg13g2_decap_8
XFILLER_32_738 VPWR VGND sg13g2_decap_4
XFILLER_13_974 VPWR VGND sg13g2_decap_8
XFILLER_40_793 VPWR VGND sg13g2_decap_4
XFILLER_9_956 VPWR VGND sg13g2_decap_8
XFILLER_8_433 VPWR VGND sg13g2_decap_8
X_1560_ _0893_ _0867_ _0890_ VPWR VGND sg13g2_xnor2_1
XFILLER_4_672 VPWR VGND sg13g2_decap_8
X_3230_ net510 VGND VPWR net259 mac1.sum_lvl3_ff\[5\] clknet_leaf_35_clk sg13g2_dfrbpq_2
X_3161_ net521 VGND VPWR net94 mac1.sum_lvl2_ff\[19\] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_2112_ _1396_ _1389_ _1394_ _1395_ VPWR VGND sg13g2_and3_1
X_3092_ net541 VGND VPWR _0071_ mac1.products_ff\[79\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_2043_ _1334_ mac1.sum_lvl3_ff\[14\] mac1.sum_lvl3_ff\[34\] VPWR VGND sg13g2_nand2_1
XFILLER_35_521 VPWR VGND sg13g2_fill_2
XFILLER_35_554 VPWR VGND sg13g2_decap_8
X_2945_ _0761_ _0757_ _0827_ VPWR VGND sg13g2_xor2_1
X_2876_ DP_1.Q_range.out_data\[4\] DP_1.Q_range.out_data\[6\] _0766_ VPWR VGND sg13g2_nor2_1
X_1827_ _1153_ net462 net401 VPWR VGND sg13g2_nand2_1
XFILLER_30_292 VPWR VGND sg13g2_decap_8
X_1758_ _1086_ _1044_ _1084_ VPWR VGND sg13g2_xnor2_1
X_1689_ _1008_ _1016_ _1018_ _1019_ VPWR VGND sg13g2_or3_1
XFILLER_16_1002 VPWR VGND sg13g2_decap_8
XFILLER_41_579 VPWR VGND sg13g2_decap_8
XFILLER_9_219 VPWR VGND sg13g2_decap_8
XFILLER_22_771 VPWR VGND sg13g2_decap_8
XFILLER_10_922 VPWR VGND sg13g2_decap_8
XFILLER_6_937 VPWR VGND sg13g2_decap_8
XFILLER_10_999 VPWR VGND sg13g2_decap_8
XFILLER_1_653 VPWR VGND sg13g2_decap_8
XFILLER_49_657 VPWR VGND sg13g2_decap_8
XFILLER_49_635 VPWR VGND sg13g2_fill_1
XFILLER_23_1017 VPWR VGND sg13g2_decap_8
XFILLER_23_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_679 VPWR VGND sg13g2_decap_8
XFILLER_48_167 VPWR VGND sg13g2_decap_8
XFILLER_45_830 VPWR VGND sg13g2_decap_8
XFILLER_29_370 VPWR VGND sg13g2_decap_8
X_2730_ VGND VPWR _0626_ _0624_ _0619_ sg13g2_or2_1
XFILLER_9_753 VPWR VGND sg13g2_decap_8
XFILLER_8_230 VPWR VGND sg13g2_decap_4
X_2661_ _0559_ _0554_ _0558_ VPWR VGND sg13g2_xnor2_1
X_1612_ _0944_ _0919_ _0943_ VPWR VGND sg13g2_xnor2_1
X_2592_ _0478_ VPWR _0491_ VGND _0456_ _0479_ sg13g2_o21ai_1
XFILLER_5_63 VPWR VGND sg13g2_decap_8
X_1543_ _0877_ _0870_ _0875_ _0876_ VPWR VGND sg13g2_and3_1
X_3213_ net509 VGND VPWR net114 mac1.sum_lvl3_ff\[24\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_3144_ net544 VGND VPWR net85 mac1.sum_lvl1_ff\[51\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_3075_ net517 VGND VPWR _0128_ DP_2.matrix\[74\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_39_178 VPWR VGND sg13g2_decap_8
XFILLER_39_1002 VPWR VGND sg13g2_decap_8
X_2026_ _1320_ mac1.sum_lvl3_ff\[11\] mac1.sum_lvl3_ff\[31\] VPWR VGND sg13g2_nand2_1
XFILLER_35_340 VPWR VGND sg13g2_fill_1
XFILLER_23_579 VPWR VGND sg13g2_decap_8
X_2928_ _0816_ VPWR _0084_ VGND _0812_ net374 sg13g2_o21ai_1
XFILLER_31_590 VPWR VGND sg13g2_decap_8
XFILLER_40_38 VPWR VGND sg13g2_fill_2
X_2859_ _0749_ net376 _0748_ _0732_ net215 VPWR VGND sg13g2_a22oi_1
Xhold252 _1324_ VPWR VGND net292 sg13g2_dlygate4sd3_1
Xhold230 DP_2.matrix\[36\] VPWR VGND net270 sg13g2_dlygate4sd3_1
Xhold241 _0004_ VPWR VGND net281 sg13g2_dlygate4sd3_1
XFILLER_49_14 VPWR VGND sg13g2_decap_8
Xhold263 _0001_ VPWR VGND net303 sg13g2_dlygate4sd3_1
XFILLER_19_808 VPWR VGND sg13g2_fill_1
XFILLER_46_649 VPWR VGND sg13g2_fill_2
XFILLER_14_502 VPWR VGND sg13g2_decap_8
XFILLER_42_888 VPWR VGND sg13g2_decap_8
XFILLER_41_343 VPWR VGND sg13g2_decap_8
XFILLER_14_579 VPWR VGND sg13g2_decap_4
XFILLER_41_398 VPWR VGND sg13g2_fill_2
XFILLER_41_387 VPWR VGND sg13g2_decap_4
XFILLER_14_94 VPWR VGND sg13g2_decap_8
XFILLER_10_796 VPWR VGND sg13g2_decap_8
XFILLER_6_734 VPWR VGND sg13g2_decap_8
XFILLER_5_211 VPWR VGND sg13g2_decap_4
XFILLER_5_244 VPWR VGND sg13g2_fill_2
XFILLER_30_60 VPWR VGND sg13g2_decap_8
XFILLER_30_82 VPWR VGND sg13g2_decap_8
XFILLER_2_951 VPWR VGND sg13g2_decap_8
XFILLER_49_421 VPWR VGND sg13g2_decap_8
XFILLER_7_1022 VPWR VGND sg13g2_decap_8
XFILLER_49_465 VPWR VGND sg13g2_decap_8
XFILLER_36_104 VPWR VGND sg13g2_decap_8
Xinput9 uio_in[0] net9 VPWR VGND sg13g2_buf_1
XFILLER_18_874 VPWR VGND sg13g2_decap_8
XFILLER_33_811 VPWR VGND sg13g2_fill_1
XFILLER_17_395 VPWR VGND sg13g2_decap_8
XFILLER_32_332 VPWR VGND sg13g2_decap_8
XFILLER_20_516 VPWR VGND sg13g2_decap_8
X_2713_ _0573_ _0608_ _0571_ _0610_ VPWR VGND sg13g2_nand3_1
X_2644_ _0495_ _0498_ _0542_ VPWR VGND sg13g2_nor2_1
X_2575_ _0464_ _0472_ _0474_ _0475_ VPWR VGND sg13g2_or3_1
X_1526_ _0861_ _0860_ _0854_ VPWR VGND sg13g2_nand2b_1
X_3127_ net547 VGND VPWR net121 mac1.sum_lvl1_ff\[14\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_27_126 VPWR VGND sg13g2_decap_8
XFILLER_35_38 VPWR VGND sg13g2_decap_4
X_3058_ net531 VGND VPWR net222 DP_2.matrix\[1\] clknet_leaf_14_clk sg13g2_dfrbpq_2
X_2009_ net288 _1306_ _0029_ VPWR VGND sg13g2_and2_1
XFILLER_24_844 VPWR VGND sg13g2_decap_8
XFILLER_11_527 VPWR VGND sg13g2_fill_1
XFILLER_11_549 VPWR VGND sg13g2_fill_2
XFILLER_13_1016 VPWR VGND sg13g2_decap_8
XFILLER_13_1027 VPWR VGND sg13g2_fill_2
XFILLER_3_759 VPWR VGND sg13g2_decap_8
Xfanout540 net541 net540 VPWR VGND sg13g2_buf_8
XFILLER_19_616 VPWR VGND sg13g2_decap_8
XFILLER_20_1009 VPWR VGND sg13g2_decap_8
XFILLER_47_969 VPWR VGND sg13g2_decap_8
XFILLER_15_844 VPWR VGND sg13g2_decap_8
XFILLER_42_641 VPWR VGND sg13g2_decap_4
XFILLER_42_685 VPWR VGND sg13g2_decap_8
XFILLER_14_398 VPWR VGND sg13g2_decap_8
XFILLER_30_836 VPWR VGND sg13g2_decap_8
X_2360_ _0240_ VPWR _0270_ VGND _0238_ _0241_ sg13g2_o21ai_1
X_2291_ _0203_ DP_1.matrix\[74\] net502 VPWR VGND sg13g2_nand2_1
XFILLER_38_903 VPWR VGND sg13g2_decap_8
XFILLER_49_284 VPWR VGND sg13g2_decap_8
XFILLER_37_424 VPWR VGND sg13g2_decap_4
XFILLER_33_663 VPWR VGND sg13g2_decap_8
XFILLER_36_1005 VPWR VGND sg13g2_decap_8
XFILLER_21_847 VPWR VGND sg13g2_decap_8
X_2627_ _0502_ VPWR _0526_ VGND _0522_ _0524_ sg13g2_o21ai_1
X_2558_ _0458_ net489 net426 VPWR VGND sg13g2_nand2_1
X_1509_ net417 net470 net472 net412 _0846_ VPWR VGND sg13g2_and4_1
X_2489_ _0391_ _0390_ _0387_ VPWR VGND sg13g2_nand2b_1
XFILLER_28_424 VPWR VGND sg13g2_fill_1
XFILLER_46_37 VPWR VGND sg13g2_decap_8
XFILLER_29_969 VPWR VGND sg13g2_decap_8
XFILLER_43_416 VPWR VGND sg13g2_decap_8
XFILLER_37_980 VPWR VGND sg13g2_decap_8
XFILLER_15_118 VPWR VGND sg13g2_decap_8
XFILLER_24_630 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_35_clk clknet_3_1__leaf_clk clknet_leaf_35_clk VPWR VGND sg13g2_buf_8
XFILLER_12_814 VPWR VGND sg13g2_fill_2
XFILLER_23_151 VPWR VGND sg13g2_decap_8
XFILLER_24_696 VPWR VGND sg13g2_fill_2
XFILLER_3_501 VPWR VGND sg13g2_fill_1
Xfanout381 net185 net381 VPWR VGND sg13g2_buf_8
Xfanout392 net393 net392 VPWR VGND sg13g2_buf_2
XFILLER_47_766 VPWR VGND sg13g2_fill_2
XFILLER_46_276 VPWR VGND sg13g2_decap_8
XFILLER_34_438 VPWR VGND sg13g2_fill_1
XFILLER_43_950 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_26_clk clknet_3_5__leaf_clk clknet_leaf_26_clk VPWR VGND sg13g2_buf_8
XFILLER_30_655 VPWR VGND sg13g2_decap_8
X_1860_ _1185_ _1148_ _1183_ VPWR VGND sg13g2_xnor2_1
Xinput12 uio_in[3] net12 VPWR VGND sg13g2_buf_1
X_1791_ _1118_ net405 net462 VPWR VGND sg13g2_nand2_1
XFILLER_7_840 VPWR VGND sg13g2_decap_8
XFILLER_11_891 VPWR VGND sg13g2_decap_8
XFILLER_6_372 VPWR VGND sg13g2_decap_4
X_2412_ _0303_ _0295_ _0302_ _0320_ VPWR VGND sg13g2_a21o_1
X_2343_ _0243_ _0253_ _0254_ VPWR VGND sg13g2_nor2_1
X_2274_ _0187_ _0181_ _0185_ VPWR VGND sg13g2_xnor2_1
XFILLER_25_405 VPWR VGND sg13g2_fill_1
XFILLER_37_243 VPWR VGND sg13g2_decap_8
XFILLER_16_29 VPWR VGND sg13g2_decap_4
XFILLER_37_287 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_17_clk clknet_3_7__leaf_clk clknet_leaf_17_clk VPWR VGND sg13g2_buf_8
XFILLER_18_490 VPWR VGND sg13g2_decap_8
XFILLER_34_961 VPWR VGND sg13g2_decap_8
X_1989_ _1291_ mac1.sum_lvl3_ff\[3\] net200 VPWR VGND sg13g2_xnor2_1
XFILLER_0_559 VPWR VGND sg13g2_decap_8
XFILLER_29_755 VPWR VGND sg13g2_fill_2
XFILLER_17_928 VPWR VGND sg13g2_decap_8
XFILLER_28_265 VPWR VGND sg13g2_decap_8
XFILLER_12_611 VPWR VGND sg13g2_fill_2
XFILLER_25_983 VPWR VGND sg13g2_decap_8
XFILLER_40_953 VPWR VGND sg13g2_decap_8
XFILLER_12_688 VPWR VGND sg13g2_decap_4
XFILLER_7_136 VPWR VGND sg13g2_fill_2
XFILLER_4_854 VPWR VGND sg13g2_decap_8
XFILLER_21_8 VPWR VGND sg13g2_fill_1
XFILLER_47_596 VPWR VGND sg13g2_decap_8
XFILLER_35_725 VPWR VGND sg13g2_fill_2
XFILLER_34_246 VPWR VGND sg13g2_decap_8
XFILLER_34_257 VPWR VGND sg13g2_fill_2
X_2961_ _0837_ _0801_ _0803_ VPWR VGND sg13g2_xnor2_1
XFILLER_15_460 VPWR VGND sg13g2_decap_4
XFILLER_34_268 VPWR VGND sg13g2_fill_2
X_1912_ net254 mac1.sum_lvl2_ff\[21\] _1231_ VPWR VGND sg13g2_xor2_1
XFILLER_15_482 VPWR VGND sg13g2_decap_8
XFILLER_31_964 VPWR VGND sg13g2_decap_8
XFILLER_33_1008 VPWR VGND sg13g2_decap_8
X_2892_ _0781_ DP_2.I_range.out_data\[2\] DP_2.Q_range.out_data\[2\] VPWR VGND sg13g2_xnor2_1
XFILLER_8_52 VPWR VGND sg13g2_decap_8
X_1843_ VGND VPWR _1116_ _1136_ _1169_ _1138_ sg13g2_a21oi_1
X_1774_ _1100_ _1091_ _1102_ VPWR VGND sg13g2_xor2_1
Xclkbuf_leaf_6_clk clknet_3_6__leaf_clk clknet_leaf_6_clk VPWR VGND sg13g2_buf_8
X_2326_ _0220_ _0213_ _0183_ _0237_ VPWR VGND sg13g2_a21o_1
X_2257_ _0170_ _0165_ _0168_ VPWR VGND sg13g2_xnor2_1
X_2188_ VGND VPWR _1466_ _1467_ _1470_ _1448_ sg13g2_a21oi_1
XFILLER_25_224 VPWR VGND sg13g2_decap_8
XFILLER_41_706 VPWR VGND sg13g2_decap_8
XFILLER_26_758 VPWR VGND sg13g2_decap_8
XFILLER_26_769 VPWR VGND sg13g2_fill_2
XFILLER_34_780 VPWR VGND sg13g2_fill_1
XFILLER_22_931 VPWR VGND sg13g2_decap_8
XFILLER_21_463 VPWR VGND sg13g2_decap_8
XFILLER_0_312 VPWR VGND sg13g2_decap_8
XFILLER_1_835 VPWR VGND sg13g2_decap_8
XFILLER_49_839 VPWR VGND sg13g2_decap_8
XFILLER_0_356 VPWR VGND sg13g2_fill_1
XFILLER_17_703 VPWR VGND sg13g2_decap_8
XFILLER_29_541 VPWR VGND sg13g2_decap_4
XFILLER_1_1017 VPWR VGND sg13g2_decap_8
XFILLER_1_1028 VPWR VGND sg13g2_fill_1
XFILLER_29_574 VPWR VGND sg13g2_fill_1
XFILLER_17_758 VPWR VGND sg13g2_decap_4
XFILLER_44_577 VPWR VGND sg13g2_decap_8
XFILLER_12_430 VPWR VGND sg13g2_decap_4
XFILLER_13_953 VPWR VGND sg13g2_decap_8
XFILLER_9_935 VPWR VGND sg13g2_decap_8
XFILLER_8_412 VPWR VGND sg13g2_decap_8
XFILLER_8_423 VPWR VGND sg13g2_fill_1
XFILLER_8_478 VPWR VGND sg13g2_decap_4
XFILLER_4_651 VPWR VGND sg13g2_decap_8
X_3160_ net547 VGND VPWR net79 mac1.sum_lvl2_ff\[15\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_12_4 VPWR VGND sg13g2_decap_4
X_2111_ _1390_ VPWR _1395_ VGND _1391_ _1393_ sg13g2_o21ai_1
X_3091_ net542 VGND VPWR _0070_ mac1.products_ff\[78\] clknet_leaf_23_clk sg13g2_dfrbpq_1
Xhold1 mac1.sum_lvl1_ff\[87\] VPWR VGND net41 sg13g2_dlygate4sd3_1
XFILLER_39_349 VPWR VGND sg13g2_decap_8
X_2042_ VGND VPWR mac1.sum_lvl3_ff\[13\] mac1.sum_lvl3_ff\[33\] _1333_ _1331_ sg13g2_a21oi_1
XFILLER_22_216 VPWR VGND sg13g2_fill_2
XFILLER_35_599 VPWR VGND sg13g2_decap_8
X_2944_ VGND VPWR net371 _0825_ _0091_ _0826_ sg13g2_a21oi_1
X_2875_ _0765_ _0762_ _0764_ VPWR VGND sg13g2_nand2b_1
X_1826_ _1152_ net467 net494 VPWR VGND sg13g2_nand2_1
X_1757_ VGND VPWR _1085_ _1083_ _1045_ sg13g2_or2_1
X_1688_ VGND VPWR _1014_ _1015_ _1018_ _1009_ sg13g2_a21oi_1
X_2309_ _0221_ _0213_ _0220_ VPWR VGND sg13g2_xnor2_1
XFILLER_39_883 VPWR VGND sg13g2_decap_8
XFILLER_41_514 VPWR VGND sg13g2_fill_1
XFILLER_13_205 VPWR VGND sg13g2_fill_2
XFILLER_14_717 VPWR VGND sg13g2_decap_8
XFILLER_26_577 VPWR VGND sg13g2_fill_1
XFILLER_10_901 VPWR VGND sg13g2_decap_8
XFILLER_21_282 VPWR VGND sg13g2_decap_8
XFILLER_10_978 VPWR VGND sg13g2_decap_8
XFILLER_6_916 VPWR VGND sg13g2_decap_8
XFILLER_1_632 VPWR VGND sg13g2_decap_8
XFILLER_49_603 VPWR VGND sg13g2_fill_2
XFILLER_0_197 VPWR VGND sg13g2_decap_8
XFILLER_17_533 VPWR VGND sg13g2_decap_8
XFILLER_45_886 VPWR VGND sg13g2_decap_8
XFILLER_32_503 VPWR VGND sg13g2_decap_4
XFILLER_44_385 VPWR VGND sg13g2_decap_4
XFILLER_32_547 VPWR VGND sg13g2_fill_2
XFILLER_9_732 VPWR VGND sg13g2_decap_8
X_2660_ _0558_ _0505_ _0555_ VPWR VGND sg13g2_xnor2_1
X_1611_ _0940_ _0942_ _0943_ VPWR VGND sg13g2_nor2_1
X_2591_ _0066_ _0449_ _0490_ VPWR VGND sg13g2_xnor2_1
XFILLER_5_993 VPWR VGND sg13g2_decap_8
X_1542_ _0871_ VPWR _0876_ VGND _0872_ _0874_ sg13g2_o21ai_1
X_3212_ net509 VGND VPWR net141 mac1.sum_lvl3_ff\[23\] clknet_leaf_36_clk sg13g2_dfrbpq_1
XFILLER_39_124 VPWR VGND sg13g2_decap_8
X_3143_ net544 VGND VPWR net63 mac1.sum_lvl1_ff\[50\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_3074_ net518 VGND VPWR _0127_ DP_2.matrix\[73\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_2025_ mac1.sum_lvl3_ff\[11\] mac1.sum_lvl3_ff\[31\] _1319_ VPWR VGND sg13g2_nor2_1
XFILLER_36_886 VPWR VGND sg13g2_decap_8
XFILLER_23_536 VPWR VGND sg13g2_decap_4
X_2927_ _0816_ net495 net374 VPWR VGND sg13g2_nand2_1
X_2858_ net470 net488 net379 _0748_ VPWR VGND sg13g2_mux2_1
X_2789_ _0682_ _0655_ _0683_ VPWR VGND sg13g2_xor2_1
X_1809_ _1136_ _1125_ _1135_ VPWR VGND sg13g2_xnor2_1
Xhold220 DP_1.matrix\[3\] VPWR VGND net260 sg13g2_dlygate4sd3_1
Xhold242 DP_2.matrix\[5\] VPWR VGND net282 sg13g2_dlygate4sd3_1
XFILLER_2_418 VPWR VGND sg13g2_fill_2
Xhold253 _0019_ VPWR VGND net293 sg13g2_dlygate4sd3_1
Xhold231 DP_1.matrix\[73\] VPWR VGND net271 sg13g2_dlygate4sd3_1
Xhold264 mac1.sum_lvl2_ff\[7\] VPWR VGND net304 sg13g2_dlygate4sd3_1
XFILLER_45_127 VPWR VGND sg13g2_fill_2
XFILLER_45_116 VPWR VGND sg13g2_decap_8
XFILLER_27_897 VPWR VGND sg13g2_decap_8
XFILLER_41_333 VPWR VGND sg13g2_fill_1
XFILLER_41_311 VPWR VGND sg13g2_fill_2
XFILLER_42_867 VPWR VGND sg13g2_decap_8
XFILLER_14_558 VPWR VGND sg13g2_decap_8
XFILLER_22_580 VPWR VGND sg13g2_decap_8
XFILLER_14_73 VPWR VGND sg13g2_decap_8
XFILLER_10_775 VPWR VGND sg13g2_decap_8
XFILLER_6_713 VPWR VGND sg13g2_decap_8
XFILLER_5_289 VPWR VGND sg13g2_decap_8
XFILLER_2_930 VPWR VGND sg13g2_decap_8
XFILLER_49_400 VPWR VGND sg13g2_decap_8
XFILLER_7_1001 VPWR VGND sg13g2_decap_8
XFILLER_45_672 VPWR VGND sg13g2_fill_1
XFILLER_17_374 VPWR VGND sg13g2_decap_8
XFILLER_33_889 VPWR VGND sg13g2_decap_8
XFILLER_32_388 VPWR VGND sg13g2_decap_8
X_2712_ VGND VPWR _0571_ _0573_ _0609_ _0608_ sg13g2_a21oi_1
XFILLER_9_540 VPWR VGND sg13g2_decap_8
X_2643_ _0523_ VPWR _0541_ VGND _0502_ _0524_ sg13g2_o21ai_1
X_2574_ VGND VPWR _0470_ _0471_ _0474_ _0465_ sg13g2_a21oi_1
XFILLER_5_790 VPWR VGND sg13g2_decap_8
X_1525_ _0858_ _0859_ _0860_ VPWR VGND sg13g2_nor2b_1
X_3126_ net545 VGND VPWR net117 mac1.sum_lvl1_ff\[13\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_28_628 VPWR VGND sg13g2_fill_2
XFILLER_42_108 VPWR VGND sg13g2_decap_4
X_3057_ net531 VGND VPWR net199 DP_2.matrix\[0\] clknet_leaf_14_clk sg13g2_dfrbpq_2
XFILLER_36_650 VPWR VGND sg13g2_decap_8
XFILLER_36_661 VPWR VGND sg13g2_fill_2
X_2008_ _1298_ _1301_ _1304_ _1306_ VPWR VGND sg13g2_or3_1
XFILLER_24_823 VPWR VGND sg13g2_decap_8
XFILLER_23_399 VPWR VGND sg13g2_decap_8
XFILLER_2_204 VPWR VGND sg13g2_decap_8
XFILLER_3_738 VPWR VGND sg13g2_decap_8
Xfanout541 net542 net541 VPWR VGND sg13g2_buf_8
Xfanout530 net532 net530 VPWR VGND sg13g2_buf_2
XFILLER_47_948 VPWR VGND sg13g2_decap_8
XFILLER_18_149 VPWR VGND sg13g2_decap_8
XFILLER_34_609 VPWR VGND sg13g2_fill_2
XFILLER_6_510 VPWR VGND sg13g2_decap_8
XFILLER_10_583 VPWR VGND sg13g2_decap_4
X_2290_ _0177_ VPWR _0202_ VGND _0175_ _0178_ sg13g2_o21ai_1
XFILLER_2_32 VPWR VGND sg13g2_decap_4
XFILLER_49_263 VPWR VGND sg13g2_decap_8
XFILLER_2_54 VPWR VGND sg13g2_decap_8
XFILLER_38_959 VPWR VGND sg13g2_decap_8
XFILLER_46_981 VPWR VGND sg13g2_decap_8
XFILLER_21_826 VPWR VGND sg13g2_decap_8
XFILLER_32_152 VPWR VGND sg13g2_decap_4
XFILLER_36_1028 VPWR VGND sg13g2_fill_1
XFILLER_20_336 VPWR VGND sg13g2_fill_1
XFILLER_32_196 VPWR VGND sg13g2_decap_8
X_2626_ _0502_ _0522_ _0524_ _0525_ VPWR VGND sg13g2_or3_1
X_2557_ _0436_ _0426_ _0434_ _0457_ VPWR VGND sg13g2_a21o_1
X_1508_ net472 net412 _0845_ VPWR VGND sg13g2_and2_1
X_2488_ _0389_ _0366_ _0390_ VPWR VGND sg13g2_xor2_1
XFILLER_29_948 VPWR VGND sg13g2_decap_8
XFILLER_44_929 VPWR VGND sg13g2_decap_8
X_3109_ net529 VGND VPWR _0050_ mac1.products_ff\[148\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_36_480 VPWR VGND sg13g2_decap_8
XFILLER_11_52 VPWR VGND sg13g2_decap_4
XFILLER_3_535 VPWR VGND sg13g2_decap_8
XFILLER_47_712 VPWR VGND sg13g2_fill_2
XFILLER_47_701 VPWR VGND sg13g2_decap_8
Xfanout371 net372 net371 VPWR VGND sg13g2_buf_2
XFILLER_4_1015 VPWR VGND sg13g2_decap_8
Xfanout393 net395 net393 VPWR VGND sg13g2_buf_1
Xfanout382 net383 net382 VPWR VGND sg13g2_buf_8
XFILLER_35_929 VPWR VGND sg13g2_decap_8
XFILLER_30_634 VPWR VGND sg13g2_decap_8
Xinput13 uio_in[4] net13 VPWR VGND sg13g2_buf_1
XFILLER_11_870 VPWR VGND sg13g2_decap_8
X_1790_ _1099_ _1092_ _1061_ _1117_ VPWR VGND sg13g2_a21o_2
XFILLER_6_340 VPWR VGND sg13g2_decap_8
XFILLER_7_896 VPWR VGND sg13g2_decap_8
XFILLER_6_395 VPWR VGND sg13g2_decap_8
XFILLER_42_4 VPWR VGND sg13g2_decap_4
X_2411_ _0307_ _0309_ _0319_ VPWR VGND sg13g2_and2_1
X_2342_ _0251_ _0244_ _0253_ VPWR VGND sg13g2_xor2_1
XFILLER_42_1021 VPWR VGND sg13g2_decap_8
X_2273_ _0186_ _0181_ _0185_ VPWR VGND sg13g2_nand2_1
XFILLER_38_712 VPWR VGND sg13g2_decap_8
XFILLER_38_734 VPWR VGND sg13g2_fill_2
XFILLER_19_992 VPWR VGND sg13g2_decap_8
XFILLER_34_940 VPWR VGND sg13g2_decap_8
XFILLER_33_450 VPWR VGND sg13g2_decap_8
XFILLER_21_645 VPWR VGND sg13g2_fill_2
XFILLER_20_133 VPWR VGND sg13g2_decap_4
XFILLER_21_678 VPWR VGND sg13g2_decap_8
XFILLER_21_689 VPWR VGND sg13g2_fill_1
X_1988_ _1290_ mac1.sum_lvl3_ff\[3\] net200 VPWR VGND sg13g2_nand2_1
XFILLER_20_188 VPWR VGND sg13g2_decap_8
X_2609_ _0508_ _0459_ _0506_ VPWR VGND sg13g2_xnor2_1
XFILLER_0_538 VPWR VGND sg13g2_decap_8
XFILLER_17_907 VPWR VGND sg13g2_decap_8
XFILLER_28_244 VPWR VGND sg13g2_decap_8
XFILLER_16_439 VPWR VGND sg13g2_decap_8
XFILLER_25_962 VPWR VGND sg13g2_decap_8
XFILLER_12_601 VPWR VGND sg13g2_fill_2
XFILLER_40_932 VPWR VGND sg13g2_decap_8
XFILLER_11_177 VPWR VGND sg13g2_decap_8
XFILLER_4_833 VPWR VGND sg13g2_decap_8
XFILLER_22_95 VPWR VGND sg13g2_decap_8
XFILLER_3_387 VPWR VGND sg13g2_fill_1
XFILLER_3_376 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_14_8 VPWR VGND sg13g2_fill_1
XFILLER_19_211 VPWR VGND sg13g2_fill_2
XFILLER_19_222 VPWR VGND sg13g2_decap_8
XFILLER_47_575 VPWR VGND sg13g2_decap_8
XFILLER_19_277 VPWR VGND sg13g2_fill_2
X_2960_ _0836_ VPWR _0113_ VGND net374 _0835_ sg13g2_o21ai_1
XFILLER_16_995 VPWR VGND sg13g2_decap_8
X_2891_ DP_2.Q_range.out_data\[2\] DP_2.I_range.out_data\[2\] _0780_ VPWR VGND sg13g2_nor2b_1
X_1911_ mac1.sum_lvl2_ff\[21\] mac1.sum_lvl2_ff\[2\] _1230_ VPWR VGND sg13g2_and2_1
XFILLER_31_943 VPWR VGND sg13g2_decap_8
X_1842_ _1166_ _1145_ _1168_ VPWR VGND sg13g2_xor2_1
X_1773_ _1101_ _1091_ _1100_ VPWR VGND sg13g2_nand2b_1
XFILLER_7_693 VPWR VGND sg13g2_decap_8
X_2325_ _0222_ VPWR _0236_ VGND _0211_ _0223_ sg13g2_o21ai_1
XFILLER_27_18 VPWR VGND sg13g2_decap_8
X_2256_ _0169_ _0168_ _0165_ VPWR VGND sg13g2_nand2b_1
X_2187_ _1466_ _1467_ _1448_ _1469_ VPWR VGND sg13g2_nand3_1
XFILLER_25_203 VPWR VGND sg13g2_decap_8
XFILLER_22_910 VPWR VGND sg13g2_decap_8
XFILLER_22_987 VPWR VGND sg13g2_decap_8
XFILLER_21_497 VPWR VGND sg13g2_decap_8
XFILLER_4_129 VPWR VGND sg13g2_fill_2
XFILLER_1_814 VPWR VGND sg13g2_decap_8
XFILLER_0_335 VPWR VGND sg13g2_decap_8
XFILLER_49_818 VPWR VGND sg13g2_decap_8
XFILLER_44_523 VPWR VGND sg13g2_fill_1
XFILLER_17_737 VPWR VGND sg13g2_decap_8
XFILLER_17_62 VPWR VGND sg13g2_fill_1
XFILLER_17_84 VPWR VGND sg13g2_decap_8
XFILLER_13_932 VPWR VGND sg13g2_decap_8
XFILLER_9_914 VPWR VGND sg13g2_decap_8
XFILLER_12_486 VPWR VGND sg13g2_decap_8
XFILLER_4_630 VPWR VGND sg13g2_decap_8
XFILLER_3_162 VPWR VGND sg13g2_decap_8
X_3090_ net543 VGND VPWR _0079_ mac1.products_ff\[77\] clknet_leaf_24_clk sg13g2_dfrbpq_1
X_2110_ _1390_ _1391_ _1393_ _1394_ VPWR VGND sg13g2_or3_1
Xhold2 mac1.sum_lvl1_ff\[50\] VPWR VGND net42 sg13g2_dlygate4sd3_1
XFILLER_39_328 VPWR VGND sg13g2_decap_8
X_2041_ net233 _1332_ _0020_ VPWR VGND sg13g2_nor2b_1
XFILLER_48_884 VPWR VGND sg13g2_decap_8
XFILLER_47_372 VPWR VGND sg13g2_decap_8
X_2943_ net483 net371 _0826_ VPWR VGND sg13g2_nor2_1
XFILLER_22_239 VPWR VGND sg13g2_decap_4
XFILLER_31_762 VPWR VGND sg13g2_fill_1
XFILLER_31_795 VPWR VGND sg13g2_decap_8
X_2874_ _0764_ _0735_ _0763_ _0732_ net441 VPWR VGND sg13g2_a22oi_1
X_1825_ _1120_ VPWR _1151_ VGND _1118_ _1121_ sg13g2_o21ai_1
XFILLER_8_991 VPWR VGND sg13g2_decap_8
X_1756_ _1084_ net467 net404 VPWR VGND sg13g2_nand2_1
X_1687_ _1014_ _1015_ _1009_ _1017_ VPWR VGND sg13g2_nand3_1
X_2308_ _0218_ _0219_ _0220_ VPWR VGND sg13g2_nor2b_1
XFILLER_39_862 VPWR VGND sg13g2_decap_8
X_2239_ _1446_ VPWR _0153_ VGND _0149_ _0151_ sg13g2_o21ai_1
XFILLER_26_556 VPWR VGND sg13g2_decap_8
XFILLER_41_548 VPWR VGND sg13g2_decap_4
XFILLER_10_957 VPWR VGND sg13g2_decap_8
XFILLER_1_611 VPWR VGND sg13g2_decap_8
XFILLER_49_626 VPWR VGND sg13g2_decap_8
XFILLER_0_176 VPWR VGND sg13g2_decap_8
XFILLER_1_688 VPWR VGND sg13g2_decap_8
XFILLER_36_309 VPWR VGND sg13g2_decap_8
XFILLER_29_350 VPWR VGND sg13g2_fill_2
XFILLER_45_865 VPWR VGND sg13g2_decap_8
XFILLER_17_556 VPWR VGND sg13g2_decap_8
XFILLER_28_94 VPWR VGND sg13g2_fill_1
XFILLER_32_515 VPWR VGND sg13g2_decap_4
XFILLER_9_711 VPWR VGND sg13g2_decap_8
XFILLER_9_788 VPWR VGND sg13g2_decap_8
X_1610_ VGND VPWR _0938_ _0939_ _0942_ _0921_ sg13g2_a21oi_1
XFILLER_8_298 VPWR VGND sg13g2_decap_8
X_2590_ _0487_ _0489_ _0490_ VPWR VGND sg13g2_nor2_1
XFILLER_5_972 VPWR VGND sg13g2_decap_8
X_1541_ _0871_ _0872_ _0874_ _0875_ VPWR VGND sg13g2_or3_1
X_3211_ net509 VGND VPWR net115 mac1.sum_lvl3_ff\[22\] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_3142_ net540 VGND VPWR net47 mac1.sum_lvl1_ff\[49\] clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_39_158 VPWR VGND sg13g2_fill_1
X_3073_ net518 VGND VPWR _0126_ DP_2.matrix\[72\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_2024_ _1317_ _1315_ _0017_ VPWR VGND sg13g2_xor2_1
XFILLER_36_865 VPWR VGND sg13g2_decap_8
XFILLER_35_375 VPWR VGND sg13g2_fill_1
XFILLER_23_559 VPWR VGND sg13g2_decap_8
X_2926_ _0779_ _0813_ _0778_ _0815_ VPWR VGND _0814_ sg13g2_nand4_1
X_2857_ _0742_ _0746_ _0747_ VPWR VGND sg13g2_nor2b_1
X_1808_ _1135_ _1126_ _1133_ VPWR VGND sg13g2_xnor2_1
X_2788_ _0682_ net476 net424 VPWR VGND sg13g2_nand2_1
Xhold210 _0819_ VPWR VGND net250 sg13g2_dlygate4sd3_1
Xhold221 mac1.sum_lvl3_ff\[26\] VPWR VGND net261 sg13g2_dlygate4sd3_1
Xhold243 mac1.sum_lvl2_ff\[26\] VPWR VGND net283 sg13g2_dlygate4sd3_1
X_1739_ _1068_ _1052_ _1066_ VPWR VGND sg13g2_xnor2_1
Xhold232 DP_1.matrix\[76\] VPWR VGND net272 sg13g2_dlygate4sd3_1
Xhold265 _1247_ VPWR VGND net305 sg13g2_dlygate4sd3_1
Xhold254 mac1.sum_lvl2_ff\[9\] VPWR VGND net294 sg13g2_dlygate4sd3_1
XFILLER_49_49 VPWR VGND sg13g2_decap_8
XFILLER_46_629 VPWR VGND sg13g2_fill_1
XFILLER_39_681 VPWR VGND sg13g2_decap_8
XFILLER_42_802 VPWR VGND sg13g2_decap_8
XFILLER_26_342 VPWR VGND sg13g2_fill_1
XFILLER_27_876 VPWR VGND sg13g2_decap_8
XFILLER_42_846 VPWR VGND sg13g2_decap_8
XFILLER_14_537 VPWR VGND sg13g2_decap_8
XFILLER_10_754 VPWR VGND sg13g2_decap_8
XFILLER_6_769 VPWR VGND sg13g2_decap_8
XFILLER_5_246 VPWR VGND sg13g2_fill_1
XFILLER_2_986 VPWR VGND sg13g2_decap_8
XFILLER_36_128 VPWR VGND sg13g2_decap_8
XFILLER_36_139 VPWR VGND sg13g2_fill_2
XFILLER_17_353 VPWR VGND sg13g2_decap_8
XFILLER_29_191 VPWR VGND sg13g2_decap_8
XFILLER_44_172 VPWR VGND sg13g2_decap_8
XFILLER_20_529 VPWR VGND sg13g2_decap_4
XFILLER_32_378 VPWR VGND sg13g2_fill_1
X_2711_ _0606_ _0579_ _0608_ VPWR VGND sg13g2_xor2_1
XFILLER_13_581 VPWR VGND sg13g2_decap_8
X_2642_ _0500_ VPWR _0540_ VGND _0453_ _0501_ sg13g2_o21ai_1
X_2573_ _0470_ _0471_ _0465_ _0473_ VPWR VGND sg13g2_nand3_1
X_1524_ _0855_ VPWR _0859_ VGND _0856_ _0857_ sg13g2_o21ai_1
X_3125_ net545 VGND VPWR net130 mac1.sum_lvl1_ff\[12\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_3056_ net532 VGND VPWR _0109_ DP_1.matrix\[79\] clknet_leaf_11_clk sg13g2_dfrbpq_2
X_2007_ _1304_ VPWR _1305_ VGND _1298_ _1301_ sg13g2_o21ai_1
XFILLER_24_802 VPWR VGND sg13g2_decap_8
XFILLER_35_161 VPWR VGND sg13g2_decap_8
XFILLER_35_172 VPWR VGND sg13g2_fill_2
XFILLER_35_194 VPWR VGND sg13g2_fill_2
XFILLER_11_518 VPWR VGND sg13g2_decap_8
XFILLER_23_378 VPWR VGND sg13g2_decap_8
X_2909_ net410 net431 net378 _0798_ VPWR VGND sg13g2_mux2_1
XFILLER_3_717 VPWR VGND sg13g2_decap_8
Xfanout531 net532 net531 VPWR VGND sg13g2_buf_8
Xfanout520 net524 net520 VPWR VGND sg13g2_buf_8
Xfanout542 net543 net542 VPWR VGND sg13g2_buf_8
XFILLER_47_927 VPWR VGND sg13g2_decap_8
XFILLER_19_629 VPWR VGND sg13g2_decap_8
XFILLER_46_448 VPWR VGND sg13g2_decap_8
XFILLER_18_128 VPWR VGND sg13g2_decap_8
XFILLER_42_610 VPWR VGND sg13g2_decap_8
XFILLER_15_879 VPWR VGND sg13g2_decap_8
XFILLER_25_51 VPWR VGND sg13g2_fill_1
XFILLER_26_183 VPWR VGND sg13g2_fill_2
XFILLER_41_142 VPWR VGND sg13g2_fill_1
XFILLER_10_562 VPWR VGND sg13g2_fill_1
XFILLER_6_500 VPWR VGND sg13g2_fill_1
XFILLER_6_544 VPWR VGND sg13g2_fill_2
XFILLER_44_8 VPWR VGND sg13g2_decap_8
XFILLER_29_1025 VPWR VGND sg13g2_decap_4
XFILLER_2_783 VPWR VGND sg13g2_decap_8
XFILLER_49_242 VPWR VGND sg13g2_decap_8
XFILLER_2_11 VPWR VGND sg13g2_decap_8
XFILLER_38_938 VPWR VGND sg13g2_decap_8
XFILLER_37_448 VPWR VGND sg13g2_decap_8
XFILLER_46_960 VPWR VGND sg13g2_decap_8
XFILLER_17_161 VPWR VGND sg13g2_fill_2
XFILLER_18_673 VPWR VGND sg13g2_decap_8
XFILLER_21_805 VPWR VGND sg13g2_decap_8
XFILLER_33_698 VPWR VGND sg13g2_decap_8
X_2625_ VGND VPWR _0520_ _0521_ _0524_ _0503_ sg13g2_a21oi_1
X_2556_ _0456_ _0451_ _0454_ VPWR VGND sg13g2_xnor2_1
X_1507_ _0844_ net417 net472 VPWR VGND sg13g2_nand2_1
X_2487_ _0389_ net489 net429 VPWR VGND sg13g2_nand2_1
XFILLER_29_927 VPWR VGND sg13g2_decap_8
X_3108_ net519 VGND VPWR _0049_ mac1.products_ff\[147\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_44_908 VPWR VGND sg13g2_decap_8
X_3039_ net539 VGND VPWR _0092_ DP_1.matrix\[6\] clknet_leaf_14_clk sg13g2_dfrbpq_2
XFILLER_24_621 VPWR VGND sg13g2_decap_8
XFILLER_23_131 VPWR VGND sg13g2_fill_1
XFILLER_24_643 VPWR VGND sg13g2_decap_8
XFILLER_24_698 VPWR VGND sg13g2_fill_1
XFILLER_8_809 VPWR VGND sg13g2_decap_8
XFILLER_12_849 VPWR VGND sg13g2_decap_8
XFILLER_3_514 VPWR VGND sg13g2_decap_8
XFILLER_11_86 VPWR VGND sg13g2_fill_2
XFILLER_2_4 VPWR VGND sg13g2_decap_8
Xfanout383 net184 net383 VPWR VGND sg13g2_buf_8
Xfanout372 net373 net372 VPWR VGND sg13g2_buf_1
Xfanout394 net395 net394 VPWR VGND sg13g2_buf_2
XFILLER_47_768 VPWR VGND sg13g2_fill_1
XFILLER_35_908 VPWR VGND sg13g2_decap_8
XFILLER_27_481 VPWR VGND sg13g2_decap_8
XFILLER_28_993 VPWR VGND sg13g2_decap_8
XFILLER_34_429 VPWR VGND sg13g2_decap_8
XFILLER_36_50 VPWR VGND sg13g2_decap_8
XFILLER_36_83 VPWR VGND sg13g2_decap_8
XFILLER_43_985 VPWR VGND sg13g2_decap_8
XFILLER_42_473 VPWR VGND sg13g2_fill_2
XFILLER_42_495 VPWR VGND sg13g2_decap_4
Xinput14 uio_in[5] net14 VPWR VGND sg13g2_buf_1
XFILLER_7_875 VPWR VGND sg13g2_decap_8
X_2410_ _0315_ _0293_ _0317_ _0318_ VPWR VGND sg13g2_a21o_1
X_2341_ _0251_ _0244_ _0252_ VPWR VGND sg13g2_nor2b_1
XFILLER_42_1000 VPWR VGND sg13g2_decap_8
XFILLER_2_580 VPWR VGND sg13g2_decap_8
X_2272_ _0183_ _0184_ _0185_ VPWR VGND sg13g2_nor2_1
XFILLER_19_971 VPWR VGND sg13g2_decap_8
XFILLER_34_996 VPWR VGND sg13g2_decap_8
XFILLER_20_112 VPWR VGND sg13g2_decap_8
X_1987_ VGND VPWR _1286_ net175 _1289_ _1287_ sg13g2_a21oi_1
XFILLER_20_156 VPWR VGND sg13g2_decap_8
XFILLER_20_167 VPWR VGND sg13g2_fill_1
X_2608_ VGND VPWR _0507_ _0505_ _0460_ sg13g2_or2_1
XFILLER_0_517 VPWR VGND sg13g2_decap_8
X_2539_ VGND VPWR _0437_ _0438_ _0440_ _0420_ sg13g2_a21oi_1
XFILLER_28_223 VPWR VGND sg13g2_decap_8
XFILLER_29_757 VPWR VGND sg13g2_fill_1
XFILLER_44_716 VPWR VGND sg13g2_fill_2
XFILLER_16_418 VPWR VGND sg13g2_decap_4
XFILLER_43_226 VPWR VGND sg13g2_fill_1
XFILLER_25_941 VPWR VGND sg13g2_decap_8
XFILLER_40_911 VPWR VGND sg13g2_decap_8
XFILLER_12_613 VPWR VGND sg13g2_fill_1
XFILLER_19_1013 VPWR VGND sg13g2_decap_8
XFILLER_24_451 VPWR VGND sg13g2_decap_8
XFILLER_24_495 VPWR VGND sg13g2_decap_8
XFILLER_40_988 VPWR VGND sg13g2_decap_8
XFILLER_7_138 VPWR VGND sg13g2_fill_1
XFILLER_20_690 VPWR VGND sg13g2_fill_1
XFILLER_4_812 VPWR VGND sg13g2_decap_8
XFILLER_3_300 VPWR VGND sg13g2_decap_8
XFILLER_3_344 VPWR VGND sg13g2_decap_8
XFILLER_4_889 VPWR VGND sg13g2_decap_8
XFILLER_26_1028 VPWR VGND sg13g2_fill_1
XFILLER_47_521 VPWR VGND sg13g2_decap_8
XFILLER_47_82 VPWR VGND sg13g2_decap_8
XFILLER_19_256 VPWR VGND sg13g2_decap_8
XFILLER_19_289 VPWR VGND sg13g2_decap_8
XFILLER_34_215 VPWR VGND sg13g2_decap_8
XFILLER_34_226 VPWR VGND sg13g2_fill_1
XFILLER_16_974 VPWR VGND sg13g2_decap_8
X_2890_ DP_2.I_range.out_data\[3\] DP_2.Q_range.out_data\[3\] _0779_ VPWR VGND sg13g2_nor2b_1
XFILLER_43_793 VPWR VGND sg13g2_decap_8
X_1910_ _1226_ VPWR _1229_ VGND _1225_ _1227_ sg13g2_o21ai_1
XFILLER_31_922 VPWR VGND sg13g2_decap_8
XFILLER_8_32 VPWR VGND sg13g2_fill_1
X_1841_ _1166_ _1145_ _1167_ VPWR VGND sg13g2_nor2b_1
XFILLER_30_432 VPWR VGND sg13g2_decap_4
XFILLER_30_465 VPWR VGND sg13g2_decap_4
XFILLER_31_999 VPWR VGND sg13g2_decap_8
XFILLER_11_690 VPWR VGND sg13g2_fill_1
X_1772_ _1100_ _1092_ _1099_ VPWR VGND sg13g2_xnor2_1
XFILLER_7_672 VPWR VGND sg13g2_decap_8
X_2324_ _0208_ _0202_ _0210_ _0235_ VPWR VGND sg13g2_a21o_1
X_2255_ _0167_ _1483_ _0168_ VPWR VGND sg13g2_xor2_1
X_2186_ _1468_ _1448_ _1466_ _1467_ VPWR VGND sg13g2_and3_1
XFILLER_26_716 VPWR VGND sg13g2_decap_4
XFILLER_38_598 VPWR VGND sg13g2_fill_1
XFILLER_43_29 VPWR VGND sg13g2_fill_2
XFILLER_21_421 VPWR VGND sg13g2_decap_8
XFILLER_22_966 VPWR VGND sg13g2_decap_8
XFILLER_21_476 VPWR VGND sg13g2_decap_8
XFILLER_49_1028 VPWR VGND sg13g2_fill_1
XFILLER_13_911 VPWR VGND sg13g2_decap_8
XFILLER_24_270 VPWR VGND sg13g2_fill_2
XFILLER_31_229 VPWR VGND sg13g2_decap_4
XFILLER_40_763 VPWR VGND sg13g2_fill_2
XFILLER_33_40 VPWR VGND sg13g2_decap_8
XFILLER_12_465 VPWR VGND sg13g2_decap_4
XFILLER_13_988 VPWR VGND sg13g2_decap_8
XFILLER_8_447 VPWR VGND sg13g2_decap_8
XFILLER_4_686 VPWR VGND sg13g2_decap_8
XFILLER_0_881 VPWR VGND sg13g2_decap_8
Xhold3 mac1.products_ff\[75\] VPWR VGND net43 sg13g2_dlygate4sd3_1
XFILLER_48_863 VPWR VGND sg13g2_decap_8
X_2040_ _1328_ net232 _1323_ _1332_ VPWR VGND sg13g2_nand3_1
XFILLER_47_395 VPWR VGND sg13g2_decap_4
XFILLER_23_708 VPWR VGND sg13g2_decap_4
XFILLER_16_782 VPWR VGND sg13g2_decap_8
XFILLER_22_218 VPWR VGND sg13g2_fill_1
XFILLER_31_730 VPWR VGND sg13g2_decap_8
X_2942_ _0756_ _0738_ _0825_ VPWR VGND sg13g2_xor2_1
XFILLER_31_774 VPWR VGND sg13g2_decap_8
X_2873_ net461 net478 _0730_ _0763_ VPWR VGND sg13g2_mux2_1
X_1824_ _1130_ VPWR _1150_ VGND _1128_ _1131_ sg13g2_o21ai_1
XFILLER_8_970 VPWR VGND sg13g2_decap_8
X_1755_ _1083_ net467 net401 VPWR VGND sg13g2_nand2_1
X_1686_ _1016_ _1009_ _1014_ _1015_ VPWR VGND sg13g2_and3_1
X_2307_ _0214_ VPWR _0219_ VGND _0216_ _0217_ sg13g2_o21ai_1
XFILLER_38_29 VPWR VGND sg13g2_decap_8
X_2238_ _1446_ _0149_ _0151_ _0152_ VPWR VGND sg13g2_or3_1
XFILLER_38_340 VPWR VGND sg13g2_decap_8
XFILLER_38_362 VPWR VGND sg13g2_decap_4
X_2169_ _1451_ net448 net388 VPWR VGND sg13g2_nand2_1
XFILLER_26_535 VPWR VGND sg13g2_decap_8
XFILLER_38_384 VPWR VGND sg13g2_fill_2
XFILLER_26_568 VPWR VGND sg13g2_decap_8
XFILLER_41_527 VPWR VGND sg13g2_decap_8
XFILLER_16_1016 VPWR VGND sg13g2_decap_8
XFILLER_22_752 VPWR VGND sg13g2_decap_4
XFILLER_10_936 VPWR VGND sg13g2_decap_8
XFILLER_16_1027 VPWR VGND sg13g2_fill_2
XFILLER_21_262 VPWR VGND sg13g2_decap_8
XFILLER_5_417 VPWR VGND sg13g2_decap_4
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_1_667 VPWR VGND sg13g2_decap_8
XFILLER_48_104 VPWR VGND sg13g2_decap_4
XFILLER_0_155 VPWR VGND sg13g2_decap_8
XFILLER_45_844 VPWR VGND sg13g2_decap_8
XFILLER_29_384 VPWR VGND sg13g2_fill_1
XFILLER_44_61 VPWR VGND sg13g2_decap_8
XFILLER_8_200 VPWR VGND sg13g2_fill_1
XFILLER_13_785 VPWR VGND sg13g2_fill_2
XFILLER_9_767 VPWR VGND sg13g2_decap_8
XFILLER_5_951 VPWR VGND sg13g2_decap_8
X_1540_ _0874_ net466 net418 net468 net412 VPWR VGND sg13g2_a22oi_1
XFILLER_5_99 VPWR VGND sg13g2_decap_8
X_3210_ net505 VGND VPWR net89 mac1.sum_lvl3_ff\[21\] clknet_leaf_37_clk sg13g2_dfrbpq_1
X_3141_ net540 VGND VPWR net53 mac1.sum_lvl1_ff\[48\] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_3072_ net548 VGND VPWR _0125_ DP_2.matrix\[43\] clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_47_181 VPWR VGND sg13g2_decap_8
X_2023_ _1318_ _1315_ _1317_ VPWR VGND sg13g2_nand2_1
XFILLER_39_1027 VPWR VGND sg13g2_fill_2
XFILLER_39_1016 VPWR VGND sg13g2_decap_8
XFILLER_35_354 VPWR VGND sg13g2_fill_1
X_2925_ DP_2.I_range.out_data\[6\] DP_2.I_range.out_data\[5\] _0814_ VPWR VGND sg13g2_nor2b_1
X_2856_ _0743_ _0744_ _0745_ _0746_ VPWR VGND sg13g2_nor3_1
X_1807_ _1133_ _1126_ _1134_ VPWR VGND sg13g2_nor2b_1
X_2787_ _0681_ net477 net422 VPWR VGND sg13g2_nand2_1
Xhold200 _1303_ VPWR VGND net240 sg13g2_dlygate4sd3_1
Xhold211 _0088_ VPWR VGND net251 sg13g2_dlygate4sd3_1
Xhold222 _1299_ VPWR VGND net262 sg13g2_dlygate4sd3_1
Xhold244 _1246_ VPWR VGND net284 sg13g2_dlygate4sd3_1
X_1738_ _1067_ _1052_ _1066_ VPWR VGND sg13g2_nand2_1
Xhold233 DP_2.matrix\[75\] VPWR VGND net273 sg13g2_dlygate4sd3_1
XFILLER_49_28 VPWR VGND sg13g2_decap_8
XFILLER_46_1009 VPWR VGND sg13g2_decap_8
Xhold255 _1256_ VPWR VGND net295 sg13g2_dlygate4sd3_1
X_1669_ _0999_ _0991_ _0998_ VPWR VGND sg13g2_nand2_1
XFILLER_39_660 VPWR VGND sg13g2_decap_8
XFILLER_27_822 VPWR VGND sg13g2_decap_8
XFILLER_27_855 VPWR VGND sg13g2_decap_8
XFILLER_38_181 VPWR VGND sg13g2_decap_8
XFILLER_42_836 VPWR VGND sg13g2_fill_1
XFILLER_41_324 VPWR VGND sg13g2_decap_8
XFILLER_26_398 VPWR VGND sg13g2_decap_4
XFILLER_41_357 VPWR VGND sg13g2_decap_8
XFILLER_41_368 VPWR VGND sg13g2_fill_1
XFILLER_14_42 VPWR VGND sg13g2_decap_8
XFILLER_10_733 VPWR VGND sg13g2_decap_8
XFILLER_6_748 VPWR VGND sg13g2_decap_8
XFILLER_30_96 VPWR VGND sg13g2_decap_8
XFILLER_2_965 VPWR VGND sg13g2_decap_8
XFILLER_49_435 VPWR VGND sg13g2_decap_8
XFILLER_39_83 VPWR VGND sg13g2_decap_8
XFILLER_49_479 VPWR VGND sg13g2_decap_8
XFILLER_18_888 VPWR VGND sg13g2_decap_8
XFILLER_32_346 VPWR VGND sg13g2_fill_2
XFILLER_32_357 VPWR VGND sg13g2_decap_8
XFILLER_13_560 VPWR VGND sg13g2_decap_8
X_2710_ _0607_ _0606_ _0579_ VPWR VGND sg13g2_nand2b_1
X_2641_ _0528_ VPWR _0539_ VGND _0455_ _0529_ sg13g2_o21ai_1
X_2572_ _0472_ _0465_ _0470_ _0471_ VPWR VGND sg13g2_and3_1
X_1523_ _0855_ _0856_ _0857_ _0858_ VPWR VGND sg13g2_nor3_1
X_3124_ net544 VGND VPWR net45 mac1.sum_lvl1_ff\[11\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_3055_ net532 VGND VPWR _0108_ DP_1.matrix\[78\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_36_630 VPWR VGND sg13g2_decap_8
X_2006_ net239 net287 _1304_ VPWR VGND sg13g2_xor2_1
XFILLER_23_302 VPWR VGND sg13g2_fill_2
XFILLER_36_685 VPWR VGND sg13g2_decap_8
X_2908_ _0792_ _0796_ _0797_ VPWR VGND sg13g2_nor2b_1
X_2839_ _0729_ DP_1.I_range.out_data\[2\] DP_1.Q_range.out_data\[2\] VPWR VGND sg13g2_nand2b_1
XFILLER_4_8 VPWR VGND sg13g2_fill_2
Xfanout510 net513 net510 VPWR VGND sg13g2_buf_8
Xfanout521 net524 net521 VPWR VGND sg13g2_buf_8
Xfanout532 net533 net532 VPWR VGND sg13g2_buf_8
XFILLER_47_906 VPWR VGND sg13g2_decap_8
Xfanout543 net549 net543 VPWR VGND sg13g2_buf_8
XFILLER_46_405 VPWR VGND sg13g2_decap_8
XFILLER_39_490 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_38_clk clknet_3_0__leaf_clk clknet_leaf_38_clk VPWR VGND sg13g2_buf_8
XFILLER_27_641 VPWR VGND sg13g2_decap_8
XFILLER_26_173 VPWR VGND sg13g2_decap_4
XFILLER_15_858 VPWR VGND sg13g2_decap_8
XFILLER_42_699 VPWR VGND sg13g2_decap_8
XFILLER_42_666 VPWR VGND sg13g2_decap_8
XFILLER_14_368 VPWR VGND sg13g2_decap_8
XFILLER_14_379 VPWR VGND sg13g2_fill_1
XFILLER_25_74 VPWR VGND sg13g2_fill_1
XFILLER_23_891 VPWR VGND sg13g2_decap_8
XFILLER_6_556 VPWR VGND sg13g2_decap_8
XFILLER_6_589 VPWR VGND sg13g2_decap_8
XFILLER_29_1004 VPWR VGND sg13g2_decap_8
XFILLER_2_762 VPWR VGND sg13g2_decap_8
XFILLER_49_221 VPWR VGND sg13g2_decap_8
XFILLER_1_272 VPWR VGND sg13g2_fill_2
XFILLER_38_917 VPWR VGND sg13g2_decap_8
XFILLER_49_298 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_29_clk clknet_3_5__leaf_clk clknet_leaf_29_clk VPWR VGND sg13g2_buf_8
XFILLER_17_140 VPWR VGND sg13g2_fill_2
XFILLER_17_184 VPWR VGND sg13g2_decap_8
XFILLER_33_633 VPWR VGND sg13g2_decap_8
XFILLER_36_1019 VPWR VGND sg13g2_decap_8
XFILLER_14_891 VPWR VGND sg13g2_decap_8
XFILLER_32_176 VPWR VGND sg13g2_fill_2
X_2624_ _0520_ _0521_ _0503_ _0523_ VPWR VGND sg13g2_nand3_1
X_2555_ _0455_ _0451_ _0454_ VPWR VGND sg13g2_nand2_1
X_1506_ _0843_ net474 net410 VPWR VGND sg13g2_nand2_1
X_2486_ _0388_ net489 net427 VPWR VGND sg13g2_nand2_1
XFILLER_29_906 VPWR VGND sg13g2_decap_8
X_3107_ net511 VGND VPWR _0048_ mac1.products_ff\[146\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_28_438 VPWR VGND sg13g2_decap_8
X_3038_ net539 VGND VPWR _0091_ DP_1.matrix\[5\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_36_460 VPWR VGND sg13g2_fill_1
XFILLER_37_994 VPWR VGND sg13g2_decap_8
XFILLER_12_828 VPWR VGND sg13g2_decap_8
XFILLER_23_165 VPWR VGND sg13g2_decap_8
XFILLER_11_327 VPWR VGND sg13g2_fill_2
XFILLER_20_883 VPWR VGND sg13g2_decap_8
XFILLER_11_65 VPWR VGND sg13g2_decap_8
Xfanout373 _0770_ net373 VPWR VGND sg13g2_buf_2
Xfanout384 net385 net384 VPWR VGND sg13g2_buf_8
XFILLER_46_202 VPWR VGND sg13g2_decap_8
Xfanout395 net396 net395 VPWR VGND sg13g2_buf_1
XFILLER_19_449 VPWR VGND sg13g2_fill_1
XFILLER_15_600 VPWR VGND sg13g2_decap_8
XFILLER_27_460 VPWR VGND sg13g2_fill_2
XFILLER_28_972 VPWR VGND sg13g2_decap_8
XFILLER_43_964 VPWR VGND sg13g2_decap_8
XFILLER_14_143 VPWR VGND sg13g2_decap_8
XFILLER_15_655 VPWR VGND sg13g2_decap_8
Xinput15 uio_in[6] net15 VPWR VGND sg13g2_buf_1
XFILLER_7_854 VPWR VGND sg13g2_decap_8
X_2340_ _0251_ _0245_ _0250_ VPWR VGND sg13g2_xnor2_1
X_2271_ _0184_ net391 net440 net396 net496 VPWR VGND sg13g2_a22oi_1
XFILLER_28_4 VPWR VGND sg13g2_fill_2
XFILLER_19_950 VPWR VGND sg13g2_decap_8
XFILLER_26_909 VPWR VGND sg13g2_decap_8
XFILLER_37_257 VPWR VGND sg13g2_decap_8
XFILLER_33_430 VPWR VGND sg13g2_fill_1
XFILLER_34_975 VPWR VGND sg13g2_decap_8
XFILLER_21_625 VPWR VGND sg13g2_decap_8
XFILLER_21_647 VPWR VGND sg13g2_fill_1
X_1986_ net175 _1286_ _0024_ VPWR VGND sg13g2_xor2_1
Xclkbuf_leaf_9_clk clknet_3_2__leaf_clk clknet_leaf_9_clk VPWR VGND sg13g2_buf_8
XFILLER_9_191 VPWR VGND sg13g2_decap_8
X_2607_ _0506_ net482 net429 VPWR VGND sg13g2_nand2_1
X_2538_ _0437_ _0438_ _0420_ _0439_ VPWR VGND sg13g2_nand3_1
X_2469_ net439 net486 net485 net436 _0372_ VPWR VGND sg13g2_and4_1
XFILLER_29_725 VPWR VGND sg13g2_decap_8
XFILLER_43_216 VPWR VGND sg13g2_decap_4
XFILLER_25_920 VPWR VGND sg13g2_decap_8
XFILLER_28_279 VPWR VGND sg13g2_decap_8
XFILLER_37_780 VPWR VGND sg13g2_fill_2
XFILLER_43_238 VPWR VGND sg13g2_decap_8
XFILLER_24_430 VPWR VGND sg13g2_decap_8
XFILLER_11_113 VPWR VGND sg13g2_decap_8
XFILLER_25_997 VPWR VGND sg13g2_decap_8
XFILLER_40_967 VPWR VGND sg13g2_decap_8
XFILLER_8_629 VPWR VGND sg13g2_fill_2
XFILLER_8_618 VPWR VGND sg13g2_decap_8
XFILLER_22_42 VPWR VGND sg13g2_fill_2
XFILLER_4_868 VPWR VGND sg13g2_decap_8
XFILLER_26_1007 VPWR VGND sg13g2_decap_8
XFILLER_19_279 VPWR VGND sg13g2_fill_1
XFILLER_16_953 VPWR VGND sg13g2_decap_8
XFILLER_31_901 VPWR VGND sg13g2_decap_8
XFILLER_42_260 VPWR VGND sg13g2_decap_8
XFILLER_15_496 VPWR VGND sg13g2_decap_8
Xclkbuf_3_4__f_clk clknet_0_clk clknet_3_4__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_8_22 VPWR VGND sg13g2_decap_4
X_1840_ _1164_ _1163_ _1166_ VPWR VGND sg13g2_xor2_1
XFILLER_31_978 VPWR VGND sg13g2_decap_8
XFILLER_8_66 VPWR VGND sg13g2_decap_4
XFILLER_8_77 VPWR VGND sg13g2_decap_8
X_1771_ _1097_ _1098_ _1099_ VPWR VGND sg13g2_nor2b_1
XFILLER_10_190 VPWR VGND sg13g2_decap_4
X_2323_ _0233_ _0231_ _0048_ VPWR VGND sg13g2_xor2_1
X_2254_ _0167_ net451 net382 VPWR VGND sg13g2_nand2_1
XFILLER_38_500 VPWR VGND sg13g2_fill_2
X_2185_ _1455_ VPWR _1467_ VGND _1463_ _1465_ sg13g2_o21ai_1
XFILLER_38_577 VPWR VGND sg13g2_decap_8
XFILLER_25_238 VPWR VGND sg13g2_decap_4
XFILLER_40_208 VPWR VGND sg13g2_decap_8
XFILLER_21_400 VPWR VGND sg13g2_decap_8
XFILLER_22_945 VPWR VGND sg13g2_decap_8
XFILLER_34_794 VPWR VGND sg13g2_fill_1
X_1969_ VGND VPWR mac1.sum_lvl2_ff\[32\] mac1.sum_lvl2_ff\[13\] _1276_ _1274_ sg13g2_a21oi_1
XFILLER_49_1007 VPWR VGND sg13g2_decap_8
XFILLER_1_849 VPWR VGND sg13g2_decap_8
XFILLER_44_514 VPWR VGND sg13g2_decap_8
XFILLER_17_717 VPWR VGND sg13g2_decap_4
XFILLER_29_588 VPWR VGND sg13g2_decap_8
XFILLER_44_547 VPWR VGND sg13g2_decap_8
XFILLER_17_53 VPWR VGND sg13g2_decap_8
XFILLER_44_558 VPWR VGND sg13g2_fill_1
XFILLER_32_709 VPWR VGND sg13g2_fill_2
XFILLER_40_742 VPWR VGND sg13g2_decap_8
XFILLER_13_967 VPWR VGND sg13g2_decap_8
XFILLER_40_797 VPWR VGND sg13g2_fill_2
XFILLER_9_949 VPWR VGND sg13g2_decap_8
XFILLER_32_1011 VPWR VGND sg13g2_decap_8
XFILLER_4_665 VPWR VGND sg13g2_decap_8
Xhold4 mac1.sum_lvl1_ff\[6\] VPWR VGND net44 sg13g2_dlygate4sd3_1
XFILLER_0_860 VPWR VGND sg13g2_decap_8
XFILLER_48_842 VPWR VGND sg13g2_decap_8
XFILLER_47_330 VPWR VGND sg13g2_decap_8
XFILLER_35_547 VPWR VGND sg13g2_decap_8
XFILLER_16_761 VPWR VGND sg13g2_decap_8
XFILLER_43_580 VPWR VGND sg13g2_fill_2
XFILLER_16_772 VPWR VGND sg13g2_fill_1
X_2941_ VGND VPWR net371 _0824_ _0090_ _0823_ sg13g2_a21oi_1
XFILLER_43_591 VPWR VGND sg13g2_fill_2
XFILLER_31_742 VPWR VGND sg13g2_fill_1
XFILLER_30_252 VPWR VGND sg13g2_decap_8
X_2872_ _0757_ _0761_ _0762_ VPWR VGND sg13g2_nor2b_1
X_1823_ _1149_ _1148_ _1146_ VPWR VGND sg13g2_nand2b_1
X_1754_ _1082_ net471 net494 VPWR VGND sg13g2_nand2_1
X_1685_ _1010_ VPWR _1015_ VGND _1011_ _1013_ sg13g2_o21ai_1
X_2306_ _0214_ _0216_ _0217_ _0218_ VPWR VGND sg13g2_nor3_1
X_2237_ VGND VPWR _0147_ _0148_ _0151_ _1480_ sg13g2_a21oi_1
XFILLER_39_897 VPWR VGND sg13g2_decap_8
X_2168_ _1450_ net447 net386 VPWR VGND sg13g2_nand2_1
X_2099_ _1383_ net458 net384 VPWR VGND sg13g2_nand2_1
XFILLER_22_731 VPWR VGND sg13g2_decap_8
XFILLER_10_915 VPWR VGND sg13g2_decap_8
XFILLER_21_241 VPWR VGND sg13g2_decap_8
XFILLER_21_252 VPWR VGND sg13g2_fill_1
XFILLER_21_296 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_1_646 VPWR VGND sg13g2_decap_8
XFILLER_17_503 VPWR VGND sg13g2_decap_4
XFILLER_45_823 VPWR VGND sg13g2_decap_8
XFILLER_44_322 VPWR VGND sg13g2_decap_8
XFILLER_44_40 VPWR VGND sg13g2_decap_8
XFILLER_12_241 VPWR VGND sg13g2_decap_8
XFILLER_40_583 VPWR VGND sg13g2_fill_1
XFILLER_9_746 VPWR VGND sg13g2_decap_8
XFILLER_8_234 VPWR VGND sg13g2_fill_2
XFILLER_8_223 VPWR VGND sg13g2_decap_8
XFILLER_8_278 VPWR VGND sg13g2_decap_4
XFILLER_8_256 VPWR VGND sg13g2_decap_4
XFILLER_5_930 VPWR VGND sg13g2_decap_8
XFILLER_5_34 VPWR VGND sg13g2_decap_4
XFILLER_5_56 VPWR VGND sg13g2_decap_8
XFILLER_4_473 VPWR VGND sg13g2_decap_4
X_3140_ net540 VGND VPWR net67 mac1.sum_lvl1_ff\[47\] clknet_leaf_23_clk sg13g2_dfrbpq_1
XFILLER_48_661 VPWR VGND sg13g2_fill_2
X_3071_ net548 VGND VPWR _0124_ DP_2.matrix\[42\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_10_4 VPWR VGND sg13g2_decap_8
X_2022_ net213 net206 _1317_ VPWR VGND sg13g2_xor2_1
XFILLER_23_506 VPWR VGND sg13g2_fill_2
XFILLER_16_580 VPWR VGND sg13g2_fill_2
X_2924_ DP_2.I_range.out_data\[2\] DP_2.I_range.out_data\[4\] _0813_ VPWR VGND sg13g2_nor2_1
X_2855_ net490 _0728_ _0731_ _0745_ VPWR VGND sg13g2_nor3_1
X_1806_ _1133_ _1127_ _1132_ VPWR VGND sg13g2_xnor2_1
X_2786_ _0680_ net482 net495 VPWR VGND sg13g2_nand2_1
Xhold201 _1310_ VPWR VGND net241 sg13g2_dlygate4sd3_1
Xhold212 DP_2.matrix\[7\] VPWR VGND net252 sg13g2_dlygate4sd3_1
Xhold223 _1302_ VPWR VGND net263 sg13g2_dlygate4sd3_1
X_1737_ _1065_ _1058_ _1066_ VPWR VGND sg13g2_xor2_1
Xhold234 DP_1.matrix\[43\] VPWR VGND net274 sg13g2_dlygate4sd3_1
Xhold256 mac1.sum_lvl2_ff\[6\] VPWR VGND net296 sg13g2_dlygate4sd3_1
Xhold245 _0014_ VPWR VGND net285 sg13g2_dlygate4sd3_1
X_1668_ _0996_ _0992_ _0998_ VPWR VGND sg13g2_xor2_1
X_1599_ net414 net464 net419 _0931_ VPWR VGND net463 sg13g2_nand4_1
X_3269_ net516 VGND VPWR net11 DP_2.Q_range.out_data\[4\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_14_87 VPWR VGND sg13g2_decap_8
XFILLER_6_727 VPWR VGND sg13g2_decap_8
XFILLER_5_204 VPWR VGND sg13g2_decap_8
XFILLER_10_789 VPWR VGND sg13g2_decap_8
XFILLER_5_215 VPWR VGND sg13g2_fill_2
XFILLER_30_53 VPWR VGND sg13g2_decap_8
XFILLER_2_944 VPWR VGND sg13g2_decap_8
XFILLER_49_414 VPWR VGND sg13g2_decap_8
XFILLER_7_1015 VPWR VGND sg13g2_decap_8
XFILLER_39_40 VPWR VGND sg13g2_decap_4
XFILLER_49_458 VPWR VGND sg13g2_decap_8
XFILLER_39_62 VPWR VGND sg13g2_decap_8
XFILLER_18_801 VPWR VGND sg13g2_decap_8
XFILLER_45_642 VPWR VGND sg13g2_decap_4
XFILLER_18_867 VPWR VGND sg13g2_decap_8
XFILLER_33_804 VPWR VGND sg13g2_decap_8
XFILLER_17_388 VPWR VGND sg13g2_decap_8
XFILLER_20_509 VPWR VGND sg13g2_decap_8
XFILLER_41_892 VPWR VGND sg13g2_decap_8
XFILLER_40_391 VPWR VGND sg13g2_fill_2
XFILLER_9_554 VPWR VGND sg13g2_fill_2
X_2640_ _0538_ _0533_ _0537_ VPWR VGND sg13g2_nand2_1
X_2571_ _0466_ VPWR _0471_ VGND _0467_ _0469_ sg13g2_o21ai_1
X_1522_ _0857_ net468 net417 net413 net470 VPWR VGND sg13g2_a22oi_1
X_3123_ net544 VGND VPWR net151 mac1.sum_lvl1_ff\[10\] clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_27_119 VPWR VGND sg13g2_decap_8
X_3054_ net519 VGND VPWR _0107_ DP_1.matrix\[77\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2005_ _1303_ mac1.sum_lvl3_ff\[7\] net239 VPWR VGND sg13g2_nand2_1
XFILLER_24_837 VPWR VGND sg13g2_decap_8
XFILLER_35_196 VPWR VGND sg13g2_fill_1
XFILLER_32_892 VPWR VGND sg13g2_decap_8
X_2907_ _0795_ VPWR _0796_ VGND _0793_ _0794_ sg13g2_o21ai_1
XFILLER_13_1009 VPWR VGND sg13g2_decap_8
X_2838_ _0728_ DP_1.I_range.out_data\[3\] DP_1.Q_range.out_data\[3\] VPWR VGND sg13g2_xnor2_1
X_2769_ VGND VPWR _0664_ _0663_ _0651_ sg13g2_or2_1
XFILLER_2_218 VPWR VGND sg13g2_fill_2
Xfanout500 net501 net500 VPWR VGND sg13g2_buf_8
Xfanout533 rst_n net533 VPWR VGND sg13g2_buf_8
Xfanout511 net513 net511 VPWR VGND sg13g2_buf_8
Xfanout522 net524 net522 VPWR VGND sg13g2_buf_8
Xfanout544 net546 net544 VPWR VGND sg13g2_buf_8
XFILLER_27_620 VPWR VGND sg13g2_decap_8
XFILLER_15_837 VPWR VGND sg13g2_decap_8
XFILLER_25_31 VPWR VGND sg13g2_decap_8
XFILLER_23_870 VPWR VGND sg13g2_decap_8
XFILLER_30_829 VPWR VGND sg13g2_decap_8
XFILLER_6_524 VPWR VGND sg13g2_decap_4
XFILLER_6_546 VPWR VGND sg13g2_fill_1
XFILLER_2_741 VPWR VGND sg13g2_decap_8
XFILLER_49_200 VPWR VGND sg13g2_decap_8
XFILLER_49_277 VPWR VGND sg13g2_decap_8
XFILLER_37_428 VPWR VGND sg13g2_fill_2
XFILLER_46_995 VPWR VGND sg13g2_decap_8
XFILLER_17_163 VPWR VGND sg13g2_fill_1
XFILLER_45_494 VPWR VGND sg13g2_decap_8
XFILLER_33_656 VPWR VGND sg13g2_decap_8
XFILLER_33_678 VPWR VGND sg13g2_decap_8
XFILLER_14_870 VPWR VGND sg13g2_decap_8
XFILLER_13_391 VPWR VGND sg13g2_decap_8
X_2623_ _0522_ _0503_ _0520_ _0521_ VPWR VGND sg13g2_and3_1
X_2554_ _0452_ _0453_ _0454_ VPWR VGND sg13g2_nor2b_1
XFILLER_49_0 VPWR VGND sg13g2_decap_8
X_1505_ VPWR DP_1.Q_range.data_plus_4\[6\] net8 VGND sg13g2_inv_1
X_2485_ _0387_ net492 net426 VPWR VGND sg13g2_nand2_1
X_3106_ net511 VGND VPWR _0057_ mac1.products_ff\[145\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_43_409 VPWR VGND sg13g2_decap_8
X_3037_ net539 VGND VPWR _0090_ DP_1.matrix\[4\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_37_973 VPWR VGND sg13g2_decap_8
XFILLER_36_494 VPWR VGND sg13g2_fill_2
XFILLER_12_807 VPWR VGND sg13g2_decap_8
XFILLER_23_144 VPWR VGND sg13g2_decap_8
XFILLER_24_667 VPWR VGND sg13g2_fill_2
XFILLER_24_689 VPWR VGND sg13g2_decap_8
XFILLER_11_11 VPWR VGND sg13g2_fill_2
XFILLER_3_549 VPWR VGND sg13g2_decap_4
Xfanout374 _0815_ net374 VPWR VGND sg13g2_buf_8
XFILLER_47_737 VPWR VGND sg13g2_fill_2
Xfanout385 net177 net385 VPWR VGND sg13g2_buf_8
Xfanout396 DP_2.matrix\[73\] net396 VPWR VGND sg13g2_buf_8
XFILLER_28_951 VPWR VGND sg13g2_decap_8
XFILLER_43_943 VPWR VGND sg13g2_decap_8
XFILLER_14_188 VPWR VGND sg13g2_fill_2
XFILLER_30_626 VPWR VGND sg13g2_fill_2
XFILLER_35_1020 VPWR VGND sg13g2_decap_8
XFILLER_30_648 VPWR VGND sg13g2_decap_8
Xinput16 uio_in[7] net16 VPWR VGND sg13g2_buf_1
XFILLER_7_833 VPWR VGND sg13g2_decap_8
XFILLER_11_884 VPWR VGND sg13g2_decap_8
XFILLER_6_376 VPWR VGND sg13g2_fill_1
XFILLER_6_365 VPWR VGND sg13g2_decap_8
X_2270_ net440 net496 net396 net390 _0183_ VPWR VGND sg13g2_and4_1
XFILLER_18_483 VPWR VGND sg13g2_decap_8
XFILLER_34_954 VPWR VGND sg13g2_decap_8
XFILLER_33_497 VPWR VGND sg13g2_decap_8
X_1985_ net174 mac1.sum_lvl3_ff\[2\] _1288_ VPWR VGND sg13g2_xor2_1
X_2606_ _0505_ net482 net427 VPWR VGND sg13g2_nand2_2
X_2537_ _0436_ _0435_ _0426_ _0438_ VPWR VGND sg13g2_a21o_1
X_2468_ _0371_ net488 net431 VPWR VGND sg13g2_nand2_1
XFILLER_29_704 VPWR VGND sg13g2_decap_4
X_2399_ _0308_ _0281_ _0306_ VPWR VGND sg13g2_xnor2_1
XFILLER_29_748 VPWR VGND sg13g2_decap_8
XFILLER_44_718 VPWR VGND sg13g2_fill_1
XFILLER_28_258 VPWR VGND sg13g2_decap_8
XFILLER_37_792 VPWR VGND sg13g2_fill_2
XFILLER_25_976 VPWR VGND sg13g2_decap_8
XFILLER_40_946 VPWR VGND sg13g2_decap_8
XFILLER_24_475 VPWR VGND sg13g2_decap_8
XFILLER_7_129 VPWR VGND sg13g2_decap_8
XFILLER_11_158 VPWR VGND sg13g2_fill_2
XFILLER_4_847 VPWR VGND sg13g2_decap_8
XFILLER_47_545 VPWR VGND sg13g2_fill_2
XFILLER_19_236 VPWR VGND sg13g2_decap_4
XFILLER_47_589 VPWR VGND sg13g2_decap_8
XFILLER_28_770 VPWR VGND sg13g2_decap_4
XFILLER_16_932 VPWR VGND sg13g2_decap_8
XFILLER_27_280 VPWR VGND sg13g2_decap_8
XFILLER_28_792 VPWR VGND sg13g2_decap_8
XFILLER_34_239 VPWR VGND sg13g2_decap_8
XFILLER_43_762 VPWR VGND sg13g2_decap_8
XFILLER_43_740 VPWR VGND sg13g2_fill_2
XFILLER_15_464 VPWR VGND sg13g2_fill_2
XFILLER_15_475 VPWR VGND sg13g2_decap_8
XFILLER_30_401 VPWR VGND sg13g2_decap_4
XFILLER_31_957 VPWR VGND sg13g2_decap_8
XFILLER_8_45 VPWR VGND sg13g2_decap_8
X_1770_ _1093_ VPWR _1098_ VGND _1095_ _1096_ sg13g2_o21ai_1
XFILLER_6_162 VPWR VGND sg13g2_decap_8
XFILLER_40_4 VPWR VGND sg13g2_decap_4
X_2322_ _0231_ _0233_ _0234_ VPWR VGND sg13g2_nor2_1
X_2253_ _0166_ net451 net380 VPWR VGND sg13g2_nand2_1
X_2184_ _1455_ _1463_ _1465_ _1466_ VPWR VGND sg13g2_or3_1
XFILLER_25_217 VPWR VGND sg13g2_decap_8
XFILLER_18_291 VPWR VGND sg13g2_decap_8
XFILLER_34_762 VPWR VGND sg13g2_decap_8
XFILLER_22_924 VPWR VGND sg13g2_decap_8
XFILLER_33_294 VPWR VGND sg13g2_decap_8
X_1968_ _1274_ net280 _0004_ VPWR VGND sg13g2_nor2b_2
XFILLER_30_990 VPWR VGND sg13g2_decap_8
X_1899_ _1222_ _1219_ _1221_ VPWR VGND sg13g2_xnor2_1
XFILLER_0_305 VPWR VGND sg13g2_decap_8
XFILLER_1_828 VPWR VGND sg13g2_decap_8
XFILLER_0_349 VPWR VGND sg13g2_decap_8
XFILLER_29_501 VPWR VGND sg13g2_decap_8
XFILLER_29_545 VPWR VGND sg13g2_fill_2
XFILLER_29_534 VPWR VGND sg13g2_decap_8
XFILLER_17_32 VPWR VGND sg13g2_decap_8
XFILLER_29_567 VPWR VGND sg13g2_decap_8
XFILLER_17_98 VPWR VGND sg13g2_fill_1
XFILLER_12_423 VPWR VGND sg13g2_decap_8
XFILLER_12_434 VPWR VGND sg13g2_fill_2
XFILLER_13_946 VPWR VGND sg13g2_decap_8
XFILLER_40_765 VPWR VGND sg13g2_fill_1
XFILLER_9_928 VPWR VGND sg13g2_decap_8
XFILLER_33_97 VPWR VGND sg13g2_decap_8
XFILLER_4_644 VPWR VGND sg13g2_decap_8
XFILLER_3_132 VPWR VGND sg13g2_fill_2
XFILLER_48_821 VPWR VGND sg13g2_decap_8
XFILLER_12_8 VPWR VGND sg13g2_fill_1
Xhold5 mac1.products_ff\[11\] VPWR VGND net45 sg13g2_dlygate4sd3_1
XFILLER_48_898 VPWR VGND sg13g2_decap_8
XFILLER_16_740 VPWR VGND sg13g2_decap_8
XFILLER_22_209 VPWR VGND sg13g2_decap_8
X_2940_ _0755_ _0751_ _0824_ VPWR VGND sg13g2_xor2_1
X_2871_ _0758_ VPWR _0761_ VGND _0759_ _0760_ sg13g2_o21ai_1
X_1822_ VGND VPWR _1148_ _1147_ _1094_ sg13g2_or2_1
X_1753_ _1055_ VPWR _1081_ VGND _1053_ _1056_ sg13g2_o21ai_1
X_1684_ _1010_ _1011_ _1013_ _1014_ VPWR VGND sg13g2_or3_1
XFILLER_31_0 VPWR VGND sg13g2_fill_2
X_2305_ _0217_ net387 net443 net389 net441 VPWR VGND sg13g2_a22oi_1
X_2236_ _0147_ _0148_ _1480_ _0150_ VPWR VGND sg13g2_nand3_1
XFILLER_39_876 VPWR VGND sg13g2_decap_8
XFILLER_26_504 VPWR VGND sg13g2_fill_2
X_2167_ _1449_ net453 net384 VPWR VGND sg13g2_nand2_1
XFILLER_0_1021 VPWR VGND sg13g2_decap_8
X_2098_ _1373_ VPWR _1382_ VGND _1365_ _1374_ sg13g2_o21ai_1
XFILLER_22_710 VPWR VGND sg13g2_decap_8
XFILLER_34_581 VPWR VGND sg13g2_decap_8
XFILLER_6_909 VPWR VGND sg13g2_decap_8
XFILLER_1_625 VPWR VGND sg13g2_decap_8
XFILLER_28_20 VPWR VGND sg13g2_fill_2
XFILLER_45_802 VPWR VGND sg13g2_decap_8
XFILLER_28_42 VPWR VGND sg13g2_decap_8
XFILLER_17_526 VPWR VGND sg13g2_decap_8
XFILLER_45_879 VPWR VGND sg13g2_decap_8
XFILLER_32_507 VPWR VGND sg13g2_fill_1
XFILLER_40_551 VPWR VGND sg13g2_fill_2
XFILLER_9_725 VPWR VGND sg13g2_decap_8
XFILLER_12_231 VPWR VGND sg13g2_fill_1
XFILLER_13_754 VPWR VGND sg13g2_decap_4
XFILLER_13_787 VPWR VGND sg13g2_fill_1
XFILLER_5_986 VPWR VGND sg13g2_decap_8
X_3070_ net548 VGND VPWR _0123_ DP_2.matrix\[41\] clknet_leaf_21_clk sg13g2_dfrbpq_2
XFILLER_39_117 VPWR VGND sg13g2_decap_8
X_2021_ _1316_ net206 mac1.sum_lvl3_ff\[30\] VPWR VGND sg13g2_nand2_1
XFILLER_36_879 VPWR VGND sg13g2_decap_8
X_2923_ _0811_ _0809_ _0812_ VPWR VGND sg13g2_xor2_1
XFILLER_31_562 VPWR VGND sg13g2_decap_8
X_2854_ net456 net376 _0744_ VPWR VGND sg13g2_nor2_1
X_2785_ _0657_ VPWR _0679_ VGND _0654_ _0658_ sg13g2_o21ai_1
X_1805_ _1131_ _1128_ _1132_ VPWR VGND sg13g2_xor2_1
Xhold202 _0030_ VPWR VGND net242 sg13g2_dlygate4sd3_1
X_1736_ _1065_ _1059_ _1063_ VPWR VGND sg13g2_xnor2_1
Xhold213 DP_1.matrix\[8\] VPWR VGND net253 sg13g2_dlygate4sd3_1
Xhold224 _0028_ VPWR VGND net264 sg13g2_dlygate4sd3_1
Xhold235 DP_2.matrix\[76\] VPWR VGND net275 sg13g2_dlygate4sd3_1
Xhold257 _1242_ VPWR VGND net297 sg13g2_dlygate4sd3_1
X_1667_ _0992_ _0996_ _0997_ VPWR VGND sg13g2_nor2_1
Xhold246 DP_1.matrix\[77\] VPWR VGND net286 sg13g2_dlygate4sd3_1
X_1598_ net419 net414 net464 net463 _0930_ VPWR VGND sg13g2_and4_1
X_3268_ net516 VGND VPWR net10 DP_2.Q_range.out_data\[3\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_39_651 VPWR VGND sg13g2_fill_1
XFILLER_22_1022 VPWR VGND sg13g2_decap_8
XFILLER_45_109 VPWR VGND sg13g2_decap_8
X_3199_ net512 VGND VPWR net125 mac1.sum_lvl1_ff\[78\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2219_ _1500_ net442 net390 VPWR VGND sg13g2_nand2_1
XFILLER_38_150 VPWR VGND sg13g2_decap_8
XFILLER_38_194 VPWR VGND sg13g2_decap_8
XFILLER_14_66 VPWR VGND sg13g2_decap_8
XFILLER_10_768 VPWR VGND sg13g2_decap_8
XFILLER_6_706 VPWR VGND sg13g2_decap_8
XFILLER_30_32 VPWR VGND sg13g2_decap_8
XFILLER_2_923 VPWR VGND sg13g2_decap_8
XFILLER_29_150 VPWR VGND sg13g2_fill_2
XFILLER_29_172 VPWR VGND sg13g2_decap_8
XFILLER_17_334 VPWR VGND sg13g2_fill_2
XFILLER_45_665 VPWR VGND sg13g2_decap_8
XFILLER_17_367 VPWR VGND sg13g2_decap_8
XFILLER_44_186 VPWR VGND sg13g2_decap_8
XFILLER_32_315 VPWR VGND sg13g2_decap_4
XFILLER_41_871 VPWR VGND sg13g2_decap_8
XFILLER_9_533 VPWR VGND sg13g2_decap_8
XFILLER_13_595 VPWR VGND sg13g2_fill_1
XFILLER_9_599 VPWR VGND sg13g2_decap_8
X_2570_ _0466_ _0467_ _0469_ _0470_ VPWR VGND sg13g2_or3_1
XFILLER_5_783 VPWR VGND sg13g2_decap_8
XFILLER_4_260 VPWR VGND sg13g2_fill_1
X_1521_ net417 net470 net412 net468 _0856_ VPWR VGND sg13g2_and4_1
X_3122_ net541 VGND VPWR net152 mac1.sum_lvl1_ff\[9\] clknet_leaf_23_clk sg13g2_dfrbpq_1
XFILLER_49_993 VPWR VGND sg13g2_decap_8
X_3053_ net517 VGND VPWR _0106_ DP_1.matrix\[76\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_2004_ _1301_ net263 _0028_ VPWR VGND sg13g2_nor2b_1
XFILLER_24_816 VPWR VGND sg13g2_decap_8
XFILLER_32_871 VPWR VGND sg13g2_decap_8
X_2906_ net377 net416 _0795_ VPWR VGND net378 sg13g2_nand3b_1
X_2837_ _0043_ _0727_ _0844_ _0042_ _0845_ VPWR VGND sg13g2_a22oi_1
X_2768_ _0661_ _0652_ _0663_ VPWR VGND sg13g2_xor2_1
X_2699_ net479 net476 net430 net428 _0596_ VPWR VGND sg13g2_and4_1
X_1719_ _1048_ _1043_ _1046_ VPWR VGND sg13g2_xnor2_1
Xfanout501 DP_1.matrix\[8\] net501 VPWR VGND sg13g2_buf_1
Xfanout512 net513 net512 VPWR VGND sg13g2_buf_8
Xfanout523 net524 net523 VPWR VGND sg13g2_buf_8
Xfanout545 net546 net545 VPWR VGND sg13g2_buf_8
Xfanout534 net535 net534 VPWR VGND sg13g2_buf_8
XFILLER_27_610 VPWR VGND sg13g2_decap_4
XFILLER_26_131 VPWR VGND sg13g2_fill_1
XFILLER_27_687 VPWR VGND sg13g2_fill_1
XFILLER_42_624 VPWR VGND sg13g2_fill_1
XFILLER_25_43 VPWR VGND sg13g2_decap_4
XFILLER_26_197 VPWR VGND sg13g2_decap_8
XFILLER_10_587 VPWR VGND sg13g2_fill_1
XFILLER_10_576 VPWR VGND sg13g2_decap_8
XFILLER_2_720 VPWR VGND sg13g2_decap_8
XFILLER_2_25 VPWR VGND sg13g2_decap_8
XFILLER_2_797 VPWR VGND sg13g2_decap_8
XFILLER_49_256 VPWR VGND sg13g2_decap_8
XFILLER_2_36 VPWR VGND sg13g2_fill_2
XFILLER_2_47 VPWR VGND sg13g2_decap_8
XFILLER_46_974 VPWR VGND sg13g2_decap_8
XFILLER_45_451 VPWR VGND sg13g2_fill_1
XFILLER_13_370 VPWR VGND sg13g2_decap_8
XFILLER_32_189 VPWR VGND sg13g2_decap_8
XFILLER_9_341 VPWR VGND sg13g2_decap_8
XFILLER_12_1010 VPWR VGND sg13g2_decap_8
X_2622_ _0509_ VPWR _0521_ VGND _0517_ _0519_ sg13g2_o21ai_1
X_2553_ net491 net425 net493 _0453_ VPWR VGND net421 sg13g2_nand4_1
X_1504_ VPWR DP_2.Q_range.data_plus_4\[6\] net12 VGND sg13g2_inv_1
X_2484_ _0377_ VPWR _0386_ VGND _0369_ _0378_ sg13g2_o21ai_1
X_3105_ net512 VGND VPWR _0056_ mac1.products_ff\[144\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_28_407 VPWR VGND sg13g2_decap_4
XFILLER_49_790 VPWR VGND sg13g2_decap_8
X_3036_ net531 VGND VPWR _0089_ DP_1.matrix\[3\] clknet_leaf_14_clk sg13g2_dfrbpq_2
XFILLER_37_952 VPWR VGND sg13g2_decap_8
XFILLER_11_329 VPWR VGND sg13g2_fill_1
XFILLER_11_56 VPWR VGND sg13g2_fill_1
XFILLER_11_45 VPWR VGND sg13g2_decap_8
XFILLER_3_528 VPWR VGND sg13g2_decap_8
Xfanout375 _0815_ net375 VPWR VGND sg13g2_buf_8
XFILLER_4_1008 VPWR VGND sg13g2_decap_8
Xfanout397 net398 net397 VPWR VGND sg13g2_buf_2
Xfanout386 net387 net386 VPWR VGND sg13g2_buf_8
XFILLER_28_930 VPWR VGND sg13g2_decap_8
XFILLER_43_922 VPWR VGND sg13g2_decap_8
XFILLER_14_101 VPWR VGND sg13g2_decap_4
XFILLER_14_112 VPWR VGND sg13g2_decap_8
XFILLER_15_635 VPWR VGND sg13g2_fill_1
XFILLER_36_97 VPWR VGND sg13g2_decap_8
XFILLER_30_605 VPWR VGND sg13g2_fill_1
XFILLER_43_999 VPWR VGND sg13g2_decap_8
XFILLER_7_812 VPWR VGND sg13g2_decap_8
XFILLER_11_863 VPWR VGND sg13g2_decap_8
XFILLER_6_333 VPWR VGND sg13g2_decap_8
XFILLER_7_889 VPWR VGND sg13g2_decap_8
XFILLER_42_8 VPWR VGND sg13g2_fill_1
XFILLER_42_1014 VPWR VGND sg13g2_decap_8
XFILLER_2_594 VPWR VGND sg13g2_decap_8
XFILLER_38_705 VPWR VGND sg13g2_decap_8
XFILLER_18_462 VPWR VGND sg13g2_decap_8
XFILLER_19_985 VPWR VGND sg13g2_decap_8
XFILLER_45_281 VPWR VGND sg13g2_decap_8
XFILLER_33_421 VPWR VGND sg13g2_decap_4
XFILLER_34_933 VPWR VGND sg13g2_decap_8
XFILLER_33_443 VPWR VGND sg13g2_decap_8
X_1984_ mac1.sum_lvl3_ff\[2\] net174 _1287_ VPWR VGND sg13g2_and2_1
XFILLER_20_126 VPWR VGND sg13g2_decap_8
X_2605_ _0504_ net487 net426 VPWR VGND sg13g2_nand2_1
X_2536_ _0435_ _0436_ _0426_ _0437_ VPWR VGND sg13g2_nand3_1
X_2467_ _0356_ VPWR _0370_ VGND _0354_ _0357_ sg13g2_o21ai_1
X_2398_ _0307_ _0306_ _0281_ VPWR VGND sg13g2_nand2b_1
XFILLER_28_237 VPWR VGND sg13g2_decap_8
X_3019_ net547 VGND VPWR _0062_ mac1.products_ff\[13\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_37_782 VPWR VGND sg13g2_fill_1
XFILLER_19_1027 VPWR VGND sg13g2_fill_2
XFILLER_25_955 VPWR VGND sg13g2_decap_8
XFILLER_40_925 VPWR VGND sg13g2_decap_8
XFILLER_24_465 VPWR VGND sg13g2_fill_1
XFILLER_4_826 VPWR VGND sg13g2_decap_8
XFILLER_3_369 VPWR VGND sg13g2_decap_8
XFILLER_19_204 VPWR VGND sg13g2_decap_8
XFILLER_47_535 VPWR VGND sg13g2_fill_2
XFILLER_47_568 VPWR VGND sg13g2_decap_8
XFILLER_47_96 VPWR VGND sg13g2_decap_8
XFILLER_16_911 VPWR VGND sg13g2_decap_8
XFILLER_15_421 VPWR VGND sg13g2_fill_2
XFILLER_15_443 VPWR VGND sg13g2_fill_2
XFILLER_42_251 VPWR VGND sg13g2_fill_1
XFILLER_16_988 VPWR VGND sg13g2_decap_8
XFILLER_31_936 VPWR VGND sg13g2_decap_8
XFILLER_30_424 VPWR VGND sg13g2_fill_2
XFILLER_11_660 VPWR VGND sg13g2_fill_1
XFILLER_7_686 VPWR VGND sg13g2_decap_8
XFILLER_3_892 VPWR VGND sg13g2_decap_8
X_2321_ VGND VPWR _0232_ _0233_ _0198_ _0158_ sg13g2_a21oi_2
X_2252_ _0165_ net456 net502 VPWR VGND sg13g2_nand2_1
XFILLER_33_4 VPWR VGND sg13g2_decap_8
X_2183_ VGND VPWR _1461_ _1462_ _1465_ _1456_ sg13g2_a21oi_1
XFILLER_19_782 VPWR VGND sg13g2_decap_8
XFILLER_22_903 VPWR VGND sg13g2_decap_8
XFILLER_34_741 VPWR VGND sg13g2_decap_8
XFILLER_33_251 VPWR VGND sg13g2_decap_4
X_1967_ _1271_ _1273_ net279 _1275_ VPWR VGND sg13g2_nand3_1
X_1898_ _1220_ _1205_ _1221_ VPWR VGND sg13g2_xor2_1
XFILLER_1_807 VPWR VGND sg13g2_decap_8
XFILLER_0_328 VPWR VGND sg13g2_decap_8
X_2519_ _0402_ _0392_ _0400_ _0420_ VPWR VGND sg13g2_a21o_1
XFILLER_17_11 VPWR VGND sg13g2_fill_1
XFILLER_25_752 VPWR VGND sg13g2_decap_8
XFILLER_40_700 VPWR VGND sg13g2_decap_8
XFILLER_13_925 VPWR VGND sg13g2_decap_8
XFILLER_25_763 VPWR VGND sg13g2_fill_2
XFILLER_25_785 VPWR VGND sg13g2_fill_1
XFILLER_9_907 VPWR VGND sg13g2_decap_8
XFILLER_33_54 VPWR VGND sg13g2_decap_4
XFILLER_33_76 VPWR VGND sg13g2_fill_1
XFILLER_21_980 VPWR VGND sg13g2_decap_8
XFILLER_4_623 VPWR VGND sg13g2_decap_8
XFILLER_48_800 VPWR VGND sg13g2_decap_8
XFILLER_0_895 VPWR VGND sg13g2_decap_8
Xhold6 mac1.products_ff\[144\] VPWR VGND net46 sg13g2_dlygate4sd3_1
XFILLER_48_877 VPWR VGND sg13g2_decap_8
XFILLER_47_365 VPWR VGND sg13g2_decap_8
XFILLER_43_582 VPWR VGND sg13g2_fill_1
XFILLER_15_273 VPWR VGND sg13g2_fill_1
XFILLER_16_796 VPWR VGND sg13g2_decap_4
X_2870_ net376 VPWR _0760_ VGND DP_1.matrix\[6\] _0731_ sg13g2_o21ai_1
X_1821_ _1147_ net405 net498 VPWR VGND sg13g2_nand2_2
XFILLER_31_755 VPWR VGND sg13g2_decap_8
XFILLER_31_788 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_10_clk clknet_3_2__leaf_clk clknet_leaf_10_clk VPWR VGND sg13g2_buf_8
XFILLER_8_984 VPWR VGND sg13g2_decap_8
X_1752_ _1047_ VPWR _1080_ VGND _0993_ _1045_ sg13g2_o21ai_1
X_1683_ _1013_ net498 net420 net459 net414 VPWR VGND sg13g2_a22oi_1
X_2304_ net443 net441 net389 net387 _0216_ VPWR VGND sg13g2_and4_1
X_2235_ _0149_ _1480_ _0147_ _0148_ VPWR VGND sg13g2_and3_1
X_2166_ _1430_ _1420_ _1428_ _1448_ VPWR VGND sg13g2_a21o_1
XFILLER_0_1000 VPWR VGND sg13g2_decap_8
X_2097_ _1380_ _1360_ _0036_ VPWR VGND sg13g2_xor2_1
XFILLER_19_590 VPWR VGND sg13g2_decap_8
XFILLER_26_549 VPWR VGND sg13g2_fill_2
XFILLER_0_91 VPWR VGND sg13g2_decap_8
X_2999_ net394 _0127_ VPWR VGND sg13g2_buf_1
XFILLER_1_604 VPWR VGND sg13g2_decap_8
XFILLER_49_619 VPWR VGND sg13g2_decap_8
XFILLER_0_169 VPWR VGND sg13g2_decap_8
XFILLER_29_343 VPWR VGND sg13g2_decap_8
XFILLER_28_87 VPWR VGND sg13g2_decap_8
XFILLER_45_858 VPWR VGND sg13g2_decap_8
XFILLER_44_368 VPWR VGND sg13g2_decap_4
XFILLER_25_593 VPWR VGND sg13g2_fill_1
XFILLER_40_563 VPWR VGND sg13g2_fill_2
XFILLER_9_704 VPWR VGND sg13g2_decap_8
XFILLER_40_596 VPWR VGND sg13g2_decap_4
XFILLER_5_965 VPWR VGND sg13g2_decap_8
XFILLER_4_442 VPWR VGND sg13g2_decap_4
XFILLER_0_692 VPWR VGND sg13g2_decap_8
X_2020_ _1315_ _1312_ _1314_ VPWR VGND sg13g2_nand2_1
XFILLER_47_195 VPWR VGND sg13g2_decap_8
XFILLER_44_880 VPWR VGND sg13g2_decap_8
X_2922_ _0811_ _0784_ _0810_ _0783_ net502 VPWR VGND sg13g2_a22oi_1
XFILLER_16_582 VPWR VGND sg13g2_fill_1
XFILLER_43_390 VPWR VGND sg13g2_decap_8
X_2853_ VGND VPWR net472 net376 _0743_ net379 sg13g2_a21oi_1
X_2784_ _0660_ _0653_ _0662_ _0678_ VPWR VGND sg13g2_a21o_1
X_1804_ _1131_ _1083_ _1129_ VPWR VGND sg13g2_xnor2_1
XFILLER_8_781 VPWR VGND sg13g2_decap_8
X_1735_ _1064_ _1059_ _1063_ VPWR VGND sg13g2_nand2_1
Xhold225 mac1.sum_lvl2_ff\[4\] VPWR VGND net265 sg13g2_dlygate4sd3_1
Xhold214 mac1.sum_lvl2_ff\[2\] VPWR VGND net254 sg13g2_dlygate4sd3_1
Xhold203 mac1.sum_lvl2_ff\[3\] VPWR VGND net243 sg13g2_dlygate4sd3_1
Xhold247 mac1.sum_lvl3_ff\[7\] VPWR VGND net287 sg13g2_dlygate4sd3_1
Xhold258 _1245_ VPWR VGND net298 sg13g2_dlygate4sd3_1
X_1666_ VGND VPWR _0996_ _0995_ _0994_ sg13g2_or2_1
Xhold236 DP_1.matrix\[37\] VPWR VGND net276 sg13g2_dlygate4sd3_1
X_1597_ _0929_ net411 net466 VPWR VGND sg13g2_nand2_1
X_3267_ net516 VGND VPWR net9 DP_2.Q_range.out_data\[2\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_22_1001 VPWR VGND sg13g2_decap_8
XFILLER_39_674 VPWR VGND sg13g2_decap_8
X_3198_ net512 VGND VPWR net108 mac1.sum_lvl1_ff\[77\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2218_ _1459_ VPWR _1499_ VGND _1457_ _1460_ sg13g2_o21ai_1
XFILLER_27_836 VPWR VGND sg13g2_fill_2
X_2149_ _1430_ _1429_ _1420_ _1432_ VPWR VGND sg13g2_a21o_1
XFILLER_27_869 VPWR VGND sg13g2_decap_8
XFILLER_41_305 VPWR VGND sg13g2_fill_1
XFILLER_35_880 VPWR VGND sg13g2_decap_8
XFILLER_14_56 VPWR VGND sg13g2_decap_4
XFILLER_10_747 VPWR VGND sg13g2_decap_8
XFILLER_30_11 VPWR VGND sg13g2_decap_8
XFILLER_2_902 VPWR VGND sg13g2_decap_8
XFILLER_2_979 VPWR VGND sg13g2_decap_8
XFILLER_39_97 VPWR VGND sg13g2_decap_4
XFILLER_45_611 VPWR VGND sg13g2_decap_8
XFILLER_44_165 VPWR VGND sg13g2_decap_8
XFILLER_40_360 VPWR VGND sg13g2_decap_8
XFILLER_13_574 VPWR VGND sg13g2_decap_8
XFILLER_40_393 VPWR VGND sg13g2_fill_1
XFILLER_5_762 VPWR VGND sg13g2_decap_8
X_1520_ _0855_ net472 net410 VPWR VGND sg13g2_nand2_1
XFILLER_45_1012 VPWR VGND sg13g2_decap_8
X_3121_ net542 VGND VPWR net96 mac1.sum_lvl1_ff\[8\] clknet_leaf_24_clk sg13g2_dfrbpq_1
XFILLER_49_972 VPWR VGND sg13g2_decap_8
X_3052_ net517 VGND VPWR _0105_ DP_1.matrix\[75\] clknet_leaf_8_clk sg13g2_dfrbpq_2
XFILLER_36_611 VPWR VGND sg13g2_decap_8
XFILLER_48_493 VPWR VGND sg13g2_fill_1
XFILLER_48_482 VPWR VGND sg13g2_fill_2
X_2003_ net262 VPWR _1302_ VGND _1296_ _1300_ sg13g2_o21ai_1
XFILLER_35_143 VPWR VGND sg13g2_fill_1
XFILLER_23_338 VPWR VGND sg13g2_fill_1
XFILLER_35_187 VPWR VGND sg13g2_decap_8
XFILLER_36_699 VPWR VGND sg13g2_decap_8
X_2905_ net378 VPWR _0794_ VGND net433 _0782_ sg13g2_o21ai_1
X_2836_ _0727_ net474 net412 VPWR VGND sg13g2_nand2_1
XFILLER_31_393 VPWR VGND sg13g2_decap_8
X_2767_ _0661_ _0652_ _0662_ VPWR VGND sg13g2_nor2b_1
X_2698_ _0595_ net476 net428 VPWR VGND sg13g2_nand2_2
X_1718_ _1047_ _1046_ _1043_ VPWR VGND sg13g2_nand2b_1
X_1649_ _0955_ VPWR _0980_ VGND _0976_ _0978_ sg13g2_o21ai_1
Xfanout502 DP_2.matrix\[80\] net502 VPWR VGND sg13g2_buf_8
Xfanout513 net533 net513 VPWR VGND sg13g2_buf_8
Xfanout524 net533 net524 VPWR VGND sg13g2_buf_8
Xfanout546 net547 net546 VPWR VGND sg13g2_buf_8
Xfanout535 net537 net535 VPWR VGND sg13g2_buf_8
XFILLER_42_603 VPWR VGND sg13g2_decap_8
XFILLER_26_143 VPWR VGND sg13g2_fill_2
XFILLER_27_655 VPWR VGND sg13g2_fill_1
XFILLER_14_327 VPWR VGND sg13g2_decap_8
XFILLER_25_88 VPWR VGND sg13g2_fill_2
XFILLER_41_32 VPWR VGND sg13g2_decap_8
XFILLER_41_54 VPWR VGND sg13g2_fill_2
XFILLER_10_555 VPWR VGND sg13g2_decap_8
XFILLER_41_98 VPWR VGND sg13g2_decap_8
XFILLER_6_537 VPWR VGND sg13g2_decap_8
XFILLER_29_1018 VPWR VGND sg13g2_decap_8
XFILLER_2_776 VPWR VGND sg13g2_decap_8
XFILLER_49_235 VPWR VGND sg13g2_decap_8
XFILLER_46_953 VPWR VGND sg13g2_decap_8
XFILLER_45_430 VPWR VGND sg13g2_decap_8
XFILLER_17_154 VPWR VGND sg13g2_decap_8
XFILLER_17_198 VPWR VGND sg13g2_decap_8
XFILLER_33_647 VPWR VGND sg13g2_decap_4
XFILLER_9_320 VPWR VGND sg13g2_decap_8
XFILLER_9_375 VPWR VGND sg13g2_fill_2
X_2621_ _0509_ _0517_ _0519_ _0520_ VPWR VGND sg13g2_or3_1
X_2552_ _0452_ net421 net493 net425 net491 VPWR VGND sg13g2_a22oi_1
X_1503_ VPWR DP_2.I_range.data_plus_4\[6\] net16 VGND sg13g2_inv_1
XFILLER_5_592 VPWR VGND sg13g2_decap_4
X_2483_ _0384_ _0364_ _0041_ VPWR VGND sg13g2_xor2_1
X_3104_ net512 VGND VPWR _0055_ mac1.products_ff\[143\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3035_ net531 VGND VPWR net251 DP_1.matrix\[2\] clknet_leaf_14_clk sg13g2_dfrbpq_2
XFILLER_37_931 VPWR VGND sg13g2_decap_8
XFILLER_36_441 VPWR VGND sg13g2_fill_2
XFILLER_23_113 VPWR VGND sg13g2_fill_1
XFILLER_24_614 VPWR VGND sg13g2_decap_8
XFILLER_24_636 VPWR VGND sg13g2_decap_8
XFILLER_36_496 VPWR VGND sg13g2_fill_1
XFILLER_23_179 VPWR VGND sg13g2_fill_1
X_2819_ _0712_ _0705_ _0711_ VPWR VGND sg13g2_nand2_1
XFILLER_11_13 VPWR VGND sg13g2_fill_1
XFILLER_20_897 VPWR VGND sg13g2_decap_8
XFILLER_11_79 VPWR VGND sg13g2_decap_8
Xfanout398 net400 net398 VPWR VGND sg13g2_buf_1
Xfanout387 net275 net387 VPWR VGND sg13g2_buf_8
Xfanout376 _0735_ net376 VPWR VGND sg13g2_buf_8
XFILLER_46_216 VPWR VGND sg13g2_decap_4
XFILLER_43_901 VPWR VGND sg13g2_decap_8
XFILLER_28_986 VPWR VGND sg13g2_decap_8
XFILLER_36_43 VPWR VGND sg13g2_decap_8
XFILLER_15_614 VPWR VGND sg13g2_decap_4
XFILLER_27_474 VPWR VGND sg13g2_decap_8
XFILLER_36_76 VPWR VGND sg13g2_decap_8
XFILLER_43_978 VPWR VGND sg13g2_decap_8
XFILLER_15_669 VPWR VGND sg13g2_fill_1
XFILLER_42_488 VPWR VGND sg13g2_decap_8
XFILLER_14_157 VPWR VGND sg13g2_decap_4
XFILLER_42_499 VPWR VGND sg13g2_fill_1
XFILLER_11_842 VPWR VGND sg13g2_decap_8
XFILLER_7_868 VPWR VGND sg13g2_decap_8
XFILLER_2_551 VPWR VGND sg13g2_fill_2
XFILLER_37_216 VPWR VGND sg13g2_fill_1
XFILLER_19_964 VPWR VGND sg13g2_decap_8
XFILLER_45_260 VPWR VGND sg13g2_decap_8
XFILLER_34_912 VPWR VGND sg13g2_decap_8
XFILLER_20_105 VPWR VGND sg13g2_decap_8
XFILLER_34_989 VPWR VGND sg13g2_decap_8
X_1983_ _1283_ VPWR _1286_ VGND _1282_ _1284_ sg13g2_o21ai_1
XFILLER_14_680 VPWR VGND sg13g2_fill_1
XFILLER_21_639 VPWR VGND sg13g2_fill_1
XFILLER_20_149 VPWR VGND sg13g2_decap_8
X_2604_ _0473_ VPWR _0503_ VGND _0464_ _0474_ sg13g2_o21ai_1
X_2535_ _0433_ _0432_ _0427_ _0436_ VPWR VGND sg13g2_a21o_1
X_2466_ _0369_ _0368_ _0365_ VPWR VGND sg13g2_nand2b_1
X_2397_ _0304_ _0266_ _0306_ VPWR VGND sg13g2_xor2_1
XFILLER_44_709 VPWR VGND sg13g2_decap_8
X_3018_ net546 VGND VPWR _0061_ mac1.products_ff\[12\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_25_934 VPWR VGND sg13g2_decap_8
XFILLER_37_794 VPWR VGND sg13g2_fill_1
XFILLER_40_904 VPWR VGND sg13g2_decap_8
XFILLER_19_1006 VPWR VGND sg13g2_decap_8
XFILLER_24_444 VPWR VGND sg13g2_decap_8
XFILLER_11_127 VPWR VGND sg13g2_decap_4
XFILLER_20_683 VPWR VGND sg13g2_decap_8
XFILLER_4_805 VPWR VGND sg13g2_decap_8
XFILLER_3_337 VPWR VGND sg13g2_decap_8
XFILLER_47_514 VPWR VGND sg13g2_decap_8
XFILLER_47_53 VPWR VGND sg13g2_fill_2
XFILLER_47_42 VPWR VGND sg13g2_decap_8
XFILLER_47_75 VPWR VGND sg13g2_decap_8
XFILLER_19_249 VPWR VGND sg13g2_decap_8
XFILLER_35_709 VPWR VGND sg13g2_fill_2
XFILLER_34_208 VPWR VGND sg13g2_decap_8
XFILLER_16_967 VPWR VGND sg13g2_decap_8
XFILLER_43_786 VPWR VGND sg13g2_decap_8
XFILLER_31_915 VPWR VGND sg13g2_decap_8
XFILLER_42_274 VPWR VGND sg13g2_decap_4
XFILLER_30_436 VPWR VGND sg13g2_fill_1
XFILLER_30_458 VPWR VGND sg13g2_decap_8
XFILLER_30_469 VPWR VGND sg13g2_fill_2
XFILLER_7_665 VPWR VGND sg13g2_decap_8
XFILLER_3_871 VPWR VGND sg13g2_decap_8
X_2320_ VGND VPWR _0155_ _0197_ _0232_ _0196_ sg13g2_a21oi_1
X_2251_ _1496_ VPWR _0164_ VGND _1493_ _1497_ sg13g2_o21ai_1
XFILLER_26_4 VPWR VGND sg13g2_decap_8
X_2182_ _1461_ _1462_ _1456_ _1464_ VPWR VGND sg13g2_nand3_1
XFILLER_38_536 VPWR VGND sg13g2_decap_8
XFILLER_26_709 VPWR VGND sg13g2_decap_8
XFILLER_38_558 VPWR VGND sg13g2_fill_2
XFILLER_19_761 VPWR VGND sg13g2_fill_2
XFILLER_21_414 VPWR VGND sg13g2_decap_8
XFILLER_22_959 VPWR VGND sg13g2_decap_8
X_1966_ VGND VPWR net279 _1271_ _1274_ _1273_ sg13g2_a21oi_1
X_1897_ _1220_ net460 net494 VPWR VGND sg13g2_nand2_1
X_2518_ _0416_ _0415_ _0419_ VPWR VGND sg13g2_xor2_1
X_2449_ VGND VPWR _0353_ _0348_ _0346_ sg13g2_or2_1
XFILLER_25_731 VPWR VGND sg13g2_decap_8
XFILLER_13_904 VPWR VGND sg13g2_decap_8
XFILLER_24_241 VPWR VGND sg13g2_fill_2
XFILLER_33_11 VPWR VGND sg13g2_decap_8
XFILLER_40_756 VPWR VGND sg13g2_decap_8
XFILLER_12_458 VPWR VGND sg13g2_decap_8
XFILLER_12_469 VPWR VGND sg13g2_fill_2
XFILLER_32_1025 VPWR VGND sg13g2_decap_4
XFILLER_3_134 VPWR VGND sg13g2_fill_1
XFILLER_4_679 VPWR VGND sg13g2_decap_8
XFILLER_0_874 VPWR VGND sg13g2_decap_8
Xhold7 mac1.products_ff\[81\] VPWR VGND net47 sg13g2_dlygate4sd3_1
XFILLER_48_856 VPWR VGND sg13g2_decap_8
XFILLER_35_517 VPWR VGND sg13g2_decap_4
XFILLER_43_550 VPWR VGND sg13g2_fill_1
XFILLER_15_252 VPWR VGND sg13g2_decap_8
XFILLER_31_723 VPWR VGND sg13g2_decap_8
X_1820_ _1146_ net499 net406 net460 net405 VPWR VGND sg13g2_a22oi_1
XFILLER_31_767 VPWR VGND sg13g2_decap_8
XFILLER_30_266 VPWR VGND sg13g2_decap_4
XFILLER_8_963 VPWR VGND sg13g2_decap_8
X_1751_ _1067_ VPWR _1079_ VGND _1051_ _1068_ sg13g2_o21ai_1
XFILLER_30_299 VPWR VGND sg13g2_decap_8
X_1682_ net415 net459 net420 _1012_ VPWR VGND net498 sg13g2_nand4_1
XFILLER_48_1010 VPWR VGND sg13g2_decap_8
X_2303_ _0215_ net441 net387 VPWR VGND sg13g2_nand2_1
X_2234_ _1491_ VPWR _0148_ VGND _0144_ _0146_ sg13g2_o21ai_1
XFILLER_17_0 VPWR VGND sg13g2_decap_8
X_2165_ _1447_ _1442_ _1445_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_333 VPWR VGND sg13g2_decap_8
XFILLER_38_366 VPWR VGND sg13g2_fill_1
XFILLER_38_377 VPWR VGND sg13g2_decap_8
X_2096_ VGND VPWR _1381_ _1380_ _1360_ sg13g2_or2_1
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_22_745 VPWR VGND sg13g2_decap_8
XFILLER_16_1009 VPWR VGND sg13g2_decap_8
XFILLER_22_756 VPWR VGND sg13g2_fill_1
XFILLER_22_778 VPWR VGND sg13g2_decap_4
XFILLER_10_929 VPWR VGND sg13g2_decap_8
X_2998_ net399 _0126_ VPWR VGND sg13g2_buf_1
X_1949_ mac1.sum_lvl2_ff\[10\] net301 _1260_ VPWR VGND sg13g2_xor2_1
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_0_148 VPWR VGND sg13g2_decap_8
XFILLER_45_837 VPWR VGND sg13g2_decap_8
XFILLER_29_377 VPWR VGND sg13g2_decap_8
XFILLER_44_336 VPWR VGND sg13g2_decap_8
XFILLER_44_54 VPWR VGND sg13g2_decap_8
XFILLER_40_553 VPWR VGND sg13g2_fill_1
XFILLER_12_255 VPWR VGND sg13g2_decap_8
XFILLER_5_944 VPWR VGND sg13g2_decap_8
XFILLER_48_620 VPWR VGND sg13g2_decap_8
XFILLER_0_671 VPWR VGND sg13g2_decap_8
XFILLER_48_675 VPWR VGND sg13g2_fill_2
XFILLER_47_174 VPWR VGND sg13g2_decap_8
XFILLER_39_1009 VPWR VGND sg13g2_decap_8
X_2921_ DP_2.matrix\[44\] net495 _0781_ _0810_ VPWR VGND sg13g2_mux2_1
X_2852_ _0742_ net376 _0741_ _0732_ net458 VPWR VGND sg13g2_a22oi_1
X_2783_ _0677_ _0673_ _0061_ VPWR VGND sg13g2_xor2_1
X_1803_ VGND VPWR _1130_ _1129_ _1083_ sg13g2_or2_1
XFILLER_31_597 VPWR VGND sg13g2_fill_2
XFILLER_8_760 VPWR VGND sg13g2_decap_8
X_1734_ _1061_ _1062_ _1063_ VPWR VGND sg13g2_nor2_1
Xhold226 _1237_ VPWR VGND net266 sg13g2_dlygate4sd3_1
Xhold204 _1234_ VPWR VGND net244 sg13g2_dlygate4sd3_1
Xhold215 _1231_ VPWR VGND net255 sg13g2_dlygate4sd3_1
Xhold248 _1305_ VPWR VGND net288 sg13g2_dlygate4sd3_1
Xhold259 _0012_ VPWR VGND net299 sg13g2_dlygate4sd3_1
X_1665_ _0995_ net401 net473 net404 net471 VPWR VGND sg13g2_a22oi_1
Xhold237 DP_1.matrix\[72\] VPWR VGND net277 sg13g2_dlygate4sd3_1
X_1596_ _0898_ VPWR _0928_ VGND _0896_ _0899_ sg13g2_o21ai_1
X_3266_ net516 VGND VPWR net16 DP_2.I_range.out_data\[6\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_39_642 VPWR VGND sg13g2_decap_8
X_2217_ _1498_ _1493_ _1497_ VPWR VGND sg13g2_xnor2_1
X_3197_ net506 VGND VPWR net119 mac1.sum_lvl1_ff\[76\] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_2148_ _1429_ _1430_ _1420_ _1431_ VPWR VGND sg13g2_nand3_1
XFILLER_27_848 VPWR VGND sg13g2_decap_8
X_2079_ _1361_ _1363_ _1364_ VPWR VGND sg13g2_nor2_1
XFILLER_41_317 VPWR VGND sg13g2_decap_8
XFILLER_22_520 VPWR VGND sg13g2_decap_8
XFILLER_14_35 VPWR VGND sg13g2_decap_8
XFILLER_22_542 VPWR VGND sg13g2_decap_8
XFILLER_34_380 VPWR VGND sg13g2_fill_2
XFILLER_10_726 VPWR VGND sg13g2_decap_8
XFILLER_10_704 VPWR VGND sg13g2_fill_2
XFILLER_30_67 VPWR VGND sg13g2_fill_2
XFILLER_30_89 VPWR VGND sg13g2_decap_8
XFILLER_2_958 VPWR VGND sg13g2_decap_8
XFILLER_49_428 VPWR VGND sg13g2_decap_8
XFILLER_39_76 VPWR VGND sg13g2_decap_8
XFILLER_18_815 VPWR VGND sg13g2_decap_4
XFILLER_17_325 VPWR VGND sg13g2_fill_1
XFILLER_17_336 VPWR VGND sg13g2_fill_1
XFILLER_18_848 VPWR VGND sg13g2_decap_4
XFILLER_26_881 VPWR VGND sg13g2_decap_8
XFILLER_32_339 VPWR VGND sg13g2_decap_8
XFILLER_13_520 VPWR VGND sg13g2_decap_8
XFILLER_13_553 VPWR VGND sg13g2_decap_8
XFILLER_25_391 VPWR VGND sg13g2_decap_8
XFILLER_9_502 VPWR VGND sg13g2_decap_4
XFILLER_5_741 VPWR VGND sg13g2_decap_8
X_3120_ net536 VGND VPWR net106 mac1.sum_lvl1_ff\[7\] clknet_leaf_25_clk sg13g2_dfrbpq_1
XFILLER_49_951 VPWR VGND sg13g2_decap_8
X_3051_ net517 VGND VPWR _0104_ DP_1.matrix\[74\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_2002_ _1296_ net262 _1300_ _1301_ VPWR VGND sg13g2_nor3_1
X_2904_ net396 net377 _0793_ VPWR VGND sg13g2_nor2_1
X_2835_ _0064_ _0719_ _0726_ VPWR VGND sg13g2_xnor2_1
X_2766_ _0661_ _0653_ _0660_ VPWR VGND sg13g2_xnor2_1
X_2697_ _0594_ net481 net426 VPWR VGND sg13g2_nand2_1
X_1717_ _1045_ _0993_ _1046_ VPWR VGND sg13g2_xor2_1
X_1648_ _0955_ _0976_ _0978_ _0979_ VPWR VGND sg13g2_or3_1
Xfanout514 net515 net514 VPWR VGND sg13g2_buf_8
Xfanout503 net506 net503 VPWR VGND sg13g2_buf_8
Xfanout547 net548 net547 VPWR VGND sg13g2_buf_8
Xfanout525 net528 net525 VPWR VGND sg13g2_buf_8
X_1579_ _0883_ _0911_ _0912_ VPWR VGND sg13g2_nor2_1
Xfanout536 net537 net536 VPWR VGND sg13g2_buf_8
XFILLER_39_461 VPWR VGND sg13g2_fill_2
XFILLER_39_450 VPWR VGND sg13g2_decap_8
X_3249_ net504 VGND VPWR net242 net17 clknet_leaf_31_clk sg13g2_dfrbpq_2
XFILLER_39_483 VPWR VGND sg13g2_decap_8
XFILLER_26_111 VPWR VGND sg13g2_fill_1
XFILLER_27_634 VPWR VGND sg13g2_decap_8
XFILLER_26_166 VPWR VGND sg13g2_decap_8
XFILLER_26_177 VPWR VGND sg13g2_fill_2
XFILLER_23_884 VPWR VGND sg13g2_decap_8
XFILLER_41_11 VPWR VGND sg13g2_decap_8
XFILLER_2_755 VPWR VGND sg13g2_decap_8
XFILLER_49_214 VPWR VGND sg13g2_decap_8
XFILLER_18_601 VPWR VGND sg13g2_fill_1
XFILLER_46_932 VPWR VGND sg13g2_decap_8
XFILLER_18_623 VPWR VGND sg13g2_fill_1
XFILLER_18_645 VPWR VGND sg13g2_decap_4
XFILLER_17_133 VPWR VGND sg13g2_decap_8
XFILLER_17_177 VPWR VGND sg13g2_decap_8
XFILLER_41_670 VPWR VGND sg13g2_decap_8
XFILLER_14_884 VPWR VGND sg13g2_decap_8
XFILLER_32_169 VPWR VGND sg13g2_decap_8
XFILLER_41_692 VPWR VGND sg13g2_decap_8
X_2620_ VGND VPWR _0515_ _0516_ _0519_ _0510_ sg13g2_a21oi_1
X_2551_ _0425_ VPWR _0451_ VGND _0388_ _0423_ sg13g2_o21ai_1
X_1502_ VPWR DP_1.I_range.data_plus_4\[6\] net4 VGND sg13g2_inv_1
X_2482_ _0385_ _0364_ _0384_ VPWR VGND sg13g2_nand2_1
X_3103_ net512 VGND VPWR _0054_ mac1.products_ff\[142\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_37_910 VPWR VGND sg13g2_decap_8
X_3034_ net531 VGND VPWR net248 DP_1.matrix\[1\] clknet_leaf_7_clk sg13g2_dfrbpq_2
XFILLER_37_987 VPWR VGND sg13g2_decap_8
XFILLER_23_158 VPWR VGND sg13g2_fill_2
XFILLER_20_843 VPWR VGND sg13g2_decap_4
XFILLER_32_670 VPWR VGND sg13g2_decap_4
XFILLER_20_876 VPWR VGND sg13g2_decap_8
X_2818_ _0711_ _0706_ _0709_ VPWR VGND sg13g2_xnor2_1
X_2749_ _0645_ _0642_ _0644_ VPWR VGND sg13g2_nand2_1
Xfanout377 _0784_ net377 VPWR VGND sg13g2_buf_8
Xfanout399 net400 net399 VPWR VGND sg13g2_buf_2
Xfanout388 net389 net388 VPWR VGND sg13g2_buf_8
XFILLER_27_453 VPWR VGND sg13g2_decap_8
XFILLER_28_965 VPWR VGND sg13g2_decap_8
XFILLER_36_22 VPWR VGND sg13g2_decap_8
XFILLER_43_957 VPWR VGND sg13g2_decap_8
XFILLER_14_136 VPWR VGND sg13g2_decap_8
XFILLER_15_648 VPWR VGND sg13g2_decap_8
XFILLER_11_821 VPWR VGND sg13g2_decap_8
XFILLER_23_681 VPWR VGND sg13g2_fill_1
XFILLER_6_302 VPWR VGND sg13g2_fill_2
XFILLER_7_847 VPWR VGND sg13g2_decap_8
XFILLER_11_898 VPWR VGND sg13g2_decap_8
XFILLER_10_397 VPWR VGND sg13g2_decap_8
XFILLER_19_943 VPWR VGND sg13g2_decap_8
XFILLER_46_751 VPWR VGND sg13g2_decap_8
XFILLER_18_442 VPWR VGND sg13g2_decap_8
XFILLER_33_401 VPWR VGND sg13g2_decap_8
XFILLER_18_497 VPWR VGND sg13g2_decap_8
XFILLER_34_968 VPWR VGND sg13g2_decap_8
XFILLER_21_618 VPWR VGND sg13g2_decap_8
X_1982_ _0023_ _1282_ _1285_ VPWR VGND sg13g2_xnor2_1
XFILLER_13_180 VPWR VGND sg13g2_decap_8
XFILLER_9_184 VPWR VGND sg13g2_decap_8
X_2603_ _0502_ _0453_ _0501_ VPWR VGND sg13g2_xnor2_1
X_2534_ _0432_ _0433_ _0427_ _0435_ VPWR VGND sg13g2_nand3_1
XFILLER_47_0 VPWR VGND sg13g2_decap_8
X_2465_ VGND VPWR _0368_ _0366_ _0352_ sg13g2_or2_1
X_2396_ _0266_ _0304_ _0305_ VPWR VGND sg13g2_nor2_1
XFILLER_43_209 VPWR VGND sg13g2_decap_8
XFILLER_25_913 VPWR VGND sg13g2_decap_8
XFILLER_37_773 VPWR VGND sg13g2_decap_8
X_3017_ net546 VGND VPWR _0060_ mac1.products_ff\[11\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_11_106 VPWR VGND sg13g2_decap_8
XFILLER_20_673 VPWR VGND sg13g2_fill_2
XFILLER_47_21 VPWR VGND sg13g2_decap_8
XFILLER_15_423 VPWR VGND sg13g2_fill_1
XFILLER_15_445 VPWR VGND sg13g2_fill_1
XFILLER_16_946 VPWR VGND sg13g2_decap_8
XFILLER_15_489 VPWR VGND sg13g2_decap_8
XFILLER_8_26 VPWR VGND sg13g2_fill_2
XFILLER_8_59 VPWR VGND sg13g2_decap_8
XFILLER_10_194 VPWR VGND sg13g2_fill_1
XFILLER_6_176 VPWR VGND sg13g2_fill_2
XFILLER_3_850 VPWR VGND sg13g2_decap_8
X_2250_ _1484_ _1487_ _0163_ VPWR VGND sg13g2_nor2_1
XFILLER_19_4 VPWR VGND sg13g2_decap_8
X_2181_ _1463_ _1456_ _1461_ _1462_ VPWR VGND sg13g2_and3_1
XFILLER_34_710 VPWR VGND sg13g2_decap_8
XFILLER_34_776 VPWR VGND sg13g2_decap_4
XFILLER_22_938 VPWR VGND sg13g2_decap_8
X_1965_ _1273_ mac1.sum_lvl2_ff\[32\] mac1.sum_lvl2_ff\[13\] VPWR VGND sg13g2_xnor2_1
X_1896_ _1208_ VPWR _1219_ VGND _1179_ _1206_ sg13g2_o21ai_1
X_2517_ _0418_ _0415_ _0416_ VPWR VGND sg13g2_xnor2_1
X_2448_ _0352_ net492 net429 VPWR VGND sg13g2_nand2_2
XFILLER_25_1011 VPWR VGND sg13g2_decap_8
X_2379_ _0287_ _0288_ _0289_ VPWR VGND sg13g2_nor2_1
XFILLER_44_507 VPWR VGND sg13g2_decap_8
XFILLER_17_46 VPWR VGND sg13g2_decap_8
XFILLER_25_710 VPWR VGND sg13g2_decap_8
XFILLER_40_735 VPWR VGND sg13g2_decap_8
XFILLER_8_419 VPWR VGND sg13g2_decap_4
XFILLER_32_1004 VPWR VGND sg13g2_decap_8
XFILLER_4_658 VPWR VGND sg13g2_decap_8
XFILLER_0_853 VPWR VGND sg13g2_decap_8
XFILLER_48_835 VPWR VGND sg13g2_decap_8
XFILLER_47_301 VPWR VGND sg13g2_fill_2
Xhold8 mac1.products_ff\[137\] VPWR VGND net48 sg13g2_dlygate4sd3_1
XFILLER_47_323 VPWR VGND sg13g2_decap_8
XFILLER_35_529 VPWR VGND sg13g2_fill_1
XFILLER_15_231 VPWR VGND sg13g2_decap_8
XFILLER_16_754 VPWR VGND sg13g2_decap_8
XFILLER_43_573 VPWR VGND sg13g2_decap_8
XFILLER_30_245 VPWR VGND sg13g2_decap_8
XFILLER_12_982 VPWR VGND sg13g2_decap_8
X_1750_ VGND VPWR _1042_ _1048_ _1078_ _1050_ sg13g2_a21oi_1
XFILLER_8_942 VPWR VGND sg13g2_decap_8
XFILLER_11_492 VPWR VGND sg13g2_decap_4
X_1681_ net420 net414 net459 net498 _1011_ VPWR VGND sg13g2_and4_1
X_2302_ _0214_ net445 net384 VPWR VGND sg13g2_nand2_1
XFILLER_2_190 VPWR VGND sg13g2_decap_8
X_2233_ _1491_ _0144_ _0146_ _0147_ VPWR VGND sg13g2_or3_1
XFILLER_38_312 VPWR VGND sg13g2_decap_8
X_2164_ _1446_ _1442_ _1445_ VPWR VGND sg13g2_nand2_1
X_2095_ _1378_ _1377_ _1380_ VPWR VGND sg13g2_xor2_1
XFILLER_22_724 VPWR VGND sg13g2_fill_2
XFILLER_34_595 VPWR VGND sg13g2_decap_8
XFILLER_10_908 VPWR VGND sg13g2_decap_8
XFILLER_21_234 VPWR VGND sg13g2_decap_8
X_2997_ net402 _0125_ VPWR VGND sg13g2_buf_1
XFILLER_9_91 VPWR VGND sg13g2_decap_8
X_1948_ _1259_ net301 mac1.sum_lvl2_ff\[10\] VPWR VGND sg13g2_nand2_1
XFILLER_21_289 VPWR VGND sg13g2_decap_8
X_1879_ _1182_ VPWR _1203_ VGND _1153_ _1180_ sg13g2_o21ai_1
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_1_639 VPWR VGND sg13g2_decap_8
XFILLER_45_816 VPWR VGND sg13g2_decap_8
XFILLER_17_507 VPWR VGND sg13g2_fill_2
XFILLER_44_315 VPWR VGND sg13g2_decap_8
XFILLER_44_33 VPWR VGND sg13g2_decap_8
XFILLER_44_22 VPWR VGND sg13g2_decap_8
XFILLER_40_521 VPWR VGND sg13g2_decap_4
XFILLER_9_739 VPWR VGND sg13g2_decap_8
XFILLER_8_249 VPWR VGND sg13g2_decap_8
XFILLER_12_289 VPWR VGND sg13g2_fill_1
XFILLER_5_923 VPWR VGND sg13g2_decap_8
XFILLER_5_27 VPWR VGND sg13g2_decap_8
XFILLER_5_38 VPWR VGND sg13g2_fill_1
XFILLER_4_466 VPWR VGND sg13g2_decap_8
XFILLER_0_650 VPWR VGND sg13g2_decap_8
XFILLER_47_131 VPWR VGND sg13g2_decap_8
X_2920_ _0786_ _0805_ _0807_ _0809_ VPWR VGND sg13g2_nor3_1
XFILLER_16_573 VPWR VGND sg13g2_decap_8
XFILLER_31_543 VPWR VGND sg13g2_decap_8
X_2851_ net474 net492 net379 _0741_ VPWR VGND sg13g2_mux2_1
XFILLER_31_576 VPWR VGND sg13g2_fill_1
X_2782_ _0677_ _0676_ _0644_ _0675_ _0612_ VPWR VGND sg13g2_a22oi_1
X_1802_ _1129_ net465 net403 VPWR VGND sg13g2_nand2_1
X_1733_ _1062_ net498 net415 net459 net411 VPWR VGND sg13g2_a22oi_1
Xhold205 _0009_ VPWR VGND net245 sg13g2_dlygate4sd3_1
Xhold216 _0008_ VPWR VGND net256 sg13g2_dlygate4sd3_1
Xhold249 _0029_ VPWR VGND net289 sg13g2_dlygate4sd3_1
Xhold227 _0010_ VPWR VGND net267 sg13g2_dlygate4sd3_1
X_1664_ net471 net473 net403 net401 _0994_ VPWR VGND sg13g2_and4_1
Xhold238 mac1.sum_lvl2_ff\[31\] VPWR VGND net278 sg13g2_dlygate4sd3_1
X_1595_ _0927_ _0922_ _0925_ VPWR VGND sg13g2_xnor2_1
X_3265_ net516 VGND VPWR DP_2.I_range.data_plus_4\[6\] DP_2.I_range.out_data\[5\]
+ clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2216_ _1497_ _1450_ _1495_ VPWR VGND sg13g2_xnor2_1
X_3196_ net505 VGND VPWR net128 mac1.sum_lvl1_ff\[75\] clknet_leaf_37_clk sg13g2_dfrbpq_1
X_2147_ _1427_ _1426_ _1421_ _1430_ VPWR VGND sg13g2_a21o_1
XFILLER_27_838 VPWR VGND sg13g2_fill_1
X_2078_ net457 net454 net388 net386 _1363_ VPWR VGND sg13g2_and4_1
XFILLER_14_14 VPWR VGND sg13g2_fill_1
XFILLER_2_937 VPWR VGND sg13g2_decap_8
XFILLER_7_1008 VPWR VGND sg13g2_decap_8
XFILLER_39_33 VPWR VGND sg13g2_decap_8
XFILLER_49_407 VPWR VGND sg13g2_decap_8
XFILLER_39_55 VPWR VGND sg13g2_decap_8
XFILLER_45_646 VPWR VGND sg13g2_fill_1
XFILLER_25_370 VPWR VGND sg13g2_decap_8
XFILLER_41_885 VPWR VGND sg13g2_decap_8
XFILLER_40_384 VPWR VGND sg13g2_decap_8
XFILLER_9_547 VPWR VGND sg13g2_decap_8
XFILLER_5_720 VPWR VGND sg13g2_decap_8
XFILLER_5_797 VPWR VGND sg13g2_decap_8
XFILLER_4_274 VPWR VGND sg13g2_decap_4
XFILLER_49_930 VPWR VGND sg13g2_decap_8
X_3050_ net517 VGND VPWR _0103_ DP_1.matrix\[73\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2001_ VPWR VGND _1294_ _1293_ _1292_ net178 _1300_ mac1.sum_lvl3_ff\[25\] sg13g2_a221oi_1
XFILLER_48_484 VPWR VGND sg13g2_fill_1
XFILLER_36_657 VPWR VGND sg13g2_decap_4
XFILLER_17_893 VPWR VGND sg13g2_decap_8
XFILLER_32_885 VPWR VGND sg13g2_decap_8
X_2903_ _0792_ net377 _0791_ _0783_ DP_2.matrix\[72\] VPWR VGND sg13g2_a22oi_1
X_2834_ _0726_ _0720_ _0725_ VPWR VGND sg13g2_xnor2_1
X_2765_ _0660_ _0654_ _0659_ VPWR VGND sg13g2_xnor2_1
X_2696_ VGND VPWR net476 net434 _0593_ _0561_ sg13g2_a21oi_1
X_1716_ _1045_ net469 net404 VPWR VGND sg13g2_nand2_1
XFILLER_6_81 VPWR VGND sg13g2_decap_8
X_1647_ VGND VPWR _0974_ _0975_ _0978_ _0956_ sg13g2_a21oi_1
Xfanout504 net506 net504 VPWR VGND sg13g2_buf_8
Xfanout515 net518 net515 VPWR VGND sg13g2_buf_8
Xfanout526 net528 net526 VPWR VGND sg13g2_buf_8
X_1578_ _0910_ _0868_ _0911_ VPWR VGND sg13g2_xor2_1
Xfanout537 net549 net537 VPWR VGND sg13g2_buf_8
Xfanout548 net549 net548 VPWR VGND sg13g2_buf_8
X_3248_ net504 VGND VPWR net289 net32 clknet_leaf_32_clk sg13g2_dfrbpq_2
X_3179_ net506 VGND VPWR net147 mac1.sum_lvl2_ff\[40\] clknet_leaf_36_clk sg13g2_dfrbpq_1
XFILLER_26_145 VPWR VGND sg13g2_fill_1
XFILLER_23_852 VPWR VGND sg13g2_decap_8
XFILLER_23_863 VPWR VGND sg13g2_fill_2
XFILLER_41_56 VPWR VGND sg13g2_fill_1
XFILLER_6_517 VPWR VGND sg13g2_decap_8
XFILLER_41_78 VPWR VGND sg13g2_decap_8
XFILLER_6_528 VPWR VGND sg13g2_fill_1
XFILLER_2_734 VPWR VGND sg13g2_decap_8
XFILLER_46_911 VPWR VGND sg13g2_decap_8
XFILLER_46_988 VPWR VGND sg13g2_decap_8
XFILLER_45_465 VPWR VGND sg13g2_fill_2
XFILLER_14_863 VPWR VGND sg13g2_decap_8
XFILLER_13_384 VPWR VGND sg13g2_fill_1
XFILLER_40_192 VPWR VGND sg13g2_fill_1
XFILLER_9_377 VPWR VGND sg13g2_fill_1
XFILLER_9_355 VPWR VGND sg13g2_decap_8
XFILLER_12_1024 VPWR VGND sg13g2_decap_4
X_2550_ _0439_ VPWR _0450_ VGND _0419_ _0440_ sg13g2_o21ai_1
X_1501_ VPWR _0842_ DP_2.Q_range.out_data\[5\] VGND sg13g2_inv_1
XFILLER_5_572 VPWR VGND sg13g2_fill_2
X_2481_ _0384_ _0381_ _0382_ VPWR VGND sg13g2_xnor2_1
X_3102_ net507 VGND VPWR _0047_ mac1.products_ff\[141\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3033_ net531 VGND VPWR net195 DP_1.matrix\[0\] clknet_leaf_14_clk sg13g2_dfrbpq_2
XFILLER_37_966 VPWR VGND sg13g2_decap_8
XFILLER_36_487 VPWR VGND sg13g2_decap_8
XFILLER_23_137 VPWR VGND sg13g2_decap_8
XFILLER_31_192 VPWR VGND sg13g2_decap_4
X_2817_ _0710_ _0709_ _0706_ VPWR VGND sg13g2_nand2b_1
X_2748_ VPWR _0644_ _0643_ VGND sg13g2_inv_1
X_2679_ _0577_ _0539_ _0574_ VPWR VGND sg13g2_xnor2_1
XFILLER_47_708 VPWR VGND sg13g2_decap_4
Xfanout378 _0781_ net378 VPWR VGND sg13g2_buf_8
Xfanout389 net273 net389 VPWR VGND sg13g2_buf_8
XFILLER_28_944 VPWR VGND sg13g2_decap_8
XFILLER_43_936 VPWR VGND sg13g2_decap_8
XFILLER_14_126 VPWR VGND sg13g2_fill_2
XFILLER_23_660 VPWR VGND sg13g2_decap_8
XFILLER_30_619 VPWR VGND sg13g2_decap_8
XFILLER_35_1013 VPWR VGND sg13g2_decap_8
XFILLER_10_310 VPWR VGND sg13g2_decap_8
XFILLER_22_170 VPWR VGND sg13g2_fill_2
XFILLER_10_354 VPWR VGND sg13g2_decap_8
XFILLER_7_826 VPWR VGND sg13g2_decap_8
XFILLER_11_877 VPWR VGND sg13g2_decap_8
XFILLER_6_358 VPWR VGND sg13g2_decap_8
XFILLER_6_347 VPWR VGND sg13g2_fill_2
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_42_1028 VPWR VGND sg13g2_fill_1
XFILLER_38_719 VPWR VGND sg13g2_fill_2
XFILLER_19_922 VPWR VGND sg13g2_decap_8
XFILLER_46_730 VPWR VGND sg13g2_decap_8
XFILLER_18_421 VPWR VGND sg13g2_decap_8
XFILLER_18_476 VPWR VGND sg13g2_decap_8
XFILLER_19_999 VPWR VGND sg13g2_decap_8
XFILLER_45_295 VPWR VGND sg13g2_fill_2
XFILLER_34_947 VPWR VGND sg13g2_decap_8
XFILLER_33_457 VPWR VGND sg13g2_fill_2
XFILLER_33_468 VPWR VGND sg13g2_fill_2
X_1981_ mac1.sum_lvl3_ff\[21\] mac1.sum_lvl3_ff\[1\] _1285_ VPWR VGND sg13g2_xor2_1
XFILLER_14_671 VPWR VGND sg13g2_decap_8
X_2602_ _0501_ _0492_ _0499_ VPWR VGND sg13g2_xnor2_1
XFILLER_6_881 VPWR VGND sg13g2_decap_8
X_2533_ _0434_ _0427_ _0432_ _0433_ VPWR VGND sg13g2_and3_1
X_2464_ _0352_ _0366_ _0367_ VPWR VGND sg13g2_nor2_1
X_2395_ _0304_ _0295_ _0303_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_60 VPWR VGND sg13g2_fill_2
XFILLER_29_708 VPWR VGND sg13g2_fill_1
XFILLER_3_1011 VPWR VGND sg13g2_decap_8
XFILLER_37_752 VPWR VGND sg13g2_decap_8
X_3016_ net546 VGND VPWR _0059_ mac1.products_ff\[10\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_25_969 VPWR VGND sg13g2_decap_8
XFILLER_36_284 VPWR VGND sg13g2_decap_8
XFILLER_40_939 VPWR VGND sg13g2_decap_8
XFILLER_33_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_31_clk clknet_3_1__leaf_clk clknet_leaf_31_clk VPWR VGND sg13g2_buf_8
XFILLER_20_630 VPWR VGND sg13g2_fill_1
XFILLER_32_490 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_19_229 VPWR VGND sg13g2_decap_8
XFILLER_28_752 VPWR VGND sg13g2_decap_4
XFILLER_16_925 VPWR VGND sg13g2_decap_8
XFILLER_28_774 VPWR VGND sg13g2_fill_2
XFILLER_28_785 VPWR VGND sg13g2_decap_8
XFILLER_43_722 VPWR VGND sg13g2_decap_8
XFILLER_27_273 VPWR VGND sg13g2_decap_8
XFILLER_43_755 VPWR VGND sg13g2_decap_8
XFILLER_30_405 VPWR VGND sg13g2_fill_2
XFILLER_8_38 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_22_clk clknet_3_4__leaf_clk clknet_leaf_22_clk VPWR VGND sg13g2_buf_8
XFILLER_7_623 VPWR VGND sg13g2_decap_8
XFILLER_10_162 VPWR VGND sg13g2_fill_1
XFILLER_6_155 VPWR VGND sg13g2_decap_8
X_2180_ _1457_ VPWR _1462_ VGND _1458_ _1460_ sg13g2_o21ai_1
XFILLER_19_763 VPWR VGND sg13g2_fill_1
XFILLER_18_284 VPWR VGND sg13g2_decap_8
XFILLER_22_917 VPWR VGND sg13g2_decap_8
XFILLER_34_755 VPWR VGND sg13g2_decap_8
XFILLER_15_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_13_clk clknet_3_3__leaf_clk clknet_leaf_13_clk VPWR VGND sg13g2_buf_8
X_1964_ _1271_ _1272_ _0003_ VPWR VGND sg13g2_and2_1
XFILLER_30_983 VPWR VGND sg13g2_decap_8
X_1895_ VGND VPWR _1187_ _1211_ _1218_ _1213_ sg13g2_a21oi_1
X_2516_ _0417_ _0415_ _0416_ VPWR VGND sg13g2_nand2b_1
X_2447_ _0350_ _0343_ _0039_ VPWR VGND sg13g2_xor2_1
X_2378_ VGND VPWR _0236_ _0255_ _0288_ _0257_ sg13g2_a21oi_1
XFILLER_29_527 VPWR VGND sg13g2_decap_8
XFILLER_37_582 VPWR VGND sg13g2_decap_4
XFILLER_12_405 VPWR VGND sg13g2_decap_4
XFILLER_13_939 VPWR VGND sg13g2_decap_8
XFILLER_20_460 VPWR VGND sg13g2_decap_4
XFILLER_21_994 VPWR VGND sg13g2_decap_8
XFILLER_4_637 VPWR VGND sg13g2_decap_8
XFILLER_3_125 VPWR VGND sg13g2_decap_8
XFILLER_3_169 VPWR VGND sg13g2_decap_8
XFILLER_0_832 VPWR VGND sg13g2_decap_8
XFILLER_48_814 VPWR VGND sg13g2_decap_8
Xhold9 mac1.sum_lvl1_ff\[2\] VPWR VGND net49 sg13g2_dlygate4sd3_1
XFILLER_47_379 VPWR VGND sg13g2_decap_8
XFILLER_16_700 VPWR VGND sg13g2_decap_8
XFILLER_31_714 VPWR VGND sg13g2_fill_1
XFILLER_8_921 VPWR VGND sg13g2_decap_8
XFILLER_11_460 VPWR VGND sg13g2_decap_8
XFILLER_12_961 VPWR VGND sg13g2_decap_8
XFILLER_8_998 VPWR VGND sg13g2_decap_8
X_1680_ _1010_ net411 net462 VPWR VGND sg13g2_nand2_1
X_2301_ VGND VPWR net441 net396 _0213_ _0182_ sg13g2_a21oi_1
Xclkbuf_leaf_2_clk clknet_3_2__leaf_clk clknet_leaf_2_clk VPWR VGND sg13g2_buf_8
X_2232_ VGND VPWR _0142_ _0143_ _0146_ _1492_ sg13g2_a21oi_1
XFILLER_38_302 VPWR VGND sg13g2_fill_2
XFILLER_39_869 VPWR VGND sg13g2_decap_8
X_2163_ _1443_ _1444_ _1445_ VPWR VGND sg13g2_nor2b_1
XFILLER_19_560 VPWR VGND sg13g2_decap_8
X_2094_ _1377_ _1378_ _1379_ VPWR VGND sg13g2_nor2b_2
XFILLER_0_1014 VPWR VGND sg13g2_decap_8
XFILLER_22_703 VPWR VGND sg13g2_decap_8
XFILLER_34_574 VPWR VGND sg13g2_decap_8
XFILLER_21_224 VPWR VGND sg13g2_fill_1
X_2996_ net404 _0124_ VPWR VGND sg13g2_buf_1
X_1947_ _1258_ _1255_ _1257_ VPWR VGND sg13g2_nand2_1
X_1878_ _1185_ _1177_ _1184_ _1202_ VPWR VGND sg13g2_a21o_1
XFILLER_1_618 VPWR VGND sg13g2_decap_8
XFILLER_29_313 VPWR VGND sg13g2_decap_8
XFILLER_40_544 VPWR VGND sg13g2_decap_8
XFILLER_9_718 VPWR VGND sg13g2_decap_8
XFILLER_21_791 VPWR VGND sg13g2_decap_8
XFILLER_5_902 VPWR VGND sg13g2_decap_8
XFILLER_5_979 VPWR VGND sg13g2_decap_8
XFILLER_47_110 VPWR VGND sg13g2_decap_8
XFILLER_35_338 VPWR VGND sg13g2_fill_2
XFILLER_44_894 VPWR VGND sg13g2_decap_8
XFILLER_31_522 VPWR VGND sg13g2_decap_8
X_2850_ _0740_ net376 _0739_ _0732_ net220 VPWR VGND sg13g2_a22oi_1
X_1801_ _1128_ net469 net494 VPWR VGND sg13g2_nand2_1
XFILLER_31_555 VPWR VGND sg13g2_decap_8
X_2781_ _0676_ _0610_ _0642_ VPWR VGND sg13g2_nand2_1
XFILLER_31_599 VPWR VGND sg13g2_fill_1
X_1732_ net414 net410 net459 net498 _1061_ VPWR VGND sg13g2_and4_1
Xhold217 mac1.sum_lvl2_ff\[5\] VPWR VGND net257 sg13g2_dlygate4sd3_1
XFILLER_8_795 VPWR VGND sg13g2_decap_8
XFILLER_7_283 VPWR VGND sg13g2_fill_2
XFILLER_7_272 VPWR VGND sg13g2_fill_2
X_1663_ _0993_ net471 net401 VPWR VGND sg13g2_nand2_1
Xhold206 DP_1.matrix\[1\] VPWR VGND net246 sg13g2_dlygate4sd3_1
Xhold228 DP_2.matrix\[37\] VPWR VGND net268 sg13g2_dlygate4sd3_1
Xhold239 _1266_ VPWR VGND net279 sg13g2_dlygate4sd3_1
X_1594_ _0926_ _0925_ _0922_ VPWR VGND sg13g2_nand2b_1
X_3264_ net516 VGND VPWR net15 DP_2.I_range.out_data\[4\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_22_0 VPWR VGND sg13g2_fill_2
XFILLER_22_1015 VPWR VGND sg13g2_decap_8
X_2215_ VGND VPWR _1496_ _1494_ _1451_ sg13g2_or2_1
X_3195_ net505 VGND VPWR net91 mac1.sum_lvl1_ff\[74\] clknet_leaf_38_clk sg13g2_dfrbpq_1
XFILLER_39_688 VPWR VGND sg13g2_fill_2
X_2146_ _1426_ _1427_ _1421_ _1429_ VPWR VGND sg13g2_nand3_1
X_2077_ _1362_ net455 net386 VPWR VGND sg13g2_nand2_1
XFILLER_35_894 VPWR VGND sg13g2_decap_8
XFILLER_34_382 VPWR VGND sg13g2_fill_1
X_2979_ net464 _0099_ VPWR VGND sg13g2_buf_1
XFILLER_30_25 VPWR VGND sg13g2_decap_8
XFILLER_2_916 VPWR VGND sg13g2_decap_8
XFILLER_1_437 VPWR VGND sg13g2_fill_1
XFILLER_29_143 VPWR VGND sg13g2_decap_8
XFILLER_45_625 VPWR VGND sg13g2_fill_2
XFILLER_29_165 VPWR VGND sg13g2_decap_8
XFILLER_29_198 VPWR VGND sg13g2_decap_8
XFILLER_44_179 VPWR VGND sg13g2_decap_8
XFILLER_38_1022 VPWR VGND sg13g2_decap_8
XFILLER_41_864 VPWR VGND sg13g2_decap_8
XFILLER_9_526 VPWR VGND sg13g2_decap_8
XFILLER_40_374 VPWR VGND sg13g2_fill_2
XFILLER_13_588 VPWR VGND sg13g2_decap_8
XFILLER_5_776 VPWR VGND sg13g2_decap_8
XFILLER_4_253 VPWR VGND sg13g2_decap_8
XFILLER_45_1026 VPWR VGND sg13g2_fill_2
XFILLER_1_982 VPWR VGND sg13g2_decap_8
XFILLER_49_986 VPWR VGND sg13g2_decap_8
X_2000_ _1299_ mac1.sum_lvl3_ff\[6\] net261 VPWR VGND sg13g2_xnor2_1
XFILLER_36_625 VPWR VGND sg13g2_fill_1
XFILLER_24_809 VPWR VGND sg13g2_decap_8
XFILLER_17_872 VPWR VGND sg13g2_decap_8
XFILLER_35_168 VPWR VGND sg13g2_decap_4
XFILLER_44_680 VPWR VGND sg13g2_decap_8
X_2902_ net418 net437 net378 _0791_ VPWR VGND sg13g2_mux2_1
XFILLER_32_864 VPWR VGND sg13g2_decap_8
X_2833_ _0725_ _0712_ _0724_ VPWR VGND sg13g2_xnor2_1
X_2764_ _0656_ _0658_ _0659_ VPWR VGND sg13g2_nor2_1
X_1715_ _1044_ net469 net401 VPWR VGND sg13g2_nand2_1
X_2695_ _0565_ VPWR _0592_ VGND _0559_ _0566_ sg13g2_o21ai_1
XFILLER_6_71 VPWR VGND sg13g2_fill_1
X_1646_ _0974_ _0975_ _0956_ _0977_ VPWR VGND sg13g2_nand3_1
Xfanout505 net506 net505 VPWR VGND sg13g2_buf_8
X_1577_ _0910_ _0887_ _0907_ VPWR VGND sg13g2_xnor2_1
Xfanout538 net539 net538 VPWR VGND sg13g2_buf_8
Xfanout516 net517 net516 VPWR VGND sg13g2_buf_8
Xfanout527 net528 net527 VPWR VGND sg13g2_buf_8
Xfanout549 rst_n net549 VPWR VGND sg13g2_buf_8
X_3247_ net504 VGND VPWR net264 net31 clknet_leaf_35_clk sg13g2_dfrbpq_2
X_3178_ net505 VGND VPWR net70 mac1.sum_lvl2_ff\[39\] clknet_leaf_37_clk sg13g2_dfrbpq_1
XFILLER_26_102 VPWR VGND sg13g2_decap_8
X_2129_ _1412_ _1410_ _1411_ VPWR VGND sg13g2_nand2b_1
XFILLER_26_124 VPWR VGND sg13g2_decap_8
XFILLER_42_617 VPWR VGND sg13g2_decap_8
XFILLER_41_105 VPWR VGND sg13g2_fill_2
XFILLER_41_138 VPWR VGND sg13g2_decap_4
XFILLER_2_713 VPWR VGND sg13g2_decap_8
XFILLER_9_4 VPWR VGND sg13g2_decap_8
XFILLER_2_18 VPWR VGND sg13g2_decap_8
XFILLER_49_249 VPWR VGND sg13g2_decap_8
XFILLER_46_967 VPWR VGND sg13g2_decap_8
XFILLER_45_444 VPWR VGND sg13g2_decap_8
XFILLER_14_842 VPWR VGND sg13g2_decap_8
XFILLER_40_171 VPWR VGND sg13g2_decap_8
XFILLER_9_334 VPWR VGND sg13g2_decap_8
XFILLER_13_363 VPWR VGND sg13g2_decap_8
XFILLER_15_91 VPWR VGND sg13g2_decap_4
XFILLER_12_1003 VPWR VGND sg13g2_decap_8
X_2480_ _0383_ _0382_ _0381_ VPWR VGND sg13g2_nand2b_1
X_3101_ net508 VGND VPWR _0036_ mac1.products_ff\[140\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_49_783 VPWR VGND sg13g2_decap_8
X_3032_ net548 VGND VPWR _0085_ DP_2.matrix\[44\] clknet_leaf_21_clk sg13g2_dfrbpq_2
XFILLER_48_293 VPWR VGND sg13g2_decap_4
XFILLER_37_945 VPWR VGND sg13g2_decap_8
XFILLER_24_628 VPWR VGND sg13g2_fill_2
XFILLER_32_683 VPWR VGND sg13g2_fill_2
X_2816_ _0708_ _0681_ _0709_ VPWR VGND sg13g2_xor2_1
X_2747_ VGND VPWR _0605_ _0607_ _0643_ _0641_ sg13g2_a21oi_1
XFILLER_11_38 VPWR VGND sg13g2_decap_8
X_2678_ _0576_ _0539_ _0574_ VPWR VGND sg13g2_nand2_1
X_1629_ VGND VPWR _0960_ _0958_ _0924_ sg13g2_or2_1
XFILLER_28_1021 VPWR VGND sg13g2_decap_8
Xfanout379 _0730_ net379 VPWR VGND sg13g2_buf_8
XFILLER_28_923 VPWR VGND sg13g2_decap_8
XFILLER_43_915 VPWR VGND sg13g2_decap_8
XFILLER_36_57 VPWR VGND sg13g2_fill_2
XFILLER_14_105 VPWR VGND sg13g2_fill_2
XFILLER_27_488 VPWR VGND sg13g2_fill_2
XFILLER_10_300 VPWR VGND sg13g2_fill_1
XFILLER_7_805 VPWR VGND sg13g2_decap_8
XFILLER_11_856 VPWR VGND sg13g2_decap_8
XFILLER_22_182 VPWR VGND sg13g2_fill_1
XFILLER_6_304 VPWR VGND sg13g2_fill_1
XFILLER_2_521 VPWR VGND sg13g2_decap_8
XFILLER_42_1007 VPWR VGND sg13g2_decap_8
XFILLER_2_587 VPWR VGND sg13g2_decap_8
XFILLER_19_901 VPWR VGND sg13g2_decap_8
XFILLER_18_455 VPWR VGND sg13g2_decap_8
XFILLER_19_978 VPWR VGND sg13g2_decap_8
XFILLER_34_926 VPWR VGND sg13g2_decap_8
XFILLER_45_274 VPWR VGND sg13g2_decap_8
XFILLER_33_425 VPWR VGND sg13g2_fill_1
X_1980_ mac1.sum_lvl3_ff\[1\] mac1.sum_lvl3_ff\[21\] _1284_ VPWR VGND sg13g2_nor2_1
XFILLER_21_609 VPWR VGND sg13g2_decap_4
XFILLER_13_160 VPWR VGND sg13g2_fill_1
XFILLER_20_119 VPWR VGND sg13g2_decap_8
XFILLER_9_164 VPWR VGND sg13g2_decap_4
X_2601_ _0500_ _0492_ _0499_ VPWR VGND sg13g2_nand2_1
XFILLER_6_860 VPWR VGND sg13g2_decap_8
X_2532_ _0428_ VPWR _0433_ VGND _0429_ _0431_ sg13g2_o21ai_1
X_2463_ _0366_ net491 net427 VPWR VGND sg13g2_nand2_2
X_2394_ _0303_ _0267_ _0301_ VPWR VGND sg13g2_xnor2_1
X_3015_ net546 VGND VPWR _0068_ mac1.products_ff\[9\] clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_37_731 VPWR VGND sg13g2_decap_8
XFILLER_36_241 VPWR VGND sg13g2_decap_8
XFILLER_25_948 VPWR VGND sg13g2_decap_8
XFILLER_40_918 VPWR VGND sg13g2_decap_8
XFILLER_24_458 VPWR VGND sg13g2_decap_8
XFILLER_4_819 VPWR VGND sg13g2_decap_8
XFILLER_3_307 VPWR VGND sg13g2_fill_2
XFILLER_47_528 VPWR VGND sg13g2_decap_8
XFILLER_47_89 VPWR VGND sg13g2_decap_8
XFILLER_28_731 VPWR VGND sg13g2_decap_8
XFILLER_16_904 VPWR VGND sg13g2_decap_8
XFILLER_15_414 VPWR VGND sg13g2_decap_8
XFILLER_42_244 VPWR VGND sg13g2_decap_8
XFILLER_24_992 VPWR VGND sg13g2_decap_8
XFILLER_30_417 VPWR VGND sg13g2_decap_8
XFILLER_31_929 VPWR VGND sg13g2_decap_8
XFILLER_11_653 VPWR VGND sg13g2_decap_8
XFILLER_6_123 VPWR VGND sg13g2_fill_2
XFILLER_7_679 VPWR VGND sg13g2_decap_8
XFILLER_6_178 VPWR VGND sg13g2_fill_1
XFILLER_3_885 VPWR VGND sg13g2_decap_8
XFILLER_46_550 VPWR VGND sg13g2_decap_4
XFILLER_19_775 VPWR VGND sg13g2_decap_8
XFILLER_46_594 VPWR VGND sg13g2_fill_1
XFILLER_46_572 VPWR VGND sg13g2_decap_8
XFILLER_34_734 VPWR VGND sg13g2_decap_8
XFILLER_33_244 VPWR VGND sg13g2_decap_8
XFILLER_15_970 VPWR VGND sg13g2_decap_8
XFILLER_21_428 VPWR VGND sg13g2_decap_8
XFILLER_33_255 VPWR VGND sg13g2_fill_2
X_1963_ _1267_ _1268_ _1270_ _1272_ VPWR VGND sg13g2_or3_1
XFILLER_30_962 VPWR VGND sg13g2_decap_8
X_1894_ _1216_ VPWR _1217_ VGND _1201_ _1214_ sg13g2_o21ai_1
X_2515_ _0416_ net493 net425 VPWR VGND sg13g2_nand2_2
X_2446_ _0351_ _0343_ _0350_ VPWR VGND sg13g2_nand2_1
X_2377_ _0285_ _0264_ _0287_ VPWR VGND sg13g2_xor2_1
XFILLER_13_918 VPWR VGND sg13g2_decap_8
XFILLER_25_745 VPWR VGND sg13g2_decap_8
XFILLER_33_25 VPWR VGND sg13g2_fill_2
XFILLER_24_299 VPWR VGND sg13g2_fill_2
XFILLER_33_47 VPWR VGND sg13g2_decap_8
XFILLER_33_58 VPWR VGND sg13g2_fill_2
XFILLER_21_973 VPWR VGND sg13g2_decap_8
XFILLER_0_811 VPWR VGND sg13g2_decap_8
XFILLER_0_888 VPWR VGND sg13g2_decap_8
XFILLER_28_572 VPWR VGND sg13g2_decap_8
XFILLER_15_266 VPWR VGND sg13g2_decap_8
XFILLER_16_789 VPWR VGND sg13g2_decap_8
XFILLER_12_940 VPWR VGND sg13g2_decap_8
XFILLER_30_225 VPWR VGND sg13g2_decap_4
XFILLER_30_236 VPWR VGND sg13g2_fill_1
XFILLER_31_737 VPWR VGND sg13g2_fill_1
XFILLER_31_748 VPWR VGND sg13g2_decap_8
XFILLER_8_900 VPWR VGND sg13g2_decap_8
XFILLER_8_977 VPWR VGND sg13g2_decap_8
XFILLER_48_1024 VPWR VGND sg13g2_decap_4
XFILLER_3_682 VPWR VGND sg13g2_decap_8
X_2300_ _0186_ VPWR _0212_ VGND _0180_ _0187_ sg13g2_o21ai_1
X_2231_ _0142_ _0143_ _1492_ _0145_ VPWR VGND sg13g2_nand3_1
XFILLER_24_4 VPWR VGND sg13g2_decap_8
X_2162_ net455 net382 net458 _1444_ VPWR VGND net380 sg13g2_nand4_1
X_2093_ _1357_ VPWR _1378_ VGND _1348_ _1358_ sg13g2_o21ai_1
XFILLER_38_347 VPWR VGND sg13g2_fill_1
XFILLER_47_892 VPWR VGND sg13g2_decap_8
XFILLER_46_391 VPWR VGND sg13g2_decap_8
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_34_531 VPWR VGND sg13g2_decap_4
XFILLER_9_60 VPWR VGND sg13g2_fill_1
XFILLER_21_269 VPWR VGND sg13g2_decap_4
X_2995_ net158 _0123_ VPWR VGND sg13g2_buf_1
X_1946_ _0015_ _1254_ net295 VPWR VGND sg13g2_xnor2_1
X_1877_ VGND VPWR _1176_ _1190_ _1201_ _1189_ sg13g2_a21oi_1
X_2429_ VGND VPWR _0305_ _0329_ _0336_ _0331_ sg13g2_a21oi_1
XFILLER_29_336 VPWR VGND sg13g2_decap_8
XFILLER_25_531 VPWR VGND sg13g2_decap_8
XFILLER_44_68 VPWR VGND sg13g2_decap_4
XFILLER_25_586 VPWR VGND sg13g2_decap_8
XFILLER_40_589 VPWR VGND sg13g2_decap_8
XFILLER_5_958 VPWR VGND sg13g2_decap_8
XFILLER_4_435 VPWR VGND sg13g2_decap_8
XFILLER_0_685 VPWR VGND sg13g2_decap_8
XFILLER_47_188 VPWR VGND sg13g2_decap_8
XFILLER_29_892 VPWR VGND sg13g2_decap_8
XFILLER_16_531 VPWR VGND sg13g2_decap_8
XFILLER_28_380 VPWR VGND sg13g2_decap_4
XFILLER_44_873 VPWR VGND sg13g2_decap_8
XFILLER_43_383 VPWR VGND sg13g2_decap_8
XFILLER_15_1012 VPWR VGND sg13g2_decap_8
X_1800_ VGND VPWR _1127_ _1097_ _1095_ sg13g2_or2_1
X_2780_ _0613_ _0674_ _0675_ VPWR VGND sg13g2_nor2b_1
XFILLER_12_770 VPWR VGND sg13g2_decap_8
XFILLER_8_774 VPWR VGND sg13g2_decap_8
XFILLER_11_291 VPWR VGND sg13g2_fill_1
X_1731_ _1060_ net410 net498 VPWR VGND sg13g2_nand2_1
X_1662_ _0992_ net475 net494 VPWR VGND sg13g2_nand2_1
Xhold207 _0817_ VPWR VGND net247 sg13g2_dlygate4sd3_1
Xhold218 _1240_ VPWR VGND net258 sg13g2_dlygate4sd3_1
Xhold229 _0043_ VPWR VGND net269 sg13g2_dlygate4sd3_1
XFILLER_4_980 VPWR VGND sg13g2_decap_8
X_1593_ _0924_ _0889_ _0925_ VPWR VGND sg13g2_xor2_1
X_3263_ net516 VGND VPWR net14 DP_2.I_range.out_data\[3\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_3194_ net505 VGND VPWR net48 mac1.sum_lvl1_ff\[73\] clknet_leaf_37_clk sg13g2_dfrbpq_1
X_2214_ _1495_ net444 net388 VPWR VGND sg13g2_nand2_1
XFILLER_39_667 VPWR VGND sg13g2_decap_8
X_2145_ _1428_ _1421_ _1426_ _1427_ VPWR VGND sg13g2_and3_1
XFILLER_27_829 VPWR VGND sg13g2_decap_8
X_2076_ _1361_ net386 net457 net388 net454 VPWR VGND sg13g2_a22oi_1
XFILLER_35_840 VPWR VGND sg13g2_fill_2
Xclkbuf_3_5__f_clk clknet_0_clk clknet_3_5__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_34_350 VPWR VGND sg13g2_decap_8
XFILLER_35_873 VPWR VGND sg13g2_decap_8
XFILLER_22_534 VPWR VGND sg13g2_fill_2
XFILLER_14_49 VPWR VGND sg13g2_decap_8
XFILLER_22_556 VPWR VGND sg13g2_decap_4
X_2978_ net467 _0098_ VPWR VGND sg13g2_buf_1
X_1929_ _1239_ net297 _1243_ _1244_ VPWR VGND sg13g2_nor3_2
XFILLER_29_111 VPWR VGND sg13g2_decap_8
XFILLER_45_604 VPWR VGND sg13g2_decap_8
XFILLER_29_133 VPWR VGND sg13g2_decap_4
XFILLER_44_136 VPWR VGND sg13g2_fill_2
XFILLER_38_1001 VPWR VGND sg13g2_decap_8
XFILLER_13_534 VPWR VGND sg13g2_decap_4
XFILLER_26_895 VPWR VGND sg13g2_decap_8
XFILLER_13_567 VPWR VGND sg13g2_decap_8
XFILLER_5_755 VPWR VGND sg13g2_decap_8
XFILLER_45_1005 VPWR VGND sg13g2_decap_8
XFILLER_1_961 VPWR VGND sg13g2_decap_8
XFILLER_0_482 VPWR VGND sg13g2_decap_8
XFILLER_49_965 VPWR VGND sg13g2_decap_8
XFILLER_48_475 VPWR VGND sg13g2_decap_8
Xhold90 mac1.products_ff\[12\] VPWR VGND net130 sg13g2_dlygate4sd3_1
XFILLER_36_604 VPWR VGND sg13g2_decap_8
XFILLER_36_637 VPWR VGND sg13g2_decap_4
XFILLER_35_136 VPWR VGND sg13g2_decap_8
XFILLER_16_383 VPWR VGND sg13g2_fill_1
X_2901_ _0790_ net377 _0789_ _0783_ net389 VPWR VGND sg13g2_a22oi_1
X_2832_ _0724_ _0721_ _0723_ VPWR VGND sg13g2_xnor2_1
X_2763_ _0658_ net422 net482 net424 net479 VPWR VGND sg13g2_a22oi_1
XFILLER_8_582 VPWR VGND sg13g2_decap_4
X_1714_ _1043_ net473 net494 VPWR VGND sg13g2_nand2_1
X_2694_ _0589_ _0581_ _0591_ VPWR VGND sg13g2_xor2_1
X_1645_ _0976_ _0956_ _0974_ _0975_ VPWR VGND sg13g2_and3_1
Xfanout506 net508 net506 VPWR VGND sg13g2_buf_8
X_1576_ VGND VPWR _0905_ _0906_ _0909_ _0887_ sg13g2_a21oi_1
Xfanout528 net533 net528 VPWR VGND sg13g2_buf_8
Xfanout539 net549 net539 VPWR VGND sg13g2_buf_8
Xfanout517 net518 net517 VPWR VGND sg13g2_buf_8
XFILLER_6_1021 VPWR VGND sg13g2_decap_8
X_3246_ net503 VGND VPWR net180 net30 clknet_leaf_34_clk sg13g2_dfrbpq_2
XFILLER_39_431 VPWR VGND sg13g2_decap_4
X_3177_ net505 VGND VPWR net56 mac1.sum_lvl2_ff\[38\] clknet_leaf_38_clk sg13g2_dfrbpq_1
XFILLER_39_497 VPWR VGND sg13g2_decap_8
X_2128_ _1411_ net457 net382 VPWR VGND sg13g2_nand2_1
XFILLER_26_136 VPWR VGND sg13g2_decap_8
XFILLER_27_648 VPWR VGND sg13g2_decap_8
X_2059_ _1344_ _1345_ _1346_ VPWR VGND sg13g2_nor2b_1
XFILLER_23_832 VPWR VGND sg13g2_decap_4
XFILLER_23_898 VPWR VGND sg13g2_decap_8
XFILLER_41_47 VPWR VGND sg13g2_decap_8
XFILLER_41_25 VPWR VGND sg13g2_decap_8
XFILLER_1_268 VPWR VGND sg13g2_decap_4
XFILLER_2_769 VPWR VGND sg13g2_decap_8
XFILLER_49_228 VPWR VGND sg13g2_decap_8
XFILLER_17_103 VPWR VGND sg13g2_decap_4
XFILLER_46_946 VPWR VGND sg13g2_decap_8
XFILLER_45_423 VPWR VGND sg13g2_decap_8
XFILLER_45_467 VPWR VGND sg13g2_fill_1
XFILLER_14_810 VPWR VGND sg13g2_decap_8
XFILLER_14_821 VPWR VGND sg13g2_fill_1
XFILLER_41_640 VPWR VGND sg13g2_decap_4
XFILLER_13_342 VPWR VGND sg13g2_decap_8
XFILLER_41_684 VPWR VGND sg13g2_fill_2
XFILLER_14_898 VPWR VGND sg13g2_decap_8
XFILLER_5_574 VPWR VGND sg13g2_fill_1
XFILLER_5_552 VPWR VGND sg13g2_fill_2
X_3100_ net508 VGND VPWR _0035_ mac1.products_ff\[139\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_49_762 VPWR VGND sg13g2_decap_8
X_3031_ net538 VGND VPWR net228 DP_2.matrix\[8\] clknet_leaf_13_clk sg13g2_dfrbpq_2
XFILLER_37_924 VPWR VGND sg13g2_decap_8
XFILLER_48_272 VPWR VGND sg13g2_decap_8
XFILLER_24_607 VPWR VGND sg13g2_decap_8
XFILLER_36_456 VPWR VGND sg13g2_decap_4
X_2815_ _0708_ net500 net425 VPWR VGND sg13g2_nand2_1
X_2746_ _0607_ _0641_ _0605_ _0642_ VPWR VGND sg13g2_nand3_1
X_2677_ _0539_ _0574_ _0575_ VPWR VGND sg13g2_nor2_1
X_1628_ _0959_ net409 net467 VPWR VGND sg13g2_nand2_1
XFILLER_28_1000 VPWR VGND sg13g2_decap_8
X_1559_ _0867_ _0890_ _0892_ VPWR VGND sg13g2_and2_1
XFILLER_46_209 VPWR VGND sg13g2_decap_8
X_3229_ net510 VGND VPWR net267 mac1.sum_lvl3_ff\[4\] clknet_leaf_34_clk sg13g2_dfrbpq_1
XFILLER_28_902 VPWR VGND sg13g2_decap_8
XFILLER_27_423 VPWR VGND sg13g2_fill_2
XFILLER_36_36 VPWR VGND sg13g2_decap_8
XFILLER_39_294 VPWR VGND sg13g2_decap_8
XFILLER_15_607 VPWR VGND sg13g2_decap_8
XFILLER_15_618 VPWR VGND sg13g2_fill_1
XFILLER_28_979 VPWR VGND sg13g2_decap_8
XFILLER_11_835 VPWR VGND sg13g2_decap_8
XFILLER_2_544 VPWR VGND sg13g2_decap_8
XFILLER_46_721 VPWR VGND sg13g2_fill_1
XFILLER_19_957 VPWR VGND sg13g2_decap_8
XFILLER_46_765 VPWR VGND sg13g2_decap_4
XFILLER_45_253 VPWR VGND sg13g2_decap_8
XFILLER_34_905 VPWR VGND sg13g2_decap_8
XFILLER_46_798 VPWR VGND sg13g2_fill_2
XFILLER_45_297 VPWR VGND sg13g2_fill_1
XFILLER_42_993 VPWR VGND sg13g2_decap_8
XFILLER_13_194 VPWR VGND sg13g2_decap_8
XFILLER_9_198 VPWR VGND sg13g2_decap_8
X_2600_ _0497_ _0493_ _0499_ VPWR VGND sg13g2_xor2_1
X_2531_ _0428_ _0429_ _0431_ _0432_ VPWR VGND sg13g2_or3_1
X_2462_ _0365_ net427 net492 net429 net490 VPWR VGND sg13g2_a22oi_1
X_2393_ _0267_ _0301_ _0302_ VPWR VGND sg13g2_nor2b_1
XFILLER_49_592 VPWR VGND sg13g2_decap_8
X_3014_ net543 VGND VPWR _0067_ mac1.products_ff\[8\] clknet_leaf_24_clk sg13g2_dfrbpq_1
XFILLER_25_927 VPWR VGND sg13g2_decap_8
XFILLER_24_437 VPWR VGND sg13g2_decap_8
X_2729_ _0619_ _0624_ _0625_ VPWR VGND sg13g2_and2_1
XFILLER_47_507 VPWR VGND sg13g2_decap_8
XFILLER_47_35 VPWR VGND sg13g2_decap_8
XFILLER_47_68 VPWR VGND sg13g2_decap_8
XFILLER_28_710 VPWR VGND sg13g2_fill_2
XFILLER_42_201 VPWR VGND sg13g2_fill_1
XFILLER_15_404 VPWR VGND sg13g2_decap_4
XFILLER_27_297 VPWR VGND sg13g2_decap_4
XFILLER_31_908 VPWR VGND sg13g2_decap_8
XFILLER_43_779 VPWR VGND sg13g2_decap_8
XFILLER_42_278 VPWR VGND sg13g2_fill_2
XFILLER_42_267 VPWR VGND sg13g2_decap_8
XFILLER_24_971 VPWR VGND sg13g2_decap_8
XFILLER_11_632 VPWR VGND sg13g2_decap_8
XFILLER_23_492 VPWR VGND sg13g2_decap_8
XFILLER_6_102 VPWR VGND sg13g2_decap_8
XFILLER_12_71 VPWR VGND sg13g2_decap_8
XFILLER_3_864 VPWR VGND sg13g2_decap_8
XFILLER_2_385 VPWR VGND sg13g2_fill_2
XFILLER_38_529 VPWR VGND sg13g2_decap_8
XFILLER_19_754 VPWR VGND sg13g2_fill_2
XFILLER_18_1021 VPWR VGND sg13g2_decap_8
XFILLER_21_407 VPWR VGND sg13g2_decap_8
XFILLER_14_481 VPWR VGND sg13g2_decap_8
X_1962_ _1267_ VPWR _1271_ VGND _1268_ _1270_ sg13g2_o21ai_1
XFILLER_30_941 VPWR VGND sg13g2_decap_8
X_1893_ _0074_ _1200_ _1215_ VPWR VGND sg13g2_xnor2_1
X_2514_ _0391_ VPWR _0415_ VGND _0366_ _0389_ sg13g2_o21ai_1
X_2445_ _0348_ _0349_ _0350_ VPWR VGND sg13g2_nor2b_1
XFILLER_25_1025 VPWR VGND sg13g2_decap_4
X_2376_ _0285_ _0264_ _0286_ VPWR VGND sg13g2_nor2b_1
XFILLER_25_724 VPWR VGND sg13g2_decap_8
XFILLER_40_749 VPWR VGND sg13g2_decap_8
XFILLER_21_952 VPWR VGND sg13g2_decap_8
XFILLER_32_1018 VPWR VGND sg13g2_decap_8
XFILLER_0_867 VPWR VGND sg13g2_decap_8
XFILLER_48_849 VPWR VGND sg13g2_decap_8
XFILLER_47_337 VPWR VGND sg13g2_fill_1
XFILLER_43_532 VPWR VGND sg13g2_decap_8
XFILLER_16_768 VPWR VGND sg13g2_decap_4
XFILLER_15_245 VPWR VGND sg13g2_decap_8
XFILLER_30_259 VPWR VGND sg13g2_decap_8
XFILLER_8_956 VPWR VGND sg13g2_decap_8
XFILLER_12_996 VPWR VGND sg13g2_decap_8
XFILLER_7_466 VPWR VGND sg13g2_decap_8
XFILLER_48_1003 VPWR VGND sg13g2_decap_8
XFILLER_3_661 VPWR VGND sg13g2_decap_8
X_2230_ _0144_ _1492_ _0142_ _0143_ VPWR VGND sg13g2_and3_1
X_2161_ _1443_ net380 net458 net382 net455 VPWR VGND sg13g2_a22oi_1
XFILLER_38_326 VPWR VGND sg13g2_decap_8
X_2092_ _1377_ _1365_ _1376_ VPWR VGND sg13g2_xnor2_1
XFILLER_47_871 VPWR VGND sg13g2_decap_8
XFILLER_34_510 VPWR VGND sg13g2_decap_8
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_22_738 VPWR VGND sg13g2_decap_8
X_2994_ net407 _0122_ VPWR VGND sg13g2_buf_1
X_1945_ _1256_ VPWR _1257_ VGND _1250_ _1252_ sg13g2_o21ai_1
XFILLER_21_248 VPWR VGND sg13g2_decap_4
XFILLER_9_83 VPWR VGND sg13g2_fill_2
XFILLER_30_771 VPWR VGND sg13g2_decap_8
X_1876_ _1197_ _1199_ _1200_ VPWR VGND sg13g2_nor2_1
XFILLER_0_119 VPWR VGND sg13g2_decap_8
X_2428_ VGND VPWR _0318_ _0334_ _0335_ _0333_ sg13g2_a21oi_1
X_2359_ _0248_ VPWR _0269_ VGND _0246_ _0249_ sg13g2_o21ai_1
XFILLER_44_329 VPWR VGND sg13g2_decap_8
XFILLER_38_882 VPWR VGND sg13g2_decap_8
XFILLER_44_47 VPWR VGND sg13g2_decap_8
XFILLER_25_554 VPWR VGND sg13g2_decap_4
XFILLER_25_598 VPWR VGND sg13g2_decap_4
XFILLER_40_579 VPWR VGND sg13g2_decap_4
XFILLER_12_248 VPWR VGND sg13g2_decap_8
XFILLER_5_937 VPWR VGND sg13g2_decap_8
XFILLER_0_664 VPWR VGND sg13g2_decap_8
XFILLER_47_145 VPWR VGND sg13g2_fill_2
XFILLER_47_167 VPWR VGND sg13g2_decap_8
XFILLER_29_871 VPWR VGND sg13g2_decap_8
XFILLER_44_852 VPWR VGND sg13g2_decap_8
XFILLER_28_392 VPWR VGND sg13g2_fill_2
XFILLER_43_351 VPWR VGND sg13g2_fill_2
XFILLER_16_565 VPWR VGND sg13g2_decap_4
XFILLER_31_502 VPWR VGND sg13g2_decap_8
XFILLER_8_753 VPWR VGND sg13g2_decap_8
XFILLER_12_793 VPWR VGND sg13g2_decap_8
X_1730_ _1012_ VPWR _1059_ VGND _1010_ _1013_ sg13g2_o21ai_1
X_1661_ _0960_ VPWR _0991_ VGND _0957_ _0961_ sg13g2_o21ai_1
Xhold208 _0087_ VPWR VGND net248 sg13g2_dlygate4sd3_1
Xhold219 _0011_ VPWR VGND net259 sg13g2_dlygate4sd3_1
X_1592_ _0924_ net469 net408 VPWR VGND sg13g2_nand2_1
X_3262_ net516 VGND VPWR net13 DP_2.I_range.out_data\[2\] clknet_leaf_11_clk sg13g2_dfrbpq_2
XFILLER_39_602 VPWR VGND sg13g2_decap_8
XFILLER_39_635 VPWR VGND sg13g2_decap_8
X_3193_ net503 VGND VPWR net131 mac1.sum_lvl1_ff\[72\] clknet_leaf_38_clk sg13g2_dfrbpq_1
X_2213_ _1494_ net445 net386 VPWR VGND sg13g2_nand2_2
X_2144_ _1422_ VPWR _1427_ VGND _1423_ _1425_ sg13g2_o21ai_1
X_2075_ _0035_ _1347_ _1359_ VPWR VGND sg13g2_xnor2_1
XFILLER_19_381 VPWR VGND sg13g2_decap_8
XFILLER_35_852 VPWR VGND sg13g2_decap_8
XFILLER_10_719 VPWR VGND sg13g2_decap_8
X_2977_ net468 _0097_ VPWR VGND sg13g2_buf_1
X_1928_ VPWR VGND _1237_ _1236_ _1235_ mac1.sum_lvl2_ff\[24\] _1243_ net257 sg13g2_a221oi_1
X_1859_ _1148_ _1183_ _1184_ VPWR VGND sg13g2_nor2b_1
XFILLER_39_69 VPWR VGND sg13g2_decap_8
XFILLER_18_808 VPWR VGND sg13g2_decap_8
XFILLER_18_819 VPWR VGND sg13g2_fill_2
XFILLER_41_822 VPWR VGND sg13g2_decap_8
XFILLER_40_310 VPWR VGND sg13g2_decap_4
XFILLER_25_384 VPWR VGND sg13g2_decap_8
XFILLER_41_899 VPWR VGND sg13g2_decap_8
XFILLER_5_734 VPWR VGND sg13g2_decap_8
XFILLER_45_1028 VPWR VGND sg13g2_fill_1
XFILLER_1_940 VPWR VGND sg13g2_decap_8
XFILLER_49_944 VPWR VGND sg13g2_decap_8
XFILLER_0_461 VPWR VGND sg13g2_decap_8
Xhold80 mac1.sum_lvl1_ff\[14\] VPWR VGND net120 sg13g2_dlygate4sd3_1
Xhold91 mac1.products_ff\[136\] VPWR VGND net131 sg13g2_dlygate4sd3_1
XFILLER_35_104 VPWR VGND sg13g2_fill_2
XFILLER_17_841 VPWR VGND sg13g2_decap_8
XFILLER_29_690 VPWR VGND sg13g2_decap_8
XFILLER_16_351 VPWR VGND sg13g2_fill_2
XFILLER_16_362 VPWR VGND sg13g2_decap_8
XFILLER_31_310 VPWR VGND sg13g2_fill_2
XFILLER_32_822 VPWR VGND sg13g2_decap_8
X_2900_ net408 net429 net378 _0789_ VPWR VGND sg13g2_mux2_1
X_2831_ _0722_ _0707_ _0723_ VPWR VGND sg13g2_xor2_1
XFILLER_32_899 VPWR VGND sg13g2_decap_8
X_2762_ VGND VPWR _0657_ _0655_ _0631_ sg13g2_or2_1
XFILLER_8_572 VPWR VGND sg13g2_fill_2
X_1713_ _1006_ VPWR _1042_ VGND _1003_ _1007_ sg13g2_o21ai_1
X_2693_ _0589_ _0581_ _0590_ VPWR VGND sg13g2_nor2b_1
X_1644_ _0963_ VPWR _0975_ VGND _0971_ _0973_ sg13g2_o21ai_1
XFILLER_6_95 VPWR VGND sg13g2_decap_8
X_1575_ _0905_ _0906_ _0887_ _0908_ VPWR VGND sg13g2_nand3_1
Xfanout507 net508 net507 VPWR VGND sg13g2_buf_8
Xfanout529 net532 net529 VPWR VGND sg13g2_buf_8
Xfanout518 net519 net518 VPWR VGND sg13g2_buf_8
XFILLER_39_410 VPWR VGND sg13g2_decap_8
XFILLER_6_1000 VPWR VGND sg13g2_decap_8
X_3245_ net503 VGND VPWR net219 net29 clknet_leaf_34_clk sg13g2_dfrbpq_2
XFILLER_39_476 VPWR VGND sg13g2_fill_1
XFILLER_27_627 VPWR VGND sg13g2_decap_8
X_3176_ net545 VGND VPWR net149 mac1.sum_lvl2_ff\[34\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2127_ _1387_ VPWR _1410_ VGND _1362_ _1385_ sg13g2_o21ai_1
X_2058_ _1341_ VPWR _1345_ VGND _1342_ _1343_ sg13g2_o21ai_1
XFILLER_26_159 VPWR VGND sg13g2_decap_8
XFILLER_34_170 VPWR VGND sg13g2_fill_1
XFILLER_35_671 VPWR VGND sg13g2_fill_2
XFILLER_23_877 VPWR VGND sg13g2_decap_8
XFILLER_22_398 VPWR VGND sg13g2_decap_4
XFILLER_2_748 VPWR VGND sg13g2_decap_8
XFILLER_49_207 VPWR VGND sg13g2_decap_8
XFILLER_46_925 VPWR VGND sg13g2_decap_8
XFILLER_17_126 VPWR VGND sg13g2_decap_8
XFILLER_18_638 VPWR VGND sg13g2_decap_8
XFILLER_18_649 VPWR VGND sg13g2_fill_2
XFILLER_41_663 VPWR VGND sg13g2_decap_8
XFILLER_40_140 VPWR VGND sg13g2_decap_8
XFILLER_14_877 VPWR VGND sg13g2_decap_8
XFILLER_31_92 VPWR VGND sg13g2_decap_8
XFILLER_49_7 VPWR VGND sg13g2_decap_8
XFILLER_49_741 VPWR VGND sg13g2_decap_8
XFILLER_0_291 VPWR VGND sg13g2_decap_8
XFILLER_48_251 VPWR VGND sg13g2_decap_8
X_3030_ net532 VGND VPWR _0083_ DP_1.matrix\[80\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_37_903 VPWR VGND sg13g2_decap_8
XFILLER_45_991 VPWR VGND sg13g2_decap_8
XFILLER_23_129 VPWR VGND sg13g2_fill_2
XFILLER_32_630 VPWR VGND sg13g2_fill_1
XFILLER_32_674 VPWR VGND sg13g2_fill_1
X_2814_ _0707_ net500 net421 VPWR VGND sg13g2_nand2_1
XFILLER_20_836 VPWR VGND sg13g2_decap_8
XFILLER_20_847 VPWR VGND sg13g2_fill_1
XFILLER_31_162 VPWR VGND sg13g2_decap_8
XFILLER_20_869 VPWR VGND sg13g2_decap_8
X_2745_ _0639_ _0617_ _0641_ VPWR VGND sg13g2_xor2_1
X_2676_ _0574_ _0540_ _0572_ VPWR VGND sg13g2_xnor2_1
X_1627_ _0958_ net467 net406 VPWR VGND sg13g2_nand2_1
X_1558_ VGND VPWR _0891_ _0890_ _0867_ sg13g2_or2_1
X_3228_ net510 VGND VPWR net245 mac1.sum_lvl3_ff\[3\] clknet_leaf_34_clk sg13g2_dfrbpq_1
XFILLER_27_402 VPWR VGND sg13g2_decap_8
XFILLER_39_251 VPWR VGND sg13g2_decap_8
X_3159_ net545 VGND VPWR net120 mac1.sum_lvl2_ff\[14\] clknet_leaf_16_clk sg13g2_dfrbpq_2
XFILLER_28_958 VPWR VGND sg13g2_decap_8
XFILLER_36_15 VPWR VGND sg13g2_decap_8
XFILLER_39_284 VPWR VGND sg13g2_decap_4
XFILLER_27_446 VPWR VGND sg13g2_decap_8
XFILLER_36_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_34_clk clknet_3_1__leaf_clk clknet_leaf_34_clk VPWR VGND sg13g2_buf_8
XFILLER_23_674 VPWR VGND sg13g2_decap_8
XFILLER_35_1027 VPWR VGND sg13g2_fill_2
XFILLER_10_324 VPWR VGND sg13g2_fill_2
XFILLER_22_195 VPWR VGND sg13g2_decap_8
XFILLER_46_744 VPWR VGND sg13g2_decap_8
XFILLER_18_435 VPWR VGND sg13g2_fill_1
XFILLER_19_936 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_25_clk clknet_3_5__leaf_clk clknet_leaf_25_clk VPWR VGND sg13g2_buf_8
XFILLER_26_70 VPWR VGND sg13g2_decap_8
XFILLER_42_972 VPWR VGND sg13g2_decap_8
XFILLER_9_133 VPWR VGND sg13g2_decap_4
XFILLER_10_880 VPWR VGND sg13g2_decap_8
XFILLER_9_177 VPWR VGND sg13g2_decap_8
X_2530_ _0431_ net435 net481 net480 net438 VPWR VGND sg13g2_a22oi_1
XFILLER_6_895 VPWR VGND sg13g2_decap_8
X_2461_ _0363_ _0351_ _0040_ VPWR VGND sg13g2_xor2_1
X_2392_ _0301_ _0296_ _0299_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_96 VPWR VGND sg13g2_fill_2
X_3013_ net536 VGND VPWR _0066_ mac1.products_ff\[7\] clknet_leaf_26_clk sg13g2_dfrbpq_1
XFILLER_3_1025 VPWR VGND sg13g2_decap_4
XFILLER_25_906 VPWR VGND sg13g2_decap_8
XFILLER_37_766 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_16_clk clknet_3_7__leaf_clk clknet_leaf_16_clk VPWR VGND sg13g2_buf_8
XFILLER_20_600 VPWR VGND sg13g2_decap_8
XFILLER_32_471 VPWR VGND sg13g2_decap_8
XFILLER_32_482 VPWR VGND sg13g2_fill_1
XFILLER_33_994 VPWR VGND sg13g2_decap_8
XFILLER_20_666 VPWR VGND sg13g2_decap_8
X_2728_ _0623_ _0620_ _0624_ VPWR VGND sg13g2_xor2_1
XFILLER_3_309 VPWR VGND sg13g2_fill_1
X_2659_ _0505_ _0555_ _0557_ VPWR VGND sg13g2_and2_1
XFILLER_47_14 VPWR VGND sg13g2_decap_8
XFILLER_43_736 VPWR VGND sg13g2_decap_4
XFILLER_16_939 VPWR VGND sg13g2_decap_8
XFILLER_28_799 VPWR VGND sg13g2_decap_8
XFILLER_43_769 VPWR VGND sg13g2_fill_1
XFILLER_27_287 VPWR VGND sg13g2_fill_1
XFILLER_24_950 VPWR VGND sg13g2_decap_8
XFILLER_6_125 VPWR VGND sg13g2_fill_1
XFILLER_11_688 VPWR VGND sg13g2_fill_2
XFILLER_6_169 VPWR VGND sg13g2_decap_8
XFILLER_3_843 VPWR VGND sg13g2_decap_8
XFILLER_19_700 VPWR VGND sg13g2_decap_8
XFILLER_38_519 VPWR VGND sg13g2_fill_1
XFILLER_34_703 VPWR VGND sg13g2_decap_8
XFILLER_18_298 VPWR VGND sg13g2_decap_8
XFILLER_34_769 VPWR VGND sg13g2_decap_8
XFILLER_18_1000 VPWR VGND sg13g2_decap_8
X_1961_ VGND VPWR _1255_ _1257_ _1270_ _1269_ sg13g2_a21oi_1
XFILLER_30_920 VPWR VGND sg13g2_decap_8
X_1892_ _1215_ VPWR _1216_ VGND _1197_ _1199_ sg13g2_o21ai_1
XFILLER_30_997 VPWR VGND sg13g2_decap_8
X_2513_ _0405_ VPWR _0414_ VGND _0368_ _0406_ sg13g2_o21ai_1
XFILLER_6_692 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_5_clk clknet_3_4__leaf_clk clknet_leaf_5_clk VPWR VGND sg13g2_buf_8
X_2444_ _0345_ VPWR _0349_ VGND _0346_ _0347_ sg13g2_o21ai_1
XFILLER_25_1004 VPWR VGND sg13g2_decap_8
X_2375_ _0283_ _0282_ _0285_ VPWR VGND sg13g2_xor2_1
XFILLER_29_508 VPWR VGND sg13g2_decap_4
XFILLER_17_39 VPWR VGND sg13g2_decap_8
XFILLER_25_703 VPWR VGND sg13g2_decap_8
XFILLER_40_728 VPWR VGND sg13g2_decap_8
XFILLER_21_931 VPWR VGND sg13g2_decap_8
XFILLER_33_780 VPWR VGND sg13g2_decap_8
XFILLER_20_485 VPWR VGND sg13g2_decap_4
XFILLER_0_846 VPWR VGND sg13g2_decap_8
XFILLER_48_828 VPWR VGND sg13g2_decap_8
XFILLER_47_316 VPWR VGND sg13g2_decap_8
XFILLER_43_511 VPWR VGND sg13g2_decap_8
XFILLER_16_714 VPWR VGND sg13g2_decap_4
XFILLER_15_224 VPWR VGND sg13g2_decap_8
XFILLER_16_747 VPWR VGND sg13g2_decap_8
XFILLER_8_935 VPWR VGND sg13g2_decap_8
XFILLER_11_474 VPWR VGND sg13g2_fill_2
XFILLER_12_975 VPWR VGND sg13g2_decap_8
XFILLER_23_82 VPWR VGND sg13g2_fill_2
XFILLER_3_640 VPWR VGND sg13g2_decap_8
XFILLER_2_183 VPWR VGND sg13g2_decap_8
XFILLER_39_828 VPWR VGND sg13g2_decap_8
X_2160_ _1419_ VPWR _1442_ VGND _1384_ _1417_ sg13g2_o21ai_1
XFILLER_47_850 VPWR VGND sg13g2_decap_8
X_2091_ _1376_ _1373_ _1375_ VPWR VGND sg13g2_nand2_1
XFILLER_46_360 VPWR VGND sg13g2_fill_2
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_0_1028 VPWR VGND sg13g2_fill_1
XFILLER_22_717 VPWR VGND sg13g2_decap_8
XFILLER_34_555 VPWR VGND sg13g2_decap_4
X_2993_ net408 _0121_ VPWR VGND sg13g2_buf_1
XFILLER_34_588 VPWR VGND sg13g2_decap_8
X_1944_ net294 mac1.sum_lvl2_ff\[28\] _1256_ VPWR VGND sg13g2_xor2_1
XFILLER_30_761 VPWR VGND sg13g2_decap_4
X_1875_ _1199_ _1192_ _1198_ VPWR VGND sg13g2_nand2_1
X_2427_ _0334_ _0318_ _0052_ VPWR VGND sg13g2_xor2_1
XFILLER_28_16 VPWR VGND sg13g2_decap_4
X_2358_ _0268_ _0267_ _0265_ VPWR VGND sg13g2_nand2b_1
XFILLER_45_809 VPWR VGND sg13g2_decap_8
XFILLER_28_49 VPWR VGND sg13g2_decap_8
X_2289_ _0169_ VPWR _0201_ VGND _1483_ _0167_ sg13g2_o21ai_1
XFILLER_44_308 VPWR VGND sg13g2_decap_8
XFILLER_37_360 VPWR VGND sg13g2_fill_1
XFILLER_38_861 VPWR VGND sg13g2_decap_8
XFILLER_44_15 VPWR VGND sg13g2_decap_8
XFILLER_37_382 VPWR VGND sg13g2_fill_2
XFILLER_37_393 VPWR VGND sg13g2_fill_2
XFILLER_40_525 VPWR VGND sg13g2_fill_2
XFILLER_40_514 VPWR VGND sg13g2_decap_8
XFILLER_40_569 VPWR VGND sg13g2_fill_2
XFILLER_5_916 VPWR VGND sg13g2_decap_8
XFILLER_4_459 VPWR VGND sg13g2_decap_8
XFILLER_0_643 VPWR VGND sg13g2_decap_8
XFILLER_47_124 VPWR VGND sg13g2_decap_8
XFILLER_35_308 VPWR VGND sg13g2_fill_2
XFILLER_44_831 VPWR VGND sg13g2_decap_8
XFILLER_18_93 VPWR VGND sg13g2_decap_8
XFILLER_31_536 VPWR VGND sg13g2_decap_8
XFILLER_31_569 VPWR VGND sg13g2_decap_8
XFILLER_8_732 VPWR VGND sg13g2_decap_8
X_1660_ _0977_ VPWR _0990_ VGND _0955_ _0978_ sg13g2_o21ai_1
X_1591_ _0923_ net469 net406 VPWR VGND sg13g2_nand2_1
Xhold209 DP_1.matrix\[2\] VPWR VGND net249 sg13g2_dlygate4sd3_1
X_3261_ net515 VGND VPWR net8 DP_1.Q_range.out_data\[6\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2212_ _1493_ net451 net384 VPWR VGND sg13g2_nand2_1
X_3192_ net529 VGND VPWR net41 mac1.sum_lvl2_ff\[53\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2143_ _1422_ _1423_ _1425_ _1426_ VPWR VGND sg13g2_or3_1
XFILLER_38_157 VPWR VGND sg13g2_fill_2
XFILLER_47_680 VPWR VGND sg13g2_decap_8
X_2074_ _1360_ _1359_ _1347_ VPWR VGND sg13g2_nand2b_1
XFILLER_19_360 VPWR VGND sg13g2_decap_8
XFILLER_35_842 VPWR VGND sg13g2_fill_1
X_2976_ net470 _0096_ VPWR VGND sg13g2_buf_1
X_1927_ _1242_ mac1.sum_lvl2_ff\[25\] net296 VPWR VGND sg13g2_xnor2_1
X_1858_ _1183_ _1178_ _1181_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_39 VPWR VGND sg13g2_fill_1
X_1789_ _1101_ VPWR _1116_ VGND _1090_ _1102_ sg13g2_o21ai_1
XFILLER_39_48 VPWR VGND sg13g2_decap_8
XFILLER_29_179 VPWR VGND sg13g2_decap_4
XFILLER_38_691 VPWR VGND sg13g2_fill_2
XFILLER_41_878 VPWR VGND sg13g2_decap_8
XFILLER_21_580 VPWR VGND sg13g2_decap_8
XFILLER_5_713 VPWR VGND sg13g2_decap_8
XFILLER_20_50 VPWR VGND sg13g2_fill_2
XFILLER_20_61 VPWR VGND sg13g2_decap_8
XFILLER_4_278 VPWR VGND sg13g2_fill_2
XFILLER_0_440 VPWR VGND sg13g2_decap_8
XFILLER_49_923 VPWR VGND sg13g2_decap_8
XFILLER_1_996 VPWR VGND sg13g2_decap_8
Xhold81 mac1.products_ff\[14\] VPWR VGND net121 sg13g2_dlygate4sd3_1
Xhold92 mac1.sum_lvl1_ff\[84\] VPWR VGND net132 sg13g2_dlygate4sd3_1
Xhold70 mac1.products_ff\[150\] VPWR VGND net110 sg13g2_dlygate4sd3_1
XFILLER_17_820 VPWR VGND sg13g2_decap_8
XFILLER_17_886 VPWR VGND sg13g2_decap_8
X_2830_ _0722_ net477 DP_2.matrix\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_31_377 VPWR VGND sg13g2_fill_2
XFILLER_32_878 VPWR VGND sg13g2_decap_8
X_2761_ net482 net480 net424 net422 _0656_ VPWR VGND sg13g2_and4_1
X_2692_ _0589_ _0582_ _0588_ VPWR VGND sg13g2_xnor2_1
XFILLER_8_551 VPWR VGND sg13g2_decap_8
X_1712_ _0994_ _0997_ _1041_ VPWR VGND sg13g2_nor2_1
X_1643_ _0963_ _0971_ _0973_ _0974_ VPWR VGND sg13g2_or3_1
X_1574_ _0907_ _0905_ _0906_ VPWR VGND sg13g2_nand2_1
Xfanout508 net533 net508 VPWR VGND sg13g2_buf_8
Xfanout519 net533 net519 VPWR VGND sg13g2_buf_8
X_3244_ net503 VGND VPWR net202 net28 clknet_leaf_34_clk sg13g2_dfrbpq_2
X_3175_ net544 VGND VPWR net42 mac1.sum_lvl2_ff\[33\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_2126_ _1409_ _1401_ _1403_ VPWR VGND sg13g2_nand2_1
X_2057_ _1341_ _1342_ _1343_ _1344_ VPWR VGND sg13g2_nor3_1
XFILLER_19_190 VPWR VGND sg13g2_decap_8
XFILLER_22_333 VPWR VGND sg13g2_fill_2
XFILLER_23_845 VPWR VGND sg13g2_decap_8
X_2959_ _0836_ net429 net375 VPWR VGND sg13g2_nand2_1
XFILLER_2_727 VPWR VGND sg13g2_decap_8
XFILLER_46_904 VPWR VGND sg13g2_decap_8
XFILLER_26_683 VPWR VGND sg13g2_fill_1
XFILLER_14_856 VPWR VGND sg13g2_decap_8
XFILLER_41_686 VPWR VGND sg13g2_fill_1
XFILLER_13_377 VPWR VGND sg13g2_decap_8
XFILLER_40_185 VPWR VGND sg13g2_decap_8
XFILLER_9_348 VPWR VGND sg13g2_decap_8
XFILLER_12_1017 VPWR VGND sg13g2_decap_8
XFILLER_12_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_720 VPWR VGND sg13g2_decap_8
XFILLER_0_270 VPWR VGND sg13g2_decap_8
XFILLER_1_793 VPWR VGND sg13g2_decap_8
XFILLER_48_230 VPWR VGND sg13g2_decap_8
XFILLER_49_797 VPWR VGND sg13g2_decap_8
XFILLER_37_959 VPWR VGND sg13g2_decap_8
XFILLER_17_650 VPWR VGND sg13g2_decap_8
XFILLER_45_970 VPWR VGND sg13g2_decap_8
XFILLER_16_160 VPWR VGND sg13g2_decap_8
XFILLER_17_672 VPWR VGND sg13g2_decap_8
XFILLER_17_683 VPWR VGND sg13g2_fill_1
XFILLER_16_182 VPWR VGND sg13g2_fill_2
XFILLER_31_141 VPWR VGND sg13g2_decap_4
X_2813_ _0706_ net480 DP_2.matrix\[8\] VPWR VGND sg13g2_nand2_1
X_2744_ _0639_ _0617_ _0640_ VPWR VGND sg13g2_nor2b_1
XFILLER_9_893 VPWR VGND sg13g2_decap_8
X_2675_ _0573_ _0540_ _0572_ VPWR VGND sg13g2_nand2b_1
X_1626_ _0957_ net471 net405 VPWR VGND sg13g2_nand2_1
X_1557_ _0890_ net470 net408 VPWR VGND sg13g2_nand2_1
X_3227_ net509 VGND VPWR net256 mac1.sum_lvl3_ff\[2\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_3158_ net545 VGND VPWR net99 mac1.sum_lvl2_ff\[13\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_28_937 VPWR VGND sg13g2_decap_8
X_2109_ _1393_ net393 net447 net444 net398 VPWR VGND sg13g2_a22oi_1
XFILLER_43_929 VPWR VGND sg13g2_decap_8
X_3089_ net543 VGND VPWR _0078_ mac1.products_ff\[76\] clknet_leaf_25_clk sg13g2_dfrbpq_1
XFILLER_14_119 VPWR VGND sg13g2_decap_8
XFILLER_36_970 VPWR VGND sg13g2_decap_8
XFILLER_23_653 VPWR VGND sg13g2_decap_8
XFILLER_35_1006 VPWR VGND sg13g2_decap_8
XFILLER_23_686 VPWR VGND sg13g2_fill_2
XFILLER_7_819 VPWR VGND sg13g2_decap_8
XFILLER_19_915 VPWR VGND sg13g2_decap_8
XFILLER_18_414 VPWR VGND sg13g2_decap_8
XFILLER_18_469 VPWR VGND sg13g2_decap_8
XFILLER_27_981 VPWR VGND sg13g2_decap_8
XFILLER_45_288 VPWR VGND sg13g2_decap_8
XFILLER_42_951 VPWR VGND sg13g2_decap_8
XFILLER_14_664 VPWR VGND sg13g2_decap_8
XFILLER_9_112 VPWR VGND sg13g2_decap_8
XFILLER_6_874 VPWR VGND sg13g2_decap_8
X_2460_ _0351_ _0363_ _0364_ VPWR VGND sg13g2_nor2_1
X_2391_ _0300_ _0299_ _0296_ VPWR VGND sg13g2_nand2b_1
XFILLER_3_53 VPWR VGND sg13g2_decap_8
XFILLER_1_590 VPWR VGND sg13g2_decap_8
XFILLER_3_1004 VPWR VGND sg13g2_decap_8
X_3012_ net535 VGND VPWR _0065_ mac1.products_ff\[6\] clknet_leaf_29_clk sg13g2_dfrbpq_1
XFILLER_36_211 VPWR VGND sg13g2_decap_8
XFILLER_37_745 VPWR VGND sg13g2_decap_8
XFILLER_36_255 VPWR VGND sg13g2_decap_4
XFILLER_36_277 VPWR VGND sg13g2_decap_8
XFILLER_33_973 VPWR VGND sg13g2_decap_8
X_2727_ _0623_ _0595_ _0621_ VPWR VGND sg13g2_xnor2_1
X_2658_ VGND VPWR _0556_ _0555_ _0505_ sg13g2_or2_1
X_1609_ _0938_ _0939_ _0921_ _0941_ VPWR VGND sg13g2_nand3_1
X_2589_ VGND VPWR _0485_ _0486_ _0489_ _0444_ sg13g2_a21oi_1
XFILLER_27_233 VPWR VGND sg13g2_decap_4
XFILLER_28_745 VPWR VGND sg13g2_decap_8
XFILLER_28_756 VPWR VGND sg13g2_fill_1
XFILLER_43_715 VPWR VGND sg13g2_decap_8
XFILLER_16_918 VPWR VGND sg13g2_decap_8
XFILLER_42_214 VPWR VGND sg13g2_fill_2
XFILLER_6_148 VPWR VGND sg13g2_decap_8
XFILLER_3_822 VPWR VGND sg13g2_decap_8
XFILLER_3_899 VPWR VGND sg13g2_decap_8
XFILLER_19_723 VPWR VGND sg13g2_fill_2
XFILLER_46_520 VPWR VGND sg13g2_fill_2
XFILLER_46_586 VPWR VGND sg13g2_fill_2
XFILLER_18_277 VPWR VGND sg13g2_decap_8
XFILLER_19_789 VPWR VGND sg13g2_fill_2
XFILLER_34_748 VPWR VGND sg13g2_decap_8
XFILLER_15_984 VPWR VGND sg13g2_decap_8
X_1960_ _1263_ _1260_ _1269_ VPWR VGND _1262_ sg13g2_nand3b_1
X_1891_ _1214_ _1201_ _1215_ VPWR VGND sg13g2_xor2_1
XFILLER_30_976 VPWR VGND sg13g2_decap_8
XFILLER_6_671 VPWR VGND sg13g2_decap_8
X_2512_ _0408_ _0409_ _0413_ VPWR VGND _0383_ sg13g2_nand3b_1
XFILLER_5_181 VPWR VGND sg13g2_fill_2
X_2443_ _0345_ _0346_ _0347_ _0348_ VPWR VGND sg13g2_nor3_1
X_2374_ _0283_ _0282_ _0284_ VPWR VGND sg13g2_nor2b_1
XFILLER_37_575 VPWR VGND sg13g2_decap_8
XFILLER_25_759 VPWR VGND sg13g2_decap_4
XFILLER_37_586 VPWR VGND sg13g2_fill_2
XFILLER_12_409 VPWR VGND sg13g2_fill_1
XFILLER_21_910 VPWR VGND sg13g2_decap_8
XFILLER_20_453 VPWR VGND sg13g2_decap_8
XFILLER_20_464 VPWR VGND sg13g2_fill_1
XFILLER_21_987 VPWR VGND sg13g2_decap_8
XFILLER_0_825 VPWR VGND sg13g2_decap_8
XFILLER_48_807 VPWR VGND sg13g2_decap_8
XFILLER_31_707 VPWR VGND sg13g2_decap_8
XFILLER_24_781 VPWR VGND sg13g2_decap_8
XFILLER_8_914 VPWR VGND sg13g2_decap_8
XFILLER_12_954 VPWR VGND sg13g2_decap_8
XFILLER_23_291 VPWR VGND sg13g2_decap_8
XFILLER_11_453 VPWR VGND sg13g2_decap_8
XFILLER_23_50 VPWR VGND sg13g2_fill_2
XFILLER_3_696 VPWR VGND sg13g2_decap_8
X_2090_ _1372_ _1371_ _1366_ _1375_ VPWR VGND sg13g2_a21o_1
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_0_1007 VPWR VGND sg13g2_decap_8
XFILLER_19_553 VPWR VGND sg13g2_decap_8
XFILLER_19_597 VPWR VGND sg13g2_decap_8
XFILLER_0_98 VPWR VGND sg13g2_decap_8
X_2992_ net410 _0120_ VPWR VGND sg13g2_buf_1
XFILLER_9_41 VPWR VGND sg13g2_decap_4
X_1943_ _1255_ mac1.sum_lvl2_ff\[28\] mac1.sum_lvl2_ff\[9\] VPWR VGND sg13g2_nand2_1
XFILLER_9_85 VPWR VGND sg13g2_fill_1
X_1874_ _1198_ _1170_ _1193_ VPWR VGND sg13g2_nand2_1
XFILLER_31_1020 VPWR VGND sg13g2_decap_8
XFILLER_7_980 VPWR VGND sg13g2_decap_8
X_2426_ _0332_ _0319_ _0334_ VPWR VGND sg13g2_xor2_1
XFILLER_29_306 VPWR VGND sg13g2_decap_8
X_2357_ VGND VPWR _0267_ _0266_ _0215_ sg13g2_or2_1
X_2288_ _0189_ VPWR _0200_ VGND _0173_ _0190_ sg13g2_o21ai_1
XFILLER_21_784 VPWR VGND sg13g2_decap_8
XFILLER_0_622 VPWR VGND sg13g2_decap_8
XFILLER_47_103 VPWR VGND sg13g2_decap_8
XFILLER_0_699 VPWR VGND sg13g2_decap_8
XFILLER_48_648 VPWR VGND sg13g2_fill_1
XFILLER_29_840 VPWR VGND sg13g2_decap_8
XFILLER_47_147 VPWR VGND sg13g2_fill_1
XFILLER_18_72 VPWR VGND sg13g2_fill_2
XFILLER_43_353 VPWR VGND sg13g2_fill_1
XFILLER_16_545 VPWR VGND sg13g2_fill_2
XFILLER_28_394 VPWR VGND sg13g2_fill_1
XFILLER_44_887 VPWR VGND sg13g2_decap_8
XFILLER_43_364 VPWR VGND sg13g2_decap_4
XFILLER_43_397 VPWR VGND sg13g2_fill_2
XFILLER_8_711 VPWR VGND sg13g2_decap_8
XFILLER_15_1026 VPWR VGND sg13g2_fill_2
XFILLER_8_788 VPWR VGND sg13g2_decap_8
XFILLER_7_243 VPWR VGND sg13g2_decap_4
X_1590_ _0922_ net473 net405 VPWR VGND sg13g2_nand2_1
XFILLER_4_994 VPWR VGND sg13g2_decap_8
X_3260_ net515 VGND VPWR DP_1.Q_range.data_plus_4\[6\] DP_1.Q_range.out_data\[5\]
+ clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2211_ _1464_ VPWR _1492_ VGND _1455_ _1465_ sg13g2_o21ai_1
X_3191_ net530 VGND VPWR net80 mac1.sum_lvl2_ff\[52\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_22_1008 VPWR VGND sg13g2_decap_8
X_2142_ _1425_ net394 net444 net442 net399 VPWR VGND sg13g2_a22oi_1
X_2073_ _1358_ _1348_ _1359_ VPWR VGND sg13g2_xor2_1
XFILLER_35_887 VPWR VGND sg13g2_decap_8
X_2975_ net472 _0095_ VPWR VGND sg13g2_buf_1
X_1926_ mac1.sum_lvl2_ff\[25\] mac1.sum_lvl2_ff\[6\] _1241_ VPWR VGND sg13g2_and2_1
X_1857_ _1182_ _1181_ _1178_ VPWR VGND sg13g2_nand2b_1
XFILLER_30_18 VPWR VGND sg13g2_decap_8
XFILLER_2_909 VPWR VGND sg13g2_decap_8
X_1788_ _1087_ _1081_ _1089_ _1115_ VPWR VGND sg13g2_a21o_1
X_2409_ _0317_ _0311_ _0316_ VPWR VGND sg13g2_nand2_1
XFILLER_45_618 VPWR VGND sg13g2_decap_8
XFILLER_38_670 VPWR VGND sg13g2_decap_8
XFILLER_38_1015 VPWR VGND sg13g2_decap_8
XFILLER_40_323 VPWR VGND sg13g2_decap_4
XFILLER_40_367 VPWR VGND sg13g2_decap_8
XFILLER_9_519 VPWR VGND sg13g2_decap_8
XFILLER_5_769 VPWR VGND sg13g2_decap_8
XFILLER_4_246 VPWR VGND sg13g2_decap_8
XFILLER_45_1019 VPWR VGND sg13g2_decap_8
XFILLER_49_902 VPWR VGND sg13g2_decap_8
XFILLER_1_975 VPWR VGND sg13g2_decap_8
XFILLER_0_496 VPWR VGND sg13g2_decap_8
XFILLER_49_979 VPWR VGND sg13g2_decap_8
Xhold60 mac1.sum_lvl1_ff\[7\] VPWR VGND net100 sg13g2_dlygate4sd3_1
Xhold71 mac1.sum_lvl2_ff\[43\] VPWR VGND net111 sg13g2_dlygate4sd3_1
Xhold82 mac1.sum_lvl1_ff\[42\] VPWR VGND net122 sg13g2_dlygate4sd3_1
XFILLER_36_618 VPWR VGND sg13g2_decap_8
XFILLER_48_489 VPWR VGND sg13g2_decap_4
Xhold93 mac1.products_ff\[3\] VPWR VGND net133 sg13g2_dlygate4sd3_1
XFILLER_44_640 VPWR VGND sg13g2_decap_8
XFILLER_17_865 VPWR VGND sg13g2_decap_8
XFILLER_45_81 VPWR VGND sg13g2_decap_8
XFILLER_44_695 VPWR VGND sg13g2_decap_8
XFILLER_31_312 VPWR VGND sg13g2_fill_1
XFILLER_32_857 VPWR VGND sg13g2_decap_8
X_2760_ _0655_ net480 net422 VPWR VGND sg13g2_nand2_1
XFILLER_40_890 VPWR VGND sg13g2_decap_8
X_2691_ _0587_ _0583_ _0588_ VPWR VGND sg13g2_xor2_1
X_1711_ _1022_ VPWR _1040_ VGND _1001_ _1023_ sg13g2_o21ai_1
X_1642_ VGND VPWR _0969_ _0970_ _0973_ _0964_ sg13g2_a21oi_1
X_1573_ _0894_ VPWR _0906_ VGND _0902_ _0904_ sg13g2_o21ai_1
Xfanout509 net513 net509 VPWR VGND sg13g2_buf_8
XFILLER_4_791 VPWR VGND sg13g2_decap_8
X_3243_ net503 VGND VPWR net176 net27 clknet_leaf_35_clk sg13g2_dfrbpq_2
X_3174_ net540 VGND VPWR net59 mac1.sum_lvl2_ff\[32\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_2125_ _0047_ _1381_ _1408_ VPWR VGND sg13g2_xnor2_1
X_2056_ _1343_ net392 net454 net452 net397 VPWR VGND sg13g2_a22oi_1
XFILLER_22_301 VPWR VGND sg13g2_decap_4
XFILLER_41_39 VPWR VGND sg13g2_decap_4
X_2958_ _0800_ _0790_ _0835_ VPWR VGND sg13g2_xor2_1
X_1909_ _0007_ _1225_ _1228_ VPWR VGND sg13g2_xnor2_1
X_2889_ DP_2.Q_range.out_data\[2\] _0842_ DP_2.Q_range.out_data\[4\] DP_2.Q_range.out_data\[6\]
+ _0778_ VPWR VGND sg13g2_nor4_1
XFILLER_2_706 VPWR VGND sg13g2_decap_8
Xheichips25_template_40 VPWR VGND uio_oe[7] sg13g2_tiehi
XFILLER_45_437 VPWR VGND sg13g2_decap_8
XFILLER_26_662 VPWR VGND sg13g2_decap_8
XFILLER_14_835 VPWR VGND sg13g2_decap_8
XFILLER_26_695 VPWR VGND sg13g2_decap_8
XFILLER_13_356 VPWR VGND sg13g2_decap_8
XFILLER_15_84 VPWR VGND sg13g2_decap_8
XFILLER_40_164 VPWR VGND sg13g2_decap_8
XFILLER_9_327 VPWR VGND sg13g2_decap_8
XFILLER_15_95 VPWR VGND sg13g2_fill_1
XFILLER_40_197 VPWR VGND sg13g2_fill_2
XFILLER_5_500 VPWR VGND sg13g2_fill_2
XFILLER_1_772 VPWR VGND sg13g2_decap_8
XFILLER_49_776 VPWR VGND sg13g2_decap_8
XFILLER_48_286 VPWR VGND sg13g2_decap_8
XFILLER_37_938 VPWR VGND sg13g2_decap_8
XFILLER_48_297 VPWR VGND sg13g2_fill_2
XFILLER_31_120 VPWR VGND sg13g2_decap_8
X_2812_ _0684_ VPWR _0705_ VGND _0655_ _0682_ sg13g2_o21ai_1
XFILLER_13_890 VPWR VGND sg13g2_decap_8
X_2743_ _0639_ _0618_ _0638_ VPWR VGND sg13g2_xnor2_1
XFILLER_9_872 VPWR VGND sg13g2_decap_8
XFILLER_8_393 VPWR VGND sg13g2_fill_1
X_2674_ _0572_ _0541_ _0570_ VPWR VGND sg13g2_xnor2_1
X_1625_ _0937_ _0927_ _0935_ _0956_ VPWR VGND sg13g2_a21o_1
X_1556_ _0889_ net471 net406 VPWR VGND sg13g2_nand2_1
XFILLER_28_1014 VPWR VGND sg13g2_decap_8
X_3226_ net509 VGND VPWR net236 mac1.sum_lvl3_ff\[1\] clknet_leaf_36_clk sg13g2_dfrbpq_2
XFILLER_28_916 VPWR VGND sg13g2_decap_8
X_3157_ net545 VGND VPWR net97 mac1.sum_lvl2_ff\[12\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_43_908 VPWR VGND sg13g2_decap_8
X_2108_ net447 net444 net398 _1392_ VPWR VGND net393 sg13g2_nand4_1
X_3088_ net536 VGND VPWR _0077_ mac1.products_ff\[75\] clknet_leaf_29_clk sg13g2_dfrbpq_1
X_2039_ VGND VPWR _1323_ _1328_ _1331_ net232 sg13g2_a21oi_1
XFILLER_23_610 VPWR VGND sg13g2_decap_8
XFILLER_10_326 VPWR VGND sg13g2_fill_1
XFILLER_11_849 VPWR VGND sg13g2_decap_8
XFILLER_2_514 VPWR VGND sg13g2_decap_8
XFILLER_46_713 VPWR VGND sg13g2_fill_2
XFILLER_45_201 VPWR VGND sg13g2_fill_1
XFILLER_45_267 VPWR VGND sg13g2_decap_8
XFILLER_27_960 VPWR VGND sg13g2_decap_8
XFILLER_34_919 VPWR VGND sg13g2_decap_8
XFILLER_42_930 VPWR VGND sg13g2_decap_8
XFILLER_26_470 VPWR VGND sg13g2_decap_4
XFILLER_41_440 VPWR VGND sg13g2_fill_1
XFILLER_13_120 VPWR VGND sg13g2_decap_8
XFILLER_13_131 VPWR VGND sg13g2_fill_2
XFILLER_6_853 VPWR VGND sg13g2_decap_8
X_2390_ _0298_ _0272_ _0299_ VPWR VGND sg13g2_xor2_1
XFILLER_3_32 VPWR VGND sg13g2_decap_4
XFILLER_3_98 VPWR VGND sg13g2_fill_1
XFILLER_49_573 VPWR VGND sg13g2_decap_8
X_3011_ net534 VGND VPWR _0058_ mac1.products_ff\[5\] clknet_leaf_28_clk sg13g2_dfrbpq_1
XFILLER_37_702 VPWR VGND sg13g2_decap_8
XFILLER_37_724 VPWR VGND sg13g2_decap_8
XFILLER_17_470 VPWR VGND sg13g2_decap_8
XFILLER_18_993 VPWR VGND sg13g2_decap_8
XFILLER_33_952 VPWR VGND sg13g2_decap_8
XFILLER_9_680 VPWR VGND sg13g2_decap_8
X_2726_ VGND VPWR _0622_ _0621_ _0595_ sg13g2_or2_1
X_2657_ _0555_ net479 net430 VPWR VGND sg13g2_nand2_1
X_1608_ _0940_ _0921_ _0938_ _0939_ VPWR VGND sg13g2_and3_1
X_2588_ _0485_ _0486_ _0444_ _0488_ VPWR VGND sg13g2_nand3_1
X_1539_ net413 net468 net418 _0873_ VPWR VGND net466 sg13g2_nand4_1
XFILLER_41_1011 VPWR VGND sg13g2_decap_8
XFILLER_47_49 VPWR VGND sg13g2_decap_4
X_3209_ net505 VGND VPWR net50 mac1.sum_lvl3_ff\[20\] clknet_leaf_37_clk sg13g2_dfrbpq_1
XFILLER_28_724 VPWR VGND sg13g2_decap_8
XFILLER_42_237 VPWR VGND sg13g2_decap_8
XFILLER_24_985 VPWR VGND sg13g2_decap_8
XFILLER_11_646 VPWR VGND sg13g2_decap_8
XFILLER_10_145 VPWR VGND sg13g2_decap_4
XFILLER_6_116 VPWR VGND sg13g2_decap_8
XFILLER_3_801 VPWR VGND sg13g2_decap_8
XFILLER_12_85 VPWR VGND sg13g2_decap_8
XFILLER_3_878 VPWR VGND sg13g2_decap_8
Xhold190 _0113_ VPWR VGND net230 sg13g2_dlygate4sd3_1
XFILLER_46_543 VPWR VGND sg13g2_decap_8
XFILLER_46_554 VPWR VGND sg13g2_fill_2
XFILLER_18_267 VPWR VGND sg13g2_fill_1
XFILLER_19_768 VPWR VGND sg13g2_decap_8
XFILLER_34_727 VPWR VGND sg13g2_decap_8
XFILLER_14_440 VPWR VGND sg13g2_decap_8
XFILLER_15_963 VPWR VGND sg13g2_decap_8
XFILLER_42_760 VPWR VGND sg13g2_fill_1
XFILLER_14_473 VPWR VGND sg13g2_fill_2
XFILLER_41_281 VPWR VGND sg13g2_decap_8
XFILLER_14_495 VPWR VGND sg13g2_decap_8
XFILLER_30_955 VPWR VGND sg13g2_decap_8
X_1890_ _1212_ _1202_ _1214_ VPWR VGND sg13g2_xor2_1
XFILLER_6_650 VPWR VGND sg13g2_decap_8
X_2511_ _0385_ _0410_ _0412_ VPWR VGND sg13g2_nor2b_1
X_2442_ _0347_ net433 net490 net488 net437 VPWR VGND sg13g2_a22oi_1
X_2373_ VGND VPWR _0237_ _0242_ _0283_ _0254_ sg13g2_a21oi_1
XFILLER_37_532 VPWR VGND sg13g2_decap_8
XFILLER_37_543 VPWR VGND sg13g2_fill_1
XFILLER_25_738 VPWR VGND sg13g2_decap_8
XFILLER_24_237 VPWR VGND sg13g2_decap_4
XFILLER_33_18 VPWR VGND sg13g2_decap_8
XFILLER_21_966 VPWR VGND sg13g2_decap_8
X_2709_ _0604_ _0580_ _0606_ VPWR VGND sg13g2_xor2_1
XFILLER_0_804 VPWR VGND sg13g2_decap_8
XFILLER_28_532 VPWR VGND sg13g2_decap_8
XFILLER_28_543 VPWR VGND sg13g2_fill_2
XFILLER_28_565 VPWR VGND sg13g2_decap_8
XFILLER_43_546 VPWR VGND sg13g2_decap_4
XFILLER_15_259 VPWR VGND sg13g2_decap_8
XFILLER_30_218 VPWR VGND sg13g2_decap_8
XFILLER_12_933 VPWR VGND sg13g2_decap_8
XFILLER_30_229 VPWR VGND sg13g2_fill_2
XFILLER_7_425 VPWR VGND sg13g2_decap_4
XFILLER_11_476 VPWR VGND sg13g2_fill_1
XFILLER_48_1017 VPWR VGND sg13g2_decap_8
XFILLER_48_1028 VPWR VGND sg13g2_fill_1
XFILLER_3_675 VPWR VGND sg13g2_decap_8
XFILLER_2_141 VPWR VGND sg13g2_fill_2
XFILLER_2_163 VPWR VGND sg13g2_decap_4
XFILLER_17_7 VPWR VGND sg13g2_decap_4
XFILLER_19_532 VPWR VGND sg13g2_decap_8
XFILLER_46_351 VPWR VGND sg13g2_fill_1
XFILLER_47_885 VPWR VGND sg13g2_decap_8
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_34_524 VPWR VGND sg13g2_decap_8
XFILLER_34_535 VPWR VGND sg13g2_fill_1
XFILLER_34_568 VPWR VGND sg13g2_fill_1
X_2991_ net412 _0119_ VPWR VGND sg13g2_buf_1
X_1942_ _1250_ _1252_ _1254_ VPWR VGND sg13g2_nor2_1
X_1873_ VPWR VGND _1142_ _1196_ _1174_ _1111_ _1197_ _1173_ sg13g2_a221oi_1
XFILLER_43_0 VPWR VGND sg13g2_fill_2
X_2425_ _0319_ _0332_ _0333_ VPWR VGND sg13g2_nor2_1
X_2356_ _0266_ net496 net385 VPWR VGND sg13g2_nand2_2
X_2287_ VGND VPWR _0164_ _0170_ _0199_ _0172_ sg13g2_a21oi_1
XFILLER_29_329 VPWR VGND sg13g2_decap_8
XFILLER_25_524 VPWR VGND sg13g2_decap_8
XFILLER_38_896 VPWR VGND sg13g2_decap_8
XFILLER_37_395 VPWR VGND sg13g2_fill_1
XFILLER_12_229 VPWR VGND sg13g2_fill_2
XFILLER_21_763 VPWR VGND sg13g2_fill_1
Xclkbuf_3_0__f_clk clknet_0_clk clknet_3_0__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_4_428 VPWR VGND sg13g2_decap_8
XFILLER_0_601 VPWR VGND sg13g2_decap_8
XFILLER_0_678 VPWR VGND sg13g2_decap_8
XFILLER_18_51 VPWR VGND sg13g2_decap_8
XFILLER_43_310 VPWR VGND sg13g2_decap_4
XFILLER_16_513 VPWR VGND sg13g2_decap_4
XFILLER_16_524 VPWR VGND sg13g2_decap_8
XFILLER_28_373 VPWR VGND sg13g2_decap_8
XFILLER_29_885 VPWR VGND sg13g2_decap_8
XFILLER_44_866 VPWR VGND sg13g2_decap_8
XFILLER_43_376 VPWR VGND sg13g2_decap_8
XFILLER_12_763 VPWR VGND sg13g2_decap_8
XFILLER_15_1005 VPWR VGND sg13g2_decap_8
XFILLER_34_94 VPWR VGND sg13g2_decap_4
XFILLER_11_262 VPWR VGND sg13g2_decap_8
XFILLER_8_767 VPWR VGND sg13g2_decap_8
XFILLER_4_973 VPWR VGND sg13g2_decap_8
XFILLER_3_472 VPWR VGND sg13g2_decap_8
XFILLER_3_494 VPWR VGND sg13g2_decap_8
XFILLER_3_483 VPWR VGND sg13g2_fill_2
X_2210_ _1491_ _1444_ _1490_ VPWR VGND sg13g2_xnor2_1
XFILLER_39_616 VPWR VGND sg13g2_decap_8
X_3190_ net530 VGND VPWR net83 mac1.sum_lvl2_ff\[51\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_39_649 VPWR VGND sg13g2_fill_2
XFILLER_15_4 VPWR VGND sg13g2_decap_8
X_2141_ net444 net442 net399 _1424_ VPWR VGND net394 sg13g2_nand4_1
X_2072_ _1358_ _1349_ _1356_ VPWR VGND sg13g2_xnor2_1
XFILLER_35_833 VPWR VGND sg13g2_decap_8
XFILLER_46_170 VPWR VGND sg13g2_decap_4
XFILLER_34_343 VPWR VGND sg13g2_decap_8
XFILLER_35_866 VPWR VGND sg13g2_decap_8
X_2974_ net474 _0094_ VPWR VGND sg13g2_buf_1
XFILLER_22_527 VPWR VGND sg13g2_decap_8
XFILLER_22_549 VPWR VGND sg13g2_decap_8
X_1925_ _0011_ _1238_ net258 VPWR VGND sg13g2_xnor2_1
X_1856_ _1180_ _1153_ _1181_ VPWR VGND sg13g2_xor2_1
X_1787_ _1113_ _1110_ _0070_ VPWR VGND sg13g2_xor2_1
X_2408_ _0316_ _0289_ _0312_ VPWR VGND sg13g2_nand2_1
X_2339_ _0249_ _0246_ _0250_ VPWR VGND sg13g2_xor2_1
XFILLER_29_137 VPWR VGND sg13g2_fill_1
XFILLER_25_343 VPWR VGND sg13g2_fill_2
XFILLER_26_855 VPWR VGND sg13g2_decap_4
XFILLER_26_888 VPWR VGND sg13g2_decap_8
XFILLER_41_836 VPWR VGND sg13g2_fill_1
XFILLER_13_527 VPWR VGND sg13g2_decap_8
XFILLER_13_538 VPWR VGND sg13g2_fill_2
XFILLER_25_398 VPWR VGND sg13g2_decap_8
XFILLER_5_748 VPWR VGND sg13g2_decap_8
XFILLER_1_954 VPWR VGND sg13g2_decap_8
XFILLER_49_958 VPWR VGND sg13g2_decap_8
XFILLER_0_475 VPWR VGND sg13g2_decap_8
Xhold50 mac1.sum_lvl2_ff\[50\] VPWR VGND net90 sg13g2_dlygate4sd3_1
XFILLER_48_468 VPWR VGND sg13g2_decap_8
Xhold83 mac1.products_ff\[1\] VPWR VGND net123 sg13g2_dlygate4sd3_1
Xhold61 mac1.sum_lvl1_ff\[5\] VPWR VGND net101 sg13g2_dlygate4sd3_1
Xhold72 mac1.sum_lvl1_ff\[80\] VPWR VGND net112 sg13g2_dlygate4sd3_1
XFILLER_29_72 VPWR VGND sg13g2_decap_8
Xhold94 mac1.sum_lvl1_ff\[77\] VPWR VGND net134 sg13g2_dlygate4sd3_1
XFILLER_35_129 VPWR VGND sg13g2_decap_8
XFILLER_16_310 VPWR VGND sg13g2_decap_8
XFILLER_16_321 VPWR VGND sg13g2_decap_8
XFILLER_16_332 VPWR VGND sg13g2_fill_2
XFILLER_45_60 VPWR VGND sg13g2_fill_1
XFILLER_44_674 VPWR VGND sg13g2_fill_1
XFILLER_16_376 VPWR VGND sg13g2_decap_8
XFILLER_43_162 VPWR VGND sg13g2_decap_8
XFILLER_31_379 VPWR VGND sg13g2_fill_1
X_2690_ _0587_ _0545_ _0585_ VPWR VGND sg13g2_xnor2_1
X_1710_ _0999_ VPWR _1039_ VGND _0952_ _1000_ sg13g2_o21ai_1
XFILLER_6_43 VPWR VGND sg13g2_fill_1
X_1641_ _0969_ _0970_ _0964_ _0972_ VPWR VGND sg13g2_nand3_1
XFILLER_4_770 VPWR VGND sg13g2_decap_8
X_1572_ _0894_ _0902_ _0904_ _0905_ VPWR VGND sg13g2_or3_1
X_3242_ net503 VGND VPWR net167 net26 clknet_leaf_37_clk sg13g2_dfrbpq_1
XFILLER_39_435 VPWR VGND sg13g2_fill_2
XFILLER_39_424 VPWR VGND sg13g2_decap_8
XFILLER_6_1014 VPWR VGND sg13g2_decap_8
X_3173_ net541 VGND VPWR net52 mac1.sum_lvl2_ff\[31\] clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_39_468 VPWR VGND sg13g2_fill_2
XFILLER_39_457 VPWR VGND sg13g2_decap_4
X_2124_ _1405_ _1379_ _1408_ VPWR VGND sg13g2_xor2_1
X_2055_ net397 net454 net452 net392 _1342_ VPWR VGND sg13g2_and4_1
XFILLER_23_825 VPWR VGND sg13g2_decap_8
XFILLER_22_357 VPWR VGND sg13g2_fill_2
XFILLER_41_18 VPWR VGND sg13g2_decap_8
X_2957_ _0834_ VPWR _0112_ VGND net374 _0833_ sg13g2_o21ai_1
XFILLER_31_880 VPWR VGND sg13g2_decap_8
X_2888_ _0081_ _0775_ _0777_ _0774_ _0765_ VPWR VGND sg13g2_a22oi_1
X_1908_ mac1.sum_lvl2_ff\[1\] mac1.sum_lvl2_ff\[20\] _1228_ VPWR VGND sg13g2_xor2_1
X_1839_ _1164_ _1163_ _1165_ VPWR VGND sg13g2_nor2b_1
XFILLER_1_239 VPWR VGND sg13g2_fill_1
XFILLER_44_1020 VPWR VGND sg13g2_decap_8
XFILLER_46_939 VPWR VGND sg13g2_decap_8
XFILLER_45_416 VPWR VGND sg13g2_decap_8
XFILLER_17_107 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_37_clk clknet_3_0__leaf_clk clknet_leaf_37_clk VPWR VGND sg13g2_buf_8
XFILLER_26_641 VPWR VGND sg13g2_decap_8
XFILLER_14_803 VPWR VGND sg13g2_decap_8
XFILLER_41_633 VPWR VGND sg13g2_decap_8
XFILLER_25_162 VPWR VGND sg13g2_decap_8
XFILLER_25_173 VPWR VGND sg13g2_fill_2
XFILLER_41_677 VPWR VGND sg13g2_decap_8
XFILLER_41_644 VPWR VGND sg13g2_fill_1
XFILLER_13_335 VPWR VGND sg13g2_decap_8
XFILLER_41_699 VPWR VGND sg13g2_decap_8
XFILLER_40_154 VPWR VGND sg13g2_decap_4
XFILLER_5_545 VPWR VGND sg13g2_decap_8
XFILLER_1_751 VPWR VGND sg13g2_decap_8
XFILLER_49_755 VPWR VGND sg13g2_decap_8
XFILLER_37_917 VPWR VGND sg13g2_decap_8
XFILLER_48_265 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_28_clk clknet_3_4__leaf_clk clknet_leaf_28_clk VPWR VGND sg13g2_buf_8
XFILLER_17_696 VPWR VGND sg13g2_decap_8
X_2811_ _0687_ _0679_ _0686_ _0704_ VPWR VGND sg13g2_a21o_1
X_2742_ _0638_ _0627_ _0637_ VPWR VGND sg13g2_xnor2_1
XFILLER_9_851 VPWR VGND sg13g2_decap_8
XFILLER_8_372 VPWR VGND sg13g2_decap_8
X_2673_ _0571_ _0541_ _0570_ VPWR VGND sg13g2_nand2_1
X_1624_ _0955_ _0950_ _0953_ VPWR VGND sg13g2_xnor2_1
X_1555_ _0888_ net475 net405 VPWR VGND sg13g2_nand2_1
X_3225_ net505 VGND VPWR net162 mac1.sum_lvl3_ff\[0\] clknet_leaf_37_clk sg13g2_dfrbpq_1
XFILLER_27_416 VPWR VGND sg13g2_decap_8
X_3156_ net544 VGND VPWR net72 mac1.sum_lvl2_ff\[11\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_3087_ net534 VGND VPWR _0076_ mac1.products_ff\[74\] clknet_leaf_26_clk sg13g2_dfrbpq_1
X_2107_ net398 net447 net444 net393 _1391_ VPWR VGND sg13g2_and4_1
Xclkbuf_leaf_19_clk clknet_3_7__leaf_clk clknet_leaf_19_clk VPWR VGND sg13g2_buf_8
XFILLER_36_29 VPWR VGND sg13g2_decap_8
X_2038_ _1330_ mac1.sum_lvl3_ff\[13\] net231 VPWR VGND sg13g2_xnor2_1
XFILLER_35_460 VPWR VGND sg13g2_decap_8
XFILLER_35_482 VPWR VGND sg13g2_decap_8
XFILLER_11_828 VPWR VGND sg13g2_decap_8
XFILLER_22_154 VPWR VGND sg13g2_fill_2
XFILLER_2_537 VPWR VGND sg13g2_decap_8
XFILLER_46_769 VPWR VGND sg13g2_fill_2
XFILLER_46_758 VPWR VGND sg13g2_decap_8
XFILLER_45_246 VPWR VGND sg13g2_decap_8
XFILLER_33_408 VPWR VGND sg13g2_decap_8
XFILLER_14_622 VPWR VGND sg13g2_decap_8
XFILLER_26_84 VPWR VGND sg13g2_decap_4
XFILLER_26_95 VPWR VGND sg13g2_decap_8
XFILLER_42_986 VPWR VGND sg13g2_decap_8
XFILLER_41_485 VPWR VGND sg13g2_fill_1
XFILLER_41_474 VPWR VGND sg13g2_fill_2
XFILLER_42_50 VPWR VGND sg13g2_fill_2
XFILLER_13_187 VPWR VGND sg13g2_decap_8
XFILLER_42_94 VPWR VGND sg13g2_decap_8
XFILLER_10_894 VPWR VGND sg13g2_decap_8
XFILLER_6_832 VPWR VGND sg13g2_decap_8
XFILLER_47_7 VPWR VGND sg13g2_decap_8
XFILLER_3_11 VPWR VGND sg13g2_decap_8
XFILLER_49_541 VPWR VGND sg13g2_decap_8
XFILLER_49_585 VPWR VGND sg13g2_decap_8
XFILLER_49_552 VPWR VGND sg13g2_fill_2
X_3010_ net526 VGND VPWR _0041_ mac1.products_ff\[4\] clknet_leaf_28_clk sg13g2_dfrbpq_1
XFILLER_18_972 VPWR VGND sg13g2_decap_8
XFILLER_33_931 VPWR VGND sg13g2_decap_8
XFILLER_17_493 VPWR VGND sg13g2_fill_1
X_2725_ _0621_ net500 net430 VPWR VGND sg13g2_nand2_1
X_2656_ _0554_ net484 net426 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_8_clk clknet_3_2__leaf_clk clknet_leaf_8_clk VPWR VGND sg13g2_buf_8
X_1607_ _0937_ _0936_ _0927_ _0939_ VPWR VGND sg13g2_a21o_1
X_2587_ _0487_ _0444_ _0485_ _0486_ VPWR VGND sg13g2_and3_1
X_1538_ net417 net412 net468 net466 _0872_ VPWR VGND sg13g2_and4_1
XFILLER_47_28 VPWR VGND sg13g2_decap_8
X_3208_ net529 VGND VPWR net51 mac1.sum_lvl1_ff\[87\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_3139_ net542 VGND VPWR net82 mac1.sum_lvl1_ff\[46\] clknet_leaf_23_clk sg13g2_dfrbpq_1
XFILLER_15_408 VPWR VGND sg13g2_fill_2
XFILLER_24_964 VPWR VGND sg13g2_decap_8
XFILLER_11_625 VPWR VGND sg13g2_decap_8
XFILLER_23_485 VPWR VGND sg13g2_decap_8
XFILLER_10_135 VPWR VGND sg13g2_fill_1
XFILLER_12_64 VPWR VGND sg13g2_decap_8
XFILLER_12_97 VPWR VGND sg13g2_decap_8
XFILLER_3_857 VPWR VGND sg13g2_decap_8
Xhold180 DP_1.matrix\[75\] VPWR VGND net220 sg13g2_dlygate4sd3_1
XFILLER_2_378 VPWR VGND sg13g2_decap_8
Xhold191 mac1.sum_lvl3_ff\[33\] VPWR VGND net231 sg13g2_dlygate4sd3_1
XFILLER_19_714 VPWR VGND sg13g2_fill_1
XFILLER_19_736 VPWR VGND sg13g2_fill_1
XFILLER_19_747 VPWR VGND sg13g2_decap_8
XFILLER_34_717 VPWR VGND sg13g2_fill_2
XFILLER_46_588 VPWR VGND sg13g2_fill_1
XFILLER_33_216 VPWR VGND sg13g2_decap_8
XFILLER_15_942 VPWR VGND sg13g2_decap_8
XFILLER_41_260 VPWR VGND sg13g2_decap_8
XFILLER_18_1014 VPWR VGND sg13g2_decap_8
XFILLER_30_934 VPWR VGND sg13g2_decap_8
X_2510_ _0411_ _0410_ _0058_ VPWR VGND sg13g2_xor2_1
X_2441_ net437 net490 net488 net433 _0346_ VPWR VGND sg13g2_and4_1
XFILLER_45_4 VPWR VGND sg13g2_decap_4
XFILLER_5_183 VPWR VGND sg13g2_fill_1
X_2372_ _0280_ _0268_ _0282_ VPWR VGND sg13g2_xor2_1
XFILLER_25_1018 VPWR VGND sg13g2_decap_8
XFILLER_25_717 VPWR VGND sg13g2_decap_8
XFILLER_24_205 VPWR VGND sg13g2_decap_4
XFILLER_21_945 VPWR VGND sg13g2_decap_8
XFILLER_33_794 VPWR VGND sg13g2_fill_1
X_2708_ _0605_ _0580_ _0604_ VPWR VGND sg13g2_nand2_1
X_2639_ _0536_ _0535_ _0067_ VPWR VGND sg13g2_xor2_1
XFILLER_28_500 VPWR VGND sg13g2_decap_8
XFILLER_43_525 VPWR VGND sg13g2_decap_8
XFILLER_15_205 VPWR VGND sg13g2_decap_4
XFILLER_15_238 VPWR VGND sg13g2_decap_8
XFILLER_12_912 VPWR VGND sg13g2_decap_8
XFILLER_23_260 VPWR VGND sg13g2_decap_4
XFILLER_12_989 VPWR VGND sg13g2_decap_8
XFILLER_8_949 VPWR VGND sg13g2_decap_8
XFILLER_3_654 VPWR VGND sg13g2_decap_8
XFILLER_2_197 VPWR VGND sg13g2_decap_8
XFILLER_38_319 VPWR VGND sg13g2_decap_8
XFILLER_48_71 VPWR VGND sg13g2_fill_1
Xfanout490 net246 net490 VPWR VGND sg13g2_buf_8
XFILLER_47_864 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_34_503 VPWR VGND sg13g2_decap_8
XFILLER_15_772 VPWR VGND sg13g2_fill_2
X_2990_ net417 _0118_ VPWR VGND sg13g2_buf_1
X_1941_ _1252_ _1253_ _0014_ VPWR VGND sg13g2_nor2b_2
XFILLER_14_271 VPWR VGND sg13g2_decap_8
XFILLER_30_731 VPWR VGND sg13g2_fill_1
XFILLER_9_76 VPWR VGND sg13g2_decap_8
X_1872_ _1196_ _1171_ _1194_ VPWR VGND sg13g2_nand2_1
XFILLER_9_98 VPWR VGND sg13g2_decap_8
XFILLER_9_1012 VPWR VGND sg13g2_decap_8
X_2424_ _0330_ _0320_ _0332_ VPWR VGND sg13g2_xor2_1
X_2355_ _0265_ net384 net441 net387 net497 VPWR VGND sg13g2_a22oi_1
X_2286_ _0198_ _0159_ _0057_ VPWR VGND sg13g2_xor2_1
XFILLER_38_875 VPWR VGND sg13g2_decap_8
XFILLER_25_547 VPWR VGND sg13g2_decap_8
XFILLER_25_558 VPWR VGND sg13g2_fill_1
XFILLER_33_580 VPWR VGND sg13g2_decap_8
XFILLER_0_657 VPWR VGND sg13g2_decap_8
XFILLER_47_138 VPWR VGND sg13g2_decap_8
XFILLER_29_864 VPWR VGND sg13g2_decap_8
XFILLER_44_845 VPWR VGND sg13g2_decap_8
XFILLER_16_547 VPWR VGND sg13g2_fill_1
XFILLER_16_558 VPWR VGND sg13g2_decap_8
XFILLER_34_40 VPWR VGND sg13g2_fill_1
XFILLER_43_399 VPWR VGND sg13g2_fill_1
XFILLER_12_742 VPWR VGND sg13g2_decap_8
XFILLER_12_753 VPWR VGND sg13g2_fill_1
XFILLER_15_1028 VPWR VGND sg13g2_fill_1
XFILLER_8_746 VPWR VGND sg13g2_decap_8
XFILLER_4_952 VPWR VGND sg13g2_decap_8
X_2140_ net399 net444 net442 net394 _1423_ VPWR VGND sg13g2_and4_1
X_2071_ _1357_ _1349_ _1356_ VPWR VGND sg13g2_nand2_1
XFILLER_19_374 VPWR VGND sg13g2_decap_8
XFILLER_35_812 VPWR VGND sg13g2_decap_8
XFILLER_47_694 VPWR VGND sg13g2_decap_8
XFILLER_34_311 VPWR VGND sg13g2_decap_8
XFILLER_15_580 VPWR VGND sg13g2_decap_8
X_2973_ net159 _0085_ VPWR VGND sg13g2_buf_1
X_1924_ net257 mac1.sum_lvl2_ff\[24\] _1240_ VPWR VGND sg13g2_xor2_1
X_1855_ _1180_ net403 net460 VPWR VGND sg13g2_nand2_1
X_1786_ _1110_ _1113_ _1114_ VPWR VGND sg13g2_nor2_1
X_2407_ _0290_ _0313_ _0315_ VPWR VGND sg13g2_and2_1
X_2338_ _0249_ _0204_ _0247_ VPWR VGND sg13g2_xnor2_1
X_2269_ _0182_ net496 net390 VPWR VGND sg13g2_nand2_1
XFILLER_25_322 VPWR VGND sg13g2_decap_8
XFILLER_41_815 VPWR VGND sg13g2_decap_8
XFILLER_40_303 VPWR VGND sg13g2_decap_8
XFILLER_25_377 VPWR VGND sg13g2_decap_8
XFILLER_21_594 VPWR VGND sg13g2_fill_2
XFILLER_5_727 VPWR VGND sg13g2_decap_8
XFILLER_1_933 VPWR VGND sg13g2_decap_8
XFILLER_0_454 VPWR VGND sg13g2_decap_8
XFILLER_49_937 VPWR VGND sg13g2_decap_8
Xhold40 mac1.sum_lvl1_ff\[86\] VPWR VGND net80 sg13g2_dlygate4sd3_1
XFILLER_29_51 VPWR VGND sg13g2_decap_8
Xhold51 mac1.products_ff\[138\] VPWR VGND net91 sg13g2_dlygate4sd3_1
Xhold73 mac1.products_ff\[143\] VPWR VGND net113 sg13g2_dlygate4sd3_1
Xhold62 mac1.sum_lvl1_ff\[46\] VPWR VGND net102 sg13g2_dlygate4sd3_1
Xhold95 mac1.products_ff\[72\] VPWR VGND net135 sg13g2_dlygate4sd3_1
Xhold84 mac1.sum_lvl2_ff\[45\] VPWR VGND net124 sg13g2_dlygate4sd3_1
XFILLER_29_661 VPWR VGND sg13g2_decap_4
XFILLER_29_683 VPWR VGND sg13g2_decap_8
XFILLER_17_834 VPWR VGND sg13g2_decap_8
XFILLER_43_141 VPWR VGND sg13g2_decap_8
XFILLER_32_837 VPWR VGND sg13g2_fill_2
XFILLER_8_532 VPWR VGND sg13g2_fill_2
XFILLER_8_565 VPWR VGND sg13g2_decap_8
XFILLER_6_22 VPWR VGND sg13g2_decap_8
X_1640_ _0971_ _0964_ _0969_ _0970_ VPWR VGND sg13g2_and3_1
X_1571_ VGND VPWR _0900_ _0901_ _0904_ _0895_ sg13g2_a21oi_1
XFILLER_6_88 VPWR VGND sg13g2_decap_8
X_3241_ net503 VGND VPWR net154 net25 clknet_leaf_37_clk sg13g2_dfrbpq_1
XFILLER_39_403 VPWR VGND sg13g2_decap_8
X_3172_ net540 VGND VPWR net58 mac1.sum_lvl2_ff\[30\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_2123_ VGND VPWR _1403_ _1404_ _1407_ _1379_ sg13g2_a21oi_1
X_2054_ _1341_ net457 net390 VPWR VGND sg13g2_nand2_1
XFILLER_19_171 VPWR VGND sg13g2_decap_8
XFILLER_35_620 VPWR VGND sg13g2_decap_4
XFILLER_34_152 VPWR VGND sg13g2_decap_8
XFILLER_35_664 VPWR VGND sg13g2_decap_8
XFILLER_35_697 VPWR VGND sg13g2_decap_8
XFILLER_23_859 VPWR VGND sg13g2_decap_4
XFILLER_22_369 VPWR VGND sg13g2_fill_1
X_2956_ _0834_ net431 net374 VPWR VGND sg13g2_nand2_1
X_2887_ _0774_ _0776_ _0777_ VPWR VGND sg13g2_nor2_1
X_1907_ mac1.sum_lvl2_ff\[20\] mac1.sum_lvl2_ff\[1\] _1227_ VPWR VGND sg13g2_nor2_1
X_1838_ VGND VPWR _1124_ _1135_ _1164_ _1123_ sg13g2_a21oi_1
X_1769_ _1093_ _1095_ _1096_ _1097_ VPWR VGND sg13g2_nor3_1
XFILLER_46_918 VPWR VGND sg13g2_decap_8
XFILLER_39_981 VPWR VGND sg13g2_decap_8
XFILLER_25_141 VPWR VGND sg13g2_decap_4
XFILLER_41_612 VPWR VGND sg13g2_decap_8
XFILLER_41_656 VPWR VGND sg13g2_decap_8
XFILLER_40_133 VPWR VGND sg13g2_decap_8
XFILLER_15_53 VPWR VGND sg13g2_decap_8
XFILLER_25_196 VPWR VGND sg13g2_decap_8
XFILLER_31_85 VPWR VGND sg13g2_decap_8
Xoutput30 net30 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_1_730 VPWR VGND sg13g2_decap_8
XFILLER_49_734 VPWR VGND sg13g2_decap_8
XFILLER_48_244 VPWR VGND sg13g2_decap_8
XFILLER_0_284 VPWR VGND sg13g2_decap_8
XFILLER_17_631 VPWR VGND sg13g2_decap_8
XFILLER_29_480 VPWR VGND sg13g2_fill_2
XFILLER_36_428 VPWR VGND sg13g2_decap_8
XFILLER_44_450 VPWR VGND sg13g2_fill_2
XFILLER_17_642 VPWR VGND sg13g2_fill_2
XFILLER_45_984 VPWR VGND sg13g2_decap_8
XFILLER_44_483 VPWR VGND sg13g2_fill_2
XFILLER_44_472 VPWR VGND sg13g2_decap_8
XFILLER_16_152 VPWR VGND sg13g2_fill_2
X_2810_ VGND VPWR _0678_ _0692_ _0703_ _0691_ sg13g2_a21oi_1
XFILLER_31_155 VPWR VGND sg13g2_decap_8
X_2741_ _0637_ _0628_ _0635_ VPWR VGND sg13g2_xnor2_1
XFILLER_9_830 VPWR VGND sg13g2_decap_8
XFILLER_8_351 VPWR VGND sg13g2_decap_8
X_2672_ _0569_ _0552_ _0570_ VPWR VGND sg13g2_xor2_1
X_1623_ _0954_ _0950_ _0953_ VPWR VGND sg13g2_nand2_1
X_1554_ _0878_ _0869_ _0877_ _0887_ VPWR VGND sg13g2_a21o_2
X_3224_ net529 VGND VPWR net76 mac1.sum_lvl3_ff\[35\] clknet_leaf_6_clk sg13g2_dfrbpq_1
.ends

