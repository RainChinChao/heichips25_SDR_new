* NGSPICE file created from heichips25_template.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_2 abstract view
.subckt sg13g2_and3_2 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

.subckt heichips25_template VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
X_3155_ _2748_ _2746_ _2747_ VPWR VGND sg13g2_nand2_1
XFILLER_28_929 VPWR VGND sg13g2_decap_8
X_3086_ _2680_ net985 net907 VPWR VGND sg13g2_nand2_1
X_3988_ _0819_ net997 net927 VPWR VGND sg13g2_nand2_1
XFILLER_23_667 VPWR VGND sg13g2_fill_1
X_5727_ VGND VPWR _2423_ _2422_ _2420_ sg13g2_or2_1
X_5658_ _2361_ _2362_ net17 VPWR VGND sg13g2_nor2b_1
X_5589_ VGND VPWR _2309_ mac2.sum_lvl3_ff\[9\] mac2.sum_lvl3_ff\[29\] sg13g2_or2_1
X_4609_ _1412_ net900 net839 VPWR VGND sg13g2_nand2_1
Xhold340 mac1.sum_lvl2_ff\[2\] VPWR VGND net380 sg13g2_dlygate4sd3_1
Xhold351 _2164_ VPWR VGND net391 sg13g2_dlygate4sd3_1
Xhold362 _0080_ VPWR VGND net402 sg13g2_dlygate4sd3_1
Xhold373 DP_2.matrix\[74\] VPWR VGND net413 sg13g2_dlygate4sd3_1
Xhold395 _2139_ VPWR VGND net435 sg13g2_dlygate4sd3_1
Xhold384 _2304_ VPWR VGND net424 sg13g2_dlygate4sd3_1
Xfanout820 net496 net820 VPWR VGND sg13g2_buf_8
Xfanout831 net373 net831 VPWR VGND sg13g2_buf_8
Xfanout842 DP_4.matrix\[2\] net842 VPWR VGND sg13g2_buf_1
Xfanout853 DP_3.matrix\[79\] net853 VPWR VGND sg13g2_buf_1
Xfanout875 DP_3.matrix\[42\] net875 VPWR VGND sg13g2_buf_8
Xfanout864 net865 net864 VPWR VGND sg13g2_buf_1
Xfanout886 net323 net886 VPWR VGND sg13g2_buf_8
Xfanout897 net898 net897 VPWR VGND sg13g2_buf_8
XFILLER_42_954 VPWR VGND sg13g2_decap_8
XFILLER_1_582 VPWR VGND sg13g2_decap_4
XFILLER_49_564 VPWR VGND sg13g2_fill_2
XFILLER_37_726 VPWR VGND sg13g2_fill_1
XFILLER_36_236 VPWR VGND sg13g2_fill_2
X_4960_ net812 net809 net863 net861 _1749_ VPWR VGND sg13g2_and4_1
X_3911_ net937 net989 net941 _0744_ VPWR VGND net986 sg13g2_nand4_1
XFILLER_33_954 VPWR VGND sg13g2_decap_8
X_4891_ VGND VPWR _1686_ _1687_ _1685_ _1627_ sg13g2_a21oi_2
X_3842_ net939 net994 net941 _0677_ VPWR VGND net993 sg13g2_nand4_1
XFILLER_20_604 VPWR VGND sg13g2_fill_1
XFILLER_20_626 VPWR VGND sg13g2_decap_4
X_5512_ VGND VPWR _2244_ _2246_ _2249_ net491 sg13g2_a21oi_1
X_3773_ VPWR _0615_ _0614_ VGND sg13g2_inv_1
X_6492_ net1054 VGND VPWR _0033_ mac2.sum_lvl3_ff\[10\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_5443_ _2195_ net358 mac1.sum_lvl3_ff\[9\] VPWR VGND sg13g2_nand2_1
X_5374_ _2141_ mac1.sum_lvl2_ff\[29\] mac1.sum_lvl2_ff\[10\] VPWR VGND sg13g2_nand2_1
X_4325_ _1141_ net814 net884 net817 net883 VPWR VGND sg13g2_a22oi_1
X_4256_ _1073_ _1040_ _1074_ VPWR VGND sg13g2_xor2_1
X_3207_ _2781_ VPWR _2798_ VGND _2760_ _2782_ sg13g2_o21ai_1
X_4187_ net825 net882 net831 _1008_ VPWR VGND net880 sg13g2_nand4_1
X_3138_ _2726_ VPWR _2731_ VGND _2727_ _2729_ sg13g2_o21ai_1
X_3069_ _2659_ VPWR _2664_ VGND _2660_ _2662_ sg13g2_o21ai_1
XFILLER_24_954 VPWR VGND sg13g2_decap_8
XFILLER_12_76 VPWR VGND sg13g2_fill_2
Xhold170 mac1.products_ff\[0\] VPWR VGND net210 sg13g2_dlygate4sd3_1
Xhold181 mac1.products_ff\[75\] VPWR VGND net221 sg13g2_dlygate4sd3_1
Xhold192 mac2.products_ff\[143\] VPWR VGND net232 sg13g2_dlygate4sd3_1
XFILLER_33_217 VPWR VGND sg13g2_fill_1
XFILLER_14_431 VPWR VGND sg13g2_fill_1
XFILLER_15_976 VPWR VGND sg13g2_decap_8
XFILLER_30_946 VPWR VGND sg13g2_decap_8
X_4110_ _0937_ _0916_ _0938_ VPWR VGND sg13g2_nor2b_1
XFILLER_25_1019 VPWR VGND sg13g2_decap_8
X_5090_ _1874_ _1810_ _1875_ VPWR VGND sg13g2_xor2_1
X_4041_ _0866_ VPWR _0871_ VGND _0868_ _0869_ sg13g2_o21ai_1
X_5992_ net274 _0240_ VPWR VGND sg13g2_buf_1
X_4943_ _1736_ _1730_ _1735_ VPWR VGND sg13g2_xnor2_1
XFILLER_17_280 VPWR VGND sg13g2_fill_2
XFILLER_32_250 VPWR VGND sg13g2_fill_1
XFILLER_33_751 VPWR VGND sg13g2_fill_2
X_4874_ _1667_ _1669_ _1670_ VPWR VGND sg13g2_nor2_1
XFILLER_21_957 VPWR VGND sg13g2_decap_8
XFILLER_33_784 VPWR VGND sg13g2_fill_1
X_3825_ _0661_ _0658_ _0660_ VPWR VGND sg13g2_nand2_1
X_3756_ _0598_ _0597_ _0592_ _0596_ _0574_ VPWR VGND sg13g2_a22oi_1
Xclkbuf_4_12_0_clk clknet_0_clk clknet_4_12_0_clk VPWR VGND sg13g2_buf_8
X_6475_ net1121 VGND VPWR net216 mac2.sum_lvl2_ff\[28\] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_5426_ net533 net501 _2181_ VPWR VGND sg13g2_and2_1
X_3687_ _0531_ _0528_ _0532_ VPWR VGND sg13g2_xor2_1
X_5357_ _2123_ net509 _2127_ _2128_ VPWR VGND sg13g2_nor3_1
X_5288_ _2067_ _2062_ _2065_ VPWR VGND sg13g2_xnor2_1
X_4308_ _1122_ _1123_ _1104_ _1125_ VPWR VGND sg13g2_nand3_1
X_4239_ _1056_ _1055_ _1038_ _1058_ VPWR VGND sg13g2_a21o_1
XFILLER_43_526 VPWR VGND sg13g2_fill_1
XFILLER_15_239 VPWR VGND sg13g2_fill_2
XFILLER_3_633 VPWR VGND sg13g2_fill_1
XFILLER_15_762 VPWR VGND sg13g2_fill_2
XFILLER_42_581 VPWR VGND sg13g2_decap_8
XFILLER_9_77 VPWR VGND sg13g2_fill_1
X_3610_ VGND VPWR _0457_ _0456_ _0407_ sg13g2_or2_1
X_4590_ _1394_ net899 net841 VPWR VGND sg13g2_nand2_1
X_3541_ _0389_ _0325_ _0390_ VPWR VGND sg13g2_xor2_1
XFILLER_7_983 VPWR VGND sg13g2_decap_8
X_3472_ _0322_ _0314_ _0316_ VPWR VGND sg13g2_nand2_1
X_6260_ net1061 VGND VPWR net132 mac2.sum_lvl2_ff\[45\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_6191_ net1072 VGND VPWR net202 mac1.sum_lvl1_ff\[38\] clknet_leaf_56_clk sg13g2_dfrbpq_1
X_5211_ _1991_ _1964_ _1993_ VPWR VGND sg13g2_xor2_1
X_5142_ _1915_ VPWR _1925_ VGND _1844_ _1916_ sg13g2_o21ai_1
XFILLER_29_309 VPWR VGND sg13g2_fill_1
XFILLER_38_821 VPWR VGND sg13g2_decap_8
X_5073_ _1858_ net853 net813 net855 net806 VPWR VGND sg13g2_a22oi_1
X_4024_ _0829_ VPWR _0854_ VGND _0827_ _0830_ sg13g2_o21ai_1
XFILLER_38_898 VPWR VGND sg13g2_decap_8
XFILLER_37_386 VPWR VGND sg13g2_fill_1
X_5975_ net279 _0215_ VPWR VGND sg13g2_buf_1
XFILLER_12_209 VPWR VGND sg13g2_fill_1
X_4926_ _1720_ _1719_ _1716_ VPWR VGND sg13g2_nand2b_1
X_4857_ VPWR _1654_ _1653_ VGND sg13g2_inv_1
X_3808_ _0645_ _0644_ _0632_ VPWR VGND sg13g2_nand2b_1
X_4788_ _1587_ _1556_ _1585_ VPWR VGND sg13g2_xnor2_1
X_3739_ _0582_ _0577_ _0580_ VPWR VGND sg13g2_xnor2_1
X_6458_ net1103 VGND VPWR net45 mac2.sum_lvl2_ff\[8\] clknet_leaf_42_clk sg13g2_dfrbpq_1
X_5409_ _0023_ _2165_ _2168_ VPWR VGND sg13g2_xnor2_1
X_6389_ net1119 VGND VPWR _0136_ mac2.products_ff\[76\] clknet_leaf_40_clk sg13g2_dfrbpq_1
XFILLER_0_625 VPWR VGND sg13g2_fill_1
XFILLER_47_117 VPWR VGND sg13g2_decap_8
XFILLER_29_876 VPWR VGND sg13g2_decap_8
XFILLER_31_529 VPWR VGND sg13g2_fill_1
XFILLER_15_1018 VPWR VGND sg13g2_decap_8
XFILLER_4_986 VPWR VGND sg13g2_decap_8
XFILLER_3_463 VPWR VGND sg13g2_fill_2
XFILLER_35_846 VPWR VGND sg13g2_decap_8
XFILLER_34_356 VPWR VGND sg13g2_fill_1
XFILLER_43_890 VPWR VGND sg13g2_decap_8
X_5760_ VGND VPWR _2455_ _2454_ _2452_ sg13g2_or2_1
X_5691_ _2386_ VPWR _2389_ VGND _2385_ _2387_ sg13g2_o21ai_1
X_4711_ net902 net900 net834 net832 _1511_ VPWR VGND sg13g2_and4_1
X_4642_ _1444_ net898 net840 VPWR VGND sg13g2_nand2_1
X_4573_ net847 net843 net899 net897 _1378_ VPWR VGND sg13g2_and4_1
X_3524_ _0373_ net1006 net962 net1007 net957 VPWR VGND sg13g2_a22oi_1
X_6312_ net1046 VGND VPWR net84 mac1.sum_lvl3_ff\[31\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_3455_ _0306_ net1009 net962 net1011 net958 VPWR VGND sg13g2_a22oi_1
X_6243_ net1066 VGND VPWR net203 mac1.sum_lvl2_ff\[44\] clknet_leaf_64_clk sg13g2_dfrbpq_1
X_3386_ _0099_ _2954_ _2970_ VPWR VGND sg13g2_xnor2_1
X_6174_ net1121 VGND VPWR _0253_ DP_4.matrix\[37\] clknet_4_14_0_clk sg13g2_dfrbpq_1
X_5125_ _1909_ _1890_ _1907_ _1908_ VPWR VGND sg13g2_and3_1
X_5056_ _1841_ net792 net868 net795 net866 VPWR VGND sg13g2_a22oi_1
X_4007_ _0838_ _0833_ _0837_ VPWR VGND sg13g2_nand2_1
XFILLER_26_857 VPWR VGND sg13g2_decap_8
XFILLER_41_816 VPWR VGND sg13g2_decap_8
X_5958_ net980 _0190_ VPWR VGND sg13g2_buf_1
XFILLER_13_518 VPWR VGND sg13g2_fill_1
X_4909_ _1702_ _1688_ _1704_ VPWR VGND sg13g2_xor2_1
X_5889_ _2460_ _2456_ _2569_ VPWR VGND sg13g2_xor2_1
XFILLER_0_411 VPWR VGND sg13g2_fill_1
XFILLER_1_945 VPWR VGND sg13g2_decap_8
Xhold30 mac1.products_ff\[11\] VPWR VGND net70 sg13g2_dlygate4sd3_1
Xhold41 mac1.sum_lvl2_ff\[52\] VPWR VGND net81 sg13g2_dlygate4sd3_1
Xhold52 mac1.sum_lvl1_ff\[7\] VPWR VGND net92 sg13g2_dlygate4sd3_1
Xhold63 mac1.products_ff\[150\] VPWR VGND net103 sg13g2_dlygate4sd3_1
Xhold74 mac2.products_ff\[68\] VPWR VGND net114 sg13g2_dlygate4sd3_1
Xhold85 mac2.products_ff\[14\] VPWR VGND net125 sg13g2_dlygate4sd3_1
Xhold96 mac1.sum_lvl1_ff\[87\] VPWR VGND net136 sg13g2_dlygate4sd3_1
XFILLER_16_389 VPWR VGND sg13g2_fill_2
XFILLER_32_838 VPWR VGND sg13g2_decap_8
XFILLER_40_882 VPWR VGND sg13g2_decap_8
XFILLER_6_45 VPWR VGND sg13g2_fill_1
X_3240_ _2831_ _2797_ _2829_ VPWR VGND sg13g2_xnor2_1
X_3171_ _2763_ net911 net969 VPWR VGND sg13g2_nand2_2
XFILLER_6_1027 VPWR VGND sg13g2_fill_2
Xfanout1072 net1076 net1072 VPWR VGND sg13g2_buf_8
Xfanout1050 net1051 net1050 VPWR VGND sg13g2_buf_8
Xfanout1061 net1062 net1061 VPWR VGND sg13g2_buf_8
Xfanout1083 net1086 net1083 VPWR VGND sg13g2_buf_8
XFILLER_48_982 VPWR VGND sg13g2_decap_8
Xfanout1094 net1095 net1094 VPWR VGND sg13g2_buf_2
X_5812_ _2506_ net280 net775 VPWR VGND sg13g2_nand2_1
X_5743_ _2395_ net1032 _2437_ _2438_ VPWR VGND sg13g2_a21o_1
X_5674_ _2375_ mac1.total_sum\[12\] mac2.total_sum\[12\] VPWR VGND sg13g2_nand2_1
X_4625_ _1426_ _1427_ _1409_ _1428_ VPWR VGND sg13g2_nand3_1
X_4556_ _1365_ _1359_ _1364_ VPWR VGND sg13g2_xnor2_1
Xhold500 _0061_ VPWR VGND net540 sg13g2_dlygate4sd3_1
X_3507_ _0356_ net944 net1020 net946 net1017 VPWR VGND sg13g2_a22oi_1
X_4487_ _1299_ _1298_ _1295_ VPWR VGND sg13g2_nand2b_1
XFILLER_44_1000 VPWR VGND sg13g2_decap_8
X_3438_ _0290_ _0278_ _0289_ VPWR VGND sg13g2_xnor2_1
X_6226_ net1096 VGND VPWR net174 mac1.sum_lvl2_ff\[24\] clknet_leaf_54_clk sg13g2_dfrbpq_2
X_3369_ VGND VPWR _2931_ _2945_ _2955_ _2944_ sg13g2_a21oi_1
X_6157_ net1087 VGND VPWR _0240_ DP_3.matrix\[76\] clknet_leaf_25_clk sg13g2_dfrbpq_1
XFILLER_46_908 VPWR VGND sg13g2_decap_8
X_5108_ _1892_ net800 net856 VPWR VGND sg13g2_nand2_2
X_6088_ net1073 VGND VPWR _0194_ DP_1.matrix\[78\] clknet_leaf_60_clk sg13g2_dfrbpq_2
XFILLER_39_982 VPWR VGND sg13g2_decap_8
XFILLER_26_632 VPWR VGND sg13g2_fill_1
X_5039_ _1820_ VPWR _1825_ VGND _1821_ _1823_ sg13g2_o21ai_1
XFILLER_40_156 VPWR VGND sg13g2_fill_2
XFILLER_41_679 VPWR VGND sg13g2_fill_2
XFILLER_5_514 VPWR VGND sg13g2_fill_1
XFILLER_5_503 VPWR VGND sg13g2_fill_2
XFILLER_5_525 VPWR VGND sg13g2_fill_1
Xoutput31 net31 uo_out[6] VPWR VGND sg13g2_buf_1
Xoutput20 net20 uio_out[3] VPWR VGND sg13g2_buf_1
XFILLER_45_952 VPWR VGND sg13g2_decap_8
X_4410_ _1192_ VPWR _1224_ VGND _1139_ _1190_ sg13g2_o21ai_1
X_5390_ _0003_ net482 _2154_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_1006 VPWR VGND sg13g2_decap_8
X_4341_ net829 net826 net871 net1026 _1157_ VPWR VGND sg13g2_and4_1
X_4272_ VGND VPWR _1087_ _1088_ _1090_ _1070_ sg13g2_a21oi_1
X_6011_ net794 _0267_ VPWR VGND sg13g2_buf_1
X_3223_ _2763_ _2812_ _2814_ VPWR VGND sg13g2_and2_1
XFILLER_39_212 VPWR VGND sg13g2_fill_2
X_3154_ _2709_ _2708_ _2707_ _2747_ VPWR VGND sg13g2_a21o_2
XFILLER_28_908 VPWR VGND sg13g2_decap_8
X_3085_ _2656_ VPWR _2679_ VGND _2631_ _2654_ sg13g2_o21ai_1
XFILLER_35_440 VPWR VGND sg13g2_fill_2
XFILLER_36_985 VPWR VGND sg13g2_decap_8
X_3987_ _0818_ net997 net925 VPWR VGND sg13g2_nand2_1
X_5726_ _2422_ _2421_ net782 net781 net980 VPWR VGND sg13g2_a22oi_1
X_5657_ _2358_ _2360_ _2356_ _2362_ VPWR VGND sg13g2_nand3_1
X_5588_ mac2.sum_lvl3_ff\[29\] mac2.sum_lvl3_ff\[9\] _2308_ VPWR VGND sg13g2_and2_1
X_4608_ _1411_ net900 net837 VPWR VGND sg13g2_nand2_1
X_4539_ _1349_ _1344_ _1347_ VPWR VGND sg13g2_xnor2_1
Xhold341 _2115_ VPWR VGND net381 sg13g2_dlygate4sd3_1
Xhold330 mac1.sum_lvl2_ff\[3\] VPWR VGND net370 sg13g2_dlygate4sd3_1
Xhold352 _0006_ VPWR VGND net392 sg13g2_dlygate4sd3_1
Xhold374 DP_4.matrix\[4\] VPWR VGND net414 sg13g2_dlygate4sd3_1
Xhold396 _2140_ VPWR VGND net436 sg13g2_dlygate4sd3_1
Xhold363 DP_1.matrix\[44\] VPWR VGND net403 sg13g2_dlygate4sd3_1
Xhold385 _2305_ VPWR VGND net425 sg13g2_dlygate4sd3_1
Xfanout832 net366 net832 VPWR VGND sg13g2_buf_8
Xfanout821 net822 net821 VPWR VGND sg13g2_buf_8
X_6209_ net1097 VGND VPWR net118 mac1.sum_lvl2_ff\[4\] clknet_leaf_54_clk sg13g2_dfrbpq_1
Xfanout843 net404 net843 VPWR VGND sg13g2_buf_8
Xfanout810 net301 net810 VPWR VGND sg13g2_buf_1
Xfanout876 net340 net876 VPWR VGND sg13g2_buf_8
Xfanout854 net855 net854 VPWR VGND sg13g2_buf_8
Xfanout865 net521 net865 VPWR VGND sg13g2_buf_2
Xfanout887 DP_3.matrix\[36\] net887 VPWR VGND sg13g2_buf_1
Xfanout898 net525 net898 VPWR VGND sg13g2_buf_8
XFILLER_27_985 VPWR VGND sg13g2_decap_8
XFILLER_42_933 VPWR VGND sg13g2_decap_8
XFILLER_13_112 VPWR VGND sg13g2_fill_1
XFILLER_14_657 VPWR VGND sg13g2_fill_1
XFILLER_9_116 VPWR VGND sg13g2_fill_2
XFILLER_13_167 VPWR VGND sg13g2_fill_2
XFILLER_10_874 VPWR VGND sg13g2_fill_1
XFILLER_5_377 VPWR VGND sg13g2_fill_1
XFILLER_36_204 VPWR VGND sg13g2_fill_2
XFILLER_18_996 VPWR VGND sg13g2_decap_8
X_3910_ net941 net937 net989 net987 _0743_ VPWR VGND sg13g2_and4_1
XFILLER_33_933 VPWR VGND sg13g2_decap_8
X_4890_ VGND VPWR _1624_ _1653_ _1686_ _1655_ sg13g2_a21oi_1
X_3841_ net942 net939 net994 net993 _0676_ VPWR VGND sg13g2_and4_1
XFILLER_32_465 VPWR VGND sg13g2_decap_4
X_3772_ _0612_ _0599_ _0614_ VPWR VGND sg13g2_xor2_1
XFILLER_34_1021 VPWR VGND sg13g2_decap_8
X_5511_ _2248_ mac2.sum_lvl2_ff\[27\] net490 VPWR VGND sg13g2_xnor2_1
X_6491_ net1061 VGND VPWR _0047_ mac2.sum_lvl3_ff\[9\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_5442_ _2190_ _2192_ _2194_ VPWR VGND sg13g2_nor2_1
X_5373_ _0015_ _2137_ net436 VPWR VGND sg13g2_xnor2_1
X_4324_ net884 net883 net817 net814 _1140_ VPWR VGND sg13g2_and4_1
X_4255_ _1073_ net881 net822 VPWR VGND sg13g2_nand2_2
X_3206_ _2758_ VPWR _2797_ VGND _2713_ _2759_ sg13g2_o21ai_1
X_4186_ net831 net825 net882 net880 _1007_ VPWR VGND sg13g2_and4_1
X_3137_ _2726_ _2727_ _2729_ _2730_ VPWR VGND sg13g2_or3_1
X_3068_ _2659_ _2660_ _2662_ _2663_ VPWR VGND sg13g2_or3_1
XFILLER_24_933 VPWR VGND sg13g2_decap_8
X_5709_ _2397_ net790 _2405_ VPWR VGND sg13g2_and2_1
Xhold160 mac1.sum_lvl1_ff\[72\] VPWR VGND net200 sg13g2_dlygate4sd3_1
Xhold171 mac1.products_ff\[151\] VPWR VGND net211 sg13g2_dlygate4sd3_1
Xhold182 mac2.products_ff\[81\] VPWR VGND net222 sg13g2_dlygate4sd3_1
Xhold193 mac2.products_ff\[73\] VPWR VGND net233 sg13g2_dlygate4sd3_1
XFILLER_46_502 VPWR VGND sg13g2_decap_8
XFILLER_46_557 VPWR VGND sg13g2_fill_2
XFILLER_46_535 VPWR VGND sg13g2_fill_2
XFILLER_18_226 VPWR VGND sg13g2_fill_1
XFILLER_15_955 VPWR VGND sg13g2_decap_8
XFILLER_30_925 VPWR VGND sg13g2_decap_8
XFILLER_5_141 VPWR VGND sg13g2_fill_1
X_4040_ _0866_ _0868_ _0869_ _0870_ VPWR VGND sg13g2_nor3_1
XFILLER_49_384 VPWR VGND sg13g2_fill_1
XFILLER_49_362 VPWR VGND sg13g2_fill_2
XFILLER_37_502 VPWR VGND sg13g2_fill_2
X_5991_ net862 _0239_ VPWR VGND sg13g2_buf_1
X_4942_ _1735_ _1722_ _1734_ VPWR VGND sg13g2_xnor2_1
X_4873_ _1669_ net833 net893 net834 DP_3.matrix\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_21_936 VPWR VGND sg13g2_decap_8
X_3824_ _0657_ _0656_ _0651_ _0660_ VPWR VGND sg13g2_a21o_1
X_3755_ _0591_ VPWR _0597_ VGND _0568_ _0569_ sg13g2_o21ai_1
X_3686_ _0531_ _0484_ _0529_ VPWR VGND sg13g2_xnor2_1
X_6474_ net1121 VGND VPWR net239 mac2.sum_lvl2_ff\[27\] clknet_leaf_40_clk sg13g2_dfrbpq_2
X_5425_ _0027_ _2178_ net321 VPWR VGND sg13g2_xnor2_1
X_5356_ VPWR VGND _2121_ _2120_ _2119_ mac1.sum_lvl2_ff\[24\] _2127_ mac1.sum_lvl2_ff\[5\]
+ sg13g2_a221oi_1
X_5287_ _2066_ _2065_ _2062_ VPWR VGND sg13g2_nand2b_1
X_4307_ _1124_ _1104_ _1122_ _1123_ VPWR VGND sg13g2_and3_1
X_4238_ _1055_ _1056_ _1038_ _1057_ VPWR VGND sg13g2_nand3_1
X_4169_ _0994_ _0988_ _0993_ VPWR VGND sg13g2_xnor2_1
XFILLER_43_505 VPWR VGND sg13g2_fill_2
XFILLER_23_32 VPWR VGND sg13g2_fill_1
XFILLER_11_479 VPWR VGND sg13g2_fill_1
XFILLER_3_645 VPWR VGND sg13g2_fill_1
XFILLER_47_899 VPWR VGND sg13g2_decap_8
XFILLER_34_516 VPWR VGND sg13g2_decap_4
XFILLER_15_730 VPWR VGND sg13g2_fill_2
XFILLER_31_1024 VPWR VGND sg13g2_decap_4
XFILLER_7_962 VPWR VGND sg13g2_decap_8
X_3540_ _0389_ _0386_ _0388_ VPWR VGND sg13g2_nand2_1
XFILLER_6_450 VPWR VGND sg13g2_fill_1
X_3471_ _0105_ _0294_ _0321_ VPWR VGND sg13g2_xnor2_1
X_5210_ _1992_ _1991_ _1964_ VPWR VGND sg13g2_nand2b_1
X_6190_ net1070 VGND VPWR net199 mac1.sum_lvl1_ff\[37\] clknet_leaf_62_clk sg13g2_dfrbpq_1
XFILLER_9_1014 VPWR VGND sg13g2_decap_8
X_5141_ _1920_ VPWR _1924_ VGND _1877_ _1922_ sg13g2_o21ai_1
X_5072_ net806 net855 net813 _1857_ VPWR VGND net853 sg13g2_nand4_1
X_4023_ _0821_ VPWR _0853_ VGND _0768_ _0819_ sg13g2_o21ai_1
XFILLER_38_877 VPWR VGND sg13g2_decap_8
X_5974_ net916 _0214_ VPWR VGND sg13g2_buf_1
X_4925_ _1718_ _1691_ _1719_ VPWR VGND sg13g2_xor2_1
XFILLER_33_560 VPWR VGND sg13g2_fill_1
XFILLER_40_519 VPWR VGND sg13g2_decap_4
X_4856_ _1621_ _1652_ _1619_ _1653_ VPWR VGND sg13g2_nand3_1
X_3807_ _0643_ _0633_ _0644_ VPWR VGND sg13g2_xor2_1
X_4787_ _1586_ _1556_ _1585_ VPWR VGND sg13g2_nand2_1
X_3738_ _0581_ _0580_ _0577_ VPWR VGND sg13g2_nand2b_1
X_3669_ _0513_ _0511_ _0106_ VPWR VGND sg13g2_xor2_1
X_6457_ net1103 VGND VPWR net61 mac2.sum_lvl2_ff\[7\] clknet_leaf_43_clk sg13g2_dfrbpq_1
XFILLER_0_604 VPWR VGND sg13g2_fill_2
X_5408_ mac1.sum_lvl3_ff\[1\] mac1.sum_lvl3_ff\[21\] _2168_ VPWR VGND sg13g2_xor2_1
X_6388_ net1119 VGND VPWR _0135_ mac2.products_ff\[75\] clknet_leaf_41_clk sg13g2_dfrbpq_1
X_5339_ mac1.sum_lvl2_ff\[21\] mac1.sum_lvl2_ff\[2\] _2114_ VPWR VGND sg13g2_and2_1
Xclkbuf_leaf_67_clk clknet_4_0_0_clk clknet_leaf_67_clk VPWR VGND sg13g2_buf_8
XFILLER_29_855 VPWR VGND sg13g2_decap_8
XFILLER_44_825 VPWR VGND sg13g2_decap_4
XFILLER_34_42 VPWR VGND sg13g2_fill_2
XFILLER_34_97 VPWR VGND sg13g2_fill_1
XFILLER_7_269 VPWR VGND sg13g2_fill_1
XFILLER_4_921 VPWR VGND sg13g2_fill_2
XFILLER_4_965 VPWR VGND sg13g2_decap_8
XFILLER_19_332 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_58_clk clknet_4_9_0_clk clknet_leaf_58_clk VPWR VGND sg13g2_buf_8
Xclkbuf_4_11_0_clk clknet_0_clk clknet_4_11_0_clk VPWR VGND sg13g2_buf_8
XFILLER_35_825 VPWR VGND sg13g2_decap_8
X_4710_ _1510_ net900 net832 VPWR VGND sg13g2_nand2_1
X_5690_ net23 _2385_ _2388_ VPWR VGND sg13g2_xnor2_1
X_4641_ _1443_ net898 net837 VPWR VGND sg13g2_nand2_1
X_4572_ _1377_ net901 net841 VPWR VGND sg13g2_nand2_1
XFILLER_6_280 VPWR VGND sg13g2_fill_1
X_3523_ net957 net1007 net961 _0372_ VPWR VGND net1006 sg13g2_nand4_1
X_6311_ net1047 VGND VPWR net156 mac1.sum_lvl3_ff\[30\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_3454_ net958 net1011 net962 _0305_ VPWR VGND net1009 sg13g2_nand4_1
X_6242_ net1041 VGND VPWR net158 mac1.sum_lvl2_ff\[43\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3385_ VPWR _2971_ _2970_ VGND sg13g2_inv_1
X_6173_ net1106 VGND VPWR _0252_ DP_4.matrix\[36\] clknet_leaf_32_clk sg13g2_dfrbpq_2
X_5124_ _1896_ VPWR _1908_ VGND _1904_ _1906_ sg13g2_o21ai_1
Xclkbuf_leaf_49_clk clknet_4_10_0_clk clknet_leaf_49_clk VPWR VGND sg13g2_buf_8
X_5055_ _1817_ VPWR _1840_ VGND _1782_ _1815_ sg13g2_o21ai_1
X_4006_ _0835_ _0836_ _0837_ VPWR VGND sg13g2_nor2_1
XFILLER_26_836 VPWR VGND sg13g2_decap_4
XFILLER_38_685 VPWR VGND sg13g2_fill_2
X_5957_ net983 _0189_ VPWR VGND sg13g2_buf_1
X_4908_ _1703_ _1688_ _1702_ VPWR VGND sg13g2_nand2_1
X_5888_ net951 net772 _2568_ VPWR VGND sg13g2_nor2_1
X_4839_ _1635_ _1632_ _1636_ VPWR VGND sg13g2_xor2_1
XFILLER_20_33 VPWR VGND sg13g2_fill_2
X_6509_ net1044 VGND VPWR net339 mac2.total_sum\[11\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_1_924 VPWR VGND sg13g2_decap_8
XFILLER_29_42 VPWR VGND sg13g2_fill_1
Xhold31 mac2.products_ff\[137\] VPWR VGND net71 sg13g2_dlygate4sd3_1
Xhold20 mac2.sum_lvl2_ff\[52\] VPWR VGND net60 sg13g2_dlygate4sd3_1
Xhold53 mac1.sum_lvl1_ff\[75\] VPWR VGND net93 sg13g2_dlygate4sd3_1
Xhold64 mac2.products_ff\[8\] VPWR VGND net104 sg13g2_dlygate4sd3_1
Xhold42 mac2.sum_lvl1_ff\[47\] VPWR VGND net82 sg13g2_dlygate4sd3_1
Xhold75 mac2.sum_lvl1_ff\[83\] VPWR VGND net115 sg13g2_dlygate4sd3_1
Xhold97 mac2.sum_lvl2_ff\[41\] VPWR VGND net137 sg13g2_dlygate4sd3_1
Xhold86 mac2.products_ff\[72\] VPWR VGND net126 sg13g2_dlygate4sd3_1
XFILLER_17_836 VPWR VGND sg13g2_fill_2
XFILLER_45_96 VPWR VGND sg13g2_decap_4
XFILLER_40_861 VPWR VGND sg13g2_decap_8
XFILLER_6_1006 VPWR VGND sg13g2_decap_8
X_3170_ _2762_ net975 net909 VPWR VGND sg13g2_nand2_1
Xfanout1040 net1043 net1040 VPWR VGND sg13g2_buf_8
Xfanout1073 net1075 net1073 VPWR VGND sg13g2_buf_8
Xfanout1051 net1063 net1051 VPWR VGND sg13g2_buf_8
Xfanout1062 net1063 net1062 VPWR VGND sg13g2_buf_8
XFILLER_39_427 VPWR VGND sg13g2_decap_4
XFILLER_48_961 VPWR VGND sg13g2_decap_8
Xfanout1095 net1107 net1095 VPWR VGND sg13g2_buf_8
Xfanout1084 net1086 net1084 VPWR VGND sg13g2_buf_8
X_5811_ _2505_ _2486_ _2504_ VPWR VGND sg13g2_nand2b_1
XFILLER_16_880 VPWR VGND sg13g2_decap_8
XFILLER_23_839 VPWR VGND sg13g2_fill_2
X_5742_ net773 _2436_ _2437_ VPWR VGND sg13g2_and2_1
XFILLER_16_891 VPWR VGND sg13g2_fill_1
X_5673_ net20 _2373_ _2374_ VPWR VGND sg13g2_xnor2_1
X_4624_ _1415_ VPWR _1427_ VGND _1423_ _1425_ sg13g2_o21ai_1
Xhold501 DP_4.matrix\[8\] VPWR VGND net541 sg13g2_dlygate4sd3_1
X_4555_ _1364_ _1351_ _1363_ VPWR VGND sg13g2_xnor2_1
X_3506_ _0332_ VPWR _0355_ VGND _0297_ _0330_ sg13g2_o21ai_1
X_4486_ _1297_ _1270_ _1298_ VPWR VGND sg13g2_xor2_1
X_3437_ _0289_ _0286_ _0288_ VPWR VGND sg13g2_nand2_1
X_6225_ net1097 VGND VPWR net143 mac1.sum_lvl2_ff\[23\] clknet_leaf_54_clk sg13g2_dfrbpq_1
X_3368_ _2954_ _2953_ _2948_ _2952_ _2930_ VPWR VGND sg13g2_a22oi_1
X_6156_ net1112 VGND VPWR net70 mac1.sum_lvl1_ff\[11\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_5107_ _1891_ net860 net798 VPWR VGND sg13g2_nand2_1
Xheichips25_template_33 VPWR VGND uio_oe[0] sg13g2_tiehi
X_6087_ net1064 VGND VPWR _0068_ mac1.products_ff\[140\] clknet_leaf_66_clk sg13g2_dfrbpq_1
X_3299_ _2888_ _2840_ _2886_ VPWR VGND sg13g2_xnor2_1
XFILLER_39_961 VPWR VGND sg13g2_decap_8
X_5038_ _1820_ _1821_ _1823_ _1824_ VPWR VGND sg13g2_or3_1
XFILLER_25_110 VPWR VGND sg13g2_fill_2
XFILLER_14_817 VPWR VGND sg13g2_fill_2
XFILLER_26_699 VPWR VGND sg13g2_fill_2
XFILLER_13_349 VPWR VGND sg13g2_fill_2
XFILLER_31_21 VPWR VGND sg13g2_fill_1
Xoutput32 net32 uo_out[7] VPWR VGND sg13g2_buf_1
Xoutput21 net21 uio_out[4] VPWR VGND sg13g2_buf_1
XFILLER_36_408 VPWR VGND sg13g2_decap_8
XFILLER_45_931 VPWR VGND sg13g2_decap_8
XFILLER_36_419 VPWR VGND sg13g2_fill_1
XFILLER_32_647 VPWR VGND sg13g2_decap_4
XFILLER_9_876 VPWR VGND sg13g2_fill_1
X_4340_ _1156_ net823 net873 VPWR VGND sg13g2_nand2_1
X_4271_ _1087_ _1088_ _1070_ _1089_ VPWR VGND sg13g2_nand3_1
X_6010_ net797 _0266_ VPWR VGND sg13g2_buf_1
X_3222_ VGND VPWR _2813_ _2812_ _2763_ sg13g2_or2_1
X_3153_ _2745_ _2681_ _2746_ VPWR VGND sg13g2_xor2_1
X_3084_ _2678_ _2670_ _2672_ VPWR VGND sg13g2_nand2_1
XFILLER_36_964 VPWR VGND sg13g2_decap_8
XFILLER_10_308 VPWR VGND sg13g2_fill_2
X_3986_ _0817_ net1002 net1031 VPWR VGND sg13g2_nand2_1
X_5725_ net1015 net1000 net789 _2421_ VPWR VGND sg13g2_mux2_1
X_5656_ VGND VPWR _2356_ _2358_ _2361_ _2360_ sg13g2_a21oi_1
X_4607_ _1410_ net904 net836 VPWR VGND sg13g2_nand2_1
Xhold320 _0031_ VPWR VGND net360 sg13g2_dlygate4sd3_1
X_5587_ net423 net429 net425 _2307_ VPWR VGND sg13g2_a21o_1
X_4538_ _1348_ _1347_ _1344_ VPWR VGND sg13g2_nand2b_1
Xhold353 DP_2.matrix\[2\] VPWR VGND net393 sg13g2_dlygate4sd3_1
Xhold342 _0008_ VPWR VGND net382 sg13g2_dlygate4sd3_1
Xhold331 _2118_ VPWR VGND net371 sg13g2_dlygate4sd3_1
Xfanout800 net801 net800 VPWR VGND sg13g2_buf_8
Xhold375 _0248_ VPWR VGND net415 sg13g2_dlygate4sd3_1
Xhold386 _0062_ VPWR VGND net426 sg13g2_dlygate4sd3_1
Xhold364 DP_4.matrix\[1\] VPWR VGND net404 sg13g2_dlygate4sd3_1
X_4469_ _1280_ _1258_ _1282_ VPWR VGND sg13g2_xor2_1
Xfanout833 DP_4.matrix\[7\] net833 VPWR VGND sg13g2_buf_1
Xfanout822 net497 net822 VPWR VGND sg13g2_buf_8
X_6208_ net1095 VGND VPWR net120 mac1.sum_lvl2_ff\[3\] clknet_leaf_55_clk sg13g2_dfrbpq_1
Xhold397 _0015_ VPWR VGND net437 sg13g2_dlygate4sd3_1
Xfanout811 net812 net811 VPWR VGND sg13g2_buf_2
Xfanout855 DP_3.matrix\[78\] net855 VPWR VGND sg13g2_buf_8
Xfanout866 net867 net866 VPWR VGND sg13g2_buf_8
Xfanout844 DP_4.matrix\[1\] net844 VPWR VGND sg13g2_buf_1
XFILLER_46_717 VPWR VGND sg13g2_fill_2
Xfanout877 DP_3.matrix\[41\] net877 VPWR VGND sg13g2_buf_8
Xfanout888 net890 net888 VPWR VGND sg13g2_buf_2
X_6139_ net1106 VGND VPWR _0228_ DP_3.matrix\[36\] clknet_leaf_31_clk sg13g2_dfrbpq_1
Xfanout899 net476 net899 VPWR VGND sg13g2_buf_2
XFILLER_27_964 VPWR VGND sg13g2_decap_8
XFILLER_39_791 VPWR VGND sg13g2_fill_1
XFILLER_42_912 VPWR VGND sg13g2_decap_8
XFILLER_14_603 VPWR VGND sg13g2_fill_2
XFILLER_26_463 VPWR VGND sg13g2_fill_2
XFILLER_42_989 VPWR VGND sg13g2_decap_8
XFILLER_13_157 VPWR VGND sg13g2_fill_1
XFILLER_41_488 VPWR VGND sg13g2_decap_4
XFILLER_49_500 VPWR VGND sg13g2_fill_2
XFILLER_49_566 VPWR VGND sg13g2_fill_1
XFILLER_18_975 VPWR VGND sg13g2_decap_8
XFILLER_33_912 VPWR VGND sg13g2_decap_8
XFILLER_44_260 VPWR VGND sg13g2_fill_2
X_3840_ _0675_ net935 net997 VPWR VGND sg13g2_nand2_1
XFILLER_33_989 VPWR VGND sg13g2_decap_8
XFILLER_34_1000 VPWR VGND sg13g2_decap_8
X_3771_ VGND VPWR _0613_ _0612_ _0599_ sg13g2_or2_1
X_5510_ _2246_ _2247_ _0045_ VPWR VGND sg13g2_and2_1
X_6490_ net1051 VGND VPWR net493 mac2.sum_lvl3_ff\[8\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_5441_ _2192_ net421 _0030_ VPWR VGND sg13g2_nor2b_1
X_5372_ _2140_ net435 _2138_ VPWR VGND sg13g2_nand2b_1
X_4323_ _1139_ net883 net814 VPWR VGND sg13g2_nand2_1
X_4254_ _1072_ net881 net820 VPWR VGND sg13g2_nand2_1
X_3205_ _2786_ VPWR _2796_ VGND _2715_ _2787_ sg13g2_o21ai_1
X_4185_ _1006_ net885 net823 VPWR VGND sg13g2_nand2_1
XFILLER_41_1026 VPWR VGND sg13g2_fill_2
X_3136_ _2729_ net964 net921 net967 net918 VPWR VGND sg13g2_a22oi_1
X_3067_ _2662_ net969 net921 net972 net917 VPWR VGND sg13g2_a22oi_1
XFILLER_24_989 VPWR VGND sg13g2_decap_8
XFILLER_11_639 VPWR VGND sg13g2_fill_2
X_3969_ _0801_ _0765_ _0799_ _0800_ VPWR VGND sg13g2_and3_1
X_5708_ net772 _2403_ _2404_ VPWR VGND sg13g2_and2_1
X_5639_ _2347_ _2345_ net29 VPWR VGND sg13g2_xor2_1
XFILLER_12_78 VPWR VGND sg13g2_fill_1
Xhold161 mac1.products_ff\[144\] VPWR VGND net201 sg13g2_dlygate4sd3_1
Xhold150 mac1.sum_lvl1_ff\[48\] VPWR VGND net190 sg13g2_dlygate4sd3_1
Xhold172 mac1.products_ff\[149\] VPWR VGND net212 sg13g2_dlygate4sd3_1
Xhold183 mac2.products_ff\[79\] VPWR VGND net223 sg13g2_dlygate4sd3_1
Xhold194 mac2.products_ff\[7\] VPWR VGND net234 sg13g2_dlygate4sd3_1
XFILLER_46_514 VPWR VGND sg13g2_fill_1
XFILLER_26_271 VPWR VGND sg13g2_fill_1
XFILLER_18_1017 VPWR VGND sg13g2_decap_8
XFILLER_18_1028 VPWR VGND sg13g2_fill_1
XFILLER_30_904 VPWR VGND sg13g2_decap_8
XFILLER_6_632 VPWR VGND sg13g2_decap_8
XFILLER_6_676 VPWR VGND sg13g2_fill_1
X_5990_ net864 _0238_ VPWR VGND sg13g2_buf_1
X_4941_ _1734_ _1731_ _1733_ VPWR VGND sg13g2_xnor2_1
X_4872_ VGND VPWR _1668_ _1666_ _1641_ sg13g2_or2_1
XFILLER_33_742 VPWR VGND sg13g2_fill_2
XFILLER_33_753 VPWR VGND sg13g2_fill_1
X_3823_ VGND VPWR _0656_ _0657_ _0659_ _0651_ sg13g2_a21oi_1
X_3754_ VPWR _0596_ _0595_ VGND sg13g2_inv_1
X_3685_ VGND VPWR _0530_ _0529_ _0484_ sg13g2_or2_1
X_6473_ net1121 VGND VPWR net237 mac2.sum_lvl2_ff\[26\] clknet_leaf_41_clk sg13g2_dfrbpq_2
X_5424_ net320 mac1.sum_lvl3_ff\[25\] _2180_ VPWR VGND sg13g2_xor2_1
X_5355_ _2126_ mac1.sum_lvl2_ff\[25\] net508 VPWR VGND sg13g2_xnor2_1
X_5286_ _2064_ _2038_ _2065_ VPWR VGND sg13g2_xor2_1
X_4306_ _1111_ VPWR _1123_ VGND _1119_ _1121_ sg13g2_o21ai_1
X_4237_ _1044_ VPWR _1056_ VGND _1052_ _1054_ sg13g2_o21ai_1
X_4168_ _0993_ _0980_ _0992_ VPWR VGND sg13g2_xnor2_1
X_3119_ _2712_ net905 net984 net907 net982 VPWR VGND sg13g2_a22oi_1
X_4099_ _0927_ net926 net991 net928 net989 VPWR VGND sg13g2_a22oi_1
XFILLER_24_753 VPWR VGND sg13g2_fill_2
XFILLER_11_458 VPWR VGND sg13g2_fill_1
XFILLER_20_992 VPWR VGND sg13g2_decap_8
XFILLER_24_1010 VPWR VGND sg13g2_decap_8
XFILLER_47_878 VPWR VGND sg13g2_decap_8
XFILLER_31_1003 VPWR VGND sg13g2_decap_8
XFILLER_11_981 VPWR VGND sg13g2_decap_8
XFILLER_6_495 VPWR VGND sg13g2_fill_2
X_3470_ _0318_ _0292_ _0321_ VPWR VGND sg13g2_xor2_1
X_5140_ _1922_ _1877_ _0158_ VPWR VGND sg13g2_xor2_1
X_5071_ net813 net806 net855 net853 _1856_ VPWR VGND sg13g2_and4_1
X_4022_ _0841_ VPWR _0852_ VGND _0825_ _0842_ sg13g2_o21ai_1
XFILLER_38_856 VPWR VGND sg13g2_decap_8
X_5973_ net272 _0213_ VPWR VGND sg13g2_buf_1
X_4924_ _1718_ net834 net1029 VPWR VGND sg13g2_nand2_1
X_4855_ _1650_ _1629_ _1652_ VPWR VGND sg13g2_xor2_1
X_3806_ _0643_ _0634_ _0641_ VPWR VGND sg13g2_xnor2_1
X_4786_ _1584_ _1567_ _1585_ VPWR VGND sg13g2_xor2_1
X_3737_ _0579_ _0553_ _0580_ VPWR VGND sg13g2_xor2_1
X_3668_ _0511_ _0513_ _0514_ VPWR VGND sg13g2_nor2_1
X_6456_ net1104 VGND VPWR net153 mac2.sum_lvl2_ff\[6\] clknet_leaf_44_clk sg13g2_dfrbpq_1
X_5407_ mac1.sum_lvl3_ff\[21\] mac1.sum_lvl3_ff\[1\] _2167_ VPWR VGND sg13g2_nor2_1
X_3599_ _0446_ net1014 net944 VPWR VGND sg13g2_nand2_1
X_6387_ net1103 VGND VPWR _0134_ mac2.products_ff\[74\] clknet_leaf_42_clk sg13g2_dfrbpq_1
X_5338_ _2110_ VPWR _2113_ VGND _2109_ _2111_ sg13g2_o21ai_1
X_5269_ VGND VPWR _2009_ _2020_ _2049_ _2008_ sg13g2_a21oi_1
XFILLER_16_506 VPWR VGND sg13g2_decap_4
XFILLER_16_528 VPWR VGND sg13g2_decap_8
XFILLER_34_54 VPWR VGND sg13g2_fill_1
XFILLER_11_244 VPWR VGND sg13g2_fill_1
XFILLER_7_248 VPWR VGND sg13g2_fill_2
XFILLER_4_944 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_fill_2
XFILLER_3_465 VPWR VGND sg13g2_fill_1
X_4640_ _1442_ net902 DP_4.matrix\[5\] VPWR VGND sg13g2_nand2_1
X_6310_ net1051 VGND VPWR net79 mac1.sum_lvl3_ff\[29\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_4571_ VGND VPWR _1376_ _1371_ _1369_ sg13g2_or2_1
X_3522_ net961 net957 net1007 net1006 _0371_ VPWR VGND sg13g2_and4_1
X_3453_ net963 net958 net1011 net1009 _0304_ VPWR VGND sg13g2_and4_1
X_6241_ net1066 VGND VPWR net249 mac1.sum_lvl2_ff\[42\] clknet_leaf_64_clk sg13g2_dfrbpq_1
X_6172_ net1101 VGND VPWR _0251_ DP_4.matrix\[7\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_3384_ _2968_ _2955_ _2970_ VPWR VGND sg13g2_xor2_1
XFILLER_34_0 VPWR VGND sg13g2_fill_2
X_5123_ _1896_ _1904_ _1906_ _1907_ VPWR VGND sg13g2_or3_1
X_5054_ _1831_ VPWR _1839_ VGND _1811_ _1832_ sg13g2_o21ai_1
X_4005_ _0836_ net1035 net937 net986 net935 VPWR VGND sg13g2_a22oi_1
X_5956_ net273 _0188_ VPWR VGND sg13g2_buf_1
XFILLER_34_881 VPWR VGND sg13g2_decap_8
X_4907_ _1702_ _1675_ _1700_ VPWR VGND sg13g2_xnor2_1
X_5887_ VGND VPWR net772 _2567_ _0199_ _2566_ sg13g2_a21oi_1
X_4838_ _1635_ _1609_ _1633_ VPWR VGND sg13g2_xnor2_1
XFILLER_21_597 VPWR VGND sg13g2_fill_1
X_4769_ _1534_ VPWR _1568_ VGND _1525_ _1535_ sg13g2_o21ai_1
X_6508_ net1044 VGND VPWR net445 mac2.total_sum\[10\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_1_903 VPWR VGND sg13g2_decap_8
X_6439_ net1125 VGND VPWR net188 mac2.sum_lvl1_ff\[46\] clknet_leaf_39_clk sg13g2_dfrbpq_1
XFILLER_49_929 VPWR VGND sg13g2_decap_8
Xhold10 mac1.sum_lvl1_ff\[8\] VPWR VGND net50 sg13g2_dlygate4sd3_1
Xhold32 mac1.sum_lvl2_ff\[40\] VPWR VGND net72 sg13g2_dlygate4sd3_1
Xhold21 mac2.sum_lvl1_ff\[7\] VPWR VGND net61 sg13g2_dlygate4sd3_1
Xhold43 mac1.sum_lvl1_ff\[81\] VPWR VGND net83 sg13g2_dlygate4sd3_1
Xhold54 mac2.sum_lvl2_ff\[43\] VPWR VGND net94 sg13g2_dlygate4sd3_1
Xhold65 mac2.products_ff\[149\] VPWR VGND net105 sg13g2_dlygate4sd3_1
Xhold76 mac1.products_ff\[8\] VPWR VGND net116 sg13g2_dlygate4sd3_1
Xhold87 mac1.products_ff\[3\] VPWR VGND net127 sg13g2_dlygate4sd3_1
XFILLER_21_1013 VPWR VGND sg13g2_decap_8
Xhold98 mac2.products_ff\[2\] VPWR VGND net138 sg13g2_dlygate4sd3_1
XFILLER_43_133 VPWR VGND sg13g2_fill_2
XFILLER_43_155 VPWR VGND sg13g2_fill_2
XFILLER_12_564 VPWR VGND sg13g2_fill_1
XFILLER_40_840 VPWR VGND sg13g2_decap_8
Xfanout1030 DP_2.matrix\[80\] net1030 VPWR VGND sg13g2_buf_8
XFILLER_48_940 VPWR VGND sg13g2_decap_8
Xfanout1041 net1043 net1041 VPWR VGND sg13g2_buf_8
Xfanout1052 net1053 net1052 VPWR VGND sg13g2_buf_8
Xfanout1074 net1075 net1074 VPWR VGND sg13g2_buf_1
Xfanout1063 net1091 net1063 VPWR VGND sg13g2_buf_8
XFILLER_39_439 VPWR VGND sg13g2_fill_2
Xfanout1096 net1098 net1096 VPWR VGND sg13g2_buf_8
Xfanout1085 net1086 net1085 VPWR VGND sg13g2_buf_8
XFILLER_47_494 VPWR VGND sg13g2_fill_2
X_5810_ VGND VPWR _2504_ _2503_ _2501_ sg13g2_or2_1
X_5741_ _2435_ VPWR _2436_ VGND net384 net791 sg13g2_o21ai_1
XFILLER_22_328 VPWR VGND sg13g2_fill_1
X_5672_ _2374_ _2367_ _2371_ VPWR VGND sg13g2_nand2_1
XFILLER_31_884 VPWR VGND sg13g2_decap_8
X_4623_ _1415_ _1423_ _1425_ _1426_ VPWR VGND sg13g2_or3_1
Xhold502 mac2.sum_lvl2_ff\[14\] VPWR VGND net542 sg13g2_dlygate4sd3_1
X_4554_ _1363_ _1360_ _1362_ VPWR VGND sg13g2_xnor2_1
X_3505_ _0346_ VPWR _0354_ VGND _0326_ _0347_ sg13g2_o21ai_1
X_6224_ net1095 VGND VPWR net171 mac1.sum_lvl2_ff\[22\] clknet_leaf_55_clk sg13g2_dfrbpq_1
X_4485_ _1297_ net873 net816 VPWR VGND sg13g2_nand2_1
X_3436_ _0285_ _0284_ _0279_ _0288_ VPWR VGND sg13g2_a21o_1
X_3367_ _2947_ VPWR _2953_ VGND _2924_ _2925_ sg13g2_o21ai_1
X_6155_ net1082 VGND VPWR _0239_ DP_3.matrix\[75\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_6086_ net1067 VGND VPWR _0193_ DP_1.matrix\[77\] clknet_leaf_60_clk sg13g2_dfrbpq_1
X_5106_ _1862_ VPWR _1890_ VGND _1853_ _1863_ sg13g2_o21ai_1
Xheichips25_template_34 VPWR VGND uio_oe[1] sg13g2_tiehi
X_3298_ VGND VPWR _2887_ _2885_ _2841_ sg13g2_or2_1
X_5037_ _1823_ net855 net811 net857 net806 VPWR VGND sg13g2_a22oi_1
XFILLER_39_940 VPWR VGND sg13g2_decap_8
XFILLER_38_483 VPWR VGND sg13g2_decap_8
XFILLER_40_114 VPWR VGND sg13g2_fill_2
X_5939_ _2598_ VPWR _0251_ VGND _2549_ _2599_ sg13g2_o21ai_1
XFILLER_5_505 VPWR VGND sg13g2_fill_1
XFILLER_21_394 VPWR VGND sg13g2_fill_2
Xclkbuf_4_10_0_clk clknet_0_clk clknet_4_10_0_clk VPWR VGND sg13g2_buf_8
Xoutput22 net22 uio_out[5] VPWR VGND sg13g2_buf_1
XFILLER_0_254 VPWR VGND sg13g2_decap_4
XFILLER_0_287 VPWR VGND sg13g2_fill_1
XFILLER_45_910 VPWR VGND sg13g2_decap_8
XFILLER_45_987 VPWR VGND sg13g2_decap_8
XFILLER_13_840 VPWR VGND sg13g2_fill_1
XFILLER_9_844 VPWR VGND sg13g2_fill_1
XFILLER_9_899 VPWR VGND sg13g2_fill_2
X_4270_ _1086_ _1085_ _1076_ _1088_ VPWR VGND sg13g2_a21o_1
X_3221_ _2812_ net913 net967 VPWR VGND sg13g2_nand2_1
X_3152_ _2745_ _2742_ _2744_ VPWR VGND sg13g2_nand2_1
XFILLER_39_214 VPWR VGND sg13g2_fill_1
X_3083_ _0094_ _2650_ _2677_ VPWR VGND sg13g2_xnor2_1
XFILLER_36_943 VPWR VGND sg13g2_decap_8
X_3985_ _0781_ VPWR _0816_ VGND _0778_ _0782_ sg13g2_o21ai_1
X_5724_ _2420_ _2419_ _2415_ VPWR VGND sg13g2_nand2b_1
X_5655_ _2360_ mac1.total_sum\[8\] mac2.total_sum\[8\] VPWR VGND sg13g2_xnor2_1
XFILLER_11_1023 VPWR VGND sg13g2_decap_4
X_4606_ _1400_ VPWR _1409_ VGND _1392_ _1401_ sg13g2_o21ai_1
X_5586_ net425 _2306_ _0062_ VPWR VGND sg13g2_nor2b_1
Xhold310 _0017_ VPWR VGND net350 sg13g2_dlygate4sd3_1
X_4537_ _1346_ _1320_ _1347_ VPWR VGND sg13g2_xor2_1
Xhold343 DP_4.matrix\[44\] VPWR VGND net383 sg13g2_dlygate4sd3_1
Xhold321 mac1.sum_lvl3_ff\[23\] VPWR VGND net361 sg13g2_dlygate4sd3_1
Xhold332 _0009_ VPWR VGND net372 sg13g2_dlygate4sd3_1
Xhold376 DP_3.matrix\[5\] VPWR VGND net416 sg13g2_dlygate4sd3_1
Xhold365 DP_2.matrix\[36\] VPWR VGND net405 sg13g2_dlygate4sd3_1
Xhold354 _0198_ VPWR VGND net394 sg13g2_dlygate4sd3_1
Xhold387 DP_3.matrix\[1\] VPWR VGND net427 sg13g2_dlygate4sd3_1
X_4468_ _1280_ _1258_ _1281_ VPWR VGND sg13g2_nor2b_1
Xfanout834 net835 net834 VPWR VGND sg13g2_buf_8
Xfanout801 DP_4.matrix\[76\] net801 VPWR VGND sg13g2_buf_1
X_3419_ _0271_ _2989_ _0272_ VPWR VGND sg13g2_xor2_1
X_6207_ net1092 VGND VPWR net130 mac1.sum_lvl2_ff\[2\] clknet_leaf_56_clk sg13g2_dfrbpq_1
Xhold398 mac1.sum_lvl3_ff\[15\] VPWR VGND net438 sg13g2_dlygate4sd3_1
Xfanout812 net813 net812 VPWR VGND sg13g2_buf_2
Xfanout823 net319 net823 VPWR VGND sg13g2_buf_8
Xfanout856 net857 net856 VPWR VGND sg13g2_buf_8
Xfanout845 net846 net845 VPWR VGND sg13g2_buf_2
X_6138_ net1097 VGND VPWR net80 mac1.sum_lvl1_ff\[5\] clknet_leaf_55_clk sg13g2_dfrbpq_1
Xfanout867 net293 net867 VPWR VGND sg13g2_buf_8
X_4399_ _1213_ _1196_ _1214_ VPWR VGND sg13g2_xor2_1
Xfanout889 net890 net889 VPWR VGND sg13g2_buf_1
Xfanout878 net326 net878 VPWR VGND sg13g2_buf_8
X_6069_ net1108 VGND VPWR _0180_ DP_1.matrix\[36\] clknet_leaf_51_clk sg13g2_dfrbpq_1
XFILLER_45_228 VPWR VGND sg13g2_fill_1
XFILLER_27_943 VPWR VGND sg13g2_decap_8
XFILLER_26_453 VPWR VGND sg13g2_fill_1
XFILLER_42_968 VPWR VGND sg13g2_decap_8
XFILLER_41_456 VPWR VGND sg13g2_decap_8
XFILLER_9_118 VPWR VGND sg13g2_fill_1
XFILLER_6_814 VPWR VGND sg13g2_fill_2
XFILLER_6_869 VPWR VGND sg13g2_fill_1
XFILLER_49_556 VPWR VGND sg13g2_decap_4
XFILLER_49_534 VPWR VGND sg13g2_decap_8
XFILLER_18_954 VPWR VGND sg13g2_decap_8
XFILLER_33_968 VPWR VGND sg13g2_decap_8
X_3770_ _0610_ _0600_ _0612_ VPWR VGND sg13g2_xor2_1
XFILLER_9_641 VPWR VGND sg13g2_decap_8
XFILLER_9_685 VPWR VGND sg13g2_fill_2
XFILLER_8_162 VPWR VGND sg13g2_fill_2
X_5440_ _2188_ _2191_ net420 _2193_ VPWR VGND sg13g2_nand3_1
X_5371_ VGND VPWR _2139_ net434 mac1.sum_lvl2_ff\[28\] sg13g2_or2_1
X_4322_ _1138_ net887 net1022 VPWR VGND sg13g2_nand2_1
XFILLER_4_390 VPWR VGND sg13g2_fill_2
X_4253_ _1071_ net884 net818 VPWR VGND sg13g2_nand2_1
X_3204_ _2791_ VPWR _2795_ VGND _2748_ _2793_ sg13g2_o21ai_1
X_4184_ VGND VPWR _1005_ _1000_ _0998_ sg13g2_or2_1
XFILLER_41_1005 VPWR VGND sg13g2_decap_8
X_3135_ net918 net967 net922 _2728_ VPWR VGND net964 sg13g2_nand4_1
X_3066_ net917 net972 net921 _2661_ VPWR VGND net969 sg13g2_nand4_1
XFILLER_24_968 VPWR VGND sg13g2_decap_8
X_3968_ _0776_ VPWR _0800_ VGND _0796_ _0798_ sg13g2_o21ai_1
X_5707_ _2402_ VPWR _2403_ VGND net403 net791 sg13g2_o21ai_1
X_3899_ _0732_ _0727_ _0730_ VPWR VGND sg13g2_xnor2_1
X_5638_ mac2.total_sum\[4\] mac1.total_sum\[4\] _2347_ VPWR VGND sg13g2_xor2_1
X_5569_ mac2.sum_lvl3_ff\[25\] net396 _2293_ VPWR VGND sg13g2_nor2_1
Xhold162 mac1.products_ff\[70\] VPWR VGND net202 sg13g2_dlygate4sd3_1
Xhold140 mac1.sum_lvl1_ff\[84\] VPWR VGND net180 sg13g2_dlygate4sd3_1
Xhold151 mac2.products_ff\[141\] VPWR VGND net191 sg13g2_dlygate4sd3_1
Xhold195 mac2.sum_lvl1_ff\[87\] VPWR VGND net235 sg13g2_dlygate4sd3_1
Xhold184 mac1.products_ff\[76\] VPWR VGND net224 sg13g2_dlygate4sd3_1
Xhold173 mac1.products_ff\[13\] VPWR VGND net213 sg13g2_dlygate4sd3_1
XFILLER_46_537 VPWR VGND sg13g2_fill_1
XFILLER_27_751 VPWR VGND sg13g2_decap_4
XFILLER_45_8 VPWR VGND sg13g2_fill_2
XFILLER_49_364 VPWR VGND sg13g2_fill_1
XFILLER_37_537 VPWR VGND sg13g2_decap_8
X_4940_ _1733_ _1717_ _1732_ VPWR VGND sg13g2_xnor2_1
X_4871_ _1641_ _1666_ _1667_ VPWR VGND sg13g2_nor2_1
X_3822_ _0656_ _0657_ _0651_ _0658_ VPWR VGND sg13g2_nand3_1
X_3753_ _0595_ _0571_ _0593_ VPWR VGND sg13g2_nand2_1
X_3684_ _0529_ net1010 net946 VPWR VGND sg13g2_nand2_1
X_6472_ net1119 VGND VPWR net226 mac2.sum_lvl2_ff\[25\] clknet_leaf_42_clk sg13g2_dfrbpq_2
X_5423_ mac1.sum_lvl3_ff\[25\] net320 _2179_ VPWR VGND sg13g2_nor2_1
X_5354_ mac1.sum_lvl2_ff\[25\] net508 _2125_ VPWR VGND sg13g2_and2_1
X_4305_ _1111_ _1119_ _1121_ _1122_ VPWR VGND sg13g2_or3_1
X_5285_ _2064_ net796 net852 VPWR VGND sg13g2_nand2_1
X_4236_ _1044_ _1052_ _1054_ _1055_ VPWR VGND sg13g2_or3_1
X_4167_ _0992_ _0989_ _0991_ VPWR VGND sg13g2_xnor2_1
X_3118_ _2688_ VPWR _2711_ VGND _2653_ _2686_ sg13g2_o21ai_1
X_4098_ VGND VPWR _0926_ _0924_ _0899_ sg13g2_or2_1
X_3049_ _2645_ _2642_ _2644_ VPWR VGND sg13g2_nand2_1
XFILLER_36_570 VPWR VGND sg13g2_fill_1
XFILLER_20_971 VPWR VGND sg13g2_decap_8
XFILLER_48_97 VPWR VGND sg13g2_fill_1
XFILLER_9_14 VPWR VGND sg13g2_fill_2
XFILLER_14_264 VPWR VGND sg13g2_fill_1
XFILLER_11_960 VPWR VGND sg13g2_decap_8
XFILLER_7_997 VPWR VGND sg13g2_decap_8
X_5070_ _1855_ net804 net856 VPWR VGND sg13g2_nand2_1
X_4021_ VGND VPWR _0816_ _0822_ _0851_ _0824_ sg13g2_a21oi_1
XFILLER_49_183 VPWR VGND sg13g2_fill_1
XFILLER_37_323 VPWR VGND sg13g2_fill_1
XFILLER_38_835 VPWR VGND sg13g2_decap_8
X_5972_ net924 _0212_ VPWR VGND sg13g2_buf_1
X_4923_ _1717_ net833 net1029 VPWR VGND sg13g2_nand2_1
X_4854_ _1650_ _1629_ _1651_ VPWR VGND sg13g2_nor2b_1
XFILLER_20_212 VPWR VGND sg13g2_fill_1
X_3805_ _0642_ _0634_ _0641_ VPWR VGND sg13g2_nand2_1
X_4785_ _1584_ _1568_ _1582_ VPWR VGND sg13g2_xnor2_1
X_3736_ _0579_ net947 net1005 VPWR VGND sg13g2_nand2_1
X_3667_ VGND VPWR _0512_ _0513_ _0478_ _0438_ sg13g2_a21oi_2
X_6455_ net1102 VGND VPWR net109 mac2.sum_lvl2_ff\[5\] clknet_leaf_30_clk sg13g2_dfrbpq_1
XFILLER_47_1011 VPWR VGND sg13g2_decap_8
X_5406_ _2166_ mac1.sum_lvl3_ff\[21\] mac1.sum_lvl3_ff\[1\] VPWR VGND sg13g2_nand2_1
X_3598_ _0445_ DP_1.matrix\[1\] net1032 VPWR VGND sg13g2_nand2_1
X_6386_ net1102 VGND VPWR _0127_ mac2.products_ff\[73\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_5337_ _0007_ _2109_ _2112_ VPWR VGND sg13g2_xnor2_1
XFILLER_0_606 VPWR VGND sg13g2_fill_1
X_5268_ _2046_ _2034_ _2048_ VPWR VGND sg13g2_xor2_1
X_4219_ _1029_ VPWR _1038_ VGND _1021_ _1030_ sg13g2_o21ai_1
X_5199_ net802 net801 net854 net851 _1981_ VPWR VGND sg13g2_and4_1
XFILLER_34_44 VPWR VGND sg13g2_fill_1
XFILLER_4_923 VPWR VGND sg13g2_fill_1
XFILLER_19_389 VPWR VGND sg13g2_decap_8
X_4570_ _1375_ net903 net839 VPWR VGND sg13g2_nand2_1
X_3521_ _0370_ net954 net1009 VPWR VGND sg13g2_nand2_1
XFILLER_6_271 VPWR VGND sg13g2_fill_1
X_3452_ _0303_ net954 net1014 VPWR VGND sg13g2_nand2_1
X_6240_ net1050 VGND VPWR net93 mac1.sum_lvl2_ff\[41\] clknet_leaf_66_clk sg13g2_dfrbpq_1
X_6171_ net1101 VGND VPWR _0250_ DP_4.matrix\[6\] clknet_leaf_26_clk sg13g2_dfrbpq_1
X_3383_ VGND VPWR _2969_ _2968_ _2955_ sg13g2_or2_1
X_5122_ VGND VPWR _1902_ _1903_ _1906_ _1897_ sg13g2_a21oi_1
X_5053_ _1838_ _1837_ _0156_ VPWR VGND sg13g2_xor2_1
X_4004_ net937 net935 net986 net1035 _0835_ VPWR VGND sg13g2_and4_1
XFILLER_38_687 VPWR VGND sg13g2_fill_1
XFILLER_37_186 VPWR VGND sg13g2_fill_2
X_5955_ net278 _0187_ VPWR VGND sg13g2_buf_1
XFILLER_34_860 VPWR VGND sg13g2_decap_8
X_4906_ _1701_ _1700_ _1675_ VPWR VGND sg13g2_nand2b_1
X_5886_ _2567_ _2445_ _2455_ VPWR VGND sg13g2_xnor2_1
XFILLER_21_510 VPWR VGND sg13g2_fill_1
X_4837_ VGND VPWR _1634_ _1633_ _1609_ sg13g2_or2_1
X_4768_ _1567_ _1557_ _1565_ VPWR VGND sg13g2_xnor2_1
X_6507_ net1044 VGND VPWR net430 mac2.total_sum\[9\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_3719_ _0561_ _0549_ _0563_ VPWR VGND sg13g2_xor2_1
X_4699_ _1498_ _1499_ _1468_ _1500_ VPWR VGND sg13g2_nand3_1
X_6438_ net1119 VGND VPWR net225 mac2.sum_lvl1_ff\[45\] clknet_leaf_40_clk sg13g2_dfrbpq_1
XFILLER_49_908 VPWR VGND sg13g2_decap_8
XFILLER_1_959 VPWR VGND sg13g2_decap_8
X_6369_ net1099 VGND VPWR _0088_ mac2.products_ff\[4\] clknet_leaf_29_clk sg13g2_dfrbpq_1
Xhold22 mac2.products_ff\[12\] VPWR VGND net62 sg13g2_dlygate4sd3_1
XFILLER_0_447 VPWR VGND sg13g2_fill_2
Xhold11 mac2.products_ff\[1\] VPWR VGND net51 sg13g2_dlygate4sd3_1
Xhold44 mac1.sum_lvl2_ff\[49\] VPWR VGND net84 sg13g2_dlygate4sd3_1
Xhold55 mac1.sum_lvl1_ff\[12\] VPWR VGND net95 sg13g2_dlygate4sd3_1
Xhold33 mac2.sum_lvl1_ff\[39\] VPWR VGND net73 sg13g2_dlygate4sd3_1
Xhold66 mac1.sum_lvl1_ff\[38\] VPWR VGND net106 sg13g2_dlygate4sd3_1
Xhold88 mac2.sum_lvl2_ff\[45\] VPWR VGND net128 sg13g2_dlygate4sd3_1
Xhold77 mac2.sum_lvl1_ff\[80\] VPWR VGND net117 sg13g2_dlygate4sd3_1
Xhold99 mac2.products_ff\[142\] VPWR VGND net139 sg13g2_dlygate4sd3_1
XFILLER_29_632 VPWR VGND sg13g2_decap_8
XFILLER_17_838 VPWR VGND sg13g2_fill_1
XFILLER_43_123 VPWR VGND sg13g2_fill_2
XFILLER_31_329 VPWR VGND sg13g2_fill_2
XFILLER_40_896 VPWR VGND sg13g2_decap_8
XFILLER_4_753 VPWR VGND sg13g2_fill_1
XFILLER_4_731 VPWR VGND sg13g2_fill_1
Xfanout1020 DP_1.matrix\[0\] net1020 VPWR VGND sg13g2_buf_1
Xfanout1031 net384 net1031 VPWR VGND sg13g2_buf_8
Xfanout1042 net1043 net1042 VPWR VGND sg13g2_buf_1
Xfanout1064 net1065 net1064 VPWR VGND sg13g2_buf_8
Xfanout1053 net1055 net1053 VPWR VGND sg13g2_buf_8
Xfanout1097 net1098 net1097 VPWR VGND sg13g2_buf_8
Xfanout1075 net1076 net1075 VPWR VGND sg13g2_buf_8
Xfanout1086 net1090 net1086 VPWR VGND sg13g2_buf_8
XFILLER_48_996 VPWR VGND sg13g2_decap_8
XFILLER_47_473 VPWR VGND sg13g2_fill_2
XFILLER_19_142 VPWR VGND sg13g2_fill_1
X_5740_ VPWR _2435_ _2434_ VGND sg13g2_inv_1
XFILLER_31_863 VPWR VGND sg13g2_decap_8
X_5671_ _2373_ mac1.total_sum\[11\] mac2.total_sum\[11\] VPWR VGND sg13g2_xnor2_1
X_4622_ VGND VPWR _1421_ _1422_ _1425_ _1416_ sg13g2_a21oi_1
X_4553_ _1362_ _1345_ _1361_ VPWR VGND sg13g2_xnor2_1
Xhold503 _2276_ VPWR VGND net543 sg13g2_dlygate4sd3_1
X_4484_ _1296_ net873 net814 VPWR VGND sg13g2_nand2_1
XFILLER_7_591 VPWR VGND sg13g2_decap_4
X_3504_ _0353_ _0352_ _0112_ VPWR VGND sg13g2_xor2_1
X_3435_ VGND VPWR _0284_ _0285_ _0287_ _0279_ sg13g2_a21oi_1
X_6223_ net1092 VGND VPWR net106 mac1.sum_lvl2_ff\[21\] clknet_leaf_56_clk sg13g2_dfrbpq_1
XFILLER_44_1014 VPWR VGND sg13g2_decap_8
X_3366_ VPWR _2952_ _2951_ VGND sg13g2_inv_1
X_6154_ net1081 VGND VPWR _0238_ DP_3.matrix\[74\] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_6085_ net1067 VGND VPWR _0192_ DP_1.matrix\[76\] clknet_leaf_60_clk sg13g2_dfrbpq_1
X_3297_ _2886_ net970 net907 VPWR VGND sg13g2_nand2_1
X_5105_ _1889_ _1842_ _1888_ VPWR VGND sg13g2_xnor2_1
Xheichips25_template_35 VPWR VGND uio_oe[2] sg13g2_tiehi
X_5036_ net806 net856 net811 _1822_ VPWR VGND net855 sg13g2_nand4_1
XFILLER_38_451 VPWR VGND sg13g2_decap_4
XFILLER_39_996 VPWR VGND sg13g2_decap_8
XFILLER_25_112 VPWR VGND sg13g2_fill_1
X_5938_ _2545_ _2547_ _2599_ VPWR VGND sg13g2_nor2b_1
XFILLER_41_627 VPWR VGND sg13g2_fill_1
XFILLER_15_68 VPWR VGND sg13g2_fill_2
XFILLER_40_137 VPWR VGND sg13g2_fill_2
X_5869_ _2557_ _2424_ _2426_ VPWR VGND sg13g2_xnor2_1
Xoutput23 net23 uio_out[6] VPWR VGND sg13g2_buf_1
XFILLER_17_613 VPWR VGND sg13g2_decap_4
XFILLER_45_966 VPWR VGND sg13g2_decap_8
XFILLER_44_465 VPWR VGND sg13g2_fill_1
XFILLER_44_498 VPWR VGND sg13g2_decap_4
XFILLER_13_885 VPWR VGND sg13g2_fill_2
X_3220_ _2811_ net972 net909 VPWR VGND sg13g2_nand2_1
X_3151_ _2741_ _2740_ _2710_ _2744_ VPWR VGND sg13g2_a21o_1
X_3082_ _2674_ _2648_ _2677_ VPWR VGND sg13g2_xor2_1
XFILLER_36_922 VPWR VGND sg13g2_decap_8
XFILLER_35_421 VPWR VGND sg13g2_fill_1
XFILLER_36_999 VPWR VGND sg13g2_decap_8
X_3984_ _0769_ _0772_ _0815_ VPWR VGND sg13g2_nor2_1
XFILLER_22_126 VPWR VGND sg13g2_fill_2
X_5723_ _2419_ _2417_ _2418_ _2416_ net782 VPWR VGND sg13g2_a22oi_1
X_5654_ _2358_ _2359_ net32 VPWR VGND sg13g2_and2_1
XFILLER_11_1002 VPWR VGND sg13g2_decap_8
X_4605_ _1407_ _1387_ _0088_ VPWR VGND sg13g2_xor2_1
Xhold311 DP_3.matrix\[75\] VPWR VGND net351 sg13g2_dlygate4sd3_1
Xhold300 DP_3.matrix\[41\] VPWR VGND net340 sg13g2_dlygate4sd3_1
X_5585_ _2302_ net424 _2300_ _2306_ VPWR VGND sg13g2_nand3_1
X_4536_ _1346_ net816 net1027 VPWR VGND sg13g2_nand2_1
Xhold322 _2174_ VPWR VGND net362 sg13g2_dlygate4sd3_1
Xhold344 DP_2.matrix\[44\] VPWR VGND net384 sg13g2_dlygate4sd3_1
Xhold333 DP_4.matrix\[36\] VPWR VGND net373 sg13g2_dlygate4sd3_1
Xhold377 _0225_ VPWR VGND net417 sg13g2_dlygate4sd3_1
Xhold355 DP_1.matrix\[36\] VPWR VGND net395 sg13g2_dlygate4sd3_1
Xhold366 mac1.sum_lvl3_ff\[24\] VPWR VGND net406 sg13g2_dlygate4sd3_1
X_4467_ _1280_ _1259_ _1279_ VPWR VGND sg13g2_xnor2_1
Xhold388 DP_3.matrix\[6\] VPWR VGND net428 sg13g2_dlygate4sd3_1
Xfanout802 net803 net802 VPWR VGND sg13g2_buf_8
X_3418_ _0271_ _2990_ _0269_ VPWR VGND sg13g2_xnor2_1
X_6206_ net1070 VGND VPWR net148 mac1.sum_lvl2_ff\[1\] clknet_leaf_62_clk sg13g2_dfrbpq_1
Xhold399 _2222_ VPWR VGND net439 sg13g2_dlygate4sd3_1
X_4398_ _1213_ _1197_ _1211_ VPWR VGND sg13g2_xnor2_1
Xfanout824 DP_4.matrix\[38\] net824 VPWR VGND sg13g2_buf_1
Xfanout813 net282 net813 VPWR VGND sg13g2_buf_2
Xfanout835 net386 net835 VPWR VGND sg13g2_buf_8
X_6137_ net1101 VGND VPWR _0227_ DP_3.matrix\[7\] clknet_leaf_26_clk sg13g2_dfrbpq_1
Xfanout857 DP_3.matrix\[77\] net857 VPWR VGND sg13g2_buf_8
X_3349_ _2935_ _2910_ _2936_ VPWR VGND sg13g2_xor2_1
Xfanout846 DP_4.matrix\[1\] net846 VPWR VGND sg13g2_buf_2
Xfanout868 net869 net868 VPWR VGND sg13g2_buf_8
Xfanout879 DP_3.matrix\[40\] net879 VPWR VGND sg13g2_buf_8
X_6068_ net1094 VGND VPWR _0179_ DP_1.matrix\[7\] clknet_leaf_58_clk sg13g2_dfrbpq_2
XFILLER_39_760 VPWR VGND sg13g2_fill_2
XFILLER_27_922 VPWR VGND sg13g2_decap_8
X_5019_ _1803_ _1777_ _1806_ VPWR VGND sg13g2_xor2_1
XFILLER_42_947 VPWR VGND sg13g2_decap_8
XFILLER_27_999 VPWR VGND sg13g2_decap_8
XFILLER_41_424 VPWR VGND sg13g2_fill_2
XFILLER_14_649 VPWR VGND sg13g2_fill_1
XFILLER_41_468 VPWR VGND sg13g2_fill_2
XFILLER_42_33 VPWR VGND sg13g2_fill_2
XFILLER_6_848 VPWR VGND sg13g2_fill_1
XFILLER_5_347 VPWR VGND sg13g2_fill_1
XFILLER_27_1020 VPWR VGND sg13g2_decap_8
XFILLER_1_586 VPWR VGND sg13g2_fill_2
XFILLER_44_262 VPWR VGND sg13g2_fill_1
XFILLER_33_947 VPWR VGND sg13g2_decap_8
XFILLER_32_479 VPWR VGND sg13g2_decap_4
XFILLER_41_991 VPWR VGND sg13g2_decap_8
XFILLER_9_675 VPWR VGND sg13g2_fill_2
X_5370_ mac1.sum_lvl2_ff\[28\] net434 _2138_ VPWR VGND sg13g2_and2_1
X_4321_ _1108_ VPWR _1137_ VGND _1105_ _1109_ sg13g2_o21ai_1
X_4252_ _1053_ VPWR _1070_ VGND _1044_ _1054_ sg13g2_o21ai_1
X_3203_ _2793_ _2748_ _0103_ VPWR VGND sg13g2_xor2_1
X_4183_ _1004_ net886 net822 VPWR VGND sg13g2_nand2_1
XFILLER_41_1028 VPWR VGND sg13g2_fill_1
X_3134_ net921 net918 net967 net964 _2727_ VPWR VGND sg13g2_and4_1
X_3065_ net921 net917 net972 net969 _2660_ VPWR VGND sg13g2_and4_1
XFILLER_24_947 VPWR VGND sg13g2_decap_8
X_3967_ _0776_ _0796_ _0798_ _0799_ VPWR VGND sg13g2_or3_1
X_5706_ VPWR _2402_ _2401_ VGND sg13g2_inv_1
X_3898_ _0731_ _0727_ _0730_ VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_30_clk clknet_4_12_0_clk clknet_leaf_30_clk VPWR VGND sg13g2_buf_8
X_5637_ mac1.total_sum\[4\] mac2.total_sum\[4\] _2346_ VPWR VGND sg13g2_and2_1
X_5568_ VGND VPWR _2289_ _2291_ _2292_ _2290_ sg13g2_a21oi_1
X_4519_ _1330_ _1329_ _1304_ VPWR VGND sg13g2_nand2b_1
Xhold141 mac1.products_ff\[68\] VPWR VGND net181 sg13g2_dlygate4sd3_1
Xhold130 mac1.products_ff\[79\] VPWR VGND net170 sg13g2_dlygate4sd3_1
Xhold152 mac2.sum_lvl1_ff\[37\] VPWR VGND net192 sg13g2_dlygate4sd3_1
Xhold163 mac1.sum_lvl1_ff\[78\] VPWR VGND net203 sg13g2_dlygate4sd3_1
X_5499_ _0043_ _2236_ net388 VPWR VGND sg13g2_xnor2_1
Xhold174 mac2.sum_lvl2_ff\[40\] VPWR VGND net214 sg13g2_dlygate4sd3_1
Xhold185 mac2.products_ff\[77\] VPWR VGND net225 sg13g2_dlygate4sd3_1
Xhold196 mac2.sum_lvl2_ff\[51\] VPWR VGND net236 sg13g2_dlygate4sd3_1
XFILLER_2_1022 VPWR VGND sg13g2_decap_8
XFILLER_15_969 VPWR VGND sg13g2_decap_8
XFILLER_30_939 VPWR VGND sg13g2_decap_8
XFILLER_41_265 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_21_clk clknet_4_5_0_clk clknet_leaf_21_clk VPWR VGND sg13g2_buf_8
XFILLER_38_8 VPWR VGND sg13g2_fill_1
XFILLER_37_516 VPWR VGND sg13g2_fill_1
X_4870_ _1666_ net891 net833 VPWR VGND sg13g2_nand2_2
X_3821_ _0652_ VPWR _0657_ VGND _0653_ _0655_ sg13g2_o21ai_1
XFILLER_14_991 VPWR VGND sg13g2_decap_8
X_3752_ _0109_ _0593_ _0594_ VPWR VGND sg13g2_xnor2_1
Xclkbuf_leaf_12_clk clknet_4_12_0_clk clknet_leaf_12_clk VPWR VGND sg13g2_buf_8
X_3683_ _0528_ net1014 net1032 VPWR VGND sg13g2_nand2_1
X_6471_ net1103 VGND VPWR net252 mac2.sum_lvl2_ff\[24\] clknet_leaf_43_clk sg13g2_dfrbpq_2
X_5422_ VGND VPWR _2175_ _2177_ _2178_ _2176_ sg13g2_a21oi_1
X_5353_ _0011_ _2122_ net506 VPWR VGND sg13g2_xnor2_1
X_4304_ VGND VPWR _1117_ _1118_ _1121_ _1112_ sg13g2_a21oi_1
X_5284_ _2063_ net851 net792 VPWR VGND sg13g2_nand2_1
X_4235_ VGND VPWR _1050_ _1051_ _1054_ _1045_ sg13g2_a21oi_1
X_4166_ _0991_ _0975_ _0990_ VPWR VGND sg13g2_xnor2_1
X_3117_ _2702_ VPWR _2710_ VGND _2682_ _2703_ sg13g2_o21ai_1
X_4097_ _0899_ _0924_ _0925_ VPWR VGND sg13g2_nor2_1
X_3048_ _2641_ _2640_ _2635_ _2644_ VPWR VGND sg13g2_a21o_1
XFILLER_24_755 VPWR VGND sg13g2_fill_1
XFILLER_23_46 VPWR VGND sg13g2_fill_1
X_4999_ _1784_ _1781_ _1786_ VPWR VGND sg13g2_xor2_1
XFILLER_7_409 VPWR VGND sg13g2_fill_2
XFILLER_20_950 VPWR VGND sg13g2_decap_8
XFILLER_3_626 VPWR VGND sg13g2_decap_8
XFILLER_3_615 VPWR VGND sg13g2_fill_2
XFILLER_48_87 VPWR VGND sg13g2_fill_1
XFILLER_14_221 VPWR VGND sg13g2_fill_2
XFILLER_42_574 VPWR VGND sg13g2_decap_8
XFILLER_7_976 VPWR VGND sg13g2_decap_8
XFILLER_9_1028 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_1_clk clknet_4_0_0_clk clknet_leaf_1_clk VPWR VGND sg13g2_buf_8
X_4020_ _0850_ _0811_ _0126_ VPWR VGND sg13g2_xor2_1
XFILLER_46_880 VPWR VGND sg13g2_decap_8
X_5971_ net281 _0211_ VPWR VGND sg13g2_buf_1
X_4922_ _1716_ net892 DP_4.matrix\[8\] VPWR VGND sg13g2_nand2_1
X_4853_ _1650_ _1630_ _1649_ VPWR VGND sg13g2_xnor2_1
X_3804_ _0639_ _0640_ _0641_ VPWR VGND sg13g2_nor2b_1
X_4784_ _1583_ _1568_ _1582_ VPWR VGND sg13g2_nand2_1
X_6523_ net1057 VGND VPWR net16 DP_3.I_range.out_data\[6\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_3735_ _0578_ net1005 net944 VPWR VGND sg13g2_nand2_1
X_6454_ net1100 VGND VPWR net85 mac2.sum_lvl2_ff\[4\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_5405_ _2165_ net288 net265 VPWR VGND sg13g2_nand2_1
X_3666_ VGND VPWR _0435_ _0477_ _0512_ _0476_ sg13g2_a21oi_1
X_3597_ _0409_ VPWR _0444_ VGND _0406_ _0410_ sg13g2_o21ai_1
X_6385_ net1100 VGND VPWR _0083_ mac2.products_ff\[72\] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_5336_ mac1.sum_lvl2_ff\[1\] mac1.sum_lvl2_ff\[20\] _2112_ VPWR VGND sg13g2_xor2_1
X_5267_ VGND VPWR _2047_ _2046_ _2034_ sg13g2_or2_1
X_4218_ _1036_ _1016_ _0083_ VPWR VGND sg13g2_xor2_1
X_5198_ _1980_ net800 net852 VPWR VGND sg13g2_nand2_1
X_4149_ _0975_ net926 net1035 VPWR VGND sg13g2_nand2_1
XFILLER_29_869 VPWR VGND sg13g2_decap_8
XFILLER_43_338 VPWR VGND sg13g2_fill_1
XFILLER_43_327 VPWR VGND sg13g2_fill_2
XFILLER_8_707 VPWR VGND sg13g2_fill_1
Xclkload0 clknet_4_1_0_clk clkload0/X VPWR VGND sg13g2_buf_8
XFILLER_4_979 VPWR VGND sg13g2_decap_8
XFILLER_1_2 VPWR VGND sg13g2_fill_1
XFILLER_19_357 VPWR VGND sg13g2_decap_8
XFILLER_35_839 VPWR VGND sg13g2_decap_8
XFILLER_28_880 VPWR VGND sg13g2_decap_8
XFILLER_43_883 VPWR VGND sg13g2_decap_8
X_3520_ _0337_ VPWR _0369_ VGND _0335_ _0338_ sg13g2_o21ai_1
X_3451_ _0282_ VPWR _0302_ VGND _0280_ _0283_ sg13g2_o21ai_1
X_6170_ net1089 VGND VPWR _0249_ DP_4.matrix\[5\] clknet_leaf_26_clk sg13g2_dfrbpq_2
X_3382_ _2966_ _2956_ _2968_ VPWR VGND sg13g2_xor2_1
X_5121_ _1902_ _1903_ _1897_ _1905_ VPWR VGND sg13g2_nand3_1
X_5052_ _1804_ VPWR _1838_ VGND _1779_ _1805_ sg13g2_o21ai_1
X_4003_ _0834_ net935 net1035 VPWR VGND sg13g2_nand2_1
XFILLER_37_132 VPWR VGND sg13g2_fill_2
X_5954_ net990 _0186_ VPWR VGND sg13g2_buf_1
X_4905_ _1698_ _1660_ _1700_ VPWR VGND sg13g2_xor2_1
X_5885_ net952 net772 _2566_ VPWR VGND sg13g2_nor2_1
X_4836_ _1633_ net840 net1028 VPWR VGND sg13g2_nand2_1
X_6506_ net1044 VGND VPWR net426 mac2.total_sum\[8\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_4767_ _1557_ _1565_ _1566_ VPWR VGND sg13g2_nor2_1
X_3718_ VGND VPWR _0562_ _0561_ _0549_ sg13g2_or2_1
X_4698_ _1474_ VPWR _1499_ VGND _1495_ _1497_ sg13g2_o21ai_1
X_3649_ _0495_ net950 DP_1.matrix\[7\] VPWR VGND sg13g2_nand2_1
X_6437_ net1120 VGND VPWR net98 mac2.sum_lvl1_ff\[44\] clknet_leaf_41_clk sg13g2_dfrbpq_1
X_6368_ net1085 VGND VPWR _0087_ mac2.products_ff\[3\] clknet_leaf_29_clk sg13g2_dfrbpq_1
X_5319_ _2095_ _2085_ _2097_ VPWR VGND sg13g2_xor2_1
XFILLER_1_938 VPWR VGND sg13g2_decap_8
X_6299_ net1057 VGND VPWR net173 mac2.sum_lvl1_ff\[86\] clknet_leaf_23_clk sg13g2_dfrbpq_1
Xhold23 mac2.sum_lvl1_ff\[38\] VPWR VGND net63 sg13g2_dlygate4sd3_1
Xhold12 mac2.sum_lvl1_ff\[10\] VPWR VGND net52 sg13g2_dlygate4sd3_1
Xhold45 mac2.sum_lvl1_ff\[4\] VPWR VGND net85 sg13g2_dlygate4sd3_1
Xhold56 mac2.products_ff\[6\] VPWR VGND net96 sg13g2_dlygate4sd3_1
Xhold34 mac2.products_ff\[136\] VPWR VGND net74 sg13g2_dlygate4sd3_1
Xhold67 mac1.sum_lvl2_ff\[38\] VPWR VGND net107 sg13g2_dlygate4sd3_1
Xhold78 mac1.sum_lvl1_ff\[4\] VPWR VGND net118 sg13g2_dlygate4sd3_1
Xhold89 mac2.sum_lvl2_ff\[50\] VPWR VGND net129 sg13g2_dlygate4sd3_1
XFILLER_17_817 VPWR VGND sg13g2_fill_1
XFILLER_43_168 VPWR VGND sg13g2_fill_2
XFILLER_43_135 VPWR VGND sg13g2_fill_1
XFILLER_40_875 VPWR VGND sg13g2_decap_8
Xfanout1021 DP_4.matrix\[80\] net1021 VPWR VGND sg13g2_buf_8
Xfanout1010 net448 net1010 VPWR VGND sg13g2_buf_8
Xfanout1065 net1069 net1065 VPWR VGND sg13g2_buf_8
XFILLER_0_982 VPWR VGND sg13g2_decap_8
Xfanout1043 net1048 net1043 VPWR VGND sg13g2_buf_8
Xfanout1032 net535 net1032 VPWR VGND sg13g2_buf_8
Xfanout1054 net1055 net1054 VPWR VGND sg13g2_buf_8
Xfanout1087 net1088 net1087 VPWR VGND sg13g2_buf_8
Xfanout1076 net1091 net1076 VPWR VGND sg13g2_buf_8
Xfanout1098 net1107 net1098 VPWR VGND sg13g2_buf_8
XFILLER_48_975 VPWR VGND sg13g2_decap_8
XFILLER_47_452 VPWR VGND sg13g2_fill_1
XFILLER_47_496 VPWR VGND sg13g2_fill_1
XFILLER_34_146 VPWR VGND sg13g2_fill_2
XFILLER_34_157 VPWR VGND sg13g2_fill_2
XFILLER_34_179 VPWR VGND sg13g2_fill_1
X_5670_ mac1.total_sum\[11\] mac2.total_sum\[11\] _2372_ VPWR VGND sg13g2_nor2_1
XFILLER_31_842 VPWR VGND sg13g2_decap_8
X_4621_ _1421_ _1422_ _1416_ _1424_ VPWR VGND sg13g2_nand3_1
X_4552_ _1361_ net870 DP_4.matrix\[44\] VPWR VGND sg13g2_nand2_1
X_4483_ _1295_ net879 net1022 VPWR VGND sg13g2_nand2_1
X_3503_ _0319_ VPWR _0353_ VGND _0294_ _0320_ sg13g2_o21ai_1
Xhold504 DP_1.matrix\[41\] VPWR VGND net544 sg13g2_dlygate4sd3_1
X_3434_ _0284_ _0285_ _0279_ _0286_ VPWR VGND sg13g2_nand3_1
X_6222_ net1070 VGND VPWR net149 mac1.sum_lvl2_ff\[20\] clknet_leaf_62_clk sg13g2_dfrbpq_1
X_3365_ _2951_ _2927_ _2949_ VPWR VGND sg13g2_nand2_1
X_6153_ net1110 VGND VPWR net142 mac1.sum_lvl1_ff\[10\] clknet_leaf_45_clk sg13g2_dfrbpq_1
X_6084_ net1050 VGND VPWR _0067_ mac1.products_ff\[139\] clknet_leaf_66_clk sg13g2_dfrbpq_1
X_3296_ _2885_ net971 net905 VPWR VGND sg13g2_nand2_1
X_5104_ _1888_ _1879_ _1886_ VPWR VGND sg13g2_xnor2_1
Xheichips25_template_36 VPWR VGND uio_oe[3] sg13g2_tiehi
X_5035_ net811 net806 net856 net855 _1821_ VPWR VGND sg13g2_and4_1
XFILLER_39_975 VPWR VGND sg13g2_decap_8
X_5937_ _2598_ net832 net767 VPWR VGND sg13g2_nand2_1
XFILLER_22_831 VPWR VGND sg13g2_fill_2
X_5868_ net1011 net772 _2556_ VPWR VGND sg13g2_nor2_1
X_4819_ _1615_ _1606_ _1617_ VPWR VGND sg13g2_xor2_1
XFILLER_21_396 VPWR VGND sg13g2_fill_1
X_5799_ _2493_ _2469_ net786 VPWR VGND sg13g2_nand2_1
XFILLER_31_79 VPWR VGND sg13g2_fill_2
Xoutput24 net24 uio_out[7] VPWR VGND sg13g2_buf_1
XFILLER_29_463 VPWR VGND sg13g2_decap_8
XFILLER_45_945 VPWR VGND sg13g2_decap_8
XFILLER_8_312 VPWR VGND sg13g2_fill_2
XFILLER_9_857 VPWR VGND sg13g2_fill_2
XFILLER_8_345 VPWR VGND sg13g2_fill_1
XFILLER_4_584 VPWR VGND sg13g2_fill_2
X_3150_ VGND VPWR _2740_ _2741_ _2743_ _2710_ sg13g2_a21oi_1
X_3081_ VGND VPWR _2672_ _2673_ _2676_ _2648_ sg13g2_a21oi_1
XFILLER_36_901 VPWR VGND sg13g2_decap_8
XFILLER_35_466 VPWR VGND sg13g2_fill_2
XFILLER_36_978 VPWR VGND sg13g2_decap_8
X_5722_ net782 VPWR _2418_ VGND net1002 net790 sg13g2_o21ai_1
X_3983_ _0797_ VPWR _0814_ VGND _0776_ _0798_ sg13g2_o21ai_1
X_5653_ _2351_ _2354_ _2357_ _2359_ VPWR VGND sg13g2_or3_1
X_5584_ VGND VPWR _2300_ _2302_ _2305_ net424 sg13g2_a21oi_1
X_4604_ VGND VPWR _1408_ _1407_ _1387_ sg13g2_or2_1
X_4535_ _1345_ net814 net1027 VPWR VGND sg13g2_nand2_1
Xhold301 DP_2.matrix\[0\] VPWR VGND net341 sg13g2_dlygate4sd3_1
Xhold312 DP_4.matrix\[78\] VPWR VGND net352 sg13g2_dlygate4sd3_1
Xhold334 DP_4.matrix\[75\] VPWR VGND net374 sg13g2_dlygate4sd3_1
Xhold323 _0025_ VPWR VGND net363 sg13g2_dlygate4sd3_1
Xhold367 _2177_ VPWR VGND net407 sg13g2_dlygate4sd3_1
Xhold378 DP_2.matrix\[4\] VPWR VGND net418 sg13g2_dlygate4sd3_1
Xhold356 mac2.sum_lvl3_ff\[5\] VPWR VGND net396 sg13g2_dlygate4sd3_1
Xhold345 DP_3.matrix\[4\] VPWR VGND net385 sg13g2_dlygate4sd3_1
X_4466_ _1277_ _1266_ _1279_ VPWR VGND sg13g2_xor2_1
Xfanout814 net815 net814 VPWR VGND sg13g2_buf_8
X_3417_ _0270_ _2990_ _0269_ VPWR VGND sg13g2_nand2_1
X_6205_ net1070 VGND VPWR net66 mac1.sum_lvl2_ff\[0\] clknet_leaf_63_clk sg13g2_dfrbpq_1
Xhold389 mac2.sum_lvl3_ff\[28\] VPWR VGND net429 sg13g2_dlygate4sd3_1
X_4397_ _1212_ _1197_ _1211_ VPWR VGND sg13g2_nand2_1
Xfanout825 net828 net825 VPWR VGND sg13g2_buf_8
Xfanout803 net374 net803 VPWR VGND sg13g2_buf_2
X_6136_ net1089 VGND VPWR _0226_ DP_3.matrix\[6\] clknet_leaf_26_clk sg13g2_dfrbpq_2
Xfanout836 net480 net836 VPWR VGND sg13g2_buf_8
X_3348_ _2935_ net908 net965 VPWR VGND sg13g2_nand2_1
Xfanout847 net316 net847 VPWR VGND sg13g2_buf_8
Xfanout858 net859 net858 VPWR VGND sg13g2_buf_8
Xfanout869 net489 net869 VPWR VGND sg13g2_buf_8
X_3279_ VGND VPWR _2868_ _2869_ _2834_ _2794_ sg13g2_a21oi_2
X_6067_ net1093 VGND VPWR _0178_ DP_1.matrix\[6\] clknet_leaf_58_clk sg13g2_dfrbpq_2
XFILLER_27_901 VPWR VGND sg13g2_decap_8
X_5018_ VGND VPWR _1801_ _1802_ _1805_ _1777_ sg13g2_a21oi_1
XFILLER_27_978 VPWR VGND sg13g2_decap_8
XFILLER_42_926 VPWR VGND sg13g2_decap_8
XFILLER_10_823 VPWR VGND sg13g2_fill_2
XFILLER_22_683 VPWR VGND sg13g2_fill_1
XFILLER_42_89 VPWR VGND sg13g2_fill_2
XFILLER_17_466 VPWR VGND sg13g2_fill_2
XFILLER_18_989 VPWR VGND sg13g2_decap_8
XFILLER_33_926 VPWR VGND sg13g2_decap_8
XFILLER_32_469 VPWR VGND sg13g2_fill_1
XFILLER_34_1014 VPWR VGND sg13g2_decap_8
XFILLER_41_970 VPWR VGND sg13g2_decap_8
XFILLER_9_621 VPWR VGND sg13g2_fill_2
XFILLER_40_480 VPWR VGND sg13g2_fill_1
XFILLER_8_164 VPWR VGND sg13g2_fill_1
X_4320_ _1125_ VPWR _1136_ VGND _1103_ _1126_ sg13g2_o21ai_1
X_4251_ _1067_ _1066_ _1069_ VPWR VGND sg13g2_xor2_1
X_3202_ _2746_ _2747_ _2791_ _2792_ _2794_ VPWR VGND sg13g2_and4_1
X_4182_ _1002_ _0995_ _0081_ VPWR VGND sg13g2_xor2_1
X_3133_ _2726_ net915 net969 VPWR VGND sg13g2_nand2_1
X_3064_ _2659_ net915 net975 VPWR VGND sg13g2_nand2_1
XFILLER_24_926 VPWR VGND sg13g2_decap_8
X_3966_ VGND VPWR _0794_ _0795_ _0798_ _0777_ sg13g2_a21oi_1
X_5705_ net784 VPWR _2401_ VGND net1037 net789 sg13g2_o21ai_1
XFILLER_32_992 VPWR VGND sg13g2_decap_8
X_3897_ _0728_ _0729_ _0730_ VPWR VGND sg13g2_nor2b_1
X_5636_ _2343_ VPWR _2345_ VGND _2342_ _2344_ sg13g2_o21ai_1
X_5567_ net458 _2289_ _0058_ VPWR VGND sg13g2_xor2_1
X_4518_ _1327_ _1290_ _1329_ VPWR VGND sg13g2_xor2_1
Xhold142 mac1.products_ff\[1\] VPWR VGND net182 sg13g2_dlygate4sd3_1
Xhold153 mac1.products_ff\[138\] VPWR VGND net193 sg13g2_dlygate4sd3_1
Xhold131 mac1.sum_lvl1_ff\[39\] VPWR VGND net171 sg13g2_dlygate4sd3_1
XFILLER_2_329 VPWR VGND sg13g2_fill_1
X_5498_ mac2.sum_lvl2_ff\[5\] net387 _2238_ VPWR VGND sg13g2_xor2_1
Xhold120 mac2.sum_lvl2_ff\[47\] VPWR VGND net160 sg13g2_dlygate4sd3_1
X_4449_ _1262_ net821 net1026 VPWR VGND sg13g2_nand2_1
Xhold164 mac1.products_ff\[141\] VPWR VGND net204 sg13g2_dlygate4sd3_1
Xhold175 mac2.products_ff\[146\] VPWR VGND net215 sg13g2_dlygate4sd3_1
Xhold186 mac2.sum_lvl1_ff\[42\] VPWR VGND net226 sg13g2_dlygate4sd3_1
Xhold197 mac2.sum_lvl1_ff\[43\] VPWR VGND net237 sg13g2_dlygate4sd3_1
X_6119_ net1071 VGND VPWR _0215_ DP_2.matrix\[75\] clknet_leaf_60_clk sg13g2_dfrbpq_1
XFILLER_2_1001 VPWR VGND sg13g2_decap_8
XFILLER_39_591 VPWR VGND sg13g2_decap_4
XFILLER_15_926 VPWR VGND sg13g2_fill_1
XFILLER_15_937 VPWR VGND sg13g2_decap_4
XFILLER_42_767 VPWR VGND sg13g2_fill_2
XFILLER_30_918 VPWR VGND sg13g2_decap_8
XFILLER_10_620 VPWR VGND sg13g2_fill_1
XFILLER_23_992 VPWR VGND sg13g2_decap_8
XFILLER_6_646 VPWR VGND sg13g2_fill_2
XFILLER_45_550 VPWR VGND sg13g2_decap_4
XFILLER_32_222 VPWR VGND sg13g2_fill_2
X_3820_ _0652_ _0653_ _0655_ _0656_ VPWR VGND sg13g2_or3_1
XFILLER_21_929 VPWR VGND sg13g2_decap_8
XFILLER_14_970 VPWR VGND sg13g2_decap_8
X_3751_ VGND VPWR _0571_ _0574_ _0594_ _0570_ sg13g2_a21oi_1
XFILLER_13_480 VPWR VGND sg13g2_fill_1
XFILLER_9_473 VPWR VGND sg13g2_fill_1
X_3682_ VGND VPWR _0527_ _0498_ _0496_ sg13g2_or2_1
X_6470_ net1102 VGND VPWR net53 mac2.sum_lvl2_ff\[23\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_5421_ net407 _2175_ _0026_ VPWR VGND sg13g2_xor2_1
X_5352_ mac1.sum_lvl2_ff\[5\] net505 _2124_ VPWR VGND sg13g2_xor2_1
X_4303_ _1117_ _1118_ _1112_ _1120_ VPWR VGND sg13g2_nand3_1
X_5283_ _2062_ net856 net1021 VPWR VGND sg13g2_nand2_1
XFILLER_4_93 VPWR VGND sg13g2_fill_2
X_4234_ _1050_ _1051_ _1045_ _1053_ VPWR VGND sg13g2_nand3_1
X_4165_ _0990_ net988 net1031 VPWR VGND sg13g2_nand2_1
X_3116_ _2709_ _2708_ _0101_ VPWR VGND sg13g2_xor2_1
X_4096_ _0924_ net989 net925 VPWR VGND sg13g2_nand2_2
X_3047_ VGND VPWR _2640_ _2641_ _2643_ _2635_ sg13g2_a21oi_1
XFILLER_17_1020 VPWR VGND sg13g2_decap_8
X_4998_ _1785_ _1784_ _1781_ VPWR VGND sg13g2_nand2b_1
X_3949_ VGND VPWR _0781_ _0779_ _0736_ sg13g2_or2_1
X_5619_ _2330_ VPWR _2333_ VGND _2329_ _2331_ sg13g2_o21ai_1
XFILLER_24_1024 VPWR VGND sg13g2_decap_4
XFILLER_46_325 VPWR VGND sg13g2_fill_2
XFILLER_46_369 VPWR VGND sg13g2_fill_2
XFILLER_15_712 VPWR VGND sg13g2_fill_1
XFILLER_7_911 VPWR VGND sg13g2_decap_8
XFILLER_11_995 VPWR VGND sg13g2_decap_8
XFILLER_31_1017 VPWR VGND sg13g2_decap_8
XFILLER_31_1028 VPWR VGND sg13g2_fill_1
XFILLER_7_955 VPWR VGND sg13g2_decap_8
XFILLER_9_1007 VPWR VGND sg13g2_decap_8
X_5970_ net928 _0210_ VPWR VGND sg13g2_buf_1
X_4921_ _1694_ VPWR _1715_ VGND _1666_ _1692_ sg13g2_o21ai_1
X_4852_ _1647_ _1637_ _1649_ VPWR VGND sg13g2_xor2_1
X_3803_ _0635_ VPWR _0640_ VGND _0636_ _0638_ sg13g2_o21ai_1
XFILLER_21_737 VPWR VGND sg13g2_fill_2
X_4783_ _1581_ _1574_ _1582_ VPWR VGND sg13g2_xor2_1
X_6522_ net1057 VGND VPWR DP_3.I_range.data_plus_4\[6\] DP_3.I_range.out_data\[5\]
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
X_3734_ _0577_ net1010 net1032 VPWR VGND sg13g2_nand2_1
X_3665_ _0511_ _0510_ _0509_ VPWR VGND sg13g2_nand2b_1
X_6453_ net1099 VGND VPWR net157 mac2.sum_lvl2_ff\[3\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_5404_ net286 mac1.sum_lvl2_ff\[19\] _0000_ VPWR VGND sg13g2_xor2_1
X_3596_ _0397_ _0400_ _0443_ VPWR VGND sg13g2_nor2_1
X_6384_ net1099 VGND VPWR _0082_ mac2.products_ff\[71\] clknet_leaf_29_clk sg13g2_dfrbpq_1
X_5335_ mac1.sum_lvl2_ff\[20\] mac1.sum_lvl2_ff\[1\] _2111_ VPWR VGND sg13g2_nor2_1
X_5266_ _2044_ _2035_ _2046_ VPWR VGND sg13g2_xor2_1
X_4217_ VGND VPWR _1037_ _1036_ _1016_ sg13g2_or2_1
X_5197_ _1979_ net857 net798 VPWR VGND sg13g2_nand2_1
X_4148_ _0974_ net990 DP_2.matrix\[44\] VPWR VGND sg13g2_nand2_1
XFILLER_29_848 VPWR VGND sg13g2_decap_8
XFILLER_44_829 VPWR VGND sg13g2_fill_1
X_4079_ _0908_ _0888_ _0907_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_358 VPWR VGND sg13g2_fill_1
XFILLER_11_214 VPWR VGND sg13g2_fill_1
XFILLER_7_207 VPWR VGND sg13g2_fill_1
Xclkload1 clknet_4_2_0_clk clkload1/X VPWR VGND sg13g2_buf_8
XFILLER_4_958 VPWR VGND sg13g2_decap_8
XFILLER_35_818 VPWR VGND sg13g2_decap_8
XFILLER_43_862 VPWR VGND sg13g2_decap_8
X_3450_ _0299_ _0296_ _0301_ VPWR VGND sg13g2_xor2_1
X_3381_ _2966_ _2956_ _2967_ VPWR VGND sg13g2_nor2b_1
XFILLER_41_4 VPWR VGND sg13g2_fill_2
X_5120_ _1904_ _1897_ _1902_ _1903_ VPWR VGND sg13g2_and3_1
X_5051_ _1837_ _1807_ _1835_ VPWR VGND sg13g2_xnor2_1
X_4002_ _0787_ VPWR _0833_ VGND _0785_ _0788_ sg13g2_o21ai_1
XFILLER_37_111 VPWR VGND sg13g2_fill_1
XFILLER_37_122 VPWR VGND sg13g2_decap_4
XFILLER_37_188 VPWR VGND sg13g2_fill_1
X_5953_ net992 _0185_ VPWR VGND sg13g2_buf_1
X_4904_ _1660_ _1698_ _1699_ VPWR VGND sg13g2_nor2_1
X_5884_ VGND VPWR net771 _2565_ _0198_ _2564_ sg13g2_a21oi_1
XFILLER_34_895 VPWR VGND sg13g2_decap_8
X_4835_ _1632_ net836 net891 VPWR VGND sg13g2_nand2_1
XFILLER_14_1012 VPWR VGND sg13g2_decap_8
X_4766_ _1565_ _1558_ _1564_ VPWR VGND sg13g2_xnor2_1
X_6505_ net1040 VGND VPWR net540 mac2.total_sum\[7\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3717_ _0559_ _0550_ _0561_ VPWR VGND sg13g2_xor2_1
X_4697_ _1474_ _1495_ _1497_ _1498_ VPWR VGND sg13g2_or3_1
X_3648_ _0494_ net1010 DP_2.matrix\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_20_48 VPWR VGND sg13g2_fill_2
X_6436_ net1120 VGND VPWR net196 mac2.sum_lvl1_ff\[43\] clknet_leaf_41_clk sg13g2_dfrbpq_1
XFILLER_1_917 VPWR VGND sg13g2_decap_8
X_3579_ _0404_ _0424_ _0426_ _0427_ VPWR VGND sg13g2_or3_1
X_6367_ net1086 VGND VPWR _0086_ mac2.products_ff\[2\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_5318_ _2095_ _2085_ _2096_ VPWR VGND sg13g2_nor2b_1
XFILLER_0_449 VPWR VGND sg13g2_fill_1
Xhold13 mac2.sum_lvl1_ff\[40\] VPWR VGND net53 sg13g2_dlygate4sd3_1
X_6298_ net1058 VGND VPWR net105 mac2.sum_lvl1_ff\[85\] clknet_leaf_21_clk sg13g2_dfrbpq_1
Xhold24 mac2.products_ff\[82\] VPWR VGND net64 sg13g2_dlygate4sd3_1
Xhold35 mac2.products_ff\[13\] VPWR VGND net75 sg13g2_dlygate4sd3_1
Xhold46 mac1.sum_lvl2_ff\[45\] VPWR VGND net86 sg13g2_dlygate4sd3_1
X_5249_ _0151_ _2028_ _2029_ VPWR VGND sg13g2_xnor2_1
Xhold68 mac2.sum_lvl1_ff\[48\] VPWR VGND net108 sg13g2_dlygate4sd3_1
Xhold79 mac1.products_ff\[145\] VPWR VGND net119 sg13g2_dlygate4sd3_1
XFILLER_21_1027 VPWR VGND sg13g2_fill_2
Xhold57 mac2.products_ff\[11\] VPWR VGND net97 sg13g2_dlygate4sd3_1
XFILLER_44_659 VPWR VGND sg13g2_fill_2
XFILLER_40_854 VPWR VGND sg13g2_decap_8
Xfanout1022 net383 net1022 VPWR VGND sg13g2_buf_8
Xfanout1000 net495 net1000 VPWR VGND sg13g2_buf_8
Xfanout1011 net1012 net1011 VPWR VGND sg13g2_buf_8
XFILLER_0_961 VPWR VGND sg13g2_decap_8
Xfanout1033 net314 net1033 VPWR VGND sg13g2_buf_8
Xfanout1044 net1048 net1044 VPWR VGND sg13g2_buf_8
Xfanout1055 net1063 net1055 VPWR VGND sg13g2_buf_8
XFILLER_48_954 VPWR VGND sg13g2_decap_8
Xfanout1088 net1089 net1088 VPWR VGND sg13g2_buf_8
Xfanout1066 net1067 net1066 VPWR VGND sg13g2_buf_8
Xfanout1077 net1080 net1077 VPWR VGND sg13g2_buf_8
Xfanout1099 net1101 net1099 VPWR VGND sg13g2_buf_8
XFILLER_47_475 VPWR VGND sg13g2_fill_1
XFILLER_37_1012 VPWR VGND sg13g2_decap_8
X_4620_ _1423_ _1416_ _1421_ _1422_ VPWR VGND sg13g2_and3_1
XFILLER_31_898 VPWR VGND sg13g2_decap_8
X_4551_ _1348_ VPWR _1360_ VGND _1320_ _1346_ sg13g2_o21ai_1
X_4482_ _1263_ VPWR _1294_ VGND _1261_ _1264_ sg13g2_o21ai_1
X_3502_ _0352_ _0322_ _0350_ VPWR VGND sg13g2_xnor2_1
Xhold505 mac2.sum_lvl2_ff\[9\] VPWR VGND net545 sg13g2_dlygate4sd3_1
X_3433_ _0280_ VPWR _0285_ VGND _0281_ _0283_ sg13g2_o21ai_1
X_6221_ net1066 VGND VPWR net146 mac1.sum_lvl2_ff\[19\] clknet_leaf_63_clk sg13g2_dfrbpq_1
X_6152_ net1081 VGND VPWR _0237_ DP_3.matrix\[73\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_3364_ _0098_ _2949_ _2950_ VPWR VGND sg13g2_xnor2_1
X_5103_ _1887_ _1879_ _1886_ VPWR VGND sg13g2_nand2_1
X_6083_ net1067 VGND VPWR _0191_ DP_1.matrix\[75\] clknet_leaf_60_clk sg13g2_dfrbpq_1
X_3295_ _2884_ net975 net1030 VPWR VGND sg13g2_nand2_1
Xheichips25_template_37 VPWR VGND uio_oe[4] sg13g2_tiehi
XFILLER_39_954 VPWR VGND sg13g2_decap_8
X_5034_ _1820_ net804 net859 VPWR VGND sg13g2_nand2_1
X_5936_ VGND VPWR net770 _2597_ _0250_ _2596_ sg13g2_a21oi_1
XFILLER_33_180 VPWR VGND sg13g2_fill_2
XFILLER_40_128 VPWR VGND sg13g2_fill_1
X_5867_ VGND VPWR net774 _2555_ _0175_ _2554_ sg13g2_a21oi_1
XFILLER_21_364 VPWR VGND sg13g2_fill_2
X_4818_ _1616_ _1606_ _1615_ VPWR VGND sg13g2_nand2b_1
X_5798_ _2489_ VPWR _2492_ VGND _2490_ _2491_ sg13g2_o21ai_1
X_4749_ _1547_ _1548_ _1546_ _1549_ VPWR VGND sg13g2_nand3_1
Xoutput25 net25 uo_out[0] VPWR VGND sg13g2_buf_1
X_6419_ net1102 VGND VPWR net96 mac2.sum_lvl1_ff\[6\] clknet_leaf_30_clk sg13g2_dfrbpq_1
XFILLER_48_228 VPWR VGND sg13g2_fill_2
XFILLER_45_924 VPWR VGND sg13g2_decap_8
XFILLER_29_497 VPWR VGND sg13g2_decap_4
XFILLER_16_125 VPWR VGND sg13g2_fill_1
XFILLER_17_659 VPWR VGND sg13g2_fill_2
XFILLER_13_887 VPWR VGND sg13g2_fill_1
XFILLER_40_640 VPWR VGND sg13g2_fill_2
X_3080_ _2672_ _2673_ _2648_ _2675_ VPWR VGND sg13g2_nand3_1
XFILLER_35_434 VPWR VGND sg13g2_fill_1
XFILLER_36_957 VPWR VGND sg13g2_decap_8
X_3982_ _0774_ VPWR _0813_ VGND _0729_ _0775_ sg13g2_o21ai_1
X_5721_ _2417_ net983 net790 VPWR VGND sg13g2_nand2_1
XFILLER_22_128 VPWR VGND sg13g2_fill_1
X_5652_ _2357_ VPWR _2358_ VGND _2351_ _2354_ sg13g2_o21ai_1
XFILLER_31_684 VPWR VGND sg13g2_fill_2
X_5583_ _2304_ mac2.sum_lvl3_ff\[28\] net423 VPWR VGND sg13g2_xnor2_1
X_4603_ _1405_ _1404_ _1407_ VPWR VGND sg13g2_xor2_1
X_4534_ _1344_ net873 net1022 VPWR VGND sg13g2_nand2_1
Xhold302 DP_4.matrix\[43\] VPWR VGND net342 sg13g2_dlygate4sd3_1
XFILLER_8_880 VPWR VGND sg13g2_decap_4
Xhold335 mac1.sum_lvl2_ff\[8\] VPWR VGND net375 sg13g2_dlygate4sd3_1
Xhold324 mac1.sum_lvl3_ff\[10\] VPWR VGND net364 sg13g2_dlygate4sd3_1
Xhold313 mac2.sum_lvl2_ff\[3\] VPWR VGND net353 sg13g2_dlygate4sd3_1
Xhold346 DP_4.matrix\[6\] VPWR VGND net386 sg13g2_dlygate4sd3_1
Xhold368 _0026_ VPWR VGND net408 sg13g2_dlygate4sd3_1
Xhold357 _2294_ VPWR VGND net397 sg13g2_dlygate4sd3_1
X_4465_ _1266_ _1277_ _1278_ VPWR VGND sg13g2_nor2_1
Xfanout815 net342 net815 VPWR VGND sg13g2_buf_8
Xhold379 mac1.sum_lvl3_ff\[27\] VPWR VGND net419 sg13g2_dlygate4sd3_1
X_3416_ _2995_ _0268_ _0269_ VPWR VGND sg13g2_nor2b_1
X_6204_ net1114 VGND VPWR net258 mac1.sum_lvl1_ff\[51\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_4396_ _1210_ _1203_ _1211_ VPWR VGND sg13g2_xor2_1
Xfanout804 net805 net804 VPWR VGND sg13g2_buf_8
Xfanout837 net414 net837 VPWR VGND sg13g2_buf_8
X_6135_ net1092 VGND VPWR net147 mac1.sum_lvl1_ff\[4\] clknet_leaf_54_clk sg13g2_dfrbpq_1
X_3347_ _2934_ net965 net906 VPWR VGND sg13g2_nand2_1
Xfanout848 DP_4.matrix\[0\] net848 VPWR VGND sg13g2_buf_1
Xfanout826 net828 net826 VPWR VGND sg13g2_buf_8
X_6066_ net1093 VGND VPWR _0177_ DP_1.matrix\[5\] clknet_leaf_58_clk sg13g2_dfrbpq_1
Xfanout859 DP_3.matrix\[76\] net859 VPWR VGND sg13g2_buf_2
X_3278_ VGND VPWR _2791_ _2833_ _2868_ _2832_ sg13g2_a21oi_1
X_5017_ _1801_ _1802_ _1777_ _1804_ VPWR VGND sg13g2_nand3_1
XFILLER_42_905 VPWR VGND sg13g2_decap_8
XFILLER_27_957 VPWR VGND sg13g2_decap_8
XFILLER_41_426 VPWR VGND sg13g2_fill_1
X_5919_ _0244_ net847 net767 VPWR VGND sg13g2_xnor2_1
XFILLER_6_828 VPWR VGND sg13g2_fill_1
XFILLER_1_522 VPWR VGND sg13g2_fill_1
XFILLER_49_548 VPWR VGND sg13g2_fill_2
XFILLER_18_968 VPWR VGND sg13g2_decap_8
XFILLER_33_905 VPWR VGND sg13g2_decap_8
XFILLER_17_456 VPWR VGND sg13g2_fill_1
XFILLER_13_673 VPWR VGND sg13g2_decap_8
X_4250_ _1068_ _1066_ _1067_ VPWR VGND sg13g2_nand2b_1
X_3201_ _2793_ _2791_ _2792_ VPWR VGND sg13g2_nand2_1
X_4181_ _1003_ _0995_ _1002_ VPWR VGND sg13g2_nand2_1
X_3132_ _2693_ VPWR _2725_ VGND _2691_ _2694_ sg13g2_o21ai_1
XFILLER_41_1019 VPWR VGND sg13g2_decap_8
X_3063_ _2638_ VPWR _2658_ VGND _2636_ _2639_ sg13g2_o21ai_1
XFILLER_36_798 VPWR VGND sg13g2_fill_2
X_3965_ _0794_ _0795_ _0777_ _0797_ VPWR VGND sg13g2_nand3_1
X_3896_ net1001 net927 net1004 _0729_ VPWR VGND net925 sg13g2_nand4_1
X_5704_ DP_1.Q_range.out_data\[2\] DP_1.I_range.out_data\[2\] _2400_ VPWR VGND sg13g2_xor2_1
XFILLER_31_470 VPWR VGND sg13g2_fill_2
XFILLER_32_971 VPWR VGND sg13g2_decap_8
X_5635_ _2344_ _2342_ net28 VPWR VGND sg13g2_xor2_1
X_5566_ net457 mac2.sum_lvl3_ff\[24\] _2291_ VPWR VGND sg13g2_xor2_1
Xhold110 mac2.sum_lvl1_ff\[74\] VPWR VGND net150 sg13g2_dlygate4sd3_1
X_4517_ _1290_ _1327_ _1328_ VPWR VGND sg13g2_nor2_1
X_5497_ net387 mac2.sum_lvl2_ff\[5\] _2237_ VPWR VGND sg13g2_nor2_1
Xhold121 mac2.sum_lvl1_ff\[2\] VPWR VGND net161 sg13g2_dlygate4sd3_1
Xhold132 mac2.products_ff\[74\] VPWR VGND net172 sg13g2_dlygate4sd3_1
Xhold143 mac2.products_ff\[3\] VPWR VGND net183 sg13g2_dlygate4sd3_1
X_4448_ _1261_ net818 net873 VPWR VGND sg13g2_nand2_1
Xhold165 mac1.sum_lvl1_ff\[82\] VPWR VGND net205 sg13g2_dlygate4sd3_1
Xhold176 mac2.sum_lvl1_ff\[45\] VPWR VGND net216 sg13g2_dlygate4sd3_1
Xhold154 mac2.sum_lvl1_ff\[85\] VPWR VGND net194 sg13g2_dlygate4sd3_1
Xhold187 mac2.sum_lvl2_ff\[53\] VPWR VGND net227 sg13g2_dlygate4sd3_1
Xhold198 mac1.products_ff\[148\] VPWR VGND net238 sg13g2_dlygate4sd3_1
X_4379_ _1194_ _1187_ _1193_ VPWR VGND sg13g2_xnor2_1
X_6118_ net1065 VGND VPWR _0214_ DP_2.matrix\[74\] clknet_leaf_65_clk sg13g2_dfrbpq_1
X_6049_ net1093 VGND VPWR _0160_ DP_1.matrix\[8\] clknet_leaf_58_clk sg13g2_dfrbpq_1
XFILLER_15_916 VPWR VGND sg13g2_fill_1
XFILLER_42_735 VPWR VGND sg13g2_fill_2
XFILLER_42_779 VPWR VGND sg13g2_decap_4
XFILLER_23_971 VPWR VGND sg13g2_decap_8
XFILLER_22_481 VPWR VGND sg13g2_fill_1
XFILLER_49_301 VPWR VGND sg13g2_fill_1
XFILLER_17_231 VPWR VGND sg13g2_fill_2
XFILLER_18_776 VPWR VGND sg13g2_fill_2
XFILLER_45_584 VPWR VGND sg13g2_fill_1
X_3750_ _0591_ _0592_ _0593_ VPWR VGND sg13g2_and2_1
XFILLER_9_485 VPWR VGND sg13g2_fill_2
X_3681_ _0486_ VPWR _0526_ VGND _0483_ _0487_ sg13g2_o21ai_1
X_5420_ mac1.sum_lvl3_ff\[4\] net406 _2177_ VPWR VGND sg13g2_xor2_1
X_5351_ net505 mac1.sum_lvl2_ff\[5\] _2123_ VPWR VGND sg13g2_nor2_1
X_5282_ _2040_ VPWR _2061_ VGND _2037_ _2041_ sg13g2_o21ai_1
X_4302_ _1119_ _1112_ _1117_ _1118_ VPWR VGND sg13g2_and3_1
X_4233_ _1052_ _1045_ _1050_ _1051_ VPWR VGND sg13g2_and3_1
X_4164_ _0978_ VPWR _0989_ VGND _0949_ _0976_ sg13g2_o21ai_1
X_3115_ _2675_ VPWR _2709_ VGND _2650_ _2676_ sg13g2_o21ai_1
X_4095_ _0923_ net995 net1031 VPWR VGND sg13g2_nand2_1
X_3046_ _2640_ _2641_ _2635_ _2642_ VPWR VGND sg13g2_nand3_1
XFILLER_24_724 VPWR VGND sg13g2_decap_4
XFILLER_24_746 VPWR VGND sg13g2_decap_8
XFILLER_24_779 VPWR VGND sg13g2_decap_4
X_4997_ _1783_ _1760_ _1784_ VPWR VGND sg13g2_xor2_1
X_3948_ _0780_ net933 net991 VPWR VGND sg13g2_nand2_1
XFILLER_32_790 VPWR VGND sg13g2_fill_1
X_3879_ _0713_ _0706_ _0711_ _0712_ VPWR VGND sg13g2_and3_1
XFILLER_20_985 VPWR VGND sg13g2_decap_8
X_5618_ _0053_ _2329_ net329 VPWR VGND sg13g2_xnor2_1
X_5549_ _0038_ _2277_ net528 VPWR VGND sg13g2_xnor2_1
XFILLER_24_1003 VPWR VGND sg13g2_decap_8
XFILLER_42_510 VPWR VGND sg13g2_fill_2
XFILLER_14_234 VPWR VGND sg13g2_fill_1
XFILLER_7_901 VPWR VGND sg13g2_decap_4
XFILLER_11_974 VPWR VGND sg13g2_decap_8
XFILLER_6_466 VPWR VGND sg13g2_fill_2
XFILLER_43_8 VPWR VGND sg13g2_fill_1
XFILLER_2_672 VPWR VGND sg13g2_fill_1
XFILLER_38_849 VPWR VGND sg13g2_decap_8
X_4920_ _1697_ _1689_ _1696_ _1714_ VPWR VGND sg13g2_a21o_1
X_4851_ _1637_ _1647_ _1648_ VPWR VGND sg13g2_nor2_1
XFILLER_33_532 VPWR VGND sg13g2_fill_1
X_3802_ _0635_ _0636_ _0638_ _0639_ VPWR VGND sg13g2_nor3_1
X_4782_ _1581_ _1575_ _1579_ VPWR VGND sg13g2_xnor2_1
X_6521_ net1057 VGND VPWR net15 DP_3.I_range.out_data\[4\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_3733_ _0555_ VPWR _0576_ VGND _0552_ _0556_ sg13g2_o21ai_1
X_3664_ _0474_ _0508_ _0472_ _0510_ VPWR VGND sg13g2_nand3_1
X_6452_ net1099 VGND VPWR net161 mac2.sum_lvl2_ff\[2\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_5403_ _0006_ _2163_ net391 VPWR VGND sg13g2_xnor2_1
X_3595_ _0425_ VPWR _0442_ VGND _0404_ _0426_ sg13g2_o21ai_1
X_6383_ net1085 VGND VPWR _0081_ mac2.products_ff\[70\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_47_1025 VPWR VGND sg13g2_decap_4
X_5334_ _2110_ mac1.sum_lvl2_ff\[20\] mac1.sum_lvl2_ff\[1\] VPWR VGND sg13g2_nand2_1
X_5265_ _2044_ _2035_ _2045_ VPWR VGND sg13g2_nor2b_1
X_5196_ VGND VPWR net807 net851 _1978_ _1947_ sg13g2_a21oi_1
XFILLER_29_805 VPWR VGND sg13g2_decap_4
X_4216_ _1034_ _1033_ _1036_ VPWR VGND sg13g2_xor2_1
X_4147_ _0952_ VPWR _0973_ VGND _0924_ _0950_ sg13g2_o21ai_1
X_4078_ _0905_ _0895_ _0907_ VPWR VGND sg13g2_xor2_1
X_3029_ _2626_ _2618_ _2625_ VPWR VGND sg13g2_nand2_1
XFILLER_37_893 VPWR VGND sg13g2_decap_8
XFILLER_11_226 VPWR VGND sg13g2_fill_1
Xclkload2 clknet_4_3_0_clk clkload2/X VPWR VGND sg13g2_buf_8
XFILLER_4_937 VPWR VGND sg13g2_decap_8
XFILLER_46_123 VPWR VGND sg13g2_decap_8
XFILLER_46_134 VPWR VGND sg13g2_fill_2
X_3380_ _2966_ _2942_ _2965_ VPWR VGND sg13g2_xnor2_1
X_5050_ _1835_ _1807_ _1836_ VPWR VGND sg13g2_nor2b_1
X_4001_ _0832_ _0827_ _0831_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_657 VPWR VGND sg13g2_fill_2
X_5952_ net994 _0184_ VPWR VGND sg13g2_buf_1
XFILLER_25_329 VPWR VGND sg13g2_fill_1
X_4903_ _1698_ _1689_ _1697_ VPWR VGND sg13g2_xnor2_1
XFILLER_18_392 VPWR VGND sg13g2_decap_4
X_5883_ _2565_ _2452_ _2454_ VPWR VGND sg13g2_xnor2_1
XFILLER_34_874 VPWR VGND sg13g2_decap_8
X_4834_ _1614_ _1607_ _1577_ _1631_ VPWR VGND sg13g2_a21o_2
XFILLER_21_524 VPWR VGND sg13g2_fill_2
X_4765_ _1564_ _1559_ _1562_ VPWR VGND sg13g2_xnor2_1
X_6504_ net1043 VGND VPWR net466 mac2.total_sum\[6\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3716_ _0559_ _0550_ _0560_ VPWR VGND sg13g2_nor2b_1
X_4696_ VGND VPWR _1493_ _1494_ _1497_ _1475_ sg13g2_a21oi_1
X_3647_ VGND VPWR net958 net1005 _0493_ _0462_ sg13g2_a21oi_1
X_6435_ net1103 VGND VPWR net172 mac2.sum_lvl1_ff\[42\] clknet_leaf_42_clk sg13g2_dfrbpq_1
X_3578_ VGND VPWR _0422_ _0423_ _0426_ _0405_ sg13g2_a21oi_1
X_6366_ net1083 VGND VPWR _0085_ mac2.products_ff\[1\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_5317_ _2095_ _2071_ _2094_ VPWR VGND sg13g2_xnor2_1
Xhold14 mac2.products_ff\[139\] VPWR VGND net54 sg13g2_dlygate4sd3_1
X_6297_ net1052 VGND VPWR net253 mac2.sum_lvl1_ff\[84\] clknet_leaf_21_clk sg13g2_dfrbpq_1
Xhold36 mac1.sum_lvl1_ff\[6\] VPWR VGND net76 sg13g2_dlygate4sd3_1
Xhold25 mac2.products_ff\[140\] VPWR VGND net65 sg13g2_dlygate4sd3_1
Xhold47 mac2.sum_lvl1_ff\[73\] VPWR VGND net87 sg13g2_dlygate4sd3_1
X_5248_ _1994_ _1999_ _2029_ VPWR VGND sg13g2_nor2_1
XFILLER_21_1006 VPWR VGND sg13g2_decap_8
Xhold58 mac2.products_ff\[76\] VPWR VGND net98 sg13g2_dlygate4sd3_1
Xhold69 mac2.sum_lvl1_ff\[5\] VPWR VGND net109 sg13g2_dlygate4sd3_1
X_5179_ _1962_ _1925_ _1960_ VPWR VGND sg13g2_nand2_1
XFILLER_43_104 VPWR VGND sg13g2_fill_1
XFILLER_43_148 VPWR VGND sg13g2_fill_2
XFILLER_25_852 VPWR VGND sg13g2_fill_1
XFILLER_40_833 VPWR VGND sg13g2_decap_8
XFILLER_20_590 VPWR VGND sg13g2_fill_1
Xfanout1001 net1002 net1001 VPWR VGND sg13g2_buf_8
XFILLER_0_940 VPWR VGND sg13g2_decap_8
Xfanout1012 net526 net1012 VPWR VGND sg13g2_buf_8
Xfanout1023 net541 net1023 VPWR VGND sg13g2_buf_8
Xfanout1034 DP_1.matrix\[80\] net1034 VPWR VGND sg13g2_buf_1
Xfanout1045 net1048 net1045 VPWR VGND sg13g2_buf_8
Xfanout1056 net1058 net1056 VPWR VGND sg13g2_buf_8
XFILLER_48_933 VPWR VGND sg13g2_decap_8
Xfanout1089 net1090 net1089 VPWR VGND sg13g2_buf_8
Xfanout1067 net1069 net1067 VPWR VGND sg13g2_buf_8
Xfanout1078 net1080 net1078 VPWR VGND sg13g2_buf_8
XFILLER_35_605 VPWR VGND sg13g2_fill_2
XFILLER_34_115 VPWR VGND sg13g2_fill_2
XFILLER_16_852 VPWR VGND sg13g2_fill_2
XFILLER_34_148 VPWR VGND sg13g2_fill_1
XFILLER_16_874 VPWR VGND sg13g2_fill_1
XFILLER_30_343 VPWR VGND sg13g2_fill_2
XFILLER_31_877 VPWR VGND sg13g2_decap_8
XFILLER_30_398 VPWR VGND sg13g2_fill_1
X_4550_ VGND VPWR _1328_ _1352_ _1359_ _1354_ sg13g2_a21oi_1
X_4481_ _1272_ VPWR _1293_ VGND _1269_ _1273_ sg13g2_o21ai_1
X_3501_ _0350_ _0322_ _0351_ VPWR VGND sg13g2_nor2b_1
Xhold506 mac1.sum_lvl2_ff\[31\] VPWR VGND net546 sg13g2_dlygate4sd3_1
X_3432_ _0280_ _0281_ _0283_ _0284_ VPWR VGND sg13g2_or3_1
X_6220_ net1128 VGND VPWR net169 mac1.sum_lvl2_ff\[15\] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_3363_ VGND VPWR _2927_ _2930_ _2950_ _2926_ sg13g2_a21oi_1
X_6151_ net1081 VGND VPWR _0236_ DP_3.matrix\[72\] clknet_leaf_28_clk sg13g2_dfrbpq_1
XFILLER_44_1028 VPWR VGND sg13g2_fill_1
X_5102_ _1884_ _1880_ _1886_ VPWR VGND sg13g2_xor2_1
X_6082_ net1071 VGND VPWR _0190_ DP_1.matrix\[74\] clknet_leaf_61_clk sg13g2_dfrbpq_1
X_3294_ VGND VPWR _2883_ _2854_ _2852_ sg13g2_or2_1
XFILLER_25_0 VPWR VGND sg13g2_fill_1
X_5033_ _1790_ VPWR _1819_ VGND _1788_ _1791_ sg13g2_o21ai_1
XFILLER_39_933 VPWR VGND sg13g2_decap_8
Xheichips25_template_38 VPWR VGND uio_oe[5] sg13g2_tiehi
X_5935_ _2544_ _2540_ _2597_ VPWR VGND sg13g2_xor2_1
X_5866_ _2555_ _2413_ _2423_ VPWR VGND sg13g2_xnor2_1
X_4817_ _1615_ _1607_ _1614_ VPWR VGND sg13g2_xnor2_1
Xclkbuf_leaf_60_clk clknet_4_2_0_clk clknet_leaf_60_clk VPWR VGND sg13g2_buf_8
X_5797_ net777 VPWR _2491_ VGND net903 net785 sg13g2_o21ai_1
X_4748_ _1500_ VPWR _1548_ VGND _1439_ _1501_ sg13g2_o21ai_1
X_4679_ _1443_ _1478_ _1480_ VPWR VGND sg13g2_and2_1
X_6418_ net1100 VGND VPWR net111 mac2.sum_lvl1_ff\[5\] clknet_leaf_29_clk sg13g2_dfrbpq_1
Xoutput26 net26 uo_out[1] VPWR VGND sg13g2_buf_1
X_6349_ net1039 VGND VPWR net266 mac1.total_sum\[0\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_0_247 VPWR VGND sg13g2_decap_8
XFILLER_45_903 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_51_clk clknet_4_10_0_clk clknet_leaf_51_clk VPWR VGND sg13g2_buf_8
XFILLER_8_325 VPWR VGND sg13g2_fill_2
XFILLER_8_314 VPWR VGND sg13g2_fill_1
XFILLER_39_229 VPWR VGND sg13g2_fill_1
XFILLER_36_936 VPWR VGND sg13g2_decap_8
X_3981_ _0802_ VPWR _0812_ VGND _0731_ _0803_ sg13g2_o21ai_1
XFILLER_16_660 VPWR VGND sg13g2_fill_1
XFILLER_23_608 VPWR VGND sg13g2_decap_8
XFILLER_35_468 VPWR VGND sg13g2_fill_1
XFILLER_35_479 VPWR VGND sg13g2_fill_2
X_5720_ net1018 net789 _2416_ VPWR VGND sg13g2_nor2_1
XFILLER_16_682 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_42_clk clknet_4_12_0_clk clknet_leaf_42_clk VPWR VGND sg13g2_buf_8
X_5651_ mac2.total_sum\[7\] mac1.total_sum\[7\] _2357_ VPWR VGND sg13g2_xor2_1
XFILLER_30_173 VPWR VGND sg13g2_fill_2
X_5582_ net539 _2303_ _0061_ VPWR VGND sg13g2_and2_1
X_4602_ _1404_ _1405_ _1406_ VPWR VGND sg13g2_nor2b_2
X_4533_ _1326_ _1318_ _1325_ _1343_ VPWR VGND sg13g2_a21o_1
XFILLER_11_1016 VPWR VGND sg13g2_decap_8
XFILLER_11_1027 VPWR VGND sg13g2_fill_2
Xhold303 mac2.sum_lvl3_ff\[15\] VPWR VGND net343 sg13g2_dlygate4sd3_1
Xhold325 _0018_ VPWR VGND net365 sg13g2_dlygate4sd3_1
Xhold314 _2232_ VPWR VGND net354 sg13g2_dlygate4sd3_1
Xhold369 DP_4.matrix\[3\] VPWR VGND net409 sg13g2_dlygate4sd3_1
Xhold336 _2134_ VPWR VGND net376 sg13g2_dlygate4sd3_1
Xhold358 _0059_ VPWR VGND net398 sg13g2_dlygate4sd3_1
X_6203_ net1114 VGND VPWR net141 mac1.sum_lvl1_ff\[50\] clknet_leaf_47_clk sg13g2_dfrbpq_1
Xhold347 mac2.sum_lvl2_ff\[24\] VPWR VGND net387 sg13g2_dlygate4sd3_1
X_4464_ _1275_ _1267_ _1277_ VPWR VGND sg13g2_xor2_1
Xfanout816 net817 net816 VPWR VGND sg13g2_buf_8
X_3415_ _2991_ VPWR _0268_ VGND _2992_ _2994_ sg13g2_o21ai_1
X_4395_ _1210_ _1204_ _1208_ VPWR VGND sg13g2_xnor2_1
Xfanout805 net308 net805 VPWR VGND sg13g2_buf_2
X_6134_ net1089 VGND VPWR net417 DP_3.matrix\[5\] clknet_leaf_25_clk sg13g2_dfrbpq_1
Xfanout838 DP_4.matrix\[4\] net838 VPWR VGND sg13g2_buf_1
X_3346_ _2933_ net971 net1030 VPWR VGND sg13g2_nand2_1
Xfanout827 net828 net827 VPWR VGND sg13g2_buf_2
Xfanout849 net850 net849 VPWR VGND sg13g2_buf_2
X_6065_ net1075 VGND VPWR _0176_ DP_1.matrix\[4\] clknet_leaf_57_clk sg13g2_dfrbpq_1
X_3277_ _2867_ _2866_ _2865_ VPWR VGND sg13g2_nand2b_1
X_5016_ _1801_ _1802_ _1803_ VPWR VGND sg13g2_and2_1
XFILLER_27_936 VPWR VGND sg13g2_decap_8
XFILLER_41_405 VPWR VGND sg13g2_fill_2
X_5918_ net325 VPWR _0227_ VGND _2514_ _2586_ sg13g2_o21ai_1
Xclkbuf_leaf_33_clk clknet_4_13_0_clk clknet_leaf_33_clk VPWR VGND sg13g2_buf_8
X_5849_ net817 net787 _2542_ VPWR VGND sg13g2_nor2_1
XFILLER_10_825 VPWR VGND sg13g2_fill_1
XFILLER_10_869 VPWR VGND sg13g2_fill_1
XFILLER_49_527 VPWR VGND sg13g2_decap_8
XFILLER_17_402 VPWR VGND sg13g2_decap_4
XFILLER_32_405 VPWR VGND sg13g2_fill_1
XFILLER_44_298 VPWR VGND sg13g2_fill_2
XFILLER_26_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_24_clk clknet_4_5_0_clk clknet_leaf_24_clk VPWR VGND sg13g2_buf_8
XFILLER_9_623 VPWR VGND sg13g2_fill_1
XFILLER_4_372 VPWR VGND sg13g2_fill_1
X_3200_ _2789_ _2788_ _2790_ _2792_ VPWR VGND sg13g2_a21o_1
X_4180_ _1000_ _1001_ _1002_ VPWR VGND sg13g2_nor2b_1
X_3131_ _2724_ _2718_ _2723_ VPWR VGND sg13g2_xnor2_1
X_3062_ _2655_ _2652_ _2657_ VPWR VGND sg13g2_xor2_1
XFILLER_36_766 VPWR VGND sg13g2_fill_2
X_3964_ _0796_ _0777_ _0794_ _0795_ VPWR VGND sg13g2_and3_1
XFILLER_32_950 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_15_clk clknet_4_6_0_clk clknet_leaf_15_clk VPWR VGND sg13g2_buf_8
X_3895_ _0728_ net925 net1004 net927 net1001 VPWR VGND sg13g2_a22oi_1
X_5703_ _2399_ DP_1.I_range.out_data\[2\] DP_1.Q_range.out_data\[2\] VPWR VGND sg13g2_xnor2_1
X_5634_ _2344_ mac1.total_sum\[3\] mac2.total_sum\[3\] VPWR VGND sg13g2_xnor2_1
Xhold100 mac1.sum_lvl1_ff\[5\] VPWR VGND net140 sg13g2_dlygate4sd3_1
X_5565_ mac2.sum_lvl3_ff\[24\] net457 _2290_ VPWR VGND sg13g2_and2_1
Xhold111 mac2.products_ff\[83\] VPWR VGND net151 sg13g2_dlygate4sd3_1
Xhold133 mac2.products_ff\[150\] VPWR VGND net173 sg13g2_dlygate4sd3_1
X_4516_ _1327_ _1318_ _1326_ VPWR VGND sg13g2_xnor2_1
Xhold144 mac1.sum_lvl1_ff\[43\] VPWR VGND net184 sg13g2_dlygate4sd3_1
Xhold122 mac1.products_ff\[80\] VPWR VGND net162 sg13g2_dlygate4sd3_1
X_5496_ VGND VPWR _2233_ _2235_ _2236_ _2234_ sg13g2_a21oi_1
Xhold177 mac1.sum_lvl2_ff\[44\] VPWR VGND net217 sg13g2_dlygate4sd3_1
Xhold166 mac1.products_ff\[78\] VPWR VGND net206 sg13g2_dlygate4sd3_1
Xhold155 mac2.sum_lvl1_ff\[78\] VPWR VGND net195 sg13g2_dlygate4sd3_1
X_4447_ _1243_ _1236_ _1206_ _1260_ VPWR VGND sg13g2_a21o_1
Xhold188 mac1.products_ff\[71\] VPWR VGND net228 sg13g2_dlygate4sd3_1
Xhold199 mac2.sum_lvl1_ff\[44\] VPWR VGND net239 sg13g2_dlygate4sd3_1
X_6117_ net1068 VGND VPWR _0099_ mac1.products_ff\[150\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_4378_ _1193_ _1188_ _1191_ VPWR VGND sg13g2_xnor2_1
X_3329_ _2915_ _2907_ _2917_ VPWR VGND sg13g2_xor2_1
X_6048_ net1116 VGND VPWR _0122_ mac1.products_ff\[83\] clknet_leaf_47_clk sg13g2_dfrbpq_1
XFILLER_26_221 VPWR VGND sg13g2_fill_2
XFILLER_41_202 VPWR VGND sg13g2_fill_1
XFILLER_23_950 VPWR VGND sg13g2_decap_8
XFILLER_6_648 VPWR VGND sg13g2_fill_1
XFILLER_18_700 VPWR VGND sg13g2_fill_2
XFILLER_45_574 VPWR VGND sg13g2_fill_2
XFILLER_18_799 VPWR VGND sg13g2_fill_1
XFILLER_14_950 VPWR VGND sg13g2_decap_4
XFILLER_32_224 VPWR VGND sg13g2_fill_1
X_3680_ _0525_ _0517_ _0522_ VPWR VGND sg13g2_xnor2_1
X_5350_ VGND VPWR _2119_ _2121_ _2122_ _2120_ sg13g2_a21oi_1
X_5281_ _2043_ _2036_ _2045_ _2060_ VPWR VGND sg13g2_a21o_1
X_4301_ _1113_ VPWR _1118_ VGND _1114_ _1116_ sg13g2_o21ai_1
X_4232_ _1046_ VPWR _1051_ VGND _1047_ _1049_ sg13g2_o21ai_1
Xclkbuf_leaf_4_clk clknet_4_1_0_clk clknet_leaf_4_clk VPWR VGND sg13g2_buf_8
X_4163_ VGND VPWR _0957_ _0981_ _0988_ _0983_ sg13g2_a21oi_1
X_3114_ _2708_ _2678_ _2706_ VPWR VGND sg13g2_xnor2_1
X_4094_ _0892_ VPWR _0922_ VGND _0890_ _0893_ sg13g2_o21ai_1
XFILLER_49_880 VPWR VGND sg13g2_decap_8
X_3045_ _2636_ VPWR _2641_ VGND _2637_ _2639_ sg13g2_o21ai_1
XFILLER_36_552 VPWR VGND sg13g2_decap_8
X_4996_ _1783_ net863 net802 VPWR VGND sg13g2_nand2_1
X_3947_ _0779_ net931 net991 VPWR VGND sg13g2_nand2_2
XFILLER_23_268 VPWR VGND sg13g2_fill_2
X_3878_ _0707_ VPWR _0712_ VGND _0708_ _0710_ sg13g2_o21ai_1
XFILLER_20_964 VPWR VGND sg13g2_decap_8
X_5617_ net328 mac2.sum_lvl3_ff\[34\] _2332_ VPWR VGND sg13g2_xor2_1
X_5548_ _2278_ mac2.sum_lvl2_ff\[34\] net527 VPWR VGND sg13g2_xnor2_1
X_5479_ _2223_ net284 net267 VPWR VGND sg13g2_nand2_1
XFILLER_42_533 VPWR VGND sg13g2_fill_1
XFILLER_42_588 VPWR VGND sg13g2_decap_8
XFILLER_6_423 VPWR VGND sg13g2_fill_2
XFILLER_6_489 VPWR VGND sg13g2_fill_1
XFILLER_38_828 VPWR VGND sg13g2_decap_8
XFILLER_46_894 VPWR VGND sg13g2_decap_8
X_4850_ _1645_ _1638_ _1647_ VPWR VGND sg13g2_xor2_1
X_3801_ _0638_ net998 net943 net1000 net940 VPWR VGND sg13g2_a22oi_1
X_4781_ _1580_ _1575_ _1579_ VPWR VGND sg13g2_nand2_1
XFILLER_21_739 VPWR VGND sg13g2_fill_1
XFILLER_33_599 VPWR VGND sg13g2_fill_1
X_6520_ net1056 VGND VPWR net14 DP_3.I_range.out_data\[3\] clknet_leaf_22_clk sg13g2_dfrbpq_1
X_3732_ _0558_ _0551_ _0560_ _0575_ VPWR VGND sg13g2_a21o_1
Xclkload20 VPWR clkload20/Y clknet_leaf_35_clk VGND sg13g2_inv_1
X_3663_ VGND VPWR _0472_ _0474_ _0509_ _0508_ sg13g2_a21oi_1
X_6451_ net1086 VGND VPWR net101 mac2.sum_lvl2_ff\[1\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_5402_ _2164_ mac1.sum_lvl2_ff\[34\] net390 VPWR VGND sg13g2_xnor2_1
X_6382_ net1084 VGND VPWR net402 mac2.products_ff\[69\] clknet_leaf_28_clk sg13g2_dfrbpq_1
XFILLER_47_1004 VPWR VGND sg13g2_decap_8
X_5333_ _2109_ net356 net286 VPWR VGND sg13g2_nand2_1
X_3594_ _0402_ VPWR _0441_ VGND _0357_ _0403_ sg13g2_o21ai_1
X_5264_ _2044_ _2036_ _2043_ VPWR VGND sg13g2_xnor2_1
X_5195_ _1951_ VPWR _1977_ VGND _1945_ _1952_ sg13g2_o21ai_1
X_4215_ _1033_ _1034_ _1035_ VPWR VGND sg13g2_nor2b_2
X_4146_ _0955_ _0947_ _0954_ _0972_ VPWR VGND sg13g2_a21o_1
XFILLER_18_27 VPWR VGND sg13g2_fill_2
X_4077_ _0895_ _0905_ _0906_ VPWR VGND sg13g2_nor2_1
X_3028_ _2623_ _2624_ _2625_ VPWR VGND sg13g2_nor2b_2
XFILLER_36_371 VPWR VGND sg13g2_fill_2
XFILLER_37_872 VPWR VGND sg13g2_decap_8
XFILLER_24_555 VPWR VGND sg13g2_fill_1
X_4979_ net808 net861 net812 _1767_ VPWR VGND net859 sg13g2_nand4_1
Xclkload3 clknet_4_5_0_clk clkload3/X VPWR VGND sg13g2_buf_8
XFILLER_46_113 VPWR VGND sg13g2_fill_1
XFILLER_19_349 VPWR VGND sg13g2_fill_2
XFILLER_46_179 VPWR VGND sg13g2_fill_2
XFILLER_15_500 VPWR VGND sg13g2_fill_2
XFILLER_28_894 VPWR VGND sg13g2_decap_8
XFILLER_43_897 VPWR VGND sg13g2_decap_8
XFILLER_6_297 VPWR VGND sg13g2_fill_2
XFILLER_3_982 VPWR VGND sg13g2_decap_8
XFILLER_2_470 VPWR VGND sg13g2_fill_2
X_4000_ _0831_ _0779_ _0828_ VPWR VGND sg13g2_xnor2_1
X_5951_ net997 _0183_ VPWR VGND sg13g2_buf_1
X_4902_ _1697_ _1661_ _1695_ VPWR VGND sg13g2_xnor2_1
XFILLER_34_853 VPWR VGND sg13g2_decap_8
X_5882_ net954 net771 _2564_ VPWR VGND sg13g2_nor2_1
X_4833_ _1616_ VPWR _1630_ VGND _1605_ _1617_ sg13g2_o21ai_1
X_4764_ _1563_ _1562_ _1559_ VPWR VGND sg13g2_nand2b_1
X_6503_ net1043 VGND VPWR net398 mac2.total_sum\[5\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_3715_ _0559_ _0551_ _0558_ VPWR VGND sg13g2_xnor2_1
X_6434_ net1102 VGND VPWR net233 mac2.sum_lvl1_ff\[41\] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_4695_ _1493_ _1494_ _1475_ _1496_ VPWR VGND sg13g2_nand3_1
X_3646_ _0466_ VPWR _0492_ VGND _0460_ _0467_ sg13g2_o21ai_1
X_3577_ _0422_ _0423_ _0405_ _0425_ VPWR VGND sg13g2_nand3_1
X_6365_ net1078 VGND VPWR _0084_ mac2.products_ff\[0\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_5316_ _2092_ _2086_ _2094_ VPWR VGND sg13g2_xor2_1
X_6296_ net1053 VGND VPWR net261 mac2.sum_lvl1_ff\[83\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_5247_ _2026_ _2027_ _2028_ VPWR VGND sg13g2_nor2_1
Xhold26 mac1.sum_lvl1_ff\[0\] VPWR VGND net66 sg13g2_dlygate4sd3_1
Xhold37 mac1.sum_lvl1_ff\[11\] VPWR VGND net77 sg13g2_dlygate4sd3_1
Xhold15 mac1.sum_lvl1_ff\[49\] VPWR VGND net55 sg13g2_dlygate4sd3_1
Xhold48 mac1.products_ff\[7\] VPWR VGND net88 sg13g2_dlygate4sd3_1
Xhold59 mac1.sum_lvl2_ff\[51\] VPWR VGND net99 sg13g2_dlygate4sd3_1
X_5178_ _1925_ _1960_ _1961_ VPWR VGND sg13g2_nor2_1
X_4129_ _0956_ _0947_ _0955_ VPWR VGND sg13g2_xnor2_1
XFILLER_16_308 VPWR VGND sg13g2_fill_1
XFILLER_28_179 VPWR VGND sg13g2_fill_1
XFILLER_12_514 VPWR VGND sg13g2_fill_2
XFILLER_8_518 VPWR VGND sg13g2_fill_2
XFILLER_40_889 VPWR VGND sg13g2_decap_8
XFILLER_3_267 VPWR VGND sg13g2_fill_2
Xfanout1013 net1014 net1013 VPWR VGND sg13g2_buf_8
Xfanout1002 net515 net1002 VPWR VGND sg13g2_buf_8
XFILLER_48_912 VPWR VGND sg13g2_decap_8
Xfanout1024 net317 net1024 VPWR VGND sg13g2_buf_8
Xfanout1035 net1036 net1035 VPWR VGND sg13g2_buf_8
Xfanout1046 net1047 net1046 VPWR VGND sg13g2_buf_8
XFILLER_0_996 VPWR VGND sg13g2_decap_8
Xfanout1068 net1069 net1068 VPWR VGND sg13g2_buf_8
Xfanout1079 net1080 net1079 VPWR VGND sg13g2_buf_1
Xfanout1057 net1058 net1057 VPWR VGND sg13g2_buf_8
XFILLER_48_989 VPWR VGND sg13g2_decap_8
XFILLER_47_466 VPWR VGND sg13g2_fill_1
XFILLER_31_856 VPWR VGND sg13g2_decap_8
X_3500_ _0350_ _0326_ _0349_ VPWR VGND sg13g2_xnor2_1
X_4480_ _1292_ _1291_ _1289_ VPWR VGND sg13g2_nand2b_1
X_3431_ _0283_ net1011 net963 net1013 net959 VPWR VGND sg13g2_a22oi_1
X_6150_ net1098 VGND VPWR net168 mac1.sum_lvl1_ff\[9\] clknet_leaf_52_clk sg13g2_dfrbpq_1
X_3362_ _2947_ _2948_ _2949_ VPWR VGND sg13g2_and2_1
XFILLER_44_1007 VPWR VGND sg13g2_decap_8
X_5101_ _1880_ _1884_ _1885_ VPWR VGND sg13g2_nor2_1
X_6081_ net1050 VGND VPWR _0066_ mac1.products_ff\[138\] clknet_leaf_66_clk sg13g2_dfrbpq_1
X_3293_ _2842_ VPWR _2882_ VGND _2839_ _2843_ sg13g2_o21ai_1
XFILLER_39_912 VPWR VGND sg13g2_decap_8
X_5032_ _1818_ _1813_ _1816_ VPWR VGND sg13g2_xnor2_1
Xheichips25_template_39 VPWR VGND uio_oe[6] sg13g2_tiehi
XFILLER_39_989 VPWR VGND sg13g2_decap_8
XFILLER_34_661 VPWR VGND sg13g2_fill_1
XFILLER_40_108 VPWR VGND sg13g2_fill_2
X_5934_ net835 net770 _2596_ VPWR VGND sg13g2_nor2_1
XFILLER_41_609 VPWR VGND sg13g2_fill_1
X_5865_ net1013 net774 _2554_ VPWR VGND sg13g2_nor2_1
X_4816_ _1612_ _1613_ _1614_ VPWR VGND sg13g2_nor2b_1
XFILLER_33_182 VPWR VGND sg13g2_fill_1
XFILLER_21_366 VPWR VGND sg13g2_fill_1
X_5796_ net886 net786 _2490_ VPWR VGND sg13g2_nor2_1
X_4747_ _1473_ VPWR _1547_ VGND _1543_ _1545_ sg13g2_o21ai_1
X_4678_ VGND VPWR _1479_ _1477_ _1444_ sg13g2_or2_1
X_3629_ _0440_ _0475_ _0476_ VPWR VGND sg13g2_nor2_1
X_6417_ net1100 VGND VPWR net240 mac2.sum_lvl1_ff\[4\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_6348_ net1059 VGND VPWR net227 mac2.sum_lvl3_ff\[35\] clknet_leaf_23_clk sg13g2_dfrbpq_1
Xoutput27 net27 uo_out[2] VPWR VGND sg13g2_buf_1
X_6279_ net1045 VGND VPWR net250 mac1.sum_lvl1_ff\[82\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_5_1023 VPWR VGND sg13g2_decap_4
XFILLER_44_403 VPWR VGND sg13g2_fill_2
XFILLER_17_617 VPWR VGND sg13g2_fill_2
XFILLER_45_959 VPWR VGND sg13g2_decap_8
XFILLER_13_812 VPWR VGND sg13g2_fill_2
XFILLER_12_333 VPWR VGND sg13g2_fill_2
XFILLER_4_510 VPWR VGND sg13g2_fill_2
XFILLER_47_230 VPWR VGND sg13g2_fill_2
XFILLER_36_915 VPWR VGND sg13g2_decap_8
XFILLER_47_285 VPWR VGND sg13g2_fill_2
X_3980_ _0807_ VPWR _0811_ VGND _0764_ _0809_ sg13g2_o21ai_1
XFILLER_43_491 VPWR VGND sg13g2_fill_2
X_5650_ _2356_ mac1.total_sum\[7\] mac2.total_sum\[7\] VPWR VGND sg13g2_nand2_1
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
XFILLER_31_675 VPWR VGND sg13g2_fill_1
X_4601_ _1384_ VPWR _1405_ VGND _1375_ _1385_ sg13g2_o21ai_1
X_5581_ _2295_ _2298_ net538 _2303_ VPWR VGND sg13g2_or3_1
X_4532_ _1330_ _1332_ _1342_ VPWR VGND sg13g2_and2_1
Xhold326 DP_4.matrix\[7\] VPWR VGND net366 sg13g2_dlygate4sd3_1
Xhold315 _0041_ VPWR VGND net355 sg13g2_dlygate4sd3_1
X_4463_ _1275_ _1267_ _1276_ VPWR VGND sg13g2_nor2b_1
Xhold304 _2334_ VPWR VGND net344 sg13g2_dlygate4sd3_1
Xhold337 _2135_ VPWR VGND net377 sg13g2_dlygate4sd3_1
X_3414_ _2991_ _2992_ _2994_ _2995_ VPWR VGND sg13g2_nor3_1
Xhold359 DP_2.matrix\[3\] VPWR VGND net399 sg13g2_dlygate4sd3_1
Xhold348 _2238_ VPWR VGND net388 sg13g2_dlygate4sd3_1
X_6202_ net1114 VGND VPWR net78 mac1.sum_lvl1_ff\[49\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_4394_ _1209_ _1204_ _1208_ VPWR VGND sg13g2_nand2_1
Xfanout806 net808 net806 VPWR VGND sg13g2_buf_2
Xfanout817 net500 net817 VPWR VGND sg13g2_buf_8
Xfanout839 net409 net839 VPWR VGND sg13g2_buf_8
X_3345_ _2913_ VPWR _2932_ VGND _2885_ _2911_ sg13g2_o21ai_1
Xfanout828 net400 net828 VPWR VGND sg13g2_buf_8
X_6133_ net1087 VGND VPWR _0224_ DP_3.matrix\[4\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_6064_ net1075 VGND VPWR _0175_ DP_1.matrix\[3\] clknet_leaf_56_clk sg13g2_dfrbpq_1
X_3276_ _2830_ _2864_ _2828_ _2866_ VPWR VGND sg13g2_nand3_1
X_5015_ _1800_ _1799_ _1761_ _1802_ VPWR VGND sg13g2_a21o_1
XFILLER_27_915 VPWR VGND sg13g2_decap_8
X_5917_ _2510_ _2512_ _2586_ VPWR VGND sg13g2_nor2b_1
X_5848_ _2541_ net797 net776 VPWR VGND sg13g2_nand2_1
XFILLER_42_48 VPWR VGND sg13g2_fill_1
X_5779_ DP_3.Q_range.out_data\[2\] DP_3.I_range.out_data\[2\] _2473_ VPWR VGND sg13g2_xor2_1
XFILLER_27_1013 VPWR VGND sg13g2_decap_8
XFILLER_29_252 VPWR VGND sg13g2_decap_4
XFILLER_44_211 VPWR VGND sg13g2_fill_2
XFILLER_17_425 VPWR VGND sg13g2_fill_1
XFILLER_32_417 VPWR VGND sg13g2_fill_2
XFILLER_12_152 VPWR VGND sg13g2_fill_2
XFILLER_34_1028 VPWR VGND sg13g2_fill_1
XFILLER_41_984 VPWR VGND sg13g2_decap_8
XFILLER_9_668 VPWR VGND sg13g2_fill_2
XFILLER_8_123 VPWR VGND sg13g2_fill_1
XFILLER_40_494 VPWR VGND sg13g2_fill_1
XFILLER_32_70 VPWR VGND sg13g2_fill_1
X_3130_ _2723_ _2685_ _2720_ VPWR VGND sg13g2_xnor2_1
X_3061_ _2656_ _2655_ _2652_ VPWR VGND sg13g2_nand2b_1
XFILLER_36_712 VPWR VGND sg13g2_fill_1
XFILLER_17_992 VPWR VGND sg13g2_decap_8
X_3963_ _0783_ VPWR _0795_ VGND _0791_ _0793_ sg13g2_o21ai_1
X_3894_ _0704_ VPWR _0727_ VGND _0669_ _0702_ sg13g2_o21ai_1
X_5702_ _2398_ _2396_ _2397_ VPWR VGND sg13g2_xnor2_1
X_5633_ _2343_ mac1.total_sum\[3\] mac2.total_sum\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_31_472 VPWR VGND sg13g2_fill_1
X_5564_ _2287_ VPWR _2289_ VGND _2286_ _2288_ sg13g2_o21ai_1
X_4515_ _1326_ _1291_ _1324_ VPWR VGND sg13g2_xnor2_1
Xhold101 mac1.products_ff\[82\] VPWR VGND net141 sg13g2_dlygate4sd3_1
Xhold112 mac1.products_ff\[142\] VPWR VGND net152 sg13g2_dlygate4sd3_1
Xhold134 mac1.sum_lvl1_ff\[41\] VPWR VGND net174 sg13g2_dlygate4sd3_1
Xhold123 mac2.products_ff\[70\] VPWR VGND net163 sg13g2_dlygate4sd3_1
X_5495_ net452 _2233_ _0042_ VPWR VGND sg13g2_xor2_1
Xhold145 mac1.sum_lvl2_ff\[53\] VPWR VGND net185 sg13g2_dlygate4sd3_1
Xhold156 mac2.products_ff\[75\] VPWR VGND net196 sg13g2_dlygate4sd3_1
Xhold167 mac2.products_ff\[69\] VPWR VGND net207 sg13g2_dlygate4sd3_1
X_4446_ _1245_ VPWR _1259_ VGND _1234_ _1246_ sg13g2_o21ai_1
Xhold178 mac1.sum_lvl1_ff\[50\] VPWR VGND net218 sg13g2_dlygate4sd3_1
Xhold189 mac2.sum_lvl1_ff\[76\] VPWR VGND net229 sg13g2_dlygate4sd3_1
X_4377_ _1192_ _1191_ _1188_ VPWR VGND sg13g2_nand2b_1
X_6116_ net1069 VGND VPWR _0213_ DP_2.matrix\[73\] clknet_leaf_65_clk sg13g2_dfrbpq_1
X_3328_ _2915_ _2907_ _2916_ VPWR VGND sg13g2_nor2b_1
X_3259_ VGND VPWR net920 net965 _2849_ _2818_ sg13g2_a21oi_1
X_6047_ net1114 VGND VPWR _0121_ mac1.products_ff\[82\] clknet_leaf_47_clk sg13g2_dfrbpq_1
XFILLER_2_1015 VPWR VGND sg13g2_decap_8
XFILLER_15_907 VPWR VGND sg13g2_fill_1
XFILLER_42_737 VPWR VGND sg13g2_fill_1
XFILLER_10_645 VPWR VGND sg13g2_decap_4
XFILLER_6_616 VPWR VGND sg13g2_fill_2
XFILLER_6_605 VPWR VGND sg13g2_decap_4
XFILLER_5_115 VPWR VGND sg13g2_fill_1
XFILLER_2_844 VPWR VGND sg13g2_fill_2
XFILLER_1_354 VPWR VGND sg13g2_fill_1
XFILLER_37_509 VPWR VGND sg13g2_decap_8
XFILLER_45_564 VPWR VGND sg13g2_fill_2
XFILLER_14_984 VPWR VGND sg13g2_decap_8
XFILLER_41_770 VPWR VGND sg13g2_fill_2
XFILLER_9_487 VPWR VGND sg13g2_fill_1
X_5280_ _2059_ _2056_ _0152_ VPWR VGND sg13g2_xor2_1
X_4300_ _1113_ _1114_ _1116_ _1117_ VPWR VGND sg13g2_or3_1
X_4231_ _1046_ _1047_ _1049_ _1050_ VPWR VGND sg13g2_or3_1
X_4162_ VGND VPWR _0970_ _0986_ _0987_ _0985_ sg13g2_a21oi_1
X_3113_ _2706_ _2678_ _2707_ VPWR VGND sg13g2_nor2b_1
X_4093_ _0900_ VPWR _0921_ VGND _0898_ _0901_ sg13g2_o21ai_1
X_3044_ _2636_ _2637_ _2639_ _2640_ VPWR VGND sg13g2_or3_1
XFILLER_36_542 VPWR VGND sg13g2_decap_4
X_4995_ _1782_ net863 net800 VPWR VGND sg13g2_nand2_1
X_3946_ _0778_ net997 net929 VPWR VGND sg13g2_nand2_1
XFILLER_20_943 VPWR VGND sg13g2_decap_8
X_3877_ _0707_ _0708_ _0710_ _0711_ VPWR VGND sg13g2_or3_1
X_5616_ mac2.sum_lvl3_ff\[34\] net328 _2331_ VPWR VGND sg13g2_nor2_1
X_5547_ _2274_ VPWR _2277_ VGND _2273_ _2275_ sg13g2_o21ai_1
X_5478_ net265 mac1.sum_lvl3_ff\[20\] _0016_ VPWR VGND sg13g2_xor2_1
X_4429_ _1241_ _1242_ _1243_ VPWR VGND sg13g2_nor2b_1
XFILLER_48_58 VPWR VGND sg13g2_fill_2
XFILLER_42_512 VPWR VGND sg13g2_fill_1
XFILLER_42_567 VPWR VGND sg13g2_decap_8
XFILLER_30_718 VPWR VGND sg13g2_fill_2
XFILLER_30_729 VPWR VGND sg13g2_decap_4
XFILLER_7_969 VPWR VGND sg13g2_decap_8
XFILLER_6_468 VPWR VGND sg13g2_fill_1
XFILLER_49_122 VPWR VGND sg13g2_decap_4
XFILLER_49_100 VPWR VGND sg13g2_decap_4
XFILLER_46_873 VPWR VGND sg13g2_decap_8
X_4780_ _1577_ _1578_ _1579_ VPWR VGND sg13g2_nor2_1
X_3800_ net940 net1000 net943 _0637_ VPWR VGND net998 sg13g2_nand4_1
XFILLER_33_556 VPWR VGND sg13g2_decap_4
X_3731_ _0574_ _0571_ _0108_ VPWR VGND sg13g2_xor2_1
X_3662_ _0506_ _0479_ _0508_ VPWR VGND sg13g2_xor2_1
X_6450_ net1084 VGND VPWR net59 mac2.sum_lvl2_ff\[0\] clknet_leaf_13_clk sg13g2_dfrbpq_1
Xclkload10 clknet_4_14_0_clk clkload10/Y VPWR VGND sg13g2_inv_4
Xclkload21 clknet_leaf_37_clk clkload21/Y VPWR VGND sg13g2_inv_4
X_3593_ _0430_ VPWR _0440_ VGND _0359_ _0431_ sg13g2_o21ai_1
X_5401_ _2160_ VPWR _2163_ VGND _2159_ _2161_ sg13g2_o21ai_1
X_6381_ net1079 VGND VPWR _0079_ mac2.products_ff\[68\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_5332_ _0155_ _2101_ _2108_ VPWR VGND sg13g2_xnor2_1
XFILLER_48_0 VPWR VGND sg13g2_fill_2
X_5263_ _2043_ _2037_ _2042_ VPWR VGND sg13g2_xnor2_1
X_5194_ _1974_ _1966_ _1976_ VPWR VGND sg13g2_xor2_1
X_4214_ _1013_ VPWR _1034_ VGND _1004_ _1014_ sg13g2_o21ai_1
X_4145_ _0959_ _0961_ _0971_ VPWR VGND sg13g2_and2_1
X_4076_ _0903_ _0896_ _0905_ VPWR VGND sg13g2_xor2_1
XFILLER_37_851 VPWR VGND sg13g2_decap_8
X_3027_ _2619_ VPWR _2624_ VGND _2620_ _2622_ sg13g2_o21ai_1
XFILLER_36_350 VPWR VGND sg13g2_fill_1
X_4978_ net811 net808 net861 net859 _1766_ VPWR VGND sg13g2_and4_1
X_3929_ _0761_ _0697_ _0762_ VPWR VGND sg13g2_xor2_1
Xclkload4 clknet_4_6_0_clk clkload4/X VPWR VGND sg13g2_buf_8
XFILLER_46_136 VPWR VGND sg13g2_fill_1
XFILLER_15_512 VPWR VGND sg13g2_decap_8
XFILLER_28_873 VPWR VGND sg13g2_decap_8
XFILLER_43_876 VPWR VGND sg13g2_decap_8
XFILLER_3_961 VPWR VGND sg13g2_decap_8
X_5950_ net999 _0182_ VPWR VGND sg13g2_buf_1
X_4901_ _1661_ _1695_ _1696_ VPWR VGND sg13g2_nor2b_1
XFILLER_34_832 VPWR VGND sg13g2_decap_8
X_5881_ VGND VPWR net771 _2563_ _0197_ _2562_ sg13g2_a21oi_1
X_4832_ _1602_ _1596_ _1604_ _1629_ VPWR VGND sg13g2_a21o_1
X_4763_ _1561_ _1510_ _1562_ VPWR VGND sg13g2_xor2_1
X_6502_ net1040 VGND VPWR net459 mac2.total_sum\[4\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_14_1026 VPWR VGND sg13g2_fill_2
X_3714_ _0558_ _0552_ _0557_ VPWR VGND sg13g2_xnor2_1
X_4694_ _1495_ _1475_ _1493_ _1494_ VPWR VGND sg13g2_and3_1
X_6433_ net1100 VGND VPWR net126 mac2.sum_lvl1_ff\[40\] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_3645_ _0489_ _0481_ _0491_ VPWR VGND sg13g2_xor2_1
X_3576_ _0424_ _0405_ _0422_ _0423_ VPWR VGND sg13g2_and3_1
X_6364_ net1046 VGND VPWR net440 mac1.total_sum\[15\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_5315_ _2093_ _2086_ _2092_ VPWR VGND sg13g2_nand2_1
X_6295_ net1052 VGND VPWR net215 mac2.sum_lvl1_ff\[82\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_5246_ VGND VPWR _1990_ _1992_ _2027_ _2024_ sg13g2_a21oi_1
Xhold27 mac1.products_ff\[137\] VPWR VGND net67 sg13g2_dlygate4sd3_1
Xhold38 mac1.products_ff\[81\] VPWR VGND net78 sg13g2_dlygate4sd3_1
Xhold16 mac2.sum_lvl1_ff\[11\] VPWR VGND net56 sg13g2_dlygate4sd3_1
Xhold49 mac1.sum_lvl2_ff\[41\] VPWR VGND net89 sg13g2_dlygate4sd3_1
X_5177_ _1960_ _1926_ _1958_ VPWR VGND sg13g2_xnor2_1
X_4128_ _0955_ _0919_ _0953_ VPWR VGND sg13g2_xnor2_1
XFILLER_45_37 VPWR VGND sg13g2_fill_2
X_4059_ _0874_ VPWR _0888_ VGND _0863_ _0875_ sg13g2_o21ai_1
XFILLER_12_548 VPWR VGND sg13g2_fill_2
XFILLER_40_868 VPWR VGND sg13g2_decap_8
Xfanout1003 net395 net1003 VPWR VGND sg13g2_buf_8
Xfanout1025 DP_3.matrix\[80\] net1025 VPWR VGND sg13g2_buf_1
Xfanout1014 net524 net1014 VPWR VGND sg13g2_buf_8
XFILLER_0_975 VPWR VGND sg13g2_decap_8
Xfanout1047 net1048 net1047 VPWR VGND sg13g2_buf_8
Xfanout1036 net403 net1036 VPWR VGND sg13g2_buf_2
Xfanout1069 net1091 net1069 VPWR VGND sg13g2_buf_8
Xfanout1058 net1059 net1058 VPWR VGND sg13g2_buf_8
XFILLER_48_968 VPWR VGND sg13g2_decap_8
XFILLER_34_117 VPWR VGND sg13g2_fill_1
XFILLER_16_887 VPWR VGND sg13g2_decap_4
XFILLER_31_835 VPWR VGND sg13g2_decap_8
XFILLER_37_1026 VPWR VGND sg13g2_fill_2
XFILLER_30_345 VPWR VGND sg13g2_fill_1
X_3430_ net958 net1013 net963 _0282_ VPWR VGND net1011 sg13g2_nand4_1
X_3361_ _2921_ _2923_ _2946_ _2948_ VPWR VGND sg13g2_or3_1
X_6080_ net1071 VGND VPWR _0189_ DP_1.matrix\[73\] clknet_leaf_61_clk sg13g2_dfrbpq_1
X_5100_ VGND VPWR _1884_ _1883_ _1882_ sg13g2_or2_1
X_3292_ _2881_ _2873_ _2878_ VPWR VGND sg13g2_xnor2_1
X_5031_ _1817_ _1816_ _1813_ VPWR VGND sg13g2_nand2b_1
XFILLER_38_412 VPWR VGND sg13g2_fill_2
XFILLER_39_968 VPWR VGND sg13g2_decap_8
XFILLER_47_990 VPWR VGND sg13g2_decap_8
XFILLER_25_139 VPWR VGND sg13g2_fill_1
X_5933_ _2595_ net836 net767 _0249_ VPWR VGND sg13g2_mux2_1
X_5864_ VGND VPWR net771 _2553_ _0174_ _2552_ sg13g2_a21oi_1
XFILLER_22_824 VPWR VGND sg13g2_decap_8
X_4815_ _1608_ VPWR _1613_ VGND _1610_ _1611_ sg13g2_o21ai_1
XFILLER_21_345 VPWR VGND sg13g2_fill_2
X_5795_ _2489_ net869 net775 VPWR VGND sg13g2_nand2_1
XFILLER_30_890 VPWR VGND sg13g2_decap_8
X_4746_ _1473_ _1543_ _1545_ _1546_ VPWR VGND sg13g2_or3_1
X_4677_ _1478_ net840 net896 VPWR VGND sg13g2_nand2_1
X_3628_ _0475_ _0441_ _0473_ VPWR VGND sg13g2_xnor2_1
X_6416_ net1099 VGND VPWR net183 mac2.sum_lvl1_ff\[3\] clknet_leaf_30_clk sg13g2_dfrbpq_1
Xoutput17 net17 uio_out[0] VPWR VGND sg13g2_buf_1
Xoutput28 net28 uo_out[3] VPWR VGND sg13g2_buf_1
X_6347_ net1059 VGND VPWR net60 mac2.sum_lvl3_ff\[34\] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_3559_ _0407_ net950 net1010 VPWR VGND sg13g2_nand2_2
X_6278_ net1047 VGND VPWR net119 mac1.sum_lvl1_ff\[81\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_5229_ _2010_ _2002_ _2007_ VPWR VGND sg13g2_xnor2_1
XFILLER_5_1002 VPWR VGND sg13g2_decap_8
XFILLER_45_938 VPWR VGND sg13g2_decap_8
XFILLER_24_150 VPWR VGND sg13g2_fill_2
XFILLER_13_846 VPWR VGND sg13g2_fill_2
XFILLER_13_868 VPWR VGND sg13g2_fill_2
XFILLER_8_327 VPWR VGND sg13g2_fill_1
XFILLER_13_879 VPWR VGND sg13g2_fill_1
XFILLER_46_80 VPWR VGND sg13g2_fill_1
XFILLER_44_993 VPWR VGND sg13g2_decap_8
XFILLER_16_684 VPWR VGND sg13g2_fill_1
XFILLER_31_665 VPWR VGND sg13g2_fill_1
X_4600_ _1404_ _1392_ _1403_ VPWR VGND sg13g2_xnor2_1
X_5580_ net538 VPWR _2302_ VGND _2295_ _2298_ sg13g2_o21ai_1
XFILLER_30_175 VPWR VGND sg13g2_fill_1
X_4531_ _1338_ _1316_ _1340_ _1341_ VPWR VGND sg13g2_a21o_1
XFILLER_7_360 VPWR VGND sg13g2_fill_2
Xhold316 mac1.sum_lvl2_ff\[19\] VPWR VGND net356 sg13g2_dlygate4sd3_1
Xhold305 _0054_ VPWR VGND net345 sg13g2_dlygate4sd3_1
X_4462_ _1275_ _1268_ _1274_ VPWR VGND sg13g2_xnor2_1
Xhold338 _0014_ VPWR VGND net378 sg13g2_dlygate4sd3_1
X_3413_ _2994_ net1013 net960 net1015 net959 VPWR VGND sg13g2_a22oi_1
Xhold327 mac1.sum_lvl3_ff\[13\] VPWR VGND net367 sg13g2_dlygate4sd3_1
Xhold349 _0043_ VPWR VGND net389 sg13g2_dlygate4sd3_1
X_6201_ net1114 VGND VPWR net162 mac1.sum_lvl1_ff\[48\] clknet_leaf_47_clk sg13g2_dfrbpq_1
X_4393_ _1206_ _1207_ _1208_ VPWR VGND sg13g2_nor2_1
Xfanout807 net808 net807 VPWR VGND sg13g2_buf_1
X_6132_ net1092 VGND VPWR net127 mac1.sum_lvl1_ff\[3\] clknet_leaf_55_clk sg13g2_dfrbpq_1
X_3344_ _2914_ _2908_ _2916_ _2931_ VPWR VGND sg13g2_a21o_1
Xfanout829 net830 net829 VPWR VGND sg13g2_buf_8
Xfanout818 net379 net818 VPWR VGND sg13g2_buf_8
X_6063_ net1072 VGND VPWR _0174_ DP_1.matrix\[2\] clknet_leaf_56_clk sg13g2_dfrbpq_1
X_3275_ VGND VPWR _2828_ _2830_ _2865_ _2864_ sg13g2_a21oi_1
X_5014_ _1799_ _1800_ _1761_ _1801_ VPWR VGND sg13g2_nand3_1
XFILLER_39_754 VPWR VGND sg13g2_fill_1
XFILLER_38_231 VPWR VGND sg13g2_fill_2
XFILLER_42_919 VPWR VGND sg13g2_decap_8
X_5916_ _2585_ net890 _2479_ VPWR VGND sg13g2_nand2_1
XFILLER_35_993 VPWR VGND sg13g2_decap_8
XFILLER_22_632 VPWR VGND sg13g2_decap_4
X_5847_ _2540_ _2522_ _2539_ VPWR VGND sg13g2_nand2b_1
X_5778_ _2472_ DP_3.I_range.out_data\[2\] DP_3.Q_range.out_data\[2\] VPWR VGND sg13g2_xnor2_1
X_4729_ net845 net888 net849 _1529_ VPWR VGND net1028 sg13g2_nand4_1
XFILLER_45_779 VPWR VGND sg13g2_fill_1
XFILLER_33_919 VPWR VGND sg13g2_decap_8
XFILLER_25_481 VPWR VGND sg13g2_fill_2
XFILLER_34_1007 VPWR VGND sg13g2_decap_8
XFILLER_40_462 VPWR VGND sg13g2_fill_2
XFILLER_41_963 VPWR VGND sg13g2_decap_8
X_3060_ _2654_ _2631_ _2655_ VPWR VGND sg13g2_xor2_1
XFILLER_24_919 VPWR VGND sg13g2_decap_8
XFILLER_36_768 VPWR VGND sg13g2_fill_1
XFILLER_17_971 VPWR VGND sg13g2_decap_8
X_3962_ _0783_ _0791_ _0793_ _0794_ VPWR VGND sg13g2_or3_1
X_5701_ _2397_ DP_1.I_range.out_data\[3\] DP_1.Q_range.out_data\[3\] VPWR VGND sg13g2_xnor2_1
X_3893_ _0718_ VPWR _0726_ VGND _0698_ _0719_ sg13g2_o21ai_1
XFILLER_32_985 VPWR VGND sg13g2_decap_8
X_5632_ VGND VPWR _2339_ _2341_ _2342_ _2340_ sg13g2_a21oi_1
X_5563_ net485 _2286_ _0057_ VPWR VGND sg13g2_xor2_1
X_4514_ _1291_ _1324_ _1325_ VPWR VGND sg13g2_nor2b_1
Xhold102 mac1.products_ff\[10\] VPWR VGND net142 sg13g2_dlygate4sd3_1
Xhold135 mac1.products_ff\[12\] VPWR VGND net175 sg13g2_dlygate4sd3_1
X_5494_ net451 mac2.sum_lvl2_ff\[23\] _2235_ VPWR VGND sg13g2_xor2_1
Xhold113 mac2.sum_lvl1_ff\[6\] VPWR VGND net153 sg13g2_dlygate4sd3_1
Xhold124 mac2.products_ff\[138\] VPWR VGND net164 sg13g2_dlygate4sd3_1
Xhold146 mac1.products_ff\[2\] VPWR VGND net186 sg13g2_dlygate4sd3_1
Xhold157 mac2.products_ff\[71\] VPWR VGND net197 sg13g2_dlygate4sd3_1
Xhold168 mac2.sum_lvl1_ff\[77\] VPWR VGND net208 sg13g2_dlygate4sd3_1
X_4445_ _1231_ _1225_ _1233_ _1258_ VPWR VGND sg13g2_a21o_1
Xhold179 mac1.products_ff\[77\] VPWR VGND net219 sg13g2_dlygate4sd3_1
X_4376_ _1190_ _1139_ _1191_ VPWR VGND sg13g2_xor2_1
X_6115_ net1067 VGND VPWR _0212_ DP_2.matrix\[72\] clknet_leaf_63_clk sg13g2_dfrbpq_1
X_3327_ _2915_ _2908_ _2914_ VPWR VGND sg13g2_xnor2_1
X_3258_ _2822_ VPWR _2848_ VGND _2816_ _2823_ sg13g2_o21ai_1
X_6046_ net1114 VGND VPWR _0120_ mac1.products_ff\[81\] clknet_leaf_39_clk sg13g2_dfrbpq_1
XFILLER_37_49 VPWR VGND sg13g2_fill_1
XFILLER_39_540 VPWR VGND sg13g2_fill_2
X_3189_ _2778_ _2779_ _2761_ _2781_ VPWR VGND sg13g2_nand3_1
XFILLER_39_584 VPWR VGND sg13g2_decap_8
XFILLER_26_223 VPWR VGND sg13g2_fill_1
XFILLER_27_768 VPWR VGND sg13g2_decap_4
XFILLER_23_985 VPWR VGND sg13g2_decap_8
XFILLER_6_639 VPWR VGND sg13g2_decap_8
XFILLER_18_702 VPWR VGND sg13g2_fill_1
XFILLER_40_1022 VPWR VGND sg13g2_decap_8
XFILLER_45_554 VPWR VGND sg13g2_fill_2
XFILLER_26_790 VPWR VGND sg13g2_fill_1
XFILLER_14_963 VPWR VGND sg13g2_decap_8
XFILLER_41_760 VPWR VGND sg13g2_fill_2
XFILLER_13_495 VPWR VGND sg13g2_fill_1
X_4230_ _1049_ net876 net830 net878 net827 VPWR VGND sg13g2_a22oi_1
X_4161_ _0986_ _0970_ _0121_ VPWR VGND sg13g2_xor2_1
X_3112_ _2706_ _2682_ _2705_ VPWR VGND sg13g2_xnor2_1
X_4092_ _0920_ _0919_ _0917_ VPWR VGND sg13g2_nand2b_1
X_3043_ _2639_ net972 net922 net976 net919 VPWR VGND sg13g2_a22oi_1
X_4994_ _1781_ net868 net798 VPWR VGND sg13g2_nand2_1
X_3945_ _0749_ VPWR _0777_ VGND _0740_ _0750_ sg13g2_o21ai_1
XFILLER_17_1013 VPWR VGND sg13g2_decap_8
XFILLER_23_248 VPWR VGND sg13g2_fill_2
X_3876_ _0710_ net990 net941 net991 net939 VPWR VGND sg13g2_a22oi_1
X_5615_ _2330_ mac2.sum_lvl3_ff\[34\] net328 VPWR VGND sg13g2_nand2_1
XFILLER_20_999 VPWR VGND sg13g2_decap_8
X_5546_ _0037_ _2273_ net543 VPWR VGND sg13g2_xnor2_1
X_5477_ _0022_ _2221_ net439 VPWR VGND sg13g2_xnor2_1
X_4428_ _1237_ VPWR _1242_ VGND _1239_ _1240_ sg13g2_o21ai_1
XFILLER_24_1017 VPWR VGND sg13g2_decap_8
X_4359_ _1102_ _1172_ _1174_ _1175_ VPWR VGND sg13g2_or3_1
XFILLER_24_1028 VPWR VGND sg13g2_fill_1
X_6029_ net1110 VGND VPWR _0108_ mac1.products_ff\[12\] clknet_leaf_44_clk sg13g2_dfrbpq_1
XFILLER_39_392 VPWR VGND sg13g2_fill_1
XFILLER_6_425 VPWR VGND sg13g2_fill_1
XFILLER_11_988 VPWR VGND sg13g2_decap_8
Xfanout990 net346 net990 VPWR VGND sg13g2_buf_8
XFILLER_38_92 VPWR VGND sg13g2_fill_2
XFILLER_33_546 VPWR VGND sg13g2_fill_2
XFILLER_14_782 VPWR VGND sg13g2_fill_2
X_3730_ VGND VPWR _0513_ _0572_ _0574_ _0573_ sg13g2_a21oi_1
X_3661_ _0507_ _0506_ _0479_ VPWR VGND sg13g2_nand2b_1
X_6380_ net1105 VGND VPWR _0144_ mac2.products_ff\[15\] clknet_leaf_33_clk sg13g2_dfrbpq_1
X_3592_ _0435_ VPWR _0439_ VGND _0392_ _0437_ sg13g2_o21ai_1
X_5400_ _0005_ _2159_ net461 VPWR VGND sg13g2_xnor2_1
Xclkload11 clknet_4_15_0_clk clkload11/X VPWR VGND sg13g2_buf_8
X_5331_ _2108_ _2102_ _2107_ VPWR VGND sg13g2_xnor2_1
XFILLER_6_992 VPWR VGND sg13g2_decap_8
X_5262_ _2039_ _2041_ _2042_ VPWR VGND sg13g2_nor2_1
X_4213_ _1033_ _1021_ _1032_ VPWR VGND sg13g2_xnor2_1
X_5193_ _1974_ _1966_ _1975_ VPWR VGND sg13g2_nor2b_1
X_4144_ _0967_ _0945_ _0969_ _0970_ VPWR VGND sg13g2_a21o_1
XFILLER_18_29 VPWR VGND sg13g2_fill_1
X_4075_ _0903_ _0896_ _0904_ VPWR VGND sg13g2_nor2b_1
X_3026_ _2619_ _2620_ _2622_ _2623_ VPWR VGND sg13g2_nor3_1
XFILLER_36_373 VPWR VGND sg13g2_fill_1
X_4977_ _1765_ net864 net804 VPWR VGND sg13g2_nand2_1
X_3928_ _0761_ _0758_ _0760_ VPWR VGND sg13g2_nand2_1
Xclkload5 clknet_4_7_0_clk clkload5/X VPWR VGND sg13g2_buf_8
X_3859_ _0116_ _0666_ _0693_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_417 VPWR VGND sg13g2_fill_2
X_5529_ _0034_ _2261_ _2262_ VPWR VGND sg13g2_xnor2_1
XFILLER_8_1011 VPWR VGND sg13g2_decap_8
XFILLER_28_852 VPWR VGND sg13g2_decap_8
XFILLER_46_159 VPWR VGND sg13g2_fill_2
XFILLER_27_395 VPWR VGND sg13g2_fill_2
XFILLER_43_855 VPWR VGND sg13g2_decap_8
XFILLER_23_590 VPWR VGND sg13g2_fill_2
XFILLER_3_940 VPWR VGND sg13g2_decap_8
XFILLER_37_126 VPWR VGND sg13g2_fill_2
X_4900_ _1695_ _1690_ _1693_ VPWR VGND sg13g2_xnor2_1
X_5880_ _2451_ _2447_ _2563_ VPWR VGND sg13g2_xor2_1
X_4831_ _1627_ _1625_ _0139_ VPWR VGND sg13g2_xor2_1
XFILLER_34_888 VPWR VGND sg13g2_decap_8
X_4762_ _1561_ net898 net834 VPWR VGND sg13g2_nand2_1
XFILLER_14_590 VPWR VGND sg13g2_fill_1
XFILLER_14_1005 VPWR VGND sg13g2_decap_8
X_6501_ net1039 VGND VPWR net486 mac2.total_sum\[3\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3713_ _0554_ _0556_ _0557_ VPWR VGND sg13g2_nor2_1
X_4693_ _1482_ VPWR _1494_ VGND _1490_ _1492_ sg13g2_o21ai_1
X_3644_ _0489_ _0481_ _0490_ VPWR VGND sg13g2_nor2b_1
X_6432_ net1099 VGND VPWR net197 mac2.sum_lvl1_ff\[39\] clknet_leaf_29_clk sg13g2_dfrbpq_1
X_3575_ _0411_ VPWR _0423_ VGND _0419_ _0421_ sg13g2_o21ai_1
X_6363_ net1045 VGND VPWR net479 mac1.total_sum\[14\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_5314_ _2092_ _2087_ _2090_ VPWR VGND sg13g2_xnor2_1
X_6294_ net1060 VGND VPWR net198 mac2.sum_lvl1_ff\[81\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_5245_ VPWR _2026_ _2025_ VGND sg13g2_inv_1
Xhold28 mac1.sum_lvl2_ff\[43\] VPWR VGND net68 sg13g2_dlygate4sd3_1
Xhold17 mac1.products_ff\[140\] VPWR VGND net57 sg13g2_dlygate4sd3_1
Xhold39 mac1.sum_lvl2_ff\[47\] VPWR VGND net79 sg13g2_dlygate4sd3_1
X_5176_ _1959_ _1926_ _1958_ VPWR VGND sg13g2_nand2b_1
X_4127_ _0919_ _0953_ _0954_ VPWR VGND sg13g2_nor2b_1
X_4058_ _0860_ _0854_ _0862_ _0887_ VPWR VGND sg13g2_a21o_1
X_3009_ _2608_ net981 net917 _0064_ VPWR VGND sg13g2_and3_2
Xclkbuf_leaf_63_clk clknet_4_2_0_clk clknet_leaf_63_clk VPWR VGND sg13g2_buf_8
XFILLER_36_181 VPWR VGND sg13g2_fill_1
XFILLER_40_803 VPWR VGND sg13g2_fill_2
XFILLER_12_505 VPWR VGND sg13g2_fill_1
XFILLER_12_516 VPWR VGND sg13g2_fill_1
XFILLER_12_527 VPWR VGND sg13g2_decap_4
XFILLER_40_847 VPWR VGND sg13g2_decap_8
XFILLER_3_269 VPWR VGND sg13g2_fill_1
Xfanout1004 net395 net1004 VPWR VGND sg13g2_buf_1
Xfanout1026 net313 net1026 VPWR VGND sg13g2_buf_8
Xfanout1015 net471 net1015 VPWR VGND sg13g2_buf_2
XFILLER_0_954 VPWR VGND sg13g2_decap_8
Xfanout1037 net522 net1037 VPWR VGND sg13g2_buf_8
Xfanout1048 net1063 net1048 VPWR VGND sg13g2_buf_8
Xfanout1059 net1063 net1059 VPWR VGND sg13g2_buf_8
XFILLER_48_947 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_54_clk clknet_4_8_0_clk clknet_leaf_54_clk VPWR VGND sg13g2_buf_8
XFILLER_37_1005 VPWR VGND sg13g2_decap_8
XFILLER_15_376 VPWR VGND sg13g2_fill_2
XFILLER_16_899 VPWR VGND sg13g2_fill_1
XFILLER_11_593 VPWR VGND sg13g2_fill_1
X_3360_ _2946_ VPWR _2947_ VGND _2921_ _2923_ sg13g2_o21ai_1
X_3291_ VGND VPWR _2880_ _2878_ _2873_ sg13g2_or2_1
X_5030_ _1815_ _1782_ _1816_ VPWR VGND sg13g2_xor2_1
XFILLER_39_947 VPWR VGND sg13g2_decap_8
XFILLER_20_1020 VPWR VGND sg13g2_decap_8
X_5932_ _2595_ _2522_ _2539_ VPWR VGND sg13g2_xnor2_1
XFILLER_19_671 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_45_clk clknet_4_11_0_clk clknet_leaf_45_clk VPWR VGND sg13g2_buf_8
X_5863_ _2553_ _2420_ _2422_ VPWR VGND sg13g2_xnor2_1
XFILLER_34_674 VPWR VGND sg13g2_fill_1
XFILLER_34_696 VPWR VGND sg13g2_fill_2
X_4814_ _1608_ _1610_ _1611_ _1612_ VPWR VGND sg13g2_nor3_1
XFILLER_22_847 VPWR VGND sg13g2_fill_2
X_5794_ _2488_ _2487_ net777 net775 net862 VPWR VGND sg13g2_a22oi_1
X_4745_ VGND VPWR _1541_ _1542_ _1545_ _1507_ sg13g2_a21oi_1
X_4676_ _1477_ net896 net838 VPWR VGND sg13g2_nand2_1
X_3627_ _0474_ _0441_ _0473_ VPWR VGND sg13g2_nand2b_1
X_6415_ net1085 VGND VPWR net138 mac2.sum_lvl1_ff\[2\] clknet_leaf_12_clk sg13g2_dfrbpq_1
Xoutput18 net18 uio_out[1] VPWR VGND sg13g2_buf_1
X_3558_ _0406_ net1014 net949 VPWR VGND sg13g2_nand2_1
Xoutput29 net29 uo_out[4] VPWR VGND sg13g2_buf_1
X_6346_ net1059 VGND VPWR net236 mac2.sum_lvl3_ff\[33\] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_3489_ _0335_ _0336_ _0338_ _0339_ VPWR VGND sg13g2_or3_1
X_6277_ net1041 VGND VPWR net201 mac1.sum_lvl1_ff\[80\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_5228_ VGND VPWR _2009_ _2007_ _2002_ sg13g2_or2_1
X_5159_ VGND VPWR _1942_ _1941_ _1892_ sg13g2_or2_1
XFILLER_45_917 VPWR VGND sg13g2_decap_8
XFILLER_44_405 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_36_clk clknet_4_15_0_clk clknet_leaf_36_clk VPWR VGND sg13g2_buf_8
XFILLER_37_490 VPWR VGND sg13g2_decap_8
XFILLER_13_814 VPWR VGND sg13g2_fill_1
XFILLER_24_162 VPWR VGND sg13g2_fill_2
XFILLER_40_655 VPWR VGND sg13g2_fill_2
XFILLER_4_512 VPWR VGND sg13g2_fill_1
XFILLER_4_567 VPWR VGND sg13g2_fill_1
XFILLER_47_287 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_27_clk clknet_4_7_0_clk clknet_leaf_27_clk VPWR VGND sg13g2_buf_8
XFILLER_44_972 VPWR VGND sg13g2_decap_8
XFILLER_43_460 VPWR VGND sg13g2_fill_2
X_4530_ _1340_ _1334_ _1339_ VPWR VGND sg13g2_nand2_1
XFILLER_7_372 VPWR VGND sg13g2_fill_2
Xhold317 _0007_ VPWR VGND net357 sg13g2_dlygate4sd3_1
Xhold306 DP_1.matrix\[42\] VPWR VGND net346 sg13g2_dlygate4sd3_1
X_4461_ _1273_ _1269_ _1274_ VPWR VGND sg13g2_xor2_1
X_3412_ net956 net1015 net960 _2993_ VPWR VGND net1013 sg13g2_nand4_1
X_6200_ net1115 VGND VPWR net170 mac1.sum_lvl1_ff\[47\] clknet_leaf_48_clk sg13g2_dfrbpq_1
Xhold328 _2215_ VPWR VGND net368 sg13g2_dlygate4sd3_1
Xhold339 DP_4.matrix\[41\] VPWR VGND net379 sg13g2_dlygate4sd3_1
X_6131_ net1088 VGND VPWR _0223_ DP_3.matrix\[3\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_4392_ _1207_ net1027 net826 net870 net823 VPWR VGND sg13g2_a22oi_1
Xfanout819 net820 net819 VPWR VGND sg13g2_buf_8
X_3343_ _2930_ _2927_ _0097_ VPWR VGND sg13g2_xor2_1
Xfanout808 net809 net808 VPWR VGND sg13g2_buf_2
X_6062_ net1070 VGND VPWR _0173_ DP_1.matrix\[1\] clknet_leaf_62_clk sg13g2_dfrbpq_2
X_3274_ _2862_ _2835_ _2864_ VPWR VGND sg13g2_xor2_1
XFILLER_23_0 VPWR VGND sg13g2_fill_1
X_5013_ _1798_ _1797_ _1780_ _1800_ VPWR VGND sg13g2_a21o_1
XFILLER_38_210 VPWR VGND sg13g2_fill_1
XFILLER_26_416 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_18_clk clknet_4_4_0_clk clknet_leaf_18_clk VPWR VGND sg13g2_buf_8
X_5915_ VGND VPWR net770 _2584_ _0226_ _2583_ sg13g2_a21oi_1
XFILLER_34_460 VPWR VGND sg13g2_fill_2
XFILLER_35_972 VPWR VGND sg13g2_decap_8
X_5846_ _2539_ _2538_ _2534_ VPWR VGND sg13g2_nand2b_1
XFILLER_10_817 VPWR VGND sg13g2_fill_1
X_5777_ _2471_ _2469_ _2470_ VPWR VGND sg13g2_xnor2_1
X_4728_ net850 net845 net888 net1028 _1528_ VPWR VGND sg13g2_and4_1
X_4659_ VGND VPWR _1458_ _1459_ _1461_ _1441_ sg13g2_a21oi_1
X_6329_ net1075 VGND VPWR net483 mac1.sum_lvl3_ff\[12\] clknet_leaf_59_clk sg13g2_dfrbpq_2
XFILLER_26_994 VPWR VGND sg13g2_decap_8
XFILLER_32_419 VPWR VGND sg13g2_fill_1
XFILLER_41_942 VPWR VGND sg13g2_decap_8
XFILLER_5_887 VPWR VGND sg13g2_fill_2
XFILLER_48_541 VPWR VGND sg13g2_fill_1
XFILLER_36_725 VPWR VGND sg13g2_fill_1
XFILLER_17_950 VPWR VGND sg13g2_decap_8
XFILLER_35_224 VPWR VGND sg13g2_fill_2
X_3961_ VGND VPWR _0789_ _0790_ _0793_ _0784_ sg13g2_a21oi_1
X_5700_ DP_1.Q_range.out_data\[2\] DP_1.I_range.out_data\[2\] _2396_ VPWR VGND sg13g2_nor2b_1
X_3892_ _0725_ _0724_ _0123_ VPWR VGND sg13g2_xor2_1
XFILLER_32_964 VPWR VGND sg13g2_decap_8
X_5631_ _2341_ _2339_ net27 VPWR VGND sg13g2_xor2_1
X_5562_ _2288_ mac2.sum_lvl3_ff\[23\] net484 VPWR VGND sg13g2_xnor2_1
X_4513_ _1324_ _1319_ _1322_ VPWR VGND sg13g2_xnor2_1
Xhold125 mac1.sum_lvl1_ff\[79\] VPWR VGND net165 sg13g2_dlygate4sd3_1
Xhold103 mac1.sum_lvl1_ff\[40\] VPWR VGND net143 sg13g2_dlygate4sd3_1
X_5493_ mac2.sum_lvl2_ff\[23\] mac2.sum_lvl2_ff\[4\] _2234_ VPWR VGND sg13g2_and2_1
Xhold114 mac2.sum_lvl1_ff\[81\] VPWR VGND net154 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_4_1_0_clk clknet_leaf_7_clk VPWR VGND sg13g2_buf_8
Xhold147 mac2.products_ff\[144\] VPWR VGND net187 sg13g2_dlygate4sd3_1
Xhold136 mac2.products_ff\[0\] VPWR VGND net176 sg13g2_dlygate4sd3_1
Xhold158 mac2.products_ff\[145\] VPWR VGND net198 sg13g2_dlygate4sd3_1
X_4444_ _1256_ _1254_ _0128_ VPWR VGND sg13g2_xor2_1
Xhold169 mac1.sum_lvl1_ff\[46\] VPWR VGND net209 sg13g2_dlygate4sd3_1
X_4375_ _1190_ net881 net817 VPWR VGND sg13g2_nand2_1
X_3326_ _2914_ _2909_ _2912_ VPWR VGND sg13g2_xnor2_1
X_6114_ net1068 VGND VPWR _0098_ mac1.products_ff\[149\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_6045_ net1115 VGND VPWR _0119_ mac1.products_ff\[80\] clknet_leaf_47_clk sg13g2_dfrbpq_1
X_3257_ _2845_ _2837_ _2847_ VPWR VGND sg13g2_xor2_1
XFILLER_39_530 VPWR VGND sg13g2_fill_1
XFILLER_39_552 VPWR VGND sg13g2_fill_2
X_3188_ _2780_ _2761_ _2778_ _2779_ VPWR VGND sg13g2_and3_1
XFILLER_41_216 VPWR VGND sg13g2_fill_1
XFILLER_23_964 VPWR VGND sg13g2_decap_8
X_5829_ _2519_ VPWR _2522_ VGND _2520_ _2521_ sg13g2_o21ai_1
XFILLER_6_618 VPWR VGND sg13g2_fill_1
XFILLER_2_846 VPWR VGND sg13g2_fill_1
XFILLER_40_1001 VPWR VGND sg13g2_decap_8
XFILLER_32_205 VPWR VGND sg13g2_fill_1
XFILLER_25_290 VPWR VGND sg13g2_fill_2
XFILLER_9_445 VPWR VGND sg13g2_fill_1
XFILLER_4_183 VPWR VGND sg13g2_fill_1
X_4160_ _0984_ _0971_ _0986_ VPWR VGND sg13g2_xor2_1
X_3111_ _2705_ _2702_ _2704_ VPWR VGND sg13g2_nand2_1
X_4091_ VGND VPWR _0919_ _0918_ _0867_ sg13g2_or2_1
XFILLER_49_894 VPWR VGND sg13g2_decap_8
X_3042_ net919 net975 net922 _2638_ VPWR VGND net972 sg13g2_nand4_1
XFILLER_17_791 VPWR VGND sg13g2_fill_1
X_4993_ _1771_ VPWR _1780_ VGND _1763_ _1772_ sg13g2_o21ai_1
X_3944_ _0776_ _0729_ _0775_ VPWR VGND sg13g2_xnor2_1
X_3875_ net938 net991 net941 _0709_ VPWR VGND net990 sg13g2_nand4_1
X_5614_ VGND VPWR _2325_ _2327_ _2329_ _2326_ sg13g2_a21oi_1
XFILLER_20_978 VPWR VGND sg13g2_decap_8
X_5545_ net542 mac2.sum_lvl2_ff\[33\] _2276_ VPWR VGND sg13g2_xor2_1
X_5476_ _2222_ mac1.sum_lvl3_ff\[35\] net438 VPWR VGND sg13g2_xnor2_1
X_4427_ _1237_ _1239_ _1240_ _1241_ VPWR VGND sg13g2_nor3_1
X_4358_ VGND VPWR _1170_ _1171_ _1174_ _1136_ sg13g2_a21oi_1
X_3309_ VPWR _2898_ _2897_ VGND sg13g2_inv_1
X_4289_ _1106_ net879 net820 VPWR VGND sg13g2_nand2_1
X_6028_ net1098 VGND VPWR _0107_ mac1.products_ff\[11\] clknet_leaf_45_clk sg13g2_dfrbpq_1
XFILLER_42_547 VPWR VGND sg13g2_decap_4
XFILLER_23_761 VPWR VGND sg13g2_fill_2
XFILLER_7_905 VPWR VGND sg13g2_fill_1
XFILLER_11_967 VPWR VGND sg13g2_decap_8
XFILLER_6_448 VPWR VGND sg13g2_fill_2
XFILLER_2_654 VPWR VGND sg13g2_decap_4
Xfanout980 net309 net980 VPWR VGND sg13g2_buf_2
Xfanout991 net992 net991 VPWR VGND sg13g2_buf_8
XFILLER_18_511 VPWR VGND sg13g2_fill_2
XFILLER_9_286 VPWR VGND sg13g2_fill_1
X_3660_ _0504_ _0480_ _0506_ VPWR VGND sg13g2_xor2_1
X_3591_ _0437_ _0392_ _0114_ VPWR VGND sg13g2_xor2_1
Xclkload12 clkload12/Y clknet_leaf_65_clk VPWR VGND sg13g2_inv_2
X_5330_ _2107_ _2093_ _2106_ VPWR VGND sg13g2_xnor2_1
XFILLER_6_971 VPWR VGND sg13g2_decap_8
XFILLER_47_1018 VPWR VGND sg13g2_decap_8
X_5261_ _2041_ net793 net857 net796 net855 VPWR VGND sg13g2_a22oi_1
XFILLER_48_2 VPWR VGND sg13g2_fill_1
X_4212_ _1032_ _1029_ _1031_ VPWR VGND sg13g2_nand2_1
X_5192_ _1974_ _1967_ _1973_ VPWR VGND sg13g2_xnor2_1
X_4143_ _0969_ _0963_ _0968_ VPWR VGND sg13g2_nand2_1
XFILLER_29_809 VPWR VGND sg13g2_fill_2
X_4074_ _0903_ _0897_ _0902_ VPWR VGND sg13g2_xnor2_1
X_3025_ _2622_ net976 net924 net980 net920 VPWR VGND sg13g2_a22oi_1
XFILLER_37_820 VPWR VGND sg13g2_fill_2
XFILLER_37_886 VPWR VGND sg13g2_decap_8
X_4976_ _1750_ VPWR _1764_ VGND _1748_ _1751_ sg13g2_o21ai_1
X_3927_ _0757_ _0756_ _0726_ _0760_ VPWR VGND sg13g2_a21o_1
X_3858_ _0690_ _0664_ _0693_ VPWR VGND sg13g2_xor2_1
Xclkload6 clknet_4_9_0_clk clkload6/X VPWR VGND sg13g2_buf_8
X_3789_ net943 net1002 net940 net1000 _0627_ VPWR VGND sg13g2_and4_1
X_5528_ _2262_ _2255_ _2259_ VPWR VGND sg13g2_nand2_1
X_5459_ _2203_ VPWR _2208_ VGND _2199_ _2202_ sg13g2_o21ai_1
XFILLER_15_536 VPWR VGND sg13g2_fill_1
XFILLER_15_547 VPWR VGND sg13g2_decap_4
XFILLER_6_278 VPWR VGND sg13g2_fill_2
XFILLER_3_996 VPWR VGND sg13g2_decap_8
XFILLER_34_867 VPWR VGND sg13g2_decap_8
X_4830_ _1625_ _1627_ _1628_ VPWR VGND sg13g2_nor2_1
X_4761_ _1560_ net898 net832 VPWR VGND sg13g2_nand2_1
X_6500_ net1039 VGND VPWR net475 mac2.total_sum\[2\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_14_1028 VPWR VGND sg13g2_fill_1
X_3712_ _0556_ net945 DP_1.matrix\[5\] net947 net1008 VPWR VGND sg13g2_a22oi_1
X_4692_ _1482_ _1490_ _1492_ _1493_ VPWR VGND sg13g2_or3_1
X_3643_ _0489_ _0482_ _0488_ VPWR VGND sg13g2_xnor2_1
X_6431_ net1085 VGND VPWR net163 mac2.sum_lvl1_ff\[38\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_6362_ net1045 VGND VPWR net369 mac1.total_sum\[13\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_5313_ _2091_ _2090_ _2087_ VPWR VGND sg13g2_nand2b_1
X_3574_ _0411_ _0419_ _0421_ _0422_ VPWR VGND sg13g2_or3_1
X_6293_ net1060 VGND VPWR net187 mac2.sum_lvl1_ff\[80\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_5244_ _1992_ _2024_ _1990_ _2025_ VPWR VGND sg13g2_nand3_1
Xhold18 mac1.sum_lvl1_ff\[13\] VPWR VGND net58 sg13g2_dlygate4sd3_1
Xhold29 mac2.sum_lvl2_ff\[48\] VPWR VGND net69 sg13g2_dlygate4sd3_1
X_5175_ _1958_ _1927_ _1956_ VPWR VGND sg13g2_xnor2_1
X_4126_ _0953_ _0948_ _0951_ VPWR VGND sg13g2_xnor2_1
XFILLER_29_639 VPWR VGND sg13g2_fill_2
X_4057_ _0885_ _0883_ _0117_ VPWR VGND sg13g2_xor2_1
X_3008_ net984 net923 _0064_ VPWR VGND sg13g2_and2_1
XFILLER_40_826 VPWR VGND sg13g2_decap_8
X_4959_ _1748_ net867 net805 VPWR VGND sg13g2_nand2_1
Xfanout1027 DP_3.matrix\[44\] net1027 VPWR VGND sg13g2_buf_1
Xfanout1016 DP_1.matrix\[2\] net1016 VPWR VGND sg13g2_buf_8
XFILLER_0_933 VPWR VGND sg13g2_decap_8
Xfanout1038 DP_1.matrix\[8\] net1038 VPWR VGND sg13g2_buf_1
Xfanout1005 net1006 net1005 VPWR VGND sg13g2_buf_8
XFILLER_48_926 VPWR VGND sg13g2_decap_8
Xfanout1049 net1050 net1049 VPWR VGND sg13g2_buf_8
XFILLER_15_311 VPWR VGND sg13g2_fill_2
XFILLER_27_160 VPWR VGND sg13g2_fill_1
XFILLER_37_1028 VPWR VGND sg13g2_fill_1
XFILLER_42_163 VPWR VGND sg13g2_fill_2
XFILLER_15_388 VPWR VGND sg13g2_fill_2
X_3290_ _2873_ _2878_ _2879_ VPWR VGND sg13g2_and2_1
XFILLER_39_926 VPWR VGND sg13g2_decap_8
X_5931_ VGND VPWR _2478_ _2594_ _0248_ _2593_ sg13g2_a21oi_1
X_5862_ net1015 net771 _2552_ VPWR VGND sg13g2_nor2_1
X_4813_ _1611_ net888 net840 net891 net838 VPWR VGND sg13g2_a22oi_1
X_5793_ net880 net897 net786 _2487_ VPWR VGND sg13g2_mux2_1
XFILLER_21_347 VPWR VGND sg13g2_fill_1
X_4744_ _1541_ _1542_ _1507_ _1544_ VPWR VGND sg13g2_nand3_1
XFILLER_31_19 VPWR VGND sg13g2_fill_2
X_4675_ _1476_ net900 net836 VPWR VGND sg13g2_nand2_1
X_3626_ _0473_ _0442_ _0471_ VPWR VGND sg13g2_xnor2_1
X_6414_ net1084 VGND VPWR net51 mac2.sum_lvl1_ff\[1\] clknet_leaf_12_clk sg13g2_dfrbpq_1
Xoutput19 net19 uio_out[2] VPWR VGND sg13g2_buf_1
X_3557_ _0377_ VPWR _0405_ VGND _0368_ _0378_ sg13g2_o21ai_1
X_6345_ net1055 VGND VPWR net129 mac2.sum_lvl3_ff\[32\] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_6276_ net1042 VGND VPWR net145 mac1.sum_lvl1_ff\[79\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_5227_ _2002_ _2007_ _2008_ VPWR VGND sg13g2_and2_1
X_3488_ _0338_ net1007 net961 net1009 net958 VPWR VGND sg13g2_a22oi_1
X_5158_ _1941_ net802 net854 VPWR VGND sg13g2_nand2_1
XFILLER_29_425 VPWR VGND sg13g2_fill_2
X_4109_ _0935_ _0934_ _0937_ VPWR VGND sg13g2_xor2_1
X_5089_ _1874_ _1871_ _1873_ VPWR VGND sg13g2_nand2_1
XFILLER_24_152 VPWR VGND sg13g2_fill_1
XFILLER_25_686 VPWR VGND sg13g2_decap_8
XFILLER_12_325 VPWR VGND sg13g2_fill_2
XFILLER_0_763 VPWR VGND sg13g2_fill_2
XFILLER_29_981 VPWR VGND sg13g2_decap_8
XFILLER_36_929 VPWR VGND sg13g2_decap_8
XFILLER_44_951 VPWR VGND sg13g2_decap_8
XFILLER_15_174 VPWR VGND sg13g2_fill_1
XFILLER_11_1009 VPWR VGND sg13g2_decap_8
XFILLER_8_896 VPWR VGND sg13g2_fill_2
XFILLER_7_362 VPWR VGND sg13g2_fill_1
Xhold307 DP_2.matrix\[77\] VPWR VGND net347 sg13g2_dlygate4sd3_1
X_4460_ _1273_ _1227_ _1271_ VPWR VGND sg13g2_xnor2_1
X_3411_ DP_2.matrix\[0\] net956 net1015 net1013 _2992_ VPWR VGND sg13g2_and4_1
Xhold318 mac1.sum_lvl3_ff\[29\] VPWR VGND net358 sg13g2_dlygate4sd3_1
Xhold329 _0020_ VPWR VGND net369 sg13g2_dlygate4sd3_1
X_4391_ net826 net824 net870 net1026 _1206_ VPWR VGND sg13g2_and4_1
X_3342_ VGND VPWR _2869_ _2928_ _2930_ _2929_ sg13g2_a21oi_1
X_6130_ net1088 VGND VPWR _0222_ DP_3.matrix\[2\] clknet_leaf_28_clk sg13g2_dfrbpq_1
Xfanout809 net810 net809 VPWR VGND sg13g2_buf_1
X_6061_ net1073 VGND VPWR _0172_ DP_1.matrix\[0\] clknet_leaf_61_clk sg13g2_dfrbpq_1
X_3273_ _2863_ _2862_ _2835_ VPWR VGND sg13g2_nand2b_1
X_5012_ _1797_ _1798_ _1780_ _1799_ VPWR VGND sg13g2_nand3_1
XFILLER_16_0 VPWR VGND sg13g2_fill_1
XFILLER_38_233 VPWR VGND sg13g2_fill_1
XFILLER_38_244 VPWR VGND sg13g2_fill_2
XFILLER_27_929 VPWR VGND sg13g2_decap_8
XFILLER_35_951 VPWR VGND sg13g2_decap_8
X_5914_ _2509_ _2505_ _2584_ VPWR VGND sg13g2_xor2_1
X_5845_ _2535_ VPWR _2538_ VGND _2536_ _2537_ sg13g2_o21ai_1
XFILLER_21_111 VPWR VGND sg13g2_fill_1
XFILLER_42_29 VPWR VGND sg13g2_decap_4
X_5776_ _2470_ DP_3.I_range.out_data\[2\] DP_3.Q_range.out_data\[2\] VPWR VGND sg13g2_nand2b_1
X_4727_ _1527_ net842 net891 VPWR VGND sg13g2_nand2_1
X_4658_ _1458_ _1459_ _1441_ _1460_ VPWR VGND sg13g2_nand3_1
X_3609_ _0456_ net952 net1008 VPWR VGND sg13g2_nand2_1
X_4589_ _1379_ VPWR _1393_ VGND _1377_ _1380_ sg13g2_o21ai_1
X_6328_ net1046 VGND VPWR _0002_ mac1.sum_lvl3_ff\[11\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_27_1027 VPWR VGND sg13g2_fill_2
X_6259_ net1061 VGND VPWR net195 mac2.sum_lvl2_ff\[44\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_17_406 VPWR VGND sg13g2_fill_2
XFILLER_17_439 VPWR VGND sg13g2_fill_2
XFILLER_16_30 VPWR VGND sg13g2_fill_1
XFILLER_26_973 VPWR VGND sg13g2_decap_8
XFILLER_41_921 VPWR VGND sg13g2_decap_8
XFILLER_12_133 VPWR VGND sg13g2_fill_2
XFILLER_32_40 VPWR VGND sg13g2_fill_1
XFILLER_41_998 VPWR VGND sg13g2_decap_8
XFILLER_5_866 VPWR VGND sg13g2_fill_1
XFILLER_35_214 VPWR VGND sg13g2_fill_2
X_3960_ _0789_ _0790_ _0784_ _0792_ VPWR VGND sg13g2_nand3_1
XFILLER_16_461 VPWR VGND sg13g2_fill_2
XFILLER_32_943 VPWR VGND sg13g2_decap_8
X_3891_ _0691_ VPWR _0725_ VGND _0666_ _0692_ sg13g2_o21ai_1
X_5630_ mac2.total_sum\[2\] mac1.total_sum\[2\] _2341_ VPWR VGND sg13g2_xor2_1
XFILLER_31_486 VPWR VGND sg13g2_fill_2
X_5561_ _2287_ mac2.sum_lvl3_ff\[23\] mac2.sum_lvl3_ff\[3\] VPWR VGND sg13g2_nand2_1
X_4512_ _1323_ _1322_ _1319_ VPWR VGND sg13g2_nand2b_1
X_5492_ _2231_ VPWR _2233_ VGND _2230_ _2232_ sg13g2_o21ai_1
Xhold104 mac1.products_ff\[6\] VPWR VGND net144 sg13g2_dlygate4sd3_1
Xhold115 mac1.products_ff\[136\] VPWR VGND net155 sg13g2_dlygate4sd3_1
Xhold126 mac1.products_ff\[147\] VPWR VGND net166 sg13g2_dlygate4sd3_1
Xhold137 mac1.sum_lvl1_ff\[80\] VPWR VGND net177 sg13g2_dlygate4sd3_1
Xhold159 mac1.products_ff\[69\] VPWR VGND net199 sg13g2_dlygate4sd3_1
X_4443_ _1254_ _1256_ _1257_ VPWR VGND sg13g2_nor2_1
Xhold148 mac2.products_ff\[78\] VPWR VGND net188 sg13g2_dlygate4sd3_1
X_4374_ _1189_ net881 net815 VPWR VGND sg13g2_nand2_1
X_3325_ _2913_ _2912_ _2909_ VPWR VGND sg13g2_nand2b_1
X_6113_ net1110 VGND VPWR _0211_ DP_2.matrix\[43\] clknet_leaf_45_clk sg13g2_dfrbpq_2
X_3256_ _2845_ _2837_ _2846_ VPWR VGND sg13g2_nor2b_1
X_6044_ net1113 VGND VPWR _0118_ mac1.products_ff\[79\] clknet_leaf_48_clk sg13g2_dfrbpq_1
X_3187_ _2767_ VPWR _2779_ VGND _2775_ _2777_ sg13g2_o21ai_1
XFILLER_26_269 VPWR VGND sg13g2_fill_2
XFILLER_23_943 VPWR VGND sg13g2_decap_8
XFILLER_22_431 VPWR VGND sg13g2_fill_1
X_5828_ net779 VPWR _2521_ VGND net836 net785 sg13g2_o21ai_1
X_5759_ _2454_ _2453_ net782 net781 DP_2.matrix\[74\] VPWR VGND sg13g2_a22oi_1
XFILLER_14_943 VPWR VGND sg13g2_decap_8
XFILLER_41_751 VPWR VGND sg13g2_fill_1
XFILLER_14_998 VPWR VGND sg13g2_decap_8
XFILLER_5_674 VPWR VGND sg13g2_fill_2
XFILLER_4_173 VPWR VGND sg13g2_fill_2
XFILLER_4_195 VPWR VGND sg13g2_fill_2
X_3110_ _2701_ _2700_ _2683_ _2704_ VPWR VGND sg13g2_a21o_1
X_4090_ _0918_ net929 net1036 VPWR VGND sg13g2_nand2_1
X_3041_ net922 net917 net975 net972 _2637_ VPWR VGND sg13g2_and4_1
X_4992_ _1778_ _1758_ _0093_ VPWR VGND sg13g2_xor2_1
X_3943_ _0775_ _0766_ _0773_ VPWR VGND sg13g2_xnor2_1
X_3874_ net941 DP_2.matrix\[37\] net992 net990 _0708_ VPWR VGND sg13g2_and4_1
XFILLER_20_957 VPWR VGND sg13g2_decap_8
X_5613_ _0052_ _2325_ net469 VPWR VGND sg13g2_xnor2_1
X_5544_ mac2.sum_lvl2_ff\[33\] mac2.sum_lvl2_ff\[14\] _2275_ VPWR VGND sg13g2_nor2_1
X_5475_ _2216_ VPWR _2221_ VGND _2217_ _2220_ sg13g2_o21ai_1
X_4426_ _1240_ net870 net821 net874 net819 VPWR VGND sg13g2_a22oi_1
X_4357_ _1170_ _1171_ _1136_ _1173_ VPWR VGND sg13g2_nand3_1
X_3308_ _2863_ _2896_ _2861_ _2897_ VPWR VGND sg13g2_nand3_1
X_4288_ _1105_ net883 DP_4.matrix\[41\] VPWR VGND sg13g2_nand2_1
X_3239_ _2830_ _2797_ _2829_ VPWR VGND sg13g2_nand2b_1
X_6027_ net1098 VGND VPWR _0106_ mac1.products_ff\[10\] clknet_leaf_45_clk sg13g2_dfrbpq_1
XFILLER_42_504 VPWR VGND sg13g2_fill_2
XFILLER_42_526 VPWR VGND sg13g2_decap_8
XFILLER_14_228 VPWR VGND sg13g2_fill_1
Xhold490 _2131_ VPWR VGND net530 sg13g2_dlygate4sd3_1
XFILLER_49_114 VPWR VGND sg13g2_decap_4
Xfanout970 net971 net970 VPWR VGND sg13g2_buf_1
XFILLER_49_158 VPWR VGND sg13g2_fill_2
Xfanout981 net983 net981 VPWR VGND sg13g2_buf_8
Xfanout992 net993 net992 VPWR VGND sg13g2_buf_1
XFILLER_46_887 VPWR VGND sg13g2_decap_8
XFILLER_14_784 VPWR VGND sg13g2_fill_1
XFILLER_9_232 VPWR VGND sg13g2_fill_1
XFILLER_13_283 VPWR VGND sg13g2_fill_2
X_3590_ _0390_ _0391_ _0435_ _0436_ _0438_ VPWR VGND sg13g2_and4_1
Xclkload13 VPWR clkload13/Y clknet_leaf_28_clk VGND sg13g2_inv_1
XFILLER_6_950 VPWR VGND sg13g2_decap_8
X_5260_ VGND VPWR _2040_ _2038_ _2014_ sg13g2_or2_1
XFILLER_5_493 VPWR VGND sg13g2_fill_2
X_4211_ _1028_ _1027_ _1022_ _1031_ VPWR VGND sg13g2_a21o_1
X_5191_ _1972_ _1968_ _1973_ VPWR VGND sg13g2_xor2_1
X_4142_ _0968_ _0941_ _0964_ VPWR VGND sg13g2_nand2_1
X_4073_ _0901_ _0898_ _0902_ VPWR VGND sg13g2_xor2_1
X_3024_ net920 net978 net924 _2621_ VPWR VGND net976 sg13g2_nand4_1
XFILLER_37_865 VPWR VGND sg13g2_decap_8
X_4975_ VPWR _1763_ _1762_ VGND sg13g2_inv_1
X_3926_ VGND VPWR _0756_ _0757_ _0759_ _0726_ sg13g2_a21oi_1
X_3857_ VGND VPWR _0688_ _0689_ _0692_ _0664_ sg13g2_a21oi_1
Xclkload7 clknet_4_10_0_clk clkload7/X VPWR VGND sg13g2_buf_8
X_3788_ _0626_ net1003 net936 VPWR VGND sg13g2_nand2_1
XFILLER_30_1023 VPWR VGND sg13g2_decap_4
X_5527_ _2261_ mac2.sum_lvl2_ff\[30\] mac2.sum_lvl2_ff\[11\] VPWR VGND sg13g2_xnor2_1
XFILLER_3_419 VPWR VGND sg13g2_fill_1
X_5458_ mac1.sum_lvl3_ff\[12\] mac1.sum_lvl3_ff\[32\] _2207_ VPWR VGND sg13g2_xor2_1
X_5389_ VPWR VGND _2153_ _2152_ _2144_ mac1.sum_lvl2_ff\[30\] _2154_ mac1.sum_lvl2_ff\[11\]
+ sg13g2_a221oi_1
X_4409_ _1212_ VPWR _1223_ VGND _1196_ _1213_ sg13g2_o21ai_1
XFILLER_28_887 VPWR VGND sg13g2_decap_8
XFILLER_11_710 VPWR VGND sg13g2_fill_2
XFILLER_6_224 VPWR VGND sg13g2_fill_1
XFILLER_3_975 VPWR VGND sg13g2_decap_8
XFILLER_49_93 VPWR VGND sg13g2_decap_8
XFILLER_19_876 VPWR VGND sg13g2_fill_2
XFILLER_34_846 VPWR VGND sg13g2_decap_8
X_4760_ _1559_ net902 net1023 VPWR VGND sg13g2_nand2_1
X_3711_ VGND VPWR _0555_ _0553_ _0529_ sg13g2_or2_1
X_4691_ VGND VPWR _1488_ _1489_ _1492_ _1483_ sg13g2_a21oi_1
X_3642_ _0487_ _0483_ _0488_ VPWR VGND sg13g2_xor2_1
X_6430_ net1083 VGND VPWR net207 mac2.sum_lvl1_ff\[37\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_6361_ net1045 VGND VPWR _0019_ mac1.total_sum\[12\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_5312_ _2089_ _2063_ _2090_ VPWR VGND sg13g2_xor2_1
X_3573_ VGND VPWR _0417_ _0418_ _0421_ _0412_ sg13g2_a21oi_1
XFILLER_46_0 VPWR VGND sg13g2_decap_8
X_6292_ net1060 VGND VPWR net232 mac2.sum_lvl1_ff\[79\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_5243_ _2022_ _2000_ _2024_ VPWR VGND sg13g2_xor2_1
Xhold19 mac2.sum_lvl1_ff\[0\] VPWR VGND net59 sg13g2_dlygate4sd3_1
X_5174_ _1957_ _1927_ _1956_ VPWR VGND sg13g2_nand2_1
X_4125_ _0952_ _0951_ _0948_ VPWR VGND sg13g2_nand2b_1
X_4056_ _0883_ _0885_ _0886_ VPWR VGND sg13g2_nor2_1
XFILLER_37_640 VPWR VGND sg13g2_fill_2
X_3007_ VPWR _2607_ net1026 VGND sg13g2_inv_1
XFILLER_25_824 VPWR VGND sg13g2_fill_1
XFILLER_40_805 VPWR VGND sg13g2_fill_1
X_4958_ VGND VPWR _1747_ _1742_ _1740_ sg13g2_or2_1
X_3909_ _0742_ net935 net991 VPWR VGND sg13g2_nand2_1
X_4889_ VGND VPWR _1623_ _1653_ _1685_ _1655_ sg13g2_a21oi_1
XFILLER_0_912 VPWR VGND sg13g2_decap_8
Xfanout1028 net536 net1028 VPWR VGND sg13g2_buf_8
Xfanout1017 net1018 net1017 VPWR VGND sg13g2_buf_8
Xfanout1006 net447 net1006 VPWR VGND sg13g2_buf_8
XFILLER_48_905 VPWR VGND sg13g2_decap_8
XFILLER_47_404 VPWR VGND sg13g2_fill_2
Xfanout1039 net1040 net1039 VPWR VGND sg13g2_buf_8
XFILLER_0_989 VPWR VGND sg13g2_decap_8
XFILLER_19_96 VPWR VGND sg13g2_fill_2
XFILLER_28_684 VPWR VGND sg13g2_fill_2
XFILLER_15_334 VPWR VGND sg13g2_fill_2
XFILLER_31_849 VPWR VGND sg13g2_decap_8
XFILLER_39_905 VPWR VGND sg13g2_decap_8
X_5930_ _2538_ _2534_ _2594_ VPWR VGND sg13g2_xor2_1
X_5861_ VGND VPWR net771 _2551_ _0173_ _2550_ sg13g2_a21oi_1
X_5792_ _2483_ VPWR _2486_ VGND _2484_ _2485_ sg13g2_o21ai_1
X_4812_ net840 net837 net891 net888 _1610_ VPWR VGND sg13g2_and4_1
XFILLER_22_849 VPWR VGND sg13g2_fill_1
X_4743_ _1543_ _1507_ _1541_ _1542_ VPWR VGND sg13g2_and3_1
X_6413_ net1084 VGND VPWR net176 mac2.sum_lvl1_ff\[0\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_4674_ _1457_ _1447_ _1455_ _1475_ VPWR VGND sg13g2_a21o_1
X_3625_ _0472_ _0442_ _0471_ VPWR VGND sg13g2_nand2_1
X_3556_ _0404_ _0357_ _0403_ VPWR VGND sg13g2_xnor2_1
X_6344_ net1054 VGND VPWR net110 mac2.sum_lvl3_ff\[31\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_6275_ net1064 VGND VPWR net152 mac1.sum_lvl1_ff\[78\] clknet_leaf_65_clk sg13g2_dfrbpq_1
X_5226_ _2006_ _2003_ _2007_ VPWR VGND sg13g2_xor2_1
X_3487_ net957 net1009 net961 _0337_ VPWR VGND net1007 sg13g2_nand4_1
X_5157_ _1940_ net858 net798 VPWR VGND sg13g2_nand2_1
XFILLER_5_1027 VPWR VGND sg13g2_fill_2
XFILLER_5_1016 VPWR VGND sg13g2_decap_8
X_4108_ _0935_ _0934_ _0936_ VPWR VGND sg13g2_nor2b_1
X_5088_ _1870_ _1869_ _1839_ _1873_ VPWR VGND sg13g2_a21o_1
X_4039_ _0869_ net986 net934 net990 net931 VPWR VGND sg13g2_a22oi_1
XFILLER_38_982 VPWR VGND sg13g2_decap_8
XFILLER_13_838 VPWR VGND sg13g2_fill_2
XFILLER_12_348 VPWR VGND sg13g2_fill_1
XFILLER_40_657 VPWR VGND sg13g2_fill_1
XFILLER_36_908 VPWR VGND sg13g2_decap_8
XFILLER_29_960 VPWR VGND sg13g2_decap_8
XFILLER_44_930 VPWR VGND sg13g2_decap_8
XFILLER_15_142 VPWR VGND sg13g2_fill_2
Xhold308 mac1.sum_lvl3_ff\[30\] VPWR VGND net348 sg13g2_dlygate4sd3_1
X_3410_ _2991_ net1018 net954 VPWR VGND sg13g2_nand2_1
Xhold319 _2196_ VPWR VGND net359 sg13g2_dlygate4sd3_1
X_4390_ _1205_ net823 net1027 VPWR VGND sg13g2_nand2_1
X_3341_ VGND VPWR _2866_ _2897_ _2929_ _2899_ sg13g2_a21oi_1
X_6060_ net1062 VGND VPWR _0171_ DP_4.matrix\[80\] clknet_leaf_24_clk sg13g2_dfrbpq_1
X_3272_ _2860_ _2836_ _2862_ VPWR VGND sg13g2_xor2_1
X_5011_ _1786_ VPWR _1798_ VGND _1794_ _1796_ sg13g2_o21ai_1
XFILLER_27_908 VPWR VGND sg13g2_decap_8
XFILLER_39_779 VPWR VGND sg13g2_decap_4
XFILLER_35_930 VPWR VGND sg13g2_decap_8
X_5913_ net892 net770 _2583_ VPWR VGND sg13g2_nor2_1
X_5844_ net778 VPWR _2537_ VGND net837 net785 sg13g2_o21ai_1
XFILLER_34_484 VPWR VGND sg13g2_fill_2
XFILLER_22_657 VPWR VGND sg13g2_fill_2
X_5775_ DP_3.Q_range.out_data\[3\] DP_3.I_range.out_data\[3\] _2469_ VPWR VGND sg13g2_xor2_1
X_4726_ _1486_ VPWR _1526_ VGND _1484_ _1487_ sg13g2_o21ai_1
X_4657_ _1457_ _1456_ _1447_ _1459_ VPWR VGND sg13g2_a21o_1
X_3608_ _0455_ net1012 net949 VPWR VGND sg13g2_nand2_1
X_6327_ net1046 VGND VPWR _0001_ mac1.sum_lvl3_ff\[10\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_4588_ VPWR _1392_ _1391_ VGND sg13g2_inv_1
X_3539_ _0385_ _0384_ _0354_ _0388_ VPWR VGND sg13g2_a21o_1
XFILLER_27_1006 VPWR VGND sg13g2_decap_8
X_6258_ net1077 VGND VPWR net208 mac2.sum_lvl2_ff\[43\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_6189_ net1066 VGND VPWR net181 mac1.sum_lvl1_ff\[36\] clknet_leaf_63_clk sg13g2_dfrbpq_1
X_5209_ _1989_ _1965_ _1991_ VPWR VGND sg13g2_xor2_1
XFILLER_29_256 VPWR VGND sg13g2_fill_2
XFILLER_26_952 VPWR VGND sg13g2_decap_8
XFILLER_41_900 VPWR VGND sg13g2_decap_8
XFILLER_41_977 VPWR VGND sg13g2_decap_8
XFILLER_21_690 VPWR VGND sg13g2_fill_2
XFILLER_5_812 VPWR VGND sg13g2_fill_2
XFILLER_5_889 VPWR VGND sg13g2_fill_1
XFILLER_44_760 VPWR VGND sg13g2_fill_1
XFILLER_17_985 VPWR VGND sg13g2_decap_8
XFILLER_32_922 VPWR VGND sg13g2_decap_8
X_3890_ _0724_ _0694_ _0722_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_421 VPWR VGND sg13g2_decap_4
XFILLER_32_999 VPWR VGND sg13g2_decap_8
X_5560_ VGND VPWR _2283_ _2285_ _2286_ _2284_ sg13g2_a21oi_1
X_4511_ _1321_ _1296_ _1322_ VPWR VGND sg13g2_xor2_1
X_5491_ net354 _2230_ _0041_ VPWR VGND sg13g2_xor2_1
Xhold105 mac1.products_ff\[143\] VPWR VGND net145 sg13g2_dlygate4sd3_1
Xhold116 mac1.sum_lvl2_ff\[48\] VPWR VGND net156 sg13g2_dlygate4sd3_1
X_4442_ VGND VPWR _1255_ _1256_ _1221_ _1181_ sg13g2_a21oi_2
Xhold138 mac1.sum_lvl1_ff\[42\] VPWR VGND net178 sg13g2_dlygate4sd3_1
Xhold127 mac1.sum_lvl1_ff\[83\] VPWR VGND net167 sg13g2_dlygate4sd3_1
Xhold149 mac2.sum_lvl1_ff\[9\] VPWR VGND net189 sg13g2_dlygate4sd3_1
X_4373_ _1188_ net885 net1022 VPWR VGND sg13g2_nand2_1
X_3324_ _2911_ _2885_ _2912_ VPWR VGND sg13g2_xor2_1
X_6112_ net1110 VGND VPWR _0210_ DP_2.matrix\[42\] clknet_leaf_45_clk sg13g2_dfrbpq_2
X_3255_ _2845_ _2838_ _2844_ VPWR VGND sg13g2_xnor2_1
X_6043_ net1113 VGND VPWR _0117_ mac1.products_ff\[78\] clknet_leaf_48_clk sg13g2_dfrbpq_1
X_3186_ _2767_ _2775_ _2777_ _2778_ VPWR VGND sg13g2_or3_1
XFILLER_2_1008 VPWR VGND sg13g2_decap_8
X_5827_ net818 net787 _2520_ VPWR VGND sg13g2_nor2_1
XFILLER_23_999 VPWR VGND sg13g2_decap_8
XFILLER_33_1010 VPWR VGND sg13g2_decap_8
XFILLER_10_649 VPWR VGND sg13g2_fill_2
X_5758_ net954 net936 net789 _2453_ VPWR VGND sg13g2_mux2_1
XFILLER_6_609 VPWR VGND sg13g2_fill_2
X_4709_ _1509_ net904 net1023 VPWR VGND sg13g2_nand2_1
X_5689_ mac2.total_sum\[14\] mac1.total_sum\[14\] _2388_ VPWR VGND sg13g2_xor2_1
XFILLER_2_826 VPWR VGND sg13g2_fill_2
XFILLER_27_74 VPWR VGND sg13g2_fill_2
XFILLER_33_719 VPWR VGND sg13g2_fill_2
XFILLER_25_292 VPWR VGND sg13g2_fill_1
XFILLER_14_977 VPWR VGND sg13g2_decap_8
XFILLER_5_664 VPWR VGND sg13g2_fill_1
XFILLER_5_686 VPWR VGND sg13g2_fill_1
XFILLER_49_841 VPWR VGND sg13g2_fill_2
X_3040_ _2636_ net978 net915 VPWR VGND sg13g2_nand2_1
XFILLER_36_513 VPWR VGND sg13g2_decap_8
XFILLER_36_546 VPWR VGND sg13g2_fill_2
XFILLER_36_568 VPWR VGND sg13g2_fill_2
X_4991_ VGND VPWR _1779_ _1778_ _1758_ sg13g2_or2_1
X_3942_ _0774_ _0766_ _0773_ VPWR VGND sg13g2_nand2_1
X_3873_ _0707_ net936 net995 VPWR VGND sg13g2_nand2_1
XFILLER_17_1027 VPWR VGND sg13g2_fill_2
XFILLER_20_936 VPWR VGND sg13g2_decap_8
X_5612_ _2328_ net468 _2326_ VPWR VGND sg13g2_nand2b_1
X_5543_ _2274_ mac2.sum_lvl2_ff\[33\] mac2.sum_lvl2_ff\[14\] VPWR VGND sg13g2_nand2_1
X_5474_ _0021_ net478 _2220_ VPWR VGND sg13g2_xnor2_1
X_4425_ net821 net819 net873 net870 _1239_ VPWR VGND sg13g2_and4_1
X_4356_ _1172_ _1136_ _1170_ _1171_ VPWR VGND sg13g2_and3_1
X_3307_ _2894_ _2871_ _2896_ VPWR VGND sg13g2_xor2_1
X_4287_ _1086_ _1076_ _1084_ _1104_ VPWR VGND sg13g2_a21o_1
X_6026_ net1098 VGND VPWR _0115_ mac1.products_ff\[9\] clknet_leaf_57_clk sg13g2_dfrbpq_1
X_3238_ _2829_ _2798_ _2827_ VPWR VGND sg13g2_xnor2_1
X_3169_ _2733_ VPWR _2761_ VGND _2724_ _2734_ sg13g2_o21ai_1
XFILLER_27_568 VPWR VGND sg13g2_decap_4
XFILLER_11_903 VPWR VGND sg13g2_fill_1
XFILLER_11_914 VPWR VGND sg13g2_fill_2
XFILLER_23_763 VPWR VGND sg13g2_fill_1
Xhold480 _0044_ VPWR VGND net520 sg13g2_dlygate4sd3_1
XFILLER_49_104 VPWR VGND sg13g2_fill_2
Xhold491 _2133_ VPWR VGND net531 sg13g2_dlygate4sd3_1
Xfanout960 net341 net960 VPWR VGND sg13g2_buf_8
Xfanout993 net544 net993 VPWR VGND sg13g2_buf_1
Xfanout982 net983 net982 VPWR VGND sg13g2_buf_1
Xfanout971 net327 net971 VPWR VGND sg13g2_buf_1
XFILLER_10_980 VPWR VGND sg13g2_decap_8
Xclkload14 clknet_leaf_44_clk clkload14/Y VPWR VGND sg13g2_inv_4
XFILLER_5_450 VPWR VGND sg13g2_fill_2
X_4210_ VGND VPWR _1027_ _1028_ _1030_ _1022_ sg13g2_a21oi_1
X_5190_ _1972_ _1931_ _1970_ VPWR VGND sg13g2_xnor2_1
X_4141_ _0942_ _0965_ _0967_ VPWR VGND sg13g2_and2_1
X_4072_ _0901_ _0856_ _0899_ VPWR VGND sg13g2_xnor2_1
XFILLER_23_1020 VPWR VGND sg13g2_decap_8
X_3023_ net923 net920 net978 net976 _2620_ VPWR VGND sg13g2_and4_1
XFILLER_37_844 VPWR VGND sg13g2_decap_8
X_4974_ _1759_ _1761_ _1762_ VPWR VGND sg13g2_nor2_1
X_3925_ _0756_ _0757_ _0726_ _0758_ VPWR VGND sg13g2_nand3_1
X_3856_ _0688_ _0689_ _0664_ _0691_ VPWR VGND sg13g2_nand3_1
Xclkload8 clknet_4_11_0_clk clkload8/X VPWR VGND sg13g2_buf_8
X_3787_ _0624_ net432 _0075_ VPWR VGND sg13g2_nor2_1
XFILLER_30_1002 VPWR VGND sg13g2_decap_8
X_5526_ mac2.sum_lvl2_ff\[30\] mac2.sum_lvl2_ff\[11\] _2260_ VPWR VGND sg13g2_nor2_1
X_5457_ _2206_ mac1.sum_lvl3_ff\[32\] mac1.sum_lvl3_ff\[12\] VPWR VGND sg13g2_nand2_1
X_4408_ VGND VPWR _1187_ _1193_ _1222_ _1195_ sg13g2_a21oi_1
X_5388_ _2143_ _2147_ _2153_ VPWR VGND sg13g2_nor2_1
XFILLER_8_1025 VPWR VGND sg13g2_decap_4
X_4339_ _1115_ VPWR _1155_ VGND _1113_ _1116_ sg13g2_o21ai_1
X_6009_ net799 _0265_ VPWR VGND sg13g2_buf_1
Xclkbuf_leaf_66_clk clknet_4_0_0_clk clknet_leaf_66_clk VPWR VGND sg13g2_buf_8
XFILLER_28_866 VPWR VGND sg13g2_decap_8
XFILLER_43_869 VPWR VGND sg13g2_decap_8
XFILLER_10_210 VPWR VGND sg13g2_fill_2
XFILLER_11_766 VPWR VGND sg13g2_fill_2
XFILLER_6_269 VPWR VGND sg13g2_fill_2
XFILLER_6_0 VPWR VGND sg13g2_fill_2
XFILLER_3_954 VPWR VGND sg13g2_decap_8
XFILLER_46_1020 VPWR VGND sg13g2_decap_8
Xfanout790 _2399_ net790 VPWR VGND sg13g2_buf_8
Xclkbuf_leaf_57_clk clknet_4_9_0_clk clknet_leaf_57_clk VPWR VGND sg13g2_buf_8
XFILLER_34_825 VPWR VGND sg13g2_decap_8
XFILLER_21_508 VPWR VGND sg13g2_fill_2
XFILLER_42_891 VPWR VGND sg13g2_decap_8
X_3710_ net1010 DP_1.matrix\[6\] net947 net945 _0554_ VPWR VGND sg13g2_and4_1
XFILLER_14_1019 VPWR VGND sg13g2_decap_8
X_4690_ _1488_ _1489_ _1483_ _1491_ VPWR VGND sg13g2_nand3_1
X_3641_ _0487_ _0446_ _0485_ VPWR VGND sg13g2_xnor2_1
X_3572_ _0417_ _0418_ _0412_ _0420_ VPWR VGND sg13g2_nand3_1
X_6360_ net1044 VGND VPWR net365 mac1.total_sum\[11\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_5311_ _2089_ net796 net1024 VPWR VGND sg13g2_nand2_1
X_6291_ net1061 VGND VPWR net139 mac2.sum_lvl1_ff\[78\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_5242_ _2022_ _2000_ _2023_ VPWR VGND sg13g2_nor2b_1
X_5173_ _1955_ _1938_ _1956_ VPWR VGND sg13g2_xor2_1
X_4124_ _0950_ _0924_ _0951_ VPWR VGND sg13g2_xor2_1
Xinput1 ui_in[0] net1 VPWR VGND sg13g2_buf_1
X_4055_ VGND VPWR _0884_ _0885_ _0850_ _0810_ sg13g2_a21oi_2
Xclkbuf_leaf_48_clk clknet_4_11_0_clk clknet_leaf_48_clk VPWR VGND sg13g2_buf_8
X_3006_ VPWR _2606_ net292 VGND sg13g2_inv_1
XFILLER_24_368 VPWR VGND sg13g2_fill_1
XFILLER_33_891 VPWR VGND sg13g2_decap_8
X_4957_ _1746_ net868 net803 VPWR VGND sg13g2_nand2_1
X_4888_ _1682_ _1681_ _1684_ VPWR VGND sg13g2_xor2_1
X_3908_ _0709_ VPWR _0741_ VGND _0707_ _0710_ sg13g2_o21ai_1
X_3839_ _0654_ VPWR _0674_ VGND _0652_ _0655_ sg13g2_o21ai_1
XFILLER_4_729 VPWR VGND sg13g2_fill_2
X_6489_ net1077 VGND VPWR _0045_ mac2.sum_lvl3_ff\[7\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_5509_ _2239_ _2242_ _2245_ _2247_ VPWR VGND sg13g2_or3_1
Xfanout1029 DP_3.matrix\[8\] net1029 VPWR VGND sg13g2_buf_1
Xfanout1018 net441 net1018 VPWR VGND sg13g2_buf_8
Xfanout1007 net1008 net1007 VPWR VGND sg13g2_buf_2
XFILLER_0_968 VPWR VGND sg13g2_decap_8
XFILLER_47_416 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_39_clk clknet_4_14_0_clk clknet_leaf_39_clk VPWR VGND sg13g2_buf_8
XFILLER_15_313 VPWR VGND sg13g2_fill_1
XFILLER_42_110 VPWR VGND sg13g2_fill_2
XFILLER_37_1019 VPWR VGND sg13g2_decap_8
XFILLER_24_891 VPWR VGND sg13g2_fill_1
XFILLER_7_534 VPWR VGND sg13g2_fill_2
XFILLER_47_983 VPWR VGND sg13g2_decap_8
XFILLER_46_471 VPWR VGND sg13g2_fill_1
X_5860_ _2419_ _2415_ _2551_ VPWR VGND sg13g2_xor2_1
X_4811_ _1609_ net838 net889 VPWR VGND sg13g2_nand2_1
X_5791_ net778 VPWR _2485_ VGND net894 net785 sg13g2_o21ai_1
X_4742_ _1518_ VPWR _1542_ VGND _1538_ _1540_ sg13g2_o21ai_1
XFILLER_30_883 VPWR VGND sg13g2_decap_8
X_4673_ _1474_ _1469_ _1472_ VPWR VGND sg13g2_xnor2_1
X_6412_ net1057 VGND VPWR _0155_ mac2.products_ff\[151\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_3624_ _0470_ _0453_ _0471_ VPWR VGND sg13g2_xor2_1
X_3555_ _0403_ _0394_ _0401_ VPWR VGND sg13g2_xnor2_1
X_6343_ net1054 VGND VPWR net69 mac2.sum_lvl3_ff\[30\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_6274_ net1041 VGND VPWR net204 mac1.sum_lvl1_ff\[77\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3486_ net961 net958 net1009 net1007 _0336_ VPWR VGND sg13g2_and4_1
X_5225_ _2006_ _1980_ _2004_ VPWR VGND sg13g2_xnor2_1
X_5156_ _1905_ VPWR _1939_ VGND _1896_ _1906_ sg13g2_o21ai_1
X_4107_ VGND VPWR _0889_ _0894_ _0935_ _0906_ sg13g2_a21oi_1
X_5087_ VGND VPWR _1869_ _1870_ _1872_ _1839_ sg13g2_a21oi_1
X_4038_ net934 net931 net990 net987 _0868_ VPWR VGND sg13g2_and4_1
XFILLER_38_961 VPWR VGND sg13g2_decap_8
XFILLER_25_633 VPWR VGND sg13g2_fill_2
XFILLER_37_482 VPWR VGND sg13g2_fill_2
XFILLER_12_305 VPWR VGND sg13g2_fill_2
XFILLER_12_327 VPWR VGND sg13g2_fill_1
X_5989_ net867 _0237_ VPWR VGND sg13g2_buf_1
XFILLER_21_894 VPWR VGND sg13g2_decap_8
XFILLER_43_1023 VPWR VGND sg13g2_decap_4
XFILLER_46_73 VPWR VGND sg13g2_decap_8
XFILLER_44_986 VPWR VGND sg13g2_decap_8
Xhold309 _2200_ VPWR VGND net349 sg13g2_dlygate4sd3_1
X_3340_ VGND VPWR _2865_ _2897_ _2928_ _2899_ sg13g2_a21oi_1
X_3271_ _2861_ _2836_ _2860_ VPWR VGND sg13g2_nand2_1
X_5010_ _1786_ _1794_ _1796_ _1797_ VPWR VGND sg13g2_or3_1
XFILLER_39_714 VPWR VGND sg13g2_fill_2
XFILLER_19_493 VPWR VGND sg13g2_fill_2
X_5912_ _2582_ net894 _2479_ _0225_ VPWR VGND sg13g2_mux2_1
X_5843_ net820 net787 _2536_ VPWR VGND sg13g2_nor2_1
XFILLER_22_603 VPWR VGND sg13g2_fill_2
XFILLER_35_986 VPWR VGND sg13g2_decap_8
X_5774_ DP_3.I_range.out_data\[3\] DP_3.Q_range.out_data\[3\] _2468_ VPWR VGND sg13g2_nor2b_1
X_4725_ _1525_ _1520_ _1524_ VPWR VGND sg13g2_xnor2_1
X_4656_ _1456_ _1457_ _1447_ _1458_ VPWR VGND sg13g2_nand3_1
X_3607_ _0420_ VPWR _0454_ VGND _0411_ _0421_ sg13g2_o21ai_1
X_4587_ _1388_ _1390_ _1391_ VPWR VGND sg13g2_nor2_1
X_3538_ VGND VPWR _0384_ _0385_ _0387_ _0354_ sg13g2_a21oi_1
X_6326_ net1110 VGND VPWR net437 mac1.sum_lvl3_ff\[9\] clknet_leaf_57_clk sg13g2_dfrbpq_2
X_3469_ VGND VPWR _0316_ _0317_ _0320_ _0292_ sg13g2_a21oi_1
X_6257_ net1077 VGND VPWR net229 mac2.sum_lvl2_ff\[42\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_6188_ net1088 VGND VPWR _0267_ DP_4.matrix\[79\] clknet_leaf_26_clk sg13g2_dfrbpq_1
X_5208_ _1990_ _1965_ _1989_ VPWR VGND sg13g2_nand2_1
XFILLER_18_909 VPWR VGND sg13g2_fill_2
X_5139_ _1875_ _1876_ _1920_ _1921_ _1923_ VPWR VGND sg13g2_and4_1
XFILLER_26_931 VPWR VGND sg13g2_decap_8
XFILLER_38_791 VPWR VGND sg13g2_fill_1
XFILLER_41_956 VPWR VGND sg13g2_decap_8
XFILLER_8_106 VPWR VGND sg13g2_fill_2
XFILLER_32_97 VPWR VGND sg13g2_fill_1
XFILLER_10_1022 VPWR VGND sg13g2_decap_8
XFILLER_35_216 VPWR VGND sg13g2_fill_1
XFILLER_17_964 VPWR VGND sg13g2_decap_8
XFILLER_32_901 VPWR VGND sg13g2_decap_8
XFILLER_44_794 VPWR VGND sg13g2_fill_1
XFILLER_32_978 VPWR VGND sg13g2_decap_8
XFILLER_31_488 VPWR VGND sg13g2_fill_1
X_4510_ _1321_ net816 net871 VPWR VGND sg13g2_nand2_1
X_5490_ _2232_ mac2.sum_lvl2_ff\[22\] net353 VPWR VGND sg13g2_xnor2_1
Xhold106 mac1.sum_lvl1_ff\[36\] VPWR VGND net146 sg13g2_dlygate4sd3_1
Xhold117 mac2.sum_lvl1_ff\[3\] VPWR VGND net157 sg13g2_dlygate4sd3_1
X_4441_ VGND VPWR _1178_ _1220_ _1255_ _1219_ sg13g2_a21oi_1
Xhold139 mac2.sum_lvl1_ff\[51\] VPWR VGND net179 sg13g2_dlygate4sd3_1
Xhold128 mac1.products_ff\[9\] VPWR VGND net168 sg13g2_dlygate4sd3_1
X_6111_ net1051 VGND VPWR _0097_ mac1.products_ff\[148\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_4372_ _1152_ VPWR _1187_ VGND _1149_ _1153_ sg13g2_o21ai_1
X_3323_ _2911_ net968 net908 VPWR VGND sg13g2_nand2_1
X_6042_ net1113 VGND VPWR _0126_ mac1.products_ff\[77\] clknet_leaf_49_clk sg13g2_dfrbpq_1
X_3254_ _2843_ _2839_ _2844_ VPWR VGND sg13g2_xor2_1
XFILLER_39_511 VPWR VGND sg13g2_fill_2
X_3185_ VGND VPWR _2773_ _2774_ _2777_ _2768_ sg13g2_a21oi_1
X_5826_ _2519_ net799 net776 VPWR VGND sg13g2_nand2_1
XFILLER_23_978 VPWR VGND sg13g2_decap_8
X_5757_ _2452_ _2451_ _2447_ VPWR VGND sg13g2_nand2b_1
X_4708_ _1479_ VPWR _1508_ VGND _1476_ _1480_ sg13g2_o21ai_1
X_5688_ mac1.total_sum\[14\] mac2.total_sum\[14\] _2387_ VPWR VGND sg13g2_nor2_1
X_4639_ _1424_ VPWR _1441_ VGND _1415_ _1425_ sg13g2_o21ai_1
X_6309_ net1049 VGND VPWR net90 mac1.sum_lvl3_ff\[28\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_40_1015 VPWR VGND sg13g2_decap_8
XFILLER_17_238 VPWR VGND sg13g2_fill_1
XFILLER_41_742 VPWR VGND sg13g2_decap_4
XFILLER_41_797 VPWR VGND sg13g2_fill_2
XFILLER_5_676 VPWR VGND sg13g2_fill_1
XFILLER_4_175 VPWR VGND sg13g2_fill_1
XFILLER_0_370 VPWR VGND sg13g2_fill_1
XFILLER_16_260 VPWR VGND sg13g2_fill_2
X_4990_ _1776_ _1775_ _1778_ VPWR VGND sg13g2_xor2_1
X_3941_ _0771_ _0767_ _0773_ VPWR VGND sg13g2_xor2_1
XFILLER_17_1006 VPWR VGND sg13g2_decap_8
X_3872_ _0677_ VPWR _0706_ VGND _0675_ _0678_ sg13g2_o21ai_1
X_5611_ VGND VPWR _2327_ net467 mac2.sum_lvl3_ff\[33\] sg13g2_or2_1
X_5542_ VGND VPWR _2269_ _2271_ _2273_ _2270_ sg13g2_a21oi_1
XFILLER_9_993 VPWR VGND sg13g2_decap_8
X_5473_ _2219_ VPWR _2220_ VGND mac1.sum_lvl3_ff\[33\] net367 sg13g2_o21ai_1
X_4424_ _1238_ net819 net870 VPWR VGND sg13g2_nand2_1
X_4355_ _1147_ VPWR _1171_ VGND _1167_ _1169_ sg13g2_o21ai_1
X_3306_ _2894_ _2871_ _2895_ VPWR VGND sg13g2_nor2b_1
X_4286_ _1103_ _1098_ _1101_ VPWR VGND sg13g2_xnor2_1
X_6025_ net1098 VGND VPWR _0114_ mac1.products_ff\[8\] clknet_leaf_53_clk sg13g2_dfrbpq_1
X_3237_ _2828_ _2798_ _2827_ VPWR VGND sg13g2_nand2_1
X_3168_ _2760_ _2713_ _2759_ VPWR VGND sg13g2_xnor2_1
XFILLER_27_525 VPWR VGND sg13g2_fill_2
X_3099_ net918 net969 net921 _2693_ VPWR VGND net967 sg13g2_nand4_1
XFILLER_13_22 VPWR VGND sg13g2_fill_1
X_5809_ _2503_ _2502_ net777 net775 net274 VPWR VGND sg13g2_a22oi_1
Xhold470 _2129_ VPWR VGND net510 sg13g2_dlygate4sd3_1
Xhold481 DP_3.matrix\[74\] VPWR VGND net521 sg13g2_dlygate4sd3_1
Xhold492 _0013_ VPWR VGND net532 sg13g2_dlygate4sd3_1
XFILLER_49_138 VPWR VGND sg13g2_decap_8
Xfanout961 net962 net961 VPWR VGND sg13g2_buf_2
Xfanout950 net951 net950 VPWR VGND sg13g2_buf_8
Xfanout972 net973 net972 VPWR VGND sg13g2_buf_8
Xfanout994 net996 net994 VPWR VGND sg13g2_buf_8
Xfanout983 net296 net983 VPWR VGND sg13g2_buf_8
XFILLER_46_812 VPWR VGND sg13g2_decap_8
XFILLER_33_517 VPWR VGND sg13g2_fill_2
XFILLER_13_285 VPWR VGND sg13g2_fill_1
XFILLER_9_267 VPWR VGND sg13g2_fill_2
Xclkload15 clknet_leaf_57_clk clkload15/X VPWR VGND sg13g2_buf_8
XFILLER_6_985 VPWR VGND sg13g2_decap_8
XFILLER_5_484 VPWR VGND sg13g2_fill_2
X_4140_ _0120_ _0965_ _0966_ VPWR VGND sg13g2_xnor2_1
X_4071_ VGND VPWR _0900_ _0899_ _0856_ sg13g2_or2_1
X_3022_ _2619_ net983 net916 VPWR VGND sg13g2_nand2_1
X_4973_ net868 net866 net802 net800 _1761_ VPWR VGND sg13g2_and4_1
X_3924_ _0732_ VPWR _0757_ VGND _0753_ _0755_ sg13g2_o21ai_1
X_3855_ _0688_ _0689_ _0690_ VPWR VGND sg13g2_and2_1
Xclkload9 clknet_4_13_0_clk clkload9/X VPWR VGND sg13g2_buf_8
X_3786_ _0625_ net940 net1003 net1002 net943 VPWR VGND sg13g2_a22oi_1
X_5525_ _0033_ _2257_ _2258_ VPWR VGND sg13g2_xnor2_1
X_5456_ _0018_ _2204_ _2205_ VPWR VGND sg13g2_xnor2_1
X_4407_ _1221_ _1182_ _0137_ VPWR VGND sg13g2_xor2_1
XFILLER_8_1004 VPWR VGND sg13g2_decap_8
X_5387_ _2141_ _2146_ _2152_ VPWR VGND sg13g2_nor2_1
X_4338_ _1154_ _1149_ _1153_ VPWR VGND sg13g2_xnor2_1
X_4269_ _1085_ _1086_ _1076_ _1087_ VPWR VGND sg13g2_nand3_1
X_6008_ net276 _0264_ VPWR VGND sg13g2_buf_1
XFILLER_28_845 VPWR VGND sg13g2_decap_8
XFILLER_39_171 VPWR VGND sg13g2_fill_2
XFILLER_11_712 VPWR VGND sg13g2_fill_1
XFILLER_24_76 VPWR VGND sg13g2_fill_2
XFILLER_40_97 VPWR VGND sg13g2_fill_2
XFILLER_3_933 VPWR VGND sg13g2_decap_8
Xfanout780 net781 net780 VPWR VGND sg13g2_buf_8
Xfanout791 _2399_ net791 VPWR VGND sg13g2_buf_1
XFILLER_18_333 VPWR VGND sg13g2_fill_2
XFILLER_18_344 VPWR VGND sg13g2_fill_2
XFILLER_45_163 VPWR VGND sg13g2_decap_4
XFILLER_14_550 VPWR VGND sg13g2_decap_8
XFILLER_42_870 VPWR VGND sg13g2_decap_8
X_3640_ VGND VPWR _0486_ _0484_ _0447_ sg13g2_or2_1
X_3571_ _0419_ _0412_ _0417_ _0418_ VPWR VGND sg13g2_and3_1
X_5310_ _2088_ net792 net1024 VPWR VGND sg13g2_nand2_1
X_6290_ net1062 VGND VPWR net191 mac2.sum_lvl1_ff\[77\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_5241_ _2022_ _2001_ _2021_ VPWR VGND sg13g2_xnor2_1
X_5172_ _1955_ _1939_ _1953_ VPWR VGND sg13g2_xnor2_1
X_4123_ _0950_ net928 net988 VPWR VGND sg13g2_nand2_1
X_4054_ VGND VPWR _0807_ _0849_ _0884_ _0848_ sg13g2_a21oi_1
Xinput2 ui_in[1] net2 VPWR VGND sg13g2_buf_1
X_3005_ VPWR _2605_ net1006 VGND sg13g2_inv_1
X_4956_ _1744_ _1737_ _0091_ VPWR VGND sg13g2_xor2_1
XFILLER_33_870 VPWR VGND sg13g2_decap_8
X_4887_ _1681_ _1682_ _1683_ VPWR VGND sg13g2_nor2_1
X_3907_ _0740_ _0734_ _0739_ VPWR VGND sg13g2_xnor2_1
X_3838_ _0671_ _0668_ _0673_ VPWR VGND sg13g2_xor2_1
X_5508_ _2245_ VPWR _2246_ VGND _2239_ _2242_ sg13g2_o21ai_1
X_3769_ _0610_ _0600_ _0611_ VPWR VGND sg13g2_nor2b_1
X_6488_ net1077 VGND VPWR net520 mac2.sum_lvl3_ff\[6\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_5439_ VGND VPWR net420 _2188_ _2192_ _2191_ sg13g2_a21oi_1
XFILLER_0_947 VPWR VGND sg13g2_decap_8
Xfanout1019 net335 net1019 VPWR VGND sg13g2_buf_8
Xfanout1008 net446 net1008 VPWR VGND sg13g2_buf_8
XFILLER_47_406 VPWR VGND sg13g2_fill_1
XFILLER_28_653 VPWR VGND sg13g2_fill_2
XFILLER_15_303 VPWR VGND sg13g2_fill_2
XFILLER_28_686 VPWR VGND sg13g2_fill_1
XFILLER_7_513 VPWR VGND sg13g2_fill_2
XFILLER_3_763 VPWR VGND sg13g2_fill_1
XFILLER_19_642 VPWR VGND sg13g2_decap_8
XFILLER_20_1013 VPWR VGND sg13g2_decap_8
XFILLER_47_962 VPWR VGND sg13g2_decap_8
XFILLER_19_653 VPWR VGND sg13g2_fill_1
XFILLER_34_634 VPWR VGND sg13g2_fill_2
X_4810_ _1608_ net893 net836 VPWR VGND sg13g2_nand2_1
X_5790_ net876 _2472_ _2484_ VPWR VGND sg13g2_nor2_1
X_4741_ _1518_ _1538_ _1540_ _1541_ VPWR VGND sg13g2_or3_1
XFILLER_30_862 VPWR VGND sg13g2_decap_8
X_4672_ _1473_ _1469_ _1472_ VPWR VGND sg13g2_nand2_1
X_6411_ net1057 VGND VPWR _0154_ mac2.products_ff\[150\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_3623_ _0470_ _0454_ _0468_ VPWR VGND sg13g2_xnor2_1
X_3554_ _0402_ _0394_ _0401_ VPWR VGND sg13g2_nand2_1
X_6342_ net1060 VGND VPWR net160 mac2.sum_lvl3_ff\[29\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_3485_ _0335_ net954 net1012 VPWR VGND sg13g2_nand2_1
X_6273_ net1064 VGND VPWR net57 mac1.sum_lvl1_ff\[76\] clknet_leaf_65_clk sg13g2_dfrbpq_1
X_5224_ VGND VPWR _2005_ _2004_ _1980_ sg13g2_or2_1
X_5155_ _1938_ _1928_ _1936_ VPWR VGND sg13g2_xnor2_1
X_4106_ _0932_ _0920_ _0934_ VPWR VGND sg13g2_xor2_1
X_5086_ _1869_ _1870_ _1839_ _1871_ VPWR VGND sg13g2_nand3_1
XFILLER_38_940 VPWR VGND sg13g2_decap_8
X_4037_ _0867_ net931 net988 VPWR VGND sg13g2_nand2_1
XFILLER_36_1020 VPWR VGND sg13g2_decap_8
X_5988_ net868 _0236_ VPWR VGND sg13g2_buf_1
X_4939_ _1732_ net889 DP_4.matrix\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_21_884 VPWR VGND sg13g2_fill_1
XFILLER_43_1002 VPWR VGND sg13g2_decap_8
XFILLER_29_995 VPWR VGND sg13g2_decap_8
XFILLER_44_965 VPWR VGND sg13g2_decap_8
XFILLER_15_133 VPWR VGND sg13g2_fill_1
XFILLER_31_637 VPWR VGND sg13g2_fill_1
XFILLER_12_873 VPWR VGND sg13g2_fill_1
XFILLER_12_895 VPWR VGND sg13g2_fill_2
XFILLER_11_394 VPWR VGND sg13g2_fill_2
X_3270_ _2859_ _2847_ _2860_ VPWR VGND sg13g2_xor2_1
X_5911_ _2582_ _2486_ _2504_ VPWR VGND sg13g2_xnor2_1
XFILLER_35_965 VPWR VGND sg13g2_decap_8
X_5842_ _2535_ net276 net776 VPWR VGND sg13g2_nand2_1
XFILLER_34_486 VPWR VGND sg13g2_fill_1
X_5773_ VGND VPWR _2437_ _2466_ _0163_ _2467_ sg13g2_a21oi_1
X_4724_ _1524_ _1477_ _1522_ VPWR VGND sg13g2_xnor2_1
X_4655_ _1454_ _1453_ _1448_ _1457_ VPWR VGND sg13g2_a21o_1
X_3606_ _0453_ _0443_ _0451_ VPWR VGND sg13g2_xnor2_1
X_4586_ net903 net902 net839 net837 _1390_ VPWR VGND sg13g2_and4_1
X_6325_ net1109 VGND VPWR net378 mac1.sum_lvl3_ff\[8\] clknet_leaf_52_clk sg13g2_dfrbpq_2
X_3537_ _0384_ _0385_ _0354_ _0386_ VPWR VGND sg13g2_nand3_1
X_3468_ _0316_ _0317_ _0292_ _0319_ VPWR VGND sg13g2_nand3_1
X_6256_ net1078 VGND VPWR net124 mac2.sum_lvl2_ff\[41\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_6187_ net1082 VGND VPWR _0266_ DP_4.matrix\[78\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_3399_ _2980_ net442 _0070_ VPWR VGND sg13g2_nor2_1
X_5207_ _1988_ _1976_ _1989_ VPWR VGND sg13g2_xor2_1
X_5138_ _1922_ _1920_ _1921_ VPWR VGND sg13g2_nand2_1
XFILLER_26_910 VPWR VGND sg13g2_decap_8
X_5069_ _1822_ VPWR _1854_ VGND _1820_ _1823_ sg13g2_o21ai_1
XFILLER_26_987 VPWR VGND sg13g2_decap_8
XFILLER_41_935 VPWR VGND sg13g2_decap_8
XFILLER_10_1001 VPWR VGND sg13g2_decap_8
XFILLER_17_943 VPWR VGND sg13g2_decap_8
XFILLER_44_784 VPWR VGND sg13g2_fill_2
XFILLER_32_957 VPWR VGND sg13g2_decap_8
XFILLER_31_456 VPWR VGND sg13g2_fill_1
Xhold107 mac1.products_ff\[4\] VPWR VGND net147 sg13g2_dlygate4sd3_1
X_4440_ _1254_ _1253_ _1252_ VPWR VGND sg13g2_nand2b_1
Xhold118 mac1.sum_lvl1_ff\[77\] VPWR VGND net158 sg13g2_dlygate4sd3_1
Xhold129 mac1.sum_lvl1_ff\[15\] VPWR VGND net169 sg13g2_dlygate4sd3_1
X_6110_ net1110 VGND VPWR _0209_ DP_2.matrix\[41\] clknet_leaf_57_clk sg13g2_dfrbpq_1
X_4371_ _1140_ _1143_ _1186_ VPWR VGND sg13g2_nor2_1
X_3322_ _2910_ net968 net906 VPWR VGND sg13g2_nand2_1
X_6041_ net1117 VGND VPWR _0125_ mac1.products_ff\[76\] clknet_leaf_50_clk sg13g2_dfrbpq_1
X_3253_ _2843_ _2802_ _2841_ VPWR VGND sg13g2_xnor2_1
X_3184_ _2773_ _2774_ _2768_ _2776_ VPWR VGND sg13g2_nand3_1
XFILLER_14_0 VPWR VGND sg13g2_fill_1
X_5825_ _2517_ VPWR _2518_ VGND net767 _2516_ sg13g2_o21ai_1
XFILLER_23_957 VPWR VGND sg13g2_decap_8
XFILLER_10_618 VPWR VGND sg13g2_fill_2
X_5756_ _2451_ _2449_ _2450_ _2448_ net782 VPWR VGND sg13g2_a22oi_1
X_5687_ _2386_ mac1.total_sum\[14\] mac2.total_sum\[14\] VPWR VGND sg13g2_nand2_1
X_4707_ _1496_ VPWR _1507_ VGND _1474_ _1497_ sg13g2_o21ai_1
X_4638_ _1438_ _1437_ _1440_ VPWR VGND sg13g2_xor2_1
X_4569_ _1373_ _1366_ _0086_ VPWR VGND sg13g2_xor2_1
X_6308_ net1050 VGND VPWR net86 mac1.sum_lvl3_ff\[27\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_6239_ net1065 VGND VPWR net256 mac1.sum_lvl2_ff\[40\] clknet_leaf_64_clk sg13g2_dfrbpq_1
XFILLER_14_913 VPWR VGND sg13g2_fill_2
XFILLER_26_762 VPWR VGND sg13g2_fill_1
XFILLER_22_990 VPWR VGND sg13g2_decap_8
XFILLER_49_887 VPWR VGND sg13g2_decap_8
XFILLER_36_559 VPWR VGND sg13g2_fill_1
X_3940_ _0767_ _0771_ _0772_ VPWR VGND sg13g2_nor2_1
X_3871_ _0705_ _0700_ _0703_ VPWR VGND sg13g2_xnor2_1
X_5610_ mac2.sum_lvl3_ff\[33\] net467 _2326_ VPWR VGND sg13g2_and2_1
X_5541_ _0036_ _2269_ _2272_ VPWR VGND sg13g2_xnor2_1
X_5472_ _2211_ _2214_ _2206_ _2219_ VPWR VGND sg13g2_nand3_1
X_4423_ _1237_ net877 net818 VPWR VGND sg13g2_nand2_1
X_4354_ _1147_ _1167_ _1169_ _1170_ VPWR VGND sg13g2_or3_1
X_3305_ _2894_ _2872_ _2893_ VPWR VGND sg13g2_xnor2_1
X_6024_ net1097 VGND VPWR _0113_ mac1.products_ff\[7\] clknet_leaf_53_clk sg13g2_dfrbpq_1
X_4285_ _1102_ _1098_ _1101_ VPWR VGND sg13g2_nand2_1
X_3236_ _2826_ _2809_ _2827_ VPWR VGND sg13g2_xor2_1
X_3167_ _2759_ _2750_ _2757_ VPWR VGND sg13g2_xnor2_1
X_3098_ net921 net918 net969 net967 _2692_ VPWR VGND sg13g2_and4_1
X_5808_ net878 net895 net787 _2502_ VPWR VGND sg13g2_mux2_1
XFILLER_10_459 VPWR VGND sg13g2_fill_1
X_5739_ net783 VPWR _2434_ VGND net1032 net789 sg13g2_o21ai_1
Xhold460 DP_4.matrix\[42\] VPWR VGND net500 sg13g2_dlygate4sd3_1
Xhold471 _0012_ VPWR VGND net511 sg13g2_dlygate4sd3_1
Xhold493 mac1.sum_lvl3_ff\[26\] VPWR VGND net533 sg13g2_dlygate4sd3_1
Xhold482 DP_1.matrix\[8\] VPWR VGND net522 sg13g2_dlygate4sd3_1
Xfanout940 net431 net940 VPWR VGND sg13g2_buf_8
Xfanout951 net418 net951 VPWR VGND sg13g2_buf_8
Xfanout973 net974 net973 VPWR VGND sg13g2_buf_2
Xfanout995 net996 net995 VPWR VGND sg13g2_buf_1
Xfanout962 net963 net962 VPWR VGND sg13g2_buf_1
Xfanout984 net985 net984 VPWR VGND sg13g2_buf_8
XFILLER_18_504 VPWR VGND sg13g2_decap_8
XFILLER_38_86 VPWR VGND sg13g2_fill_2
XFILLER_13_264 VPWR VGND sg13g2_fill_2
XFILLER_13_275 VPWR VGND sg13g2_fill_1
XFILLER_41_562 VPWR VGND sg13g2_fill_2
XFILLER_9_246 VPWR VGND sg13g2_fill_1
Xclkload16 clknet_leaf_50_clk clkload16/Y VPWR VGND sg13g2_inv_4
XFILLER_6_964 VPWR VGND sg13g2_decap_8
XFILLER_5_463 VPWR VGND sg13g2_fill_2
XFILLER_5_452 VPWR VGND sg13g2_fill_1
X_4070_ _0899_ net991 net927 VPWR VGND sg13g2_nand2_2
X_3021_ VGND VPWR _2618_ _2613_ _2611_ sg13g2_or2_1
XFILLER_37_879 VPWR VGND sg13g2_decap_8
X_4972_ _1760_ net866 net800 VPWR VGND sg13g2_nand2_1
X_3923_ _0732_ _0753_ _0755_ _0756_ VPWR VGND sg13g2_or3_1
X_3854_ _0687_ _0686_ _0648_ _0689_ VPWR VGND sg13g2_a21o_1
X_3785_ _0624_ net1002 net940 _0074_ VPWR VGND sg13g2_and3_2
X_5524_ _2259_ _2256_ _2258_ VPWR VGND sg13g2_nand2_1
X_5455_ _2205_ _2199_ _2201_ VPWR VGND sg13g2_nand2_1
X_4406_ _1219_ _1220_ _1221_ VPWR VGND sg13g2_nor2b_2
X_5386_ net481 mac1.sum_lvl2_ff\[31\] _2151_ VPWR VGND sg13g2_xor2_1
X_4337_ _1153_ _1106_ _1151_ VPWR VGND sg13g2_xnor2_1
X_4268_ _1083_ _1082_ _1077_ _1086_ VPWR VGND sg13g2_a21o_1
X_3219_ _2776_ VPWR _2810_ VGND _2767_ _2777_ sg13g2_o21ai_1
X_6007_ net803 _0263_ VPWR VGND sg13g2_buf_1
X_4199_ net887 net884 net822 net820 _1019_ VPWR VGND sg13g2_and4_1
XFILLER_27_356 VPWR VGND sg13g2_fill_2
XFILLER_10_212 VPWR VGND sg13g2_fill_1
XFILLER_3_989 VPWR VGND sg13g2_decap_8
XFILLER_49_41 VPWR VGND sg13g2_fill_1
Xhold290 _0053_ VPWR VGND net330 sg13g2_dlygate4sd3_1
Xfanout792 net794 net792 VPWR VGND sg13g2_buf_8
Xfanout770 _2478_ net770 VPWR VGND sg13g2_buf_8
Xfanout781 _2405_ net781 VPWR VGND sg13g2_buf_8
XFILLER_18_301 VPWR VGND sg13g2_decap_4
XFILLER_33_326 VPWR VGND sg13g2_fill_1
XFILLER_14_573 VPWR VGND sg13g2_fill_2
X_3570_ _0413_ VPWR _0418_ VGND _0414_ _0416_ sg13g2_o21ai_1
X_5240_ _2021_ _2010_ _2020_ VPWR VGND sg13g2_xnor2_1
X_5171_ _1954_ _1939_ _1953_ VPWR VGND sg13g2_nand2_1
X_4122_ _0949_ net988 net926 VPWR VGND sg13g2_nand2_1
X_4053_ _0883_ _0882_ _0881_ VPWR VGND sg13g2_nand2b_1
X_3004_ VPWR DP_1.Q_range.data_plus_4\[6\] net8 VGND sg13g2_inv_1
Xinput3 ui_in[2] net3 VPWR VGND sg13g2_buf_1
X_4955_ _1745_ _1737_ _1744_ VPWR VGND sg13g2_nand2_1
XFILLER_40_819 VPWR VGND sg13g2_decap_8
X_3906_ _0739_ _0701_ _0736_ VPWR VGND sg13g2_xnor2_1
X_4886_ VGND VPWR _1630_ _1649_ _1682_ _1651_ sg13g2_a21oi_1
X_3837_ _0672_ _0671_ _0668_ VPWR VGND sg13g2_nand2b_1
X_3768_ _0610_ _0586_ _0609_ VPWR VGND sg13g2_xnor2_1
X_5507_ mac2.sum_lvl2_ff\[7\] mac2.sum_lvl2_ff\[26\] _2245_ VPWR VGND sg13g2_xor2_1
X_3699_ _0509_ _0514_ _0544_ VPWR VGND sg13g2_nor2_1
X_6487_ net1078 VGND VPWR net389 mac2.sum_lvl3_ff\[5\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_5438_ _2191_ mac1.sum_lvl3_ff\[28\] mac1.sum_lvl3_ff\[8\] VPWR VGND sg13g2_xnor2_1
X_5369_ net375 mac1.sum_lvl2_ff\[27\] net377 _2137_ VPWR VGND sg13g2_a21o_1
XFILLER_0_926 VPWR VGND sg13g2_decap_8
Xfanout1009 net1010 net1009 VPWR VGND sg13g2_buf_2
XFILLER_48_919 VPWR VGND sg13g2_decap_8
XFILLER_19_66 VPWR VGND sg13g2_fill_2
XFILLER_42_112 VPWR VGND sg13g2_fill_1
XFILLER_27_197 VPWR VGND sg13g2_fill_2
XFILLER_11_576 VPWR VGND sg13g2_fill_1
XFILLER_7_536 VPWR VGND sg13g2_fill_1
XFILLER_11_598 VPWR VGND sg13g2_fill_2
XFILLER_3_775 VPWR VGND sg13g2_fill_2
XFILLER_39_919 VPWR VGND sg13g2_decap_8
XFILLER_47_941 VPWR VGND sg13g2_decap_8
XFILLER_18_153 VPWR VGND sg13g2_fill_2
XFILLER_19_687 VPWR VGND sg13g2_fill_2
XFILLER_33_134 VPWR VGND sg13g2_decap_4
XFILLER_15_860 VPWR VGND sg13g2_fill_1
XFILLER_33_167 VPWR VGND sg13g2_fill_2
X_4740_ VGND VPWR _1536_ _1537_ _1540_ _1519_ sg13g2_a21oi_1
X_4671_ _1470_ _1471_ _1472_ VPWR VGND sg13g2_nor2b_1
X_3622_ _0469_ _0454_ _0468_ VPWR VGND sg13g2_nand2_1
X_6410_ net1058 VGND VPWR _0153_ mac2.products_ff\[149\] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_6341_ net1051 VGND VPWR net247 mac2.sum_lvl3_ff\[28\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_3553_ _0399_ _0395_ _0401_ VPWR VGND sg13g2_xor2_1
X_3484_ _0305_ VPWR _0334_ VGND _0303_ _0306_ sg13g2_o21ai_1
X_6272_ net1049 VGND VPWR net262 mac1.sum_lvl1_ff\[75\] clknet_leaf_67_clk sg13g2_dfrbpq_1
X_5223_ _2004_ net803 net1024 VPWR VGND sg13g2_nand2_1
X_5154_ _1928_ _1936_ _1937_ VPWR VGND sg13g2_nor2_1
X_4105_ VGND VPWR _0933_ _0932_ _0920_ sg13g2_or2_1
X_5085_ _1845_ VPWR _1870_ VGND _1866_ _1868_ sg13g2_o21ai_1
X_4036_ _0866_ net991 net929 VPWR VGND sg13g2_nand2_1
XFILLER_25_602 VPWR VGND sg13g2_fill_2
XFILLER_37_484 VPWR VGND sg13g2_fill_1
XFILLER_38_996 VPWR VGND sg13g2_decap_8
XFILLER_25_635 VPWR VGND sg13g2_fill_1
X_5987_ net872 _0235_ VPWR VGND sg13g2_buf_1
XFILLER_25_679 VPWR VGND sg13g2_decap_8
X_4938_ _1720_ VPWR _1731_ VGND _1691_ _1718_ sg13g2_o21ai_1
XFILLER_33_690 VPWR VGND sg13g2_decap_4
X_4869_ _1665_ net896 net1023 VPWR VGND sg13g2_nand2_1
XFILLER_29_974 VPWR VGND sg13g2_decap_8
XFILLER_44_944 VPWR VGND sg13g2_decap_8
XFILLER_12_830 VPWR VGND sg13g2_fill_1
XFILLER_30_115 VPWR VGND sg13g2_decap_4
XFILLER_8_856 VPWR VGND sg13g2_fill_2
X_5910_ VGND VPWR net769 _2581_ _0224_ _2580_ sg13g2_a21oi_1
XFILLER_19_495 VPWR VGND sg13g2_fill_1
XFILLER_35_944 VPWR VGND sg13g2_decap_8
X_5841_ _2534_ _2533_ _2524_ VPWR VGND sg13g2_nand2b_1
X_5772_ VGND VPWR net773 _2466_ _2467_ _2438_ sg13g2_a21oi_1
X_4723_ VGND VPWR _1523_ _1521_ _1478_ sg13g2_or2_1
X_4654_ _1453_ _1454_ _1448_ _1456_ VPWR VGND sg13g2_nand3_1
X_3605_ _0443_ _0451_ _0452_ VPWR VGND sg13g2_nor2_1
X_4585_ _1389_ net902 net837 VPWR VGND sg13g2_nand2_1
X_3536_ _0360_ VPWR _0385_ VGND _0381_ _0383_ sg13g2_o21ai_1
X_6324_ net1109 VGND VPWR net532 mac1.sum_lvl3_ff\[7\] clknet_leaf_52_clk sg13g2_dfrbpq_2
X_6255_ net1078 VGND VPWR net150 mac2.sum_lvl2_ff\[40\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_5206_ _1986_ _1977_ _1988_ VPWR VGND sg13g2_xor2_1
X_3467_ _0316_ _0317_ _0318_ VPWR VGND sg13g2_and2_1
X_6186_ net1088 VGND VPWR _0265_ DP_4.matrix\[77\] clknet_leaf_26_clk sg13g2_dfrbpq_1
X_3398_ _2981_ net956 net1019 net1018 net960 VPWR VGND sg13g2_a22oi_1
X_5137_ _1918_ _1917_ _1919_ _1921_ VPWR VGND sg13g2_a21o_1
X_5068_ _1853_ _1847_ _1852_ VPWR VGND sg13g2_xnor2_1
X_4019_ _0848_ _0849_ _0850_ VPWR VGND sg13g2_nor2b_1
XFILLER_26_966 VPWR VGND sg13g2_decap_8
XFILLER_16_78 VPWR VGND sg13g2_fill_2
XFILLER_41_914 VPWR VGND sg13g2_decap_8
XFILLER_40_424 VPWR VGND sg13g2_fill_1
XFILLER_9_609 VPWR VGND sg13g2_decap_8
XFILLER_8_108 VPWR VGND sg13g2_fill_1
XFILLER_5_859 VPWR VGND sg13g2_fill_2
XFILLER_16_454 VPWR VGND sg13g2_fill_1
XFILLER_17_999 VPWR VGND sg13g2_decap_8
XFILLER_32_936 VPWR VGND sg13g2_decap_8
XFILLER_12_671 VPWR VGND sg13g2_decap_4
XFILLER_40_980 VPWR VGND sg13g2_decap_8
Xhold108 mac1.sum_lvl1_ff\[1\] VPWR VGND net148 sg13g2_dlygate4sd3_1
Xhold119 mac1.sum_lvl1_ff\[44\] VPWR VGND net159 sg13g2_dlygate4sd3_1
X_4370_ _1168_ VPWR _1185_ VGND _1147_ _1169_ sg13g2_o21ai_1
X_3321_ _2909_ net974 net1030 VPWR VGND sg13g2_nand2_1
X_6040_ net1108 VGND VPWR _0124_ mac1.products_ff\[75\] clknet_leaf_51_clk sg13g2_dfrbpq_1
X_3252_ VGND VPWR _2842_ _2840_ _2803_ sg13g2_or2_1
X_3183_ _2775_ _2768_ _2773_ _2774_ VPWR VGND sg13g2_and3_1
XFILLER_39_513 VPWR VGND sg13g2_fill_1
X_5824_ _2517_ net1023 net767 VPWR VGND sg13g2_nand2_1
XFILLER_23_936 VPWR VGND sg13g2_decap_8
X_5755_ net782 VPWR _2450_ VGND net940 net790 sg13g2_o21ai_1
XFILLER_33_1024 VPWR VGND sg13g2_decap_4
X_5686_ VGND VPWR _2381_ _2383_ _2385_ _2382_ sg13g2_a21oi_1
X_4706_ _1505_ _1504_ _0146_ VPWR VGND sg13g2_xor2_1
X_4637_ _1439_ _1437_ _1438_ VPWR VGND sg13g2_nand2b_1
X_4568_ _1374_ _1366_ _1373_ VPWR VGND sg13g2_nand2_1
X_6307_ net1067 VGND VPWR net217 mac1.sum_lvl3_ff\[26\] clknet_leaf_65_clk sg13g2_dfrbpq_2
X_3519_ _0368_ _0362_ _0367_ VPWR VGND sg13g2_xnor2_1
X_4499_ VGND VPWR _1259_ _1279_ _1311_ _1281_ sg13g2_a21oi_1
X_6238_ net1049 VGND VPWR net259 mac1.sum_lvl2_ff\[39\] clknet_leaf_67_clk sg13g2_dfrbpq_1
X_6169_ net1089 VGND VPWR net415 DP_4.matrix\[4\] clknet_leaf_26_clk sg13g2_dfrbpq_1
XFILLER_45_505 VPWR VGND sg13g2_fill_2
XFILLER_45_538 VPWR VGND sg13g2_decap_8
XFILLER_14_936 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_20_clk clknet_4_4_0_clk clknet_leaf_20_clk VPWR VGND sg13g2_buf_8
XFILLER_4_133 VPWR VGND sg13g2_fill_2
XFILLER_49_1020 VPWR VGND sg13g2_decap_8
XFILLER_1_1022 VPWR VGND sg13g2_decap_8
X_3870_ _0704_ _0703_ _0700_ VPWR VGND sg13g2_nand2b_1
X_5540_ _2272_ _2271_ _2270_ VPWR VGND sg13g2_nand2b_1
XFILLER_13_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_11_clk clknet_4_12_0_clk clknet_leaf_11_clk VPWR VGND sg13g2_buf_8
X_5471_ net477 mac1.sum_lvl3_ff\[34\] _2218_ VPWR VGND sg13g2_xor2_1
X_4422_ VGND VPWR net828 net870 _1236_ _1205_ sg13g2_a21oi_1
X_4353_ VGND VPWR _1165_ _1166_ _1169_ _1148_ sg13g2_a21oi_1
X_3304_ _2893_ _2881_ _2892_ VPWR VGND sg13g2_xnor2_1
X_4284_ _1099_ _1100_ _1101_ VPWR VGND sg13g2_nor2b_1
X_6023_ net1097 VGND VPWR _0112_ mac1.products_ff\[6\] clknet_leaf_53_clk sg13g2_dfrbpq_1
X_3235_ _2826_ _2810_ _2824_ VPWR VGND sg13g2_xnor2_1
X_3166_ _2758_ _2750_ _2757_ VPWR VGND sg13g2_nand2_1
X_3097_ _2691_ net915 net972 VPWR VGND sg13g2_nand2_1
XFILLER_10_416 VPWR VGND sg13g2_fill_2
X_3999_ _0779_ _0828_ _0830_ VPWR VGND sg13g2_and2_1
X_5807_ _2501_ _2500_ _2488_ VPWR VGND sg13g2_nand2b_1
X_5738_ VGND VPWR _2404_ _2432_ _0160_ _2433_ sg13g2_a21oi_1
X_5669_ net19 _2369_ _2370_ VPWR VGND sg13g2_xnor2_1
Xhold461 mac1.sum_lvl3_ff\[6\] VPWR VGND net501 sg13g2_dlygate4sd3_1
Xhold472 mac1.sum_lvl2_ff\[4\] VPWR VGND net512 sg13g2_dlygate4sd3_1
Xhold450 mac2.sum_lvl2_ff\[8\] VPWR VGND net490 sg13g2_dlygate4sd3_1
Xhold483 DP_2.matrix\[1\] VPWR VGND net523 sg13g2_dlygate4sd3_1
Xhold494 DP_2.matrix\[40\] VPWR VGND net534 sg13g2_dlygate4sd3_1
Xfanout941 net942 net941 VPWR VGND sg13g2_buf_2
Xfanout952 net399 net952 VPWR VGND sg13g2_buf_8
Xfanout930 net494 net930 VPWR VGND sg13g2_buf_8
Xfanout963 DP_2.matrix\[0\] net963 VPWR VGND sg13g2_buf_1
Xfanout985 net273 net985 VPWR VGND sg13g2_buf_2
Xfanout974 net318 net974 VPWR VGND sg13g2_buf_1
Xfanout996 net487 net996 VPWR VGND sg13g2_buf_8
XFILLER_45_335 VPWR VGND sg13g2_fill_1
XFILLER_33_519 VPWR VGND sg13g2_fill_1
XFILLER_9_269 VPWR VGND sg13g2_fill_1
Xclkload17 VPWR clkload17/Y clknet_leaf_48_clk VGND sg13g2_inv_1
XFILLER_10_994 VPWR VGND sg13g2_decap_8
XFILLER_5_486 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_0_clk clknet_4_0_0_clk clknet_leaf_0_clk VPWR VGND sg13g2_buf_8
X_3020_ _2617_ net984 net913 VPWR VGND sg13g2_nand2_1
XFILLER_37_858 VPWR VGND sg13g2_decap_8
X_4971_ _1759_ net800 net869 net802 net867 VPWR VGND sg13g2_a22oi_1
X_3922_ VGND VPWR _0751_ _0752_ _0755_ _0733_ sg13g2_a21oi_1
X_3853_ _0686_ _0687_ _0648_ _0688_ VPWR VGND sg13g2_nand3_1
XFILLER_9_770 VPWR VGND sg13g2_fill_1
X_3784_ net1003 net943 _0074_ VPWR VGND sg13g2_and2_1
XFILLER_30_1016 VPWR VGND sg13g2_decap_8
X_5523_ _2253_ _2251_ _2252_ _2258_ VPWR VGND sg13g2_a21o_2
XFILLER_30_1027 VPWR VGND sg13g2_fill_2
X_5454_ _2204_ _2203_ _2202_ VPWR VGND sg13g2_nand2b_1
X_5385_ mac1.sum_lvl2_ff\[31\] mac1.sum_lvl2_ff\[12\] _2150_ VPWR VGND sg13g2_nor2_1
X_4405_ _1220_ _1183_ _1218_ VPWR VGND sg13g2_nand2_1
X_4336_ VGND VPWR _1152_ _1150_ _1107_ sg13g2_or2_1
X_4267_ _1082_ _1083_ _1077_ _1085_ VPWR VGND sg13g2_nand3_1
X_3218_ _2809_ _2799_ _2807_ VPWR VGND sg13g2_xnor2_1
X_4198_ _1018_ net884 net819 VPWR VGND sg13g2_nand2_1
X_6006_ net805 _0262_ VPWR VGND sg13g2_buf_1
X_3149_ _2740_ _2741_ _2710_ _2742_ VPWR VGND sg13g2_nand3_1
XFILLER_39_173 VPWR VGND sg13g2_fill_1
XFILLER_15_519 VPWR VGND sg13g2_decap_8
XFILLER_36_880 VPWR VGND sg13g2_decap_8
XFILLER_42_349 VPWR VGND sg13g2_fill_2
XFILLER_23_574 VPWR VGND sg13g2_fill_1
XFILLER_3_913 VPWR VGND sg13g2_decap_4
XFILLER_3_902 VPWR VGND sg13g2_fill_2
XFILLER_40_99 VPWR VGND sg13g2_fill_1
XFILLER_3_968 VPWR VGND sg13g2_decap_8
XFILLER_2_456 VPWR VGND sg13g2_fill_1
Xhold280 mac1.sum_lvl3_ff\[5\] VPWR VGND net320 sg13g2_dlygate4sd3_1
Xhold291 DP_3.matrix\[38\] VPWR VGND net331 sg13g2_dlygate4sd3_1
XFILLER_49_86 VPWR VGND sg13g2_decap_8
Xfanout793 net794 net793 VPWR VGND sg13g2_buf_1
Xfanout782 net784 net782 VPWR VGND sg13g2_buf_8
Xfanout771 net774 net771 VPWR VGND sg13g2_buf_2
XFILLER_46_633 VPWR VGND sg13g2_fill_1
XFILLER_18_335 VPWR VGND sg13g2_fill_1
XFILLER_19_869 VPWR VGND sg13g2_decap_8
XFILLER_27_880 VPWR VGND sg13g2_decap_8
XFILLER_34_839 VPWR VGND sg13g2_decap_8
XFILLER_14_530 VPWR VGND sg13g2_fill_2
X_5170_ _1952_ _1945_ _1953_ VPWR VGND sg13g2_xor2_1
X_4121_ _0948_ net992 net1031 VPWR VGND sg13g2_nand2_1
X_4052_ _0846_ _0880_ _0844_ _0882_ VPWR VGND sg13g2_nand3_1
XFILLER_49_493 VPWR VGND sg13g2_decap_8
Xinput4 ui_in[3] net4 VPWR VGND sg13g2_buf_1
X_3003_ VPWR DP_3.Q_range.data_plus_4\[6\] net12 VGND sg13g2_inv_1
XFILLER_25_817 VPWR VGND sg13g2_decap_8
XFILLER_24_327 VPWR VGND sg13g2_fill_1
XFILLER_37_688 VPWR VGND sg13g2_fill_2
X_4954_ _1742_ _1743_ _1744_ VPWR VGND sg13g2_nor2b_1
X_3905_ _0701_ _0736_ _0738_ VPWR VGND sg13g2_and2_1
X_4885_ _1679_ _1658_ _1681_ VPWR VGND sg13g2_xor2_1
X_3836_ _0670_ _0647_ _0671_ VPWR VGND sg13g2_xor2_1
X_3767_ _0607_ _0601_ _0609_ VPWR VGND sg13g2_xor2_1
X_5506_ _2244_ mac2.sum_lvl2_ff\[26\] mac2.sum_lvl2_ff\[7\] VPWR VGND sg13g2_nand2_1
X_3698_ _0541_ _0542_ _0543_ VPWR VGND sg13g2_nor2_1
X_6486_ net1078 VGND VPWR net453 mac2.sum_lvl3_ff\[4\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_5437_ mac1.sum_lvl3_ff\[28\] mac1.sum_lvl3_ff\[8\] _2190_ VPWR VGND sg13g2_and2_1
XFILLER_0_905 VPWR VGND sg13g2_decap_8
X_5368_ net377 _2136_ _0014_ VPWR VGND sg13g2_nor2b_1
X_5299_ _2076_ _2077_ _2078_ VPWR VGND sg13g2_and2_1
X_4319_ _1134_ _1133_ _0135_ VPWR VGND sg13g2_xor2_1
XFILLER_15_305 VPWR VGND sg13g2_fill_1
XFILLER_24_861 VPWR VGND sg13g2_fill_2
XFILLER_47_920 VPWR VGND sg13g2_decap_8
XFILLER_18_110 VPWR VGND sg13g2_fill_1
XFILLER_47_997 VPWR VGND sg13g2_decap_8
XFILLER_22_809 VPWR VGND sg13g2_fill_2
XFILLER_33_113 VPWR VGND sg13g2_decap_4
X_4670_ DP_3.matrix\[1\] net834 net904 _1471_ VPWR VGND net832 sg13g2_nand4_1
X_3621_ _0467_ _0460_ _0468_ VPWR VGND sg13g2_xor2_1
XFILLER_30_897 VPWR VGND sg13g2_decap_8
X_3552_ _0395_ _0399_ _0400_ VPWR VGND sg13g2_nor2_1
X_6340_ net1061 VGND VPWR net128 mac2.sum_lvl3_ff\[27\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_6_570 VPWR VGND sg13g2_fill_2
X_3483_ _0333_ _0328_ _0331_ VPWR VGND sg13g2_xnor2_1
X_6271_ net1064 VGND VPWR net193 mac1.sum_lvl1_ff\[74\] clknet_leaf_66_clk sg13g2_dfrbpq_1
X_5222_ _2003_ net798 net854 VPWR VGND sg13g2_nand2_1
X_5153_ _1936_ _1929_ _1935_ VPWR VGND sg13g2_xnor2_1
XFILLER_5_1009 VPWR VGND sg13g2_decap_8
X_4104_ _0930_ _0921_ _0932_ VPWR VGND sg13g2_xor2_1
X_5084_ _1845_ _1866_ _1868_ _1869_ VPWR VGND sg13g2_or3_1
X_4035_ VGND VPWR net937 net986 _0865_ _0834_ sg13g2_a21oi_1
XFILLER_38_975 VPWR VGND sg13g2_decap_8
XFILLER_37_474 VPWR VGND sg13g2_fill_2
XFILLER_24_113 VPWR VGND sg13g2_fill_2
X_5986_ net873 _0234_ VPWR VGND sg13g2_buf_1
X_4937_ VGND VPWR _1699_ _1723_ _1730_ _1725_ sg13g2_a21oi_1
X_4868_ _1634_ VPWR _1664_ VGND _1632_ _1635_ sg13g2_o21ai_1
X_3819_ _0655_ net996 net942 net997 net939 VPWR VGND sg13g2_a22oi_1
X_4799_ _1597_ net900 net1023 VPWR VGND sg13g2_nand2_1
X_6469_ net1100 VGND VPWR net73 mac2.sum_lvl2_ff\[22\] clknet_leaf_29_clk sg13g2_dfrbpq_1
XFILLER_29_953 VPWR VGND sg13g2_decap_8
XFILLER_44_923 VPWR VGND sg13g2_decap_8
XFILLER_47_761 VPWR VGND sg13g2_fill_1
XFILLER_35_923 VPWR VGND sg13g2_decap_8
XFILLER_47_794 VPWR VGND sg13g2_fill_2
X_5840_ _2526_ _2529_ _2532_ _2533_ VPWR VGND sg13g2_nor3_1
X_5771_ _2466_ _2465_ _2441_ VPWR VGND sg13g2_nand2b_1
X_4722_ _1522_ net839 net894 VPWR VGND sg13g2_nand2_1
X_4653_ _1455_ _1448_ _1453_ _1454_ VPWR VGND sg13g2_and3_1
X_3604_ _0451_ _0444_ _0450_ VPWR VGND sg13g2_xnor2_1
X_4584_ _1388_ net837 net903 net839 net901 VPWR VGND sg13g2_a22oi_1
X_3535_ _0360_ _0381_ _0383_ _0384_ VPWR VGND sg13g2_or3_1
X_6323_ net1066 VGND VPWR net511 mac1.sum_lvl3_ff\[6\] clknet_leaf_63_clk sg13g2_dfrbpq_2
X_3466_ _0315_ _0314_ _0276_ _0317_ VPWR VGND sg13g2_a21o_1
X_6254_ net1084 VGND VPWR net87 mac2.sum_lvl2_ff\[39\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_5205_ _1987_ _1977_ _1986_ VPWR VGND sg13g2_nand2b_1
X_6185_ net1087 VGND VPWR _0264_ DP_4.matrix\[76\] clknet_leaf_24_clk sg13g2_dfrbpq_1
X_3397_ _2980_ net1018 net956 _0069_ VPWR VGND sg13g2_and3_2
X_5136_ _1918_ _1919_ _1917_ _1920_ VPWR VGND sg13g2_nand3_1
X_5067_ _1852_ _1814_ _1849_ VPWR VGND sg13g2_xnor2_1
X_4018_ _0849_ _0812_ _0847_ VPWR VGND sg13g2_nand2_1
XFILLER_26_945 VPWR VGND sg13g2_decap_8
X_5969_ net929 _0209_ VPWR VGND sg13g2_buf_1
XFILLER_40_458 VPWR VGND sg13g2_decap_4
XFILLER_21_683 VPWR VGND sg13g2_decap_8
XFILLER_0_521 VPWR VGND sg13g2_fill_1
XFILLER_17_978 VPWR VGND sg13g2_decap_8
XFILLER_32_915 VPWR VGND sg13g2_decap_8
XFILLER_12_683 VPWR VGND sg13g2_fill_1
Xhold109 mac1.sum_lvl1_ff\[37\] VPWR VGND net149 sg13g2_dlygate4sd3_1
X_3320_ _2876_ VPWR _2908_ VGND _2874_ _2877_ sg13g2_o21ai_1
X_3251_ _2841_ net973 net907 VPWR VGND sg13g2_nand2_1
X_3182_ _2769_ VPWR _2774_ VGND _2770_ _2772_ sg13g2_o21ai_1
XFILLER_39_536 VPWR VGND sg13g2_decap_4
XFILLER_39_547 VPWR VGND sg13g2_fill_1
XFILLER_35_753 VPWR VGND sg13g2_fill_2
X_5823_ net778 _2515_ _2516_ VPWR VGND sg13g2_and2_1
X_5754_ _2449_ net272 net790 VPWR VGND sg13g2_nand2_1
XFILLER_22_469 VPWR VGND sg13g2_decap_4
XFILLER_33_1003 VPWR VGND sg13g2_decap_8
X_5685_ net22 _2381_ _2384_ VPWR VGND sg13g2_xnor2_1
X_4705_ _1506_ _1504_ _1505_ VPWR VGND sg13g2_nand2_1
X_4636_ _1438_ net904 net835 VPWR VGND sg13g2_nand2_1
X_6306_ net1049 VGND VPWR net68 mac1.sum_lvl3_ff\[25\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_4567_ _1371_ _1372_ _1373_ VPWR VGND sg13g2_nor2b_1
X_4498_ _1308_ _1288_ _1310_ VPWR VGND sg13g2_xor2_1
X_3518_ _0367_ _0329_ _0364_ VPWR VGND sg13g2_xnor2_1
X_3449_ _0300_ _0299_ _0296_ VPWR VGND sg13g2_nand2b_1
X_6237_ net1041 VGND VPWR net200 mac1.sum_lvl2_ff\[38\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_6168_ net1125 VGND VPWR net231 mac1.sum_lvl1_ff\[15\] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_5119_ _1898_ VPWR _1903_ VGND _1899_ _1901_ sg13g2_o21ai_1
X_6099_ net1042 VGND VPWR _0103_ mac1.products_ff\[144\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_26_720 VPWR VGND sg13g2_fill_2
XFILLER_5_635 VPWR VGND sg13g2_fill_2
XFILLER_4_156 VPWR VGND sg13g2_fill_2
XFILLER_36_506 VPWR VGND sg13g2_decap_8
XFILLER_48_399 VPWR VGND sg13g2_fill_2
XFILLER_1_1001 VPWR VGND sg13g2_decap_8
XFILLER_44_583 VPWR VGND sg13g2_fill_2
X_5470_ mac1.sum_lvl3_ff\[34\] mac1.sum_lvl3_ff\[14\] _2217_ VPWR VGND sg13g2_nor2_1
X_4421_ _1209_ VPWR _1235_ VGND _1203_ _1210_ sg13g2_o21ai_1
X_4352_ _1165_ _1166_ _1148_ _1168_ VPWR VGND sg13g2_nand3_1
X_3303_ _2892_ _2882_ _2890_ VPWR VGND sg13g2_xnor2_1
X_4283_ DP_3.matrix\[37\] net816 net887 _1100_ VPWR VGND net814 sg13g2_nand4_1
X_3234_ _2825_ _2810_ _2824_ VPWR VGND sg13g2_nand2_1
X_6022_ net1092 VGND VPWR _0105_ mac1.products_ff\[5\] clknet_leaf_55_clk sg13g2_dfrbpq_1
X_3165_ _2755_ _2751_ _2757_ VPWR VGND sg13g2_xor2_1
X_3096_ _2661_ VPWR _2690_ VGND _2659_ _2662_ sg13g2_o21ai_1
XFILLER_35_561 VPWR VGND sg13g2_fill_1
XFILLER_22_211 VPWR VGND sg13g2_fill_2
XFILLER_22_222 VPWR VGND sg13g2_fill_1
X_3998_ VGND VPWR _0829_ _0828_ _0779_ sg13g2_or2_1
X_5806_ _2499_ _2497_ _2500_ VPWR VGND sg13g2_nor2b_1
X_5737_ VGND VPWR net773 _2432_ _2433_ _2406_ sg13g2_a21oi_1
X_5668_ _2371_ _2368_ _2370_ VPWR VGND sg13g2_nand2_1
X_5599_ _2317_ mac2.sum_lvl3_ff\[31\] mac2.sum_lvl3_ff\[11\] VPWR VGND sg13g2_xnor2_1
X_4619_ _1417_ VPWR _1422_ VGND _1418_ _1420_ sg13g2_o21ai_1
Xhold440 DP_4.matrix\[5\] VPWR VGND net480 sg13g2_dlygate4sd3_1
XFILLER_1_115 VPWR VGND sg13g2_fill_2
Xhold462 _2182_ VPWR VGND net502 sg13g2_dlygate4sd3_1
Xhold451 _2248_ VPWR VGND net491 sg13g2_dlygate4sd3_1
Xhold484 DP_1.matrix\[3\] VPWR VGND net524 sg13g2_dlygate4sd3_1
Xhold473 _2121_ VPWR VGND net513 sg13g2_dlygate4sd3_1
XFILLER_1_126 VPWR VGND sg13g2_fill_1
Xhold495 DP_2.matrix\[8\] VPWR VGND net535 sg13g2_dlygate4sd3_1
Xfanout942 net405 net942 VPWR VGND sg13g2_buf_2
Xfanout920 DP_2.matrix\[73\] net920 VPWR VGND sg13g2_buf_1
Xfanout931 net932 net931 VPWR VGND sg13g2_buf_8
Xfanout975 net977 net975 VPWR VGND sg13g2_buf_8
Xfanout964 net965 net964 VPWR VGND sg13g2_buf_2
Xfanout953 DP_2.matrix\[3\] net953 VPWR VGND sg13g2_buf_1
Xfanout986 net987 net986 VPWR VGND sg13g2_buf_2
Xfanout997 net998 net997 VPWR VGND sg13g2_buf_8
XFILLER_13_222 VPWR VGND sg13g2_fill_2
XFILLER_13_266 VPWR VGND sg13g2_fill_1
XFILLER_14_767 VPWR VGND sg13g2_fill_1
XFILLER_10_973 VPWR VGND sg13g2_decap_8
Xclkload18 clkload18/Y clknet_leaf_31_clk VPWR VGND sg13g2_inv_2
XFILLER_5_465 VPWR VGND sg13g2_fill_1
XFILLER_6_999 VPWR VGND sg13g2_decap_8
XFILLER_23_1013 VPWR VGND sg13g2_decap_8
X_4970_ _0092_ _1745_ _1757_ VPWR VGND sg13g2_xnor2_1
X_3921_ _0751_ _0752_ _0733_ _0754_ VPWR VGND sg13g2_nand3_1
X_3852_ _0685_ _0684_ _0667_ _0687_ VPWR VGND sg13g2_a21o_1
X_3783_ _0111_ _0616_ _0623_ VPWR VGND sg13g2_xnor2_1
X_5522_ VPWR _2257_ _2256_ VGND sg13g2_inv_1
X_5453_ _2203_ mac1.sum_lvl3_ff\[31\] mac1.sum_lvl3_ff\[11\] VPWR VGND sg13g2_nand2_1
X_5384_ _2149_ net546 net481 VPWR VGND sg13g2_nand2_1
X_4404_ _1183_ _1218_ _1219_ VPWR VGND sg13g2_nor2_1
XFILLER_5_81 VPWR VGND sg13g2_fill_2
X_4335_ _1151_ net821 net877 VPWR VGND sg13g2_nand2_1
XFILLER_8_1018 VPWR VGND sg13g2_decap_8
X_4266_ _1084_ _1077_ _1082_ _1083_ VPWR VGND sg13g2_and3_1
X_3217_ _2799_ _2807_ _2808_ VPWR VGND sg13g2_nor2_1
X_4197_ _1017_ net820 net887 net822 net884 VPWR VGND sg13g2_a22oi_1
X_6005_ net810 _0261_ VPWR VGND sg13g2_buf_1
X_3148_ _2716_ VPWR _2741_ VGND _2737_ _2739_ sg13g2_o21ai_1
XFILLER_28_859 VPWR VGND sg13g2_decap_8
XFILLER_27_358 VPWR VGND sg13g2_fill_1
X_3079_ _2672_ _2673_ _2674_ VPWR VGND sg13g2_and2_1
XFILLER_10_269 VPWR VGND sg13g2_fill_2
XFILLER_3_947 VPWR VGND sg13g2_decap_8
XFILLER_46_1013 VPWR VGND sg13g2_decap_8
Xhold270 mac2.sum_lvl3_ff\[12\] VPWR VGND net310 sg13g2_dlygate4sd3_1
Xhold281 _2180_ VPWR VGND net321 sg13g2_dlygate4sd3_1
Xhold292 DP_3.matrix\[0\] VPWR VGND net332 sg13g2_dlygate4sd3_1
Xfanout794 net302 net794 VPWR VGND sg13g2_buf_2
Xfanout783 net784 net783 VPWR VGND sg13g2_buf_8
Xfanout772 net774 net772 VPWR VGND sg13g2_buf_8
XFILLER_45_100 VPWR VGND sg13g2_fill_1
XFILLER_34_818 VPWR VGND sg13g2_decap_8
XFILLER_42_884 VPWR VGND sg13g2_decap_8
XFILLER_14_575 VPWR VGND sg13g2_fill_1
XFILLER_6_763 VPWR VGND sg13g2_fill_1
XFILLER_5_284 VPWR VGND sg13g2_fill_2
XFILLER_2_980 VPWR VGND sg13g2_decap_8
X_4120_ _0926_ VPWR _0947_ VGND _0923_ _0927_ sg13g2_o21ai_1
X_4051_ VGND VPWR _0844_ _0846_ _0881_ _0880_ sg13g2_a21oi_1
X_3002_ VPWR DP_3.I_range.data_plus_4\[6\] net16 VGND sg13g2_inv_1
Xinput5 ui_in[4] net5 VPWR VGND sg13g2_buf_1
XFILLER_17_380 VPWR VGND sg13g2_fill_2
X_4953_ _1739_ VPWR _1743_ VGND _1740_ _1741_ sg13g2_o21ai_1
X_3904_ VGND VPWR _0737_ _0735_ _0702_ sg13g2_or2_1
X_4884_ _1679_ _1658_ _1680_ VPWR VGND sg13g2_nor2b_1
XFILLER_33_884 VPWR VGND sg13g2_decap_8
X_3835_ _0670_ net1000 net933 VPWR VGND sg13g2_nand2_1
X_3766_ _0608_ _0601_ _0607_ VPWR VGND sg13g2_nand2_1
X_6485_ net1085 VGND VPWR net355 mac2.sum_lvl3_ff\[3\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_5505_ _2242_ net519 _0044_ VPWR VGND sg13g2_nor2b_2
X_5436_ _2188_ _2189_ _0029_ VPWR VGND sg13g2_and2_1
X_3697_ VGND VPWR _0505_ _0507_ _0542_ _0539_ sg13g2_a21oi_1
X_5367_ _2132_ net376 _2130_ _2136_ VPWR VGND sg13g2_nand3_1
X_5298_ _2050_ _2052_ _2075_ _2077_ VPWR VGND sg13g2_or3_1
X_4318_ _1135_ _1133_ _1134_ VPWR VGND sg13g2_nand2_1
X_4249_ _1067_ net887 net817 VPWR VGND sg13g2_nand2_1
XFILLER_19_68 VPWR VGND sg13g2_fill_1
XFILLER_43_648 VPWR VGND sg13g2_fill_1
XFILLER_13_1012 VPWR VGND sg13g2_decap_8
XFILLER_47_976 VPWR VGND sg13g2_decap_8
XFILLER_19_667 VPWR VGND sg13g2_decap_4
XFILLER_20_1027 VPWR VGND sg13g2_fill_2
XFILLER_19_689 VPWR VGND sg13g2_fill_1
XFILLER_34_659 VPWR VGND sg13g2_fill_2
XFILLER_33_169 VPWR VGND sg13g2_fill_1
X_3620_ _0467_ _0461_ _0465_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_876 VPWR VGND sg13g2_decap_8
X_3551_ VGND VPWR _0399_ _0398_ _0397_ sg13g2_or2_1
X_3482_ _0332_ _0331_ _0328_ VPWR VGND sg13g2_nand2b_1
X_6270_ net1049 VGND VPWR net67 mac1.sum_lvl1_ff\[73\] clknet_leaf_67_clk sg13g2_dfrbpq_1
X_5221_ _1985_ _1978_ _1948_ _2002_ VPWR VGND sg13g2_a21o_2
X_5152_ _1935_ _1930_ _1933_ VPWR VGND sg13g2_xnor2_1
X_4103_ _0930_ _0921_ _0931_ VPWR VGND sg13g2_nor2b_1
X_5083_ VGND VPWR _1864_ _1865_ _1868_ _1846_ sg13g2_a21oi_1
XFILLER_49_291 VPWR VGND sg13g2_fill_1
X_4034_ _0838_ VPWR _0864_ VGND _0832_ _0839_ sg13g2_o21ai_1
XFILLER_38_954 VPWR VGND sg13g2_decap_8
XFILLER_25_604 VPWR VGND sg13g2_fill_1
X_5985_ net876 _0233_ VPWR VGND sg13g2_buf_1
X_4936_ VGND VPWR _1712_ _1728_ _1729_ _1727_ sg13g2_a21oi_1
XFILLER_33_681 VPWR VGND sg13g2_decap_4
X_4867_ _1642_ VPWR _1663_ VGND _1640_ _1643_ sg13g2_o21ai_1
XFILLER_20_331 VPWR VGND sg13g2_fill_2
X_3818_ net939 net997 net942 _0654_ VPWR VGND net994 sg13g2_nand4_1
XFILLER_20_375 VPWR VGND sg13g2_decap_4
X_4798_ _1571_ VPWR _1596_ VGND _1569_ _1572_ sg13g2_o21ai_1
X_3749_ _0565_ _0567_ _0590_ _0592_ VPWR VGND sg13g2_or3_1
X_6468_ net1099 VGND VPWR net63 mac2.sum_lvl2_ff\[21\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_5419_ net406 mac1.sum_lvl3_ff\[4\] _2176_ VPWR VGND sg13g2_and2_1
X_6399_ net1080 VGND VPWR _0091_ mac2.products_ff\[138\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_43_1027 VPWR VGND sg13g2_fill_2
XFILLER_43_1016 VPWR VGND sg13g2_decap_8
XFILLER_29_932 VPWR VGND sg13g2_decap_8
XFILLER_44_902 VPWR VGND sg13g2_decap_8
XFILLER_44_979 VPWR VGND sg13g2_decap_8
XFILLER_8_858 VPWR VGND sg13g2_fill_1
Xclkbuf_4_9_0_clk clknet_0_clk clknet_4_9_0_clk VPWR VGND sg13g2_buf_8
XFILLER_4_1021 VPWR VGND sg13g2_decap_8
XFILLER_35_902 VPWR VGND sg13g2_decap_8
XFILLER_46_261 VPWR VGND sg13g2_fill_1
XFILLER_35_979 VPWR VGND sg13g2_decap_8
X_5770_ _2464_ _2462_ _2465_ VPWR VGND sg13g2_nor2b_1
XFILLER_22_618 VPWR VGND sg13g2_fill_1
XFILLER_34_478 VPWR VGND sg13g2_fill_1
X_4721_ _1521_ net838 net893 VPWR VGND sg13g2_nand2_2
X_4652_ _1449_ VPWR _1454_ VGND _1450_ _1452_ sg13g2_o21ai_1
X_3603_ _0450_ _0445_ _0448_ VPWR VGND sg13g2_xnor2_1
X_4583_ _0087_ _1374_ _1386_ VPWR VGND sg13g2_xnor2_1
X_3534_ VGND VPWR _0379_ _0380_ _0383_ _0361_ sg13g2_a21oi_1
X_6322_ net1064 VGND VPWR net507 mac1.sum_lvl3_ff\[5\] clknet_leaf_64_clk sg13g2_dfrbpq_2
X_3465_ _0314_ _0315_ _0276_ _0316_ VPWR VGND sg13g2_nand3_1
X_6253_ net1083 VGND VPWR net242 mac2.sum_lvl2_ff\[38\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_5204_ _1986_ _1978_ _1985_ VPWR VGND sg13g2_xnor2_1
X_6184_ net1081 VGND VPWR _0263_ DP_4.matrix\[75\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_3396_ net1019 net960 _0069_ VPWR VGND sg13g2_and2_1
X_5135_ _1871_ VPWR _1919_ VGND _1810_ _1872_ sg13g2_o21ai_1
X_5066_ _1814_ _1849_ _1851_ VPWR VGND sg13g2_and2_1
X_4017_ _0812_ _0847_ _0848_ VPWR VGND sg13g2_nor2_1
XFILLER_26_924 VPWR VGND sg13g2_decap_8
XFILLER_38_773 VPWR VGND sg13g2_fill_2
XFILLER_37_261 VPWR VGND sg13g2_fill_1
X_5968_ net931 _0208_ VPWR VGND sg13g2_buf_1
XFILLER_41_949 VPWR VGND sg13g2_decap_8
X_4919_ _1701_ _1703_ _1713_ VPWR VGND sg13g2_and2_1
X_5899_ net901 net768 _2574_ VPWR VGND sg13g2_nor2_1
XFILLER_32_68 VPWR VGND sg13g2_fill_2
XFILLER_10_1015 VPWR VGND sg13g2_decap_8
XFILLER_48_537 VPWR VGND sg13g2_decap_4
XFILLER_17_957 VPWR VGND sg13g2_decap_8
XFILLER_43_253 VPWR VGND sg13g2_fill_2
XFILLER_31_404 VPWR VGND sg13g2_fill_1
XFILLER_7_187 VPWR VGND sg13g2_fill_1
XFILLER_7_176 VPWR VGND sg13g2_fill_2
X_3250_ _2840_ net973 net905 VPWR VGND sg13g2_nand2_1
XFILLER_26_1022 VPWR VGND sg13g2_decap_8
X_3181_ _2769_ _2770_ _2772_ _2773_ VPWR VGND sg13g2_or3_1
X_5822_ DP_4.matrix\[44\] net1023 net787 _2515_ VPWR VGND sg13g2_mux2_1
X_5753_ net956 net789 _2448_ VPWR VGND sg13g2_nor2_1
XFILLER_31_982 VPWR VGND sg13g2_decap_8
X_4704_ _1467_ _1466_ _1465_ _1505_ VPWR VGND sg13g2_a21o_2
X_5684_ _2384_ _2383_ _2382_ VPWR VGND sg13g2_nand2b_1
X_4635_ _1414_ VPWR _1437_ VGND _1389_ _1412_ sg13g2_o21ai_1
X_4566_ _1368_ VPWR _1372_ VGND _1369_ _1370_ sg13g2_o21ai_1
X_6305_ net1050 VGND VPWR net263 mac1.sum_lvl3_ff\[24\] clknet_leaf_66_clk sg13g2_dfrbpq_1
X_3517_ _0329_ _0364_ _0366_ VPWR VGND sg13g2_and2_1
X_4497_ _1308_ _1288_ _1309_ VPWR VGND sg13g2_nor2b_1
X_3448_ _0298_ _0275_ _0299_ VPWR VGND sg13g2_xor2_1
X_6236_ net1128 VGND VPWR net102 mac1.sum_lvl2_ff\[34\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_6167_ net1087 VGND VPWR _0247_ DP_4.matrix\[3\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_3379_ _2963_ _2962_ _2965_ VPWR VGND sg13g2_xor2_1
XFILLER_40_1008 VPWR VGND sg13g2_decap_8
X_5118_ _1898_ _1899_ _1901_ _1902_ VPWR VGND sg13g2_or3_1
X_6098_ net1093 VGND VPWR _0201_ DP_2.matrix\[5\] clknet_leaf_58_clk sg13g2_dfrbpq_2
X_5049_ _1835_ _1811_ _1834_ VPWR VGND sg13g2_xnor2_1
XFILLER_13_404 VPWR VGND sg13g2_fill_2
XFILLER_13_448 VPWR VGND sg13g2_fill_1
XFILLER_41_746 VPWR VGND sg13g2_fill_1
XFILLER_4_113 VPWR VGND sg13g2_fill_2
XFILLER_9_986 VPWR VGND sg13g2_decap_8
X_4420_ _1232_ _1224_ _1234_ VPWR VGND sg13g2_xor2_1
X_4351_ _1167_ _1148_ _1165_ _1166_ VPWR VGND sg13g2_and3_1
X_3302_ _2890_ _2882_ _2891_ VPWR VGND sg13g2_nor2b_1
X_4282_ _1099_ net814 net886 net816 net884 VPWR VGND sg13g2_a22oi_1
X_6021_ net1092 VGND VPWR _0073_ mac1.products_ff\[4\] clknet_leaf_55_clk sg13g2_dfrbpq_1
X_3233_ _2823_ _2816_ _2824_ VPWR VGND sg13g2_xor2_1
X_3164_ _2751_ _2755_ _2756_ VPWR VGND sg13g2_nor2_1
X_3095_ _2689_ _2684_ _2687_ VPWR VGND sg13g2_xnor2_1
XFILLER_35_584 VPWR VGND sg13g2_fill_1
X_3997_ _0828_ net933 net989 VPWR VGND sg13g2_nand2_1
X_5805_ _2499_ _2498_ net777 net775 net865 VPWR VGND sg13g2_a22oi_1
X_5736_ _2432_ _2431_ _2409_ VPWR VGND sg13g2_nand2b_1
X_5667_ _2365_ _2363_ _2364_ _2370_ VPWR VGND sg13g2_a21o_2
X_4618_ _1417_ _1418_ _1420_ _1421_ VPWR VGND sg13g2_or3_1
X_5598_ mac2.sum_lvl3_ff\[31\] mac2.sum_lvl3_ff\[11\] _2316_ VPWR VGND sg13g2_nor2_1
X_4549_ VGND VPWR _1341_ _1357_ _1358_ _1356_ sg13g2_a21oi_1
Xhold463 _2185_ VPWR VGND net503 sg13g2_dlygate4sd3_1
Xhold441 mac1.sum_lvl2_ff\[12\] VPWR VGND net481 sg13g2_dlygate4sd3_1
Xhold452 _2249_ VPWR VGND net492 sg13g2_dlygate4sd3_1
Xhold430 _0052_ VPWR VGND net470 sg13g2_dlygate4sd3_1
Xhold496 DP_3.matrix\[8\] VPWR VGND net536 sg13g2_dlygate4sd3_1
Xhold474 _0010_ VPWR VGND net514 sg13g2_dlygate4sd3_1
Xhold485 DP_3.matrix\[3\] VPWR VGND net525 sg13g2_dlygate4sd3_1
Xfanout932 net534 net932 VPWR VGND sg13g2_buf_2
Xfanout943 net405 net943 VPWR VGND sg13g2_buf_8
Xfanout921 net923 net921 VPWR VGND sg13g2_buf_2
Xfanout910 net347 net910 VPWR VGND sg13g2_buf_1
X_6219_ net1128 VGND VPWR net133 mac1.sum_lvl2_ff\[14\] clknet_leaf_40_clk sg13g2_dfrbpq_1
Xfanout954 net393 net954 VPWR VGND sg13g2_buf_8
Xfanout976 net977 net976 VPWR VGND sg13g2_buf_1
Xfanout965 net966 net965 VPWR VGND sg13g2_buf_8
Xfanout998 net498 net998 VPWR VGND sg13g2_buf_8
Xfanout987 net988 net987 VPWR VGND sg13g2_buf_1
XFILLER_41_576 VPWR VGND sg13g2_fill_1
Xclkload19 clkload19/Y clknet_leaf_32_clk VPWR VGND sg13g2_inv_2
XFILLER_6_978 VPWR VGND sg13g2_decap_8
XFILLER_45_882 VPWR VGND sg13g2_decap_8
X_3920_ _0753_ _0733_ _0751_ _0752_ VPWR VGND sg13g2_and3_1
XFILLER_32_521 VPWR VGND sg13g2_decap_4
X_3851_ _0684_ _0685_ _0667_ _0686_ VPWR VGND sg13g2_nand3_1
X_3782_ _0623_ _0617_ _0622_ VPWR VGND sg13g2_xnor2_1
X_5521_ mac2.sum_lvl2_ff\[10\] mac2.sum_lvl2_ff\[29\] _2256_ VPWR VGND sg13g2_xor2_1
X_5452_ mac1.sum_lvl3_ff\[31\] mac1.sum_lvl3_ff\[11\] _2202_ VPWR VGND sg13g2_nor2_1
X_5383_ _0002_ _2147_ _2148_ VPWR VGND sg13g2_xnor2_1
X_4403_ _1218_ _1184_ _1216_ VPWR VGND sg13g2_xnor2_1
X_4334_ _1150_ net819 net877 VPWR VGND sg13g2_nand2_2
X_4265_ _1078_ VPWR _1083_ VGND _1079_ _1081_ sg13g2_o21ai_1
X_6004_ net813 _0260_ VPWR VGND sg13g2_buf_1
X_3216_ _2807_ _2800_ _2806_ VPWR VGND sg13g2_xnor2_1
X_4196_ _0082_ _1003_ _1015_ VPWR VGND sg13g2_xnor2_1
X_3147_ _2716_ _2737_ _2739_ _2740_ VPWR VGND sg13g2_or3_1
XFILLER_39_164 VPWR VGND sg13g2_decap_8
XFILLER_39_197 VPWR VGND sg13g2_fill_1
X_3078_ _2671_ _2670_ _2632_ _2673_ VPWR VGND sg13g2_a21o_1
XFILLER_39_1010 VPWR VGND sg13g2_decap_8
XFILLER_24_25 VPWR VGND sg13g2_fill_2
X_5719_ _2415_ _2414_ net782 net781 net273 VPWR VGND sg13g2_a22oi_1
XFILLER_3_904 VPWR VGND sg13g2_fill_1
Xhold260 DP_2.matrix\[78\] VPWR VGND net300 sg13g2_dlygate4sd3_1
Xhold271 _2321_ VPWR VGND net311 sg13g2_dlygate4sd3_1
Xhold282 _0027_ VPWR VGND net322 sg13g2_dlygate4sd3_1
Xhold293 DP_2.matrix\[72\] VPWR VGND net333 sg13g2_dlygate4sd3_1
Xfanout784 _2398_ net784 VPWR VGND sg13g2_buf_8
Xfanout773 net774 net773 VPWR VGND sg13g2_buf_1
Xfanout795 net797 net795 VPWR VGND sg13g2_buf_8
XFILLER_45_167 VPWR VGND sg13g2_fill_2
XFILLER_42_863 VPWR VGND sg13g2_decap_8
XFILLER_6_742 VPWR VGND sg13g2_fill_2
X_4050_ _0878_ _0851_ _0880_ VPWR VGND sg13g2_xor2_1
X_3001_ VPWR DP_1.I_range.data_plus_4\[6\] net4 VGND sg13g2_inv_1
Xinput6 ui_in[5] net6 VPWR VGND sg13g2_buf_1
X_4952_ _1739_ _1740_ _1741_ _1742_ VPWR VGND sg13g2_nor3_1
X_4883_ _1677_ _1676_ _1679_ VPWR VGND sg13g2_xor2_1
X_3903_ _0736_ net933 net995 VPWR VGND sg13g2_nand2_1
XFILLER_33_863 VPWR VGND sg13g2_decap_8
X_3834_ _0669_ net999 net931 VPWR VGND sg13g2_nand2_1
XFILLER_32_373 VPWR VGND sg13g2_fill_1
X_3765_ _0607_ _0602_ _0605_ VPWR VGND sg13g2_xnor2_1
X_3696_ VPWR _0541_ _0540_ VGND sg13g2_inv_1
X_6484_ net1085 VGND VPWR net307 mac2.sum_lvl3_ff\[2\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_5504_ net518 VPWR _2243_ VGND _2237_ _2241_ sg13g2_o21ai_1
X_5435_ _2181_ _2184_ _2187_ _2189_ VPWR VGND sg13g2_or3_1
X_5366_ VGND VPWR _2130_ _2132_ _2135_ net376 sg13g2_a21oi_1
X_5297_ _2075_ VPWR _2076_ VGND _2050_ _2052_ sg13g2_o21ai_1
X_4317_ _1096_ _1095_ _1094_ _1134_ VPWR VGND sg13g2_a21o_2
XFILLER_19_14 VPWR VGND sg13g2_fill_2
X_4248_ _1043_ VPWR _1066_ VGND _1018_ _1041_ sg13g2_o21ai_1
XFILLER_27_101 VPWR VGND sg13g2_fill_1
X_4179_ _0997_ VPWR _1001_ VGND _0998_ _0999_ sg13g2_o21ai_1
XFILLER_42_104 VPWR VGND sg13g2_fill_1
XFILLER_42_126 VPWR VGND sg13g2_fill_2
XFILLER_47_955 VPWR VGND sg13g2_decap_8
XFILLER_20_1006 VPWR VGND sg13g2_decap_8
XFILLER_15_841 VPWR VGND sg13g2_fill_2
XFILLER_30_855 VPWR VGND sg13g2_decap_8
X_3550_ _0398_ net944 net1017 net946 net1016 VPWR VGND sg13g2_a22oi_1
X_3481_ _0330_ _0297_ _0331_ VPWR VGND sg13g2_xor2_1
X_5220_ _1987_ VPWR _2001_ VGND _1976_ _1988_ sg13g2_o21ai_1
X_5151_ _1934_ _1933_ _1930_ VPWR VGND sg13g2_nand2b_1
X_4102_ _0930_ _0922_ _0929_ VPWR VGND sg13g2_xnor2_1
X_5082_ _1864_ _1865_ _1846_ _1867_ VPWR VGND sg13g2_nand3_1
X_4033_ _0861_ _0853_ _0863_ VPWR VGND sg13g2_xor2_1
XFILLER_38_933 VPWR VGND sg13g2_decap_8
XFILLER_37_454 VPWR VGND sg13g2_fill_2
XFILLER_37_476 VPWR VGND sg13g2_fill_1
X_5984_ net878 _0232_ VPWR VGND sg13g2_buf_1
X_4935_ _1728_ _1712_ _0143_ VPWR VGND sg13g2_xor2_1
XFILLER_36_1013 VPWR VGND sg13g2_decap_8
X_4866_ _1662_ _1661_ _1659_ VPWR VGND sg13g2_nand2b_1
X_4797_ _1563_ VPWR _1595_ VGND _1510_ _1561_ sg13g2_o21ai_1
X_3817_ net942 net939 net998 net996 _0653_ VPWR VGND sg13g2_and4_1
X_3748_ _0590_ VPWR _0591_ VGND _0565_ _0567_ sg13g2_o21ai_1
X_3679_ VGND VPWR _0524_ _0522_ _0517_ sg13g2_or2_1
X_6467_ net1085 VGND VPWR net192 mac2.sum_lvl2_ff\[20\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_5418_ _2173_ VPWR _2175_ VGND _2172_ _2174_ sg13g2_o21ai_1
X_6398_ net1080 VGND VPWR net295 mac2.products_ff\[137\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_5349_ net513 _2119_ _0010_ VPWR VGND sg13g2_xor2_1
XFILLER_29_911 VPWR VGND sg13g2_decap_8
XFILLER_29_988 VPWR VGND sg13g2_decap_8
XFILLER_44_958 VPWR VGND sg13g2_decap_8
XFILLER_16_649 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_50_clk clknet_4_10_0_clk clknet_leaf_50_clk VPWR VGND sg13g2_buf_8
XFILLER_7_303 VPWR VGND sg13g2_fill_2
XFILLER_4_1000 VPWR VGND sg13g2_decap_8
XFILLER_47_796 VPWR VGND sg13g2_fill_1
XFILLER_19_476 VPWR VGND sg13g2_fill_1
XFILLER_35_958 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_41_clk clknet_4_14_0_clk clknet_leaf_41_clk VPWR VGND sg13g2_buf_8
X_4720_ _1520_ net898 net836 VPWR VGND sg13g2_nand2_1
X_4651_ _1449_ _1450_ _1452_ _1453_ VPWR VGND sg13g2_or3_1
X_3602_ _0449_ _0448_ _0445_ VPWR VGND sg13g2_nand2b_1
X_4582_ _1387_ _1386_ _1374_ VPWR VGND sg13g2_nand2b_1
X_6321_ net1064 VGND VPWR net514 mac1.sum_lvl3_ff\[4\] clknet_leaf_64_clk sg13g2_dfrbpq_2
X_3533_ _0379_ _0380_ _0361_ _0382_ VPWR VGND sg13g2_nand3_1
X_3464_ _0313_ _0312_ _0295_ _0315_ VPWR VGND sg13g2_a21o_1
X_6252_ net1075 VGND VPWR net136 mac1.sum_lvl2_ff\[53\] clknet_leaf_59_clk sg13g2_dfrbpq_1
XFILLER_42_0 VPWR VGND sg13g2_fill_1
X_5203_ _1983_ _1984_ _1985_ VPWR VGND sg13g2_nor2b_1
X_6183_ net1082 VGND VPWR _0262_ DP_4.matrix\[74\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_3395_ _0100_ _2972_ _2979_ VPWR VGND sg13g2_xnor2_1
X_5134_ _1844_ VPWR _1918_ VGND _1914_ _1916_ sg13g2_o21ai_1
X_5065_ VGND VPWR _1850_ _1848_ _1815_ sg13g2_or2_1
X_4016_ _0847_ _0813_ _0845_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_903 VPWR VGND sg13g2_decap_8
X_5967_ net933 _0207_ VPWR VGND sg13g2_buf_1
XFILLER_41_928 VPWR VGND sg13g2_decap_8
X_4918_ _1709_ _1687_ _1711_ _1712_ VPWR VGND sg13g2_a21o_1
Xclkbuf_leaf_32_clk clknet_4_13_0_clk clknet_leaf_32_clk VPWR VGND sg13g2_buf_8
X_5898_ _0220_ net903 net767 VPWR VGND sg13g2_xnor2_1
X_4849_ _1645_ _1638_ _1646_ VPWR VGND sg13g2_nor2b_1
XFILLER_4_339 VPWR VGND sg13g2_fill_1
X_6519_ net1056 VGND VPWR net13 DP_3.I_range.out_data\[2\] clknet_leaf_22_clk sg13g2_dfrbpq_2
XFILLER_28_284 VPWR VGND sg13g2_decap_8
XFILLER_44_777 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_23_clk clknet_4_5_0_clk clknet_leaf_23_clk VPWR VGND sg13g2_buf_8
XFILLER_25_991 VPWR VGND sg13g2_decap_8
XFILLER_40_994 VPWR VGND sg13g2_decap_8
XFILLER_7_166 VPWR VGND sg13g2_fill_1
XFILLER_26_1001 VPWR VGND sg13g2_decap_8
X_3180_ _2772_ net1033 net922 net964 net919 VPWR VGND sg13g2_a22oi_1
XFILLER_47_582 VPWR VGND sg13g2_decap_4
X_5821_ _2475_ _2481_ _2514_ _0166_ VPWR VGND sg13g2_mux2_1
XFILLER_16_980 VPWR VGND sg13g2_decap_8
X_5752_ _2447_ _2446_ net782 net781 net924 VPWR VGND sg13g2_a22oi_1
Xclkbuf_leaf_14_clk clknet_4_6_0_clk clknet_leaf_14_clk VPWR VGND sg13g2_buf_8
XFILLER_31_961 VPWR VGND sg13g2_decap_8
X_4703_ _1503_ _1439_ _1504_ VPWR VGND sg13g2_xor2_1
X_5683_ VGND VPWR _2383_ mac2.total_sum\[13\] mac1.total_sum\[13\] sg13g2_or2_1
X_4634_ _1436_ _1428_ _1430_ VPWR VGND sg13g2_nand2_1
X_4565_ _1368_ _1369_ _1370_ _1371_ VPWR VGND sg13g2_nor3_1
X_6304_ net1050 VGND VPWR net89 mac1.sum_lvl3_ff\[23\] clknet_leaf_66_clk sg13g2_dfrbpq_1
X_3516_ VGND VPWR _0365_ _0363_ _0330_ sg13g2_or2_1
X_4496_ _1306_ _1305_ _1308_ VPWR VGND sg13g2_xor2_1
X_3447_ _0298_ net1016 net952 VPWR VGND sg13g2_nand2_1
X_6235_ net1115 VGND VPWR net218 mac1.sum_lvl2_ff\[33\] clknet_leaf_47_clk sg13g2_dfrbpq_2
X_3378_ _2964_ _2962_ _2963_ VPWR VGND sg13g2_nand2_1
X_6166_ net1087 VGND VPWR _0246_ DP_4.matrix\[2\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_5117_ _1901_ net1025 net813 net853 net807 VPWR VGND sg13g2_a22oi_1
X_6097_ net1093 VGND VPWR _0200_ DP_2.matrix\[4\] clknet_leaf_59_clk sg13g2_dfrbpq_1
X_5048_ _1834_ _1831_ _1833_ VPWR VGND sg13g2_nand2_1
Xclkbuf_4_8_0_clk clknet_0_clk clknet_4_8_0_clk VPWR VGND sg13g2_buf_8
XFILLER_43_68 VPWR VGND sg13g2_fill_2
XFILLER_22_983 VPWR VGND sg13g2_decap_8
XFILLER_48_302 VPWR VGND sg13g2_fill_2
XFILLER_0_342 VPWR VGND sg13g2_fill_1
XFILLER_44_574 VPWR VGND sg13g2_decap_4
XFILLER_44_563 VPWR VGND sg13g2_fill_2
XFILLER_17_80 VPWR VGND sg13g2_fill_1
XFILLER_16_287 VPWR VGND sg13g2_fill_2
X_4350_ _1154_ VPWR _1166_ VGND _1162_ _1164_ sg13g2_o21ai_1
X_3301_ _2890_ _2883_ _2889_ VPWR VGND sg13g2_xnor2_1
X_4281_ _1075_ VPWR _1098_ VGND _1040_ _1073_ sg13g2_o21ai_1
X_3232_ _2823_ _2817_ _2821_ VPWR VGND sg13g2_xnor2_1
X_6020_ net1092 VGND VPWR _0072_ mac1.products_ff\[3\] clknet_leaf_55_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_3_clk clknet_4_3_0_clk clknet_leaf_3_clk VPWR VGND sg13g2_buf_8
X_3163_ VGND VPWR _2755_ _2754_ _2753_ sg13g2_or2_1
XFILLER_39_346 VPWR VGND sg13g2_fill_2
XFILLER_48_891 VPWR VGND sg13g2_decap_8
X_3094_ _2688_ _2687_ _2684_ VPWR VGND sg13g2_nand2b_1
X_5804_ net882 net899 net786 _2498_ VPWR VGND sg13g2_mux2_1
X_3996_ _0827_ net994 net929 VPWR VGND sg13g2_nand2_1
X_5735_ _2430_ _2428_ _2431_ VPWR VGND sg13g2_nor2b_1
X_5666_ VPWR _2369_ _2368_ VGND sg13g2_inv_1
X_4617_ _1420_ net894 net850 net895 net846 VPWR VGND sg13g2_a22oi_1
X_5597_ _0049_ _2313_ _2314_ VPWR VGND sg13g2_xnor2_1
Xhold420 mac1.sum_lvl2_ff\[14\] VPWR VGND net460 sg13g2_dlygate4sd3_1
X_4548_ _1357_ _1341_ _0132_ VPWR VGND sg13g2_xor2_1
Xhold431 DP_1.matrix\[2\] VPWR VGND net471 sg13g2_dlygate4sd3_1
Xhold442 _2151_ VPWR VGND net482 sg13g2_dlygate4sd3_1
Xhold453 _0046_ VPWR VGND net493 sg13g2_dlygate4sd3_1
X_4479_ VGND VPWR _1291_ _1290_ _1238_ sg13g2_or2_1
Xhold475 DP_1.matrix\[37\] VPWR VGND net515 sg13g2_dlygate4sd3_1
Xhold464 _0028_ VPWR VGND net504 sg13g2_dlygate4sd3_1
Xhold486 DP_1.matrix\[4\] VPWR VGND net526 sg13g2_dlygate4sd3_1
Xfanout900 DP_3.matrix\[2\] net900 VPWR VGND sg13g2_buf_8
Xfanout911 net912 net911 VPWR VGND sg13g2_buf_8
Xfanout922 net923 net922 VPWR VGND sg13g2_buf_1
Xfanout933 net934 net933 VPWR VGND sg13g2_buf_8
X_6218_ net1116 VGND VPWR net58 mac1.sum_lvl2_ff\[13\] clknet_leaf_47_clk sg13g2_dfrbpq_1
Xhold497 mac2.sum_lvl3_ff\[7\] VPWR VGND net537 sg13g2_dlygate4sd3_1
Xfanout977 net303 net977 VPWR VGND sg13g2_buf_2
Xfanout955 DP_2.matrix\[2\] net955 VPWR VGND sg13g2_buf_1
Xfanout966 net304 net966 VPWR VGND sg13g2_buf_2
Xfanout944 DP_2.matrix\[7\] net944 VPWR VGND sg13g2_buf_8
X_6149_ net1123 VGND VPWR _0235_ DP_3.matrix\[43\] clknet_leaf_33_clk sg13g2_dfrbpq_1
Xfanout999 net1000 net999 VPWR VGND sg13g2_buf_8
Xfanout988 DP_1.matrix\[43\] net988 VPWR VGND sg13g2_buf_1
XFILLER_39_891 VPWR VGND sg13g2_decap_8
XFILLER_13_224 VPWR VGND sg13g2_fill_1
XFILLER_41_511 VPWR VGND sg13g2_fill_2
XFILLER_16_1022 VPWR VGND sg13g2_decap_8
XFILLER_6_957 VPWR VGND sg13g2_decap_8
XFILLER_49_611 VPWR VGND sg13g2_decap_4
XFILLER_0_194 VPWR VGND sg13g2_fill_1
XFILLER_36_305 VPWR VGND sg13g2_fill_2
X_3850_ _0673_ VPWR _0685_ VGND _0681_ _0683_ sg13g2_o21ai_1
X_3781_ _0622_ _0608_ _0621_ VPWR VGND sg13g2_xnor2_1
X_5520_ _2255_ mac2.sum_lvl2_ff\[29\] mac2.sum_lvl2_ff\[10\] VPWR VGND sg13g2_nand2_1
XFILLER_9_784 VPWR VGND sg13g2_fill_2
XFILLER_8_272 VPWR VGND sg13g2_fill_1
X_5451_ net349 _2198_ _0017_ VPWR VGND sg13g2_xor2_1
X_5382_ _2148_ _2141_ _2145_ VPWR VGND sg13g2_nand2_1
X_4402_ _1217_ _1184_ _1216_ VPWR VGND sg13g2_nand2b_1
X_4333_ _1149_ net881 DP_4.matrix\[41\] VPWR VGND sg13g2_nand2_1
X_4264_ _1078_ _1079_ _1081_ _1082_ VPWR VGND sg13g2_or3_1
X_6003_ net815 _0259_ VPWR VGND sg13g2_buf_1
X_3215_ _2806_ _2801_ _2804_ VPWR VGND sg13g2_xnor2_1
X_4195_ _1016_ _1015_ _1003_ VPWR VGND sg13g2_nand2b_1
X_3146_ VGND VPWR _2735_ _2736_ _2739_ _2717_ sg13g2_a21oi_1
XFILLER_39_154 VPWR VGND sg13g2_decap_4
X_3077_ _2670_ _2671_ _2632_ _2672_ VPWR VGND sg13g2_nand3_1
XFILLER_36_894 VPWR VGND sg13g2_decap_8
X_5718_ net1003 net1019 net790 _2414_ VPWR VGND sg13g2_mux2_1
X_3979_ _0809_ _0764_ _0125_ VPWR VGND sg13g2_xor2_1
X_5649_ _2354_ _2355_ net31 VPWR VGND sg13g2_nor2b_1
XFILLER_2_426 VPWR VGND sg13g2_fill_2
Xhold250 mac2.sum_lvl3_ff\[0\] VPWR VGND net290 sg13g2_dlygate4sd3_1
Xhold261 DP_4.matrix\[73\] VPWR VGND net301 sg13g2_dlygate4sd3_1
Xhold272 _0051_ VPWR VGND net312 sg13g2_dlygate4sd3_1
Xhold283 DP_3.matrix\[36\] VPWR VGND net323 sg13g2_dlygate4sd3_1
Xhold294 DP_3.matrix\[39\] VPWR VGND net334 sg13g2_dlygate4sd3_1
Xfanout785 _2473_ net785 VPWR VGND sg13g2_buf_8
Xfanout774 _2393_ net774 VPWR VGND sg13g2_buf_2
Xfanout796 net797 net796 VPWR VGND sg13g2_buf_1
XFILLER_27_894 VPWR VGND sg13g2_decap_8
XFILLER_42_842 VPWR VGND sg13g2_decap_8
XFILLER_14_588 VPWR VGND sg13g2_fill_2
XFILLER_46_7 VPWR VGND sg13g2_decap_8
XFILLER_5_286 VPWR VGND sg13g2_fill_1
XFILLER_1_492 VPWR VGND sg13g2_fill_2
X_3000_ VPWR _2604_ DP_3.Q_range.out_data\[5\] VGND sg13g2_inv_1
Xinput7 ui_in[6] net7 VPWR VGND sg13g2_buf_1
XFILLER_36_124 VPWR VGND sg13g2_fill_2
X_4951_ _1741_ net865 net812 net809 net867 VPWR VGND sg13g2_a22oi_1
X_4882_ _1677_ _1676_ _1678_ VPWR VGND sg13g2_nor2b_1
X_3902_ _0735_ net995 net931 VPWR VGND sg13g2_nand2_1
XFILLER_33_842 VPWR VGND sg13g2_decap_8
X_3833_ _0668_ net1003 net929 VPWR VGND sg13g2_nand2_1
X_3764_ _0606_ _0605_ _0602_ VPWR VGND sg13g2_nand2b_1
X_3695_ _0507_ _0539_ _0505_ _0540_ VPWR VGND sg13g2_nand3_1
X_5503_ _2237_ net518 _2241_ _2242_ VPWR VGND sg13g2_nor3_1
X_6483_ net1085 VGND VPWR net285 mac2.sum_lvl3_ff\[1\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_5434_ _2187_ VPWR _2188_ VGND _2181_ _2184_ sg13g2_o21ai_1
X_5365_ _2134_ mac1.sum_lvl2_ff\[27\] net375 VPWR VGND sg13g2_xnor2_1
XFILLER_0_919 VPWR VGND sg13g2_decap_8
X_5296_ _2074_ _2060_ _2075_ VPWR VGND sg13g2_xor2_1
X_4316_ _1132_ _1068_ _1133_ VPWR VGND sg13g2_xor2_1
X_4247_ _1065_ _1057_ _1059_ VPWR VGND sg13g2_nand2_1
X_4178_ _0997_ _0998_ _0999_ _1000_ VPWR VGND sg13g2_nor3_1
X_3129_ _2685_ _2720_ _2722_ VPWR VGND sg13g2_and2_1
XFILLER_24_820 VPWR VGND sg13g2_fill_1
XFILLER_46_400 VPWR VGND sg13g2_fill_2
XFILLER_47_934 VPWR VGND sg13g2_decap_8
XFILLER_30_845 VPWR VGND sg13g2_fill_1
X_3480_ _0330_ net1014 net953 VPWR VGND sg13g2_nand2_1
X_5150_ _1932_ _1881_ _1933_ VPWR VGND sg13g2_xor2_1
X_4101_ _0929_ _0923_ _0928_ VPWR VGND sg13g2_xnor2_1
X_5081_ _1866_ _1846_ _1864_ _1865_ VPWR VGND sg13g2_and3_1
X_4032_ _0861_ _0853_ _0862_ VPWR VGND sg13g2_nor2b_1
XFILLER_38_912 VPWR VGND sg13g2_decap_8
XFILLER_38_989 VPWR VGND sg13g2_decap_8
X_5983_ net880 _0231_ VPWR VGND sg13g2_buf_1
XFILLER_18_680 VPWR VGND sg13g2_fill_1
X_4934_ _1726_ _1713_ _1728_ VPWR VGND sg13g2_xor2_1
X_4865_ VGND VPWR _1661_ _1660_ _1609_ sg13g2_or2_1
XFILLER_20_333 VPWR VGND sg13g2_fill_1
X_3816_ _0652_ net999 net935 VPWR VGND sg13g2_nand2_1
X_4796_ _1583_ VPWR _1594_ VGND _1567_ _1584_ sg13g2_o21ai_1
X_3747_ _0589_ _0575_ _0590_ VPWR VGND sg13g2_xor2_1
X_3678_ _0517_ _0522_ _0523_ VPWR VGND sg13g2_and2_1
X_6466_ net1084 VGND VPWR net49 mac2.sum_lvl2_ff\[19\] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_5417_ net362 _2172_ _0025_ VPWR VGND sg13g2_xor2_1
X_6397_ net1079 VGND VPWR net283 mac2.products_ff\[136\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_5348_ net512 mac1.sum_lvl2_ff\[23\] _2121_ VPWR VGND sg13g2_xor2_1
X_5279_ VGND VPWR _2058_ _2059_ _2057_ _1998_ sg13g2_a21oi_2
XFILLER_29_967 VPWR VGND sg13g2_decap_8
XFILLER_44_937 VPWR VGND sg13g2_decap_8
XFILLER_3_576 VPWR VGND sg13g2_fill_2
XFILLER_38_208 VPWR VGND sg13g2_fill_2
XFILLER_19_433 VPWR VGND sg13g2_fill_2
XFILLER_35_937 VPWR VGND sg13g2_decap_8
XFILLER_43_981 VPWR VGND sg13g2_decap_8
XFILLER_15_683 VPWR VGND sg13g2_fill_1
XFILLER_30_664 VPWR VGND sg13g2_fill_2
X_4650_ _1452_ net892 net849 net893 net846 VPWR VGND sg13g2_a22oi_1
X_3601_ _0447_ _0396_ _0448_ VPWR VGND sg13g2_xor2_1
XFILLER_30_697 VPWR VGND sg13g2_fill_1
Xinput10 uio_in[1] net10 VPWR VGND sg13g2_buf_1
X_6320_ net1076 VGND VPWR net372 mac1.sum_lvl3_ff\[3\] clknet_leaf_62_clk sg13g2_dfrbpq_2
X_4581_ _1385_ _1375_ _1386_ VPWR VGND sg13g2_xor2_1
X_3532_ _0381_ _0361_ _0379_ _0380_ VPWR VGND sg13g2_and3_1
X_3463_ _0312_ _0313_ _0295_ _0314_ VPWR VGND sg13g2_nand3_1
X_6251_ net1074 VGND VPWR net254 mac1.sum_lvl2_ff\[52\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_5202_ _1979_ VPWR _1984_ VGND _1981_ _1982_ sg13g2_o21ai_1
X_6182_ net1082 VGND VPWR _0261_ DP_4.matrix\[73\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_3394_ _2979_ _2973_ _2978_ VPWR VGND sg13g2_xnor2_1
X_5133_ _1844_ _1914_ _1916_ _1917_ VPWR VGND sg13g2_or3_1
XFILLER_35_0 VPWR VGND sg13g2_fill_2
X_5064_ _1849_ net802 net858 VPWR VGND sg13g2_nand2_1
X_4015_ _0846_ _0813_ _0845_ VPWR VGND sg13g2_nand2b_1
XFILLER_26_959 VPWR VGND sg13g2_decap_8
XFILLER_41_907 VPWR VGND sg13g2_decap_8
X_5966_ net935 _0206_ VPWR VGND sg13g2_buf_1
X_4917_ _1711_ _1705_ _1710_ VPWR VGND sg13g2_nand2_1
X_5897_ _2573_ VPWR _0203_ VGND _2606_ net773 sg13g2_o21ai_1
XFILLER_21_631 VPWR VGND sg13g2_fill_1
X_4848_ _1645_ _1639_ _1644_ VPWR VGND sg13g2_xnor2_1
X_4779_ _1578_ net1029 net846 net888 net842 VPWR VGND sg13g2_a22oi_1
X_6518_ net1052 VGND VPWR net8 DP_1.Q_range.out_data\[6\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_6449_ net1053 VGND VPWR net4 DP_1.I_range.out_data\[6\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_0_557 VPWR VGND sg13g2_fill_2
XFILLER_25_970 VPWR VGND sg13g2_decap_8
XFILLER_32_929 VPWR VGND sg13g2_decap_8
XFILLER_40_973 VPWR VGND sg13g2_decap_8
XFILLER_11_196 VPWR VGND sg13g2_fill_1
XFILLER_39_506 VPWR VGND sg13g2_fill_1
XFILLER_39_528 VPWR VGND sg13g2_fill_2
X_5820_ _2514_ net770 _2513_ VPWR VGND sg13g2_nand2_1
XFILLER_23_929 VPWR VGND sg13g2_decap_8
X_5751_ net943 net960 net790 _2446_ VPWR VGND sg13g2_mux2_1
XFILLER_31_940 VPWR VGND sg13g2_decap_8
XFILLER_33_1017 VPWR VGND sg13g2_decap_8
X_4702_ _1503_ _1500_ _1502_ VPWR VGND sg13g2_nand2_1
X_5682_ mac1.total_sum\[13\] mac2.total_sum\[13\] _2382_ VPWR VGND sg13g2_and2_1
XFILLER_33_1028 VPWR VGND sg13g2_fill_1
X_4633_ _0138_ _1408_ _1435_ VPWR VGND sg13g2_xnor2_1
X_4564_ _1370_ net899 net847 net843 net901 VPWR VGND sg13g2_a22oi_1
X_6303_ net1066 VGND VPWR net72 mac1.sum_lvl3_ff\[22\] clknet_leaf_64_clk sg13g2_dfrbpq_1
X_3515_ _0364_ net953 net1012 VPWR VGND sg13g2_nand2_1
X_4495_ _1306_ _1305_ _1307_ VPWR VGND sg13g2_nor2b_1
X_6234_ net1114 VGND VPWR net55 mac1.sum_lvl2_ff\[32\] clknet_leaf_48_clk sg13g2_dfrbpq_1
X_3446_ _0297_ net1016 net950 VPWR VGND sg13g2_nand2_1
X_3377_ _2937_ VPWR _2963_ VGND _2910_ _2935_ sg13g2_o21ai_1
X_6165_ net1125 VGND VPWR net260 mac1.sum_lvl1_ff\[14\] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_6096_ net1042 VGND VPWR _0102_ mac1.products_ff\[143\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_5116_ net806 net851 net813 _1900_ VPWR VGND net1024 sg13g2_nand4_1
X_5047_ _1830_ _1829_ _1812_ _1833_ VPWR VGND sg13g2_a21o_1
XFILLER_26_701 VPWR VGND sg13g2_fill_1
XFILLER_38_572 VPWR VGND sg13g2_fill_2
XFILLER_38_561 VPWR VGND sg13g2_fill_2
XFILLER_13_406 VPWR VGND sg13g2_fill_1
X_5949_ net1001 _0181_ VPWR VGND sg13g2_buf_1
XFILLER_22_962 VPWR VGND sg13g2_decap_8
XFILLER_21_461 VPWR VGND sg13g2_fill_1
XFILLER_49_1013 VPWR VGND sg13g2_decap_8
XFILLER_49_837 VPWR VGND sg13g2_decap_4
XFILLER_1_1015 VPWR VGND sg13g2_decap_8
XFILLER_29_550 VPWR VGND sg13g2_decap_4
XFILLER_31_203 VPWR VGND sg13g2_fill_1
XFILLER_13_984 VPWR VGND sg13g2_decap_8
X_3300_ _2888_ _2884_ _2889_ VPWR VGND sg13g2_xor2_1
X_4280_ _1089_ VPWR _1097_ VGND _1069_ _1090_ sg13g2_o21ai_1
X_3231_ _2822_ _2817_ _2821_ VPWR VGND sg13g2_nand2_1
X_3162_ _2754_ net905 net982 net907 net979 VPWR VGND sg13g2_a22oi_1
X_3093_ _2686_ _2653_ _2687_ VPWR VGND sg13g2_xor2_1
XFILLER_47_380 VPWR VGND sg13g2_fill_1
X_5803_ _2492_ _2496_ _2497_ VPWR VGND sg13g2_and2_1
X_3995_ _0792_ VPWR _0826_ VGND _0783_ _0793_ sg13g2_o21ai_1
X_5734_ _2430_ _2429_ net783 net780 net315 VPWR VGND sg13g2_a22oi_1
X_5665_ mac2.total_sum\[10\] mac1.total_sum\[10\] _2368_ VPWR VGND sg13g2_xor2_1
X_4616_ net846 net895 net850 _1419_ VPWR VGND net894 sg13g2_nand4_1
Xhold410 _0055_ VPWR VGND net450 sg13g2_dlygate4sd3_1
X_5596_ _2315_ _2312_ _2314_ VPWR VGND sg13g2_nand2_1
X_4547_ _1355_ _1342_ _1357_ VPWR VGND sg13g2_xor2_1
Xhold454 DP_2.matrix\[41\] VPWR VGND net494 sg13g2_dlygate4sd3_1
Xhold432 DP_2.matrix\[5\] VPWR VGND net472 sg13g2_dlygate4sd3_1
Xhold443 _0003_ VPWR VGND net483 sg13g2_dlygate4sd3_1
Xhold421 _2162_ VPWR VGND net461 sg13g2_dlygate4sd3_1
Xhold487 mac2.sum_lvl2_ff\[15\] VPWR VGND net527 sg13g2_dlygate4sd3_1
X_4478_ _1290_ net818 net1027 VPWR VGND sg13g2_nand2_1
Xhold465 mac1.sum_lvl2_ff\[24\] VPWR VGND net505 sg13g2_dlygate4sd3_1
Xhold476 DP_3.matrix\[37\] VPWR VGND net516 sg13g2_dlygate4sd3_1
X_3429_ net963 net959 net1013 net1011 _0281_ VPWR VGND sg13g2_and4_1
Xfanout923 net924 net923 VPWR VGND sg13g2_buf_2
Xfanout934 net499 net934 VPWR VGND sg13g2_buf_8
Xfanout912 DP_2.matrix\[76\] net912 VPWR VGND sg13g2_buf_1
X_6217_ net1116 VGND VPWR net95 mac1.sum_lvl2_ff\[12\] clknet_leaf_46_clk sg13g2_dfrbpq_1
Xhold498 _2301_ VPWR VGND net538 sg13g2_dlygate4sd3_1
Xfanout901 net902 net901 VPWR VGND sg13g2_buf_8
X_6148_ net1123 VGND VPWR _0234_ DP_3.matrix\[42\] clknet_leaf_34_clk sg13g2_dfrbpq_1
Xfanout967 net968 net967 VPWR VGND sg13g2_buf_8
Xfanout956 net959 net956 VPWR VGND sg13g2_buf_8
Xfanout945 DP_2.matrix\[7\] net945 VPWR VGND sg13g2_buf_1
Xfanout978 net980 net978 VPWR VGND sg13g2_buf_8
Xfanout989 net990 net989 VPWR VGND sg13g2_buf_8
X_6079_ net1071 VGND VPWR _0188_ DP_1.matrix\[72\] clknet_leaf_60_clk sg13g2_dfrbpq_1
XFILLER_39_870 VPWR VGND sg13g2_decap_8
XFILLER_41_534 VPWR VGND sg13g2_fill_1
XFILLER_16_1001 VPWR VGND sg13g2_decap_8
XFILLER_10_987 VPWR VGND sg13g2_decap_8
XFILLER_23_1027 VPWR VGND sg13g2_fill_2
XFILLER_17_575 VPWR VGND sg13g2_fill_2
XFILLER_20_707 VPWR VGND sg13g2_decap_8
XFILLER_32_567 VPWR VGND sg13g2_fill_1
X_3780_ _0621_ _0618_ _0620_ VPWR VGND sg13g2_xnor2_1
X_5450_ _2201_ _2198_ net349 VPWR VGND sg13g2_nand2_1
XFILLER_30_1009 VPWR VGND sg13g2_decap_8
X_4401_ _1216_ _1185_ _1214_ VPWR VGND sg13g2_xnor2_1
X_5381_ _2147_ mac1.sum_lvl2_ff\[30\] mac1.sum_lvl2_ff\[11\] VPWR VGND sg13g2_xnor2_1
X_4332_ _1120_ VPWR _1148_ VGND _1111_ _1121_ sg13g2_o21ai_1
X_4263_ _1081_ net875 net829 net876 net827 VPWR VGND sg13g2_a22oi_1
X_6002_ net816 _0258_ VPWR VGND sg13g2_buf_1
X_3214_ _2805_ _2804_ _2801_ VPWR VGND sg13g2_nand2b_1
Xclkbuf_4_7_0_clk clknet_0_clk clknet_4_7_0_clk VPWR VGND sg13g2_buf_8
X_4194_ _1014_ _1004_ _1015_ VPWR VGND sg13g2_xor2_1
XFILLER_39_122 VPWR VGND sg13g2_decap_8
X_3145_ _2735_ _2736_ _2717_ _2738_ VPWR VGND sg13g2_nand3_1
X_3076_ _2669_ _2668_ _2651_ _2671_ VPWR VGND sg13g2_a21o_1
XFILLER_36_873 VPWR VGND sg13g2_decap_8
XFILLER_24_27 VPWR VGND sg13g2_fill_1
X_3978_ _0762_ _0763_ _0807_ _0808_ _0810_ VPWR VGND sg13g2_and4_1
X_5717_ _2413_ _2412_ net784 net780 net977 VPWR VGND sg13g2_a22oi_1
X_5648_ _2352_ VPWR _2355_ VGND _2349_ _2353_ sg13g2_o21ai_1
XFILLER_40_59 VPWR VGND sg13g2_fill_2
XFILLER_3_928 VPWR VGND sg13g2_fill_1
XFILLER_3_917 VPWR VGND sg13g2_fill_2
X_5579_ net537 mac2.sum_lvl3_ff\[27\] _2301_ VPWR VGND sg13g2_xor2_1
Xhold262 DP_4.matrix\[79\] VPWR VGND net302 sg13g2_dlygate4sd3_1
Xhold240 DP_3.matrix\[78\] VPWR VGND net280 sg13g2_dlygate4sd3_1
Xhold251 _0048_ VPWR VGND net291 sg13g2_dlygate4sd3_1
XFILLER_46_1027 VPWR VGND sg13g2_fill_2
Xhold284 DP_3.matrix\[7\] VPWR VGND net324 sg13g2_dlygate4sd3_1
Xhold273 DP_3.matrix\[44\] VPWR VGND net313 sg13g2_dlygate4sd3_1
Xhold295 DP_1.matrix\[0\] VPWR VGND net335 sg13g2_dlygate4sd3_1
Xfanout775 _2482_ net775 VPWR VGND sg13g2_buf_8
XFILLER_46_615 VPWR VGND sg13g2_fill_1
Xfanout786 net787 net786 VPWR VGND sg13g2_buf_8
Xfanout797 net352 net797 VPWR VGND sg13g2_buf_1
XFILLER_27_873 VPWR VGND sg13g2_decap_8
XFILLER_42_821 VPWR VGND sg13g2_decap_8
XFILLER_14_501 VPWR VGND sg13g2_fill_2
XFILLER_42_898 VPWR VGND sg13g2_decap_8
XFILLER_41_364 VPWR VGND sg13g2_fill_1
XFILLER_14_82 VPWR VGND sg13g2_fill_2
XFILLER_6_744 VPWR VGND sg13g2_fill_1
XFILLER_2_994 VPWR VGND sg13g2_decap_8
Xinput8 ui_in[7] net8 VPWR VGND sg13g2_buf_1
XFILLER_33_821 VPWR VGND sg13g2_decap_8
X_4950_ net812 net867 net809 net865 _1740_ VPWR VGND sg13g2_and4_1
X_4881_ VGND VPWR _1631_ _1636_ _1677_ _1648_ sg13g2_a21oi_1
X_3901_ _0734_ net999 net930 VPWR VGND sg13g2_nand2_1
X_3832_ _0658_ VPWR _0667_ VGND _0650_ _0659_ sg13g2_o21ai_1
XFILLER_33_898 VPWR VGND sg13g2_decap_8
X_3763_ _0604_ _0578_ _0605_ VPWR VGND sg13g2_xor2_1
X_5502_ VPWR VGND _2235_ _2234_ _2233_ net387 _2241_ mac2.sum_lvl2_ff\[5\] sg13g2_a221oi_1
X_3694_ _0537_ _0515_ _0539_ VPWR VGND sg13g2_xor2_1
X_6482_ net1083 VGND VPWR net268 mac2.sum_lvl3_ff\[0\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_5433_ mac1.sum_lvl3_ff\[7\] net419 _2187_ VPWR VGND sg13g2_xor2_1
X_5364_ _2132_ net531 _0013_ VPWR VGND sg13g2_and2_1
X_4315_ _1132_ _1129_ _1131_ VPWR VGND sg13g2_nand2_1
X_5295_ _2072_ _2047_ _2074_ VPWR VGND sg13g2_xor2_1
XFILLER_19_16 VPWR VGND sg13g2_fill_1
X_4246_ _0127_ _1037_ _1064_ VPWR VGND sg13g2_xnor2_1
X_4177_ _0999_ net882 net831 net825 net885 VPWR VGND sg13g2_a22oi_1
X_3128_ VGND VPWR _2721_ _2719_ _2686_ sg13g2_or2_1
X_3059_ _2654_ net978 net913 VPWR VGND sg13g2_nand2_1
XFILLER_42_128 VPWR VGND sg13g2_fill_1
XFILLER_13_1026 VPWR VGND sg13g2_fill_2
XFILLER_47_913 VPWR VGND sg13g2_decap_8
XFILLER_46_434 VPWR VGND sg13g2_fill_2
XFILLER_15_887 VPWR VGND sg13g2_decap_4
XFILLER_41_150 VPWR VGND sg13g2_decap_8
X_4100_ _0925_ _0927_ _0928_ VPWR VGND sg13g2_nor2_1
X_5080_ _1853_ VPWR _1865_ VGND _1861_ _1863_ sg13g2_o21ai_1
X_4031_ _0861_ _0854_ _0860_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_968 VPWR VGND sg13g2_decap_8
X_5982_ net882 _0230_ VPWR VGND sg13g2_buf_1
X_4933_ _1713_ _1726_ _1727_ VPWR VGND sg13g2_nor2_1
X_4864_ _1660_ DP_4.matrix\[5\] net1028 VPWR VGND sg13g2_nand2_1
XFILLER_32_161 VPWR VGND sg13g2_fill_1
X_3815_ _0637_ VPWR _0651_ VGND _0635_ _0638_ sg13g2_o21ai_1
X_4795_ VGND VPWR _1558_ _1564_ _1593_ _1566_ sg13g2_a21oi_1
X_3746_ _0587_ _0562_ _0589_ VPWR VGND sg13g2_xor2_1
X_6465_ net1122 VGND VPWR net220 mac2.sum_lvl2_ff\[15\] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_5416_ _2174_ net361 mac1.sum_lvl3_ff\[3\] VPWR VGND sg13g2_xnor2_1
X_3677_ _0521_ _0518_ _0522_ VPWR VGND sg13g2_xor2_1
X_6396_ net1126 VGND VPWR _0133_ mac2.products_ff\[83\] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_5347_ mac1.sum_lvl2_ff\[23\] mac1.sum_lvl2_ff\[4\] _2120_ VPWR VGND sg13g2_and2_1
X_5278_ VGND VPWR _1995_ _2025_ _2058_ _2027_ sg13g2_a21oi_1
X_4229_ net827 net878 net830 _1048_ VPWR VGND net876 sg13g2_nand4_1
XFILLER_29_946 VPWR VGND sg13g2_decap_8
XFILLER_44_916 VPWR VGND sg13g2_decap_8
XFILLER_24_695 VPWR VGND sg13g2_fill_2
XFILLER_7_305 VPWR VGND sg13g2_fill_1
XFILLER_11_345 VPWR VGND sg13g2_fill_2
XFILLER_35_916 VPWR VGND sg13g2_decap_8
XFILLER_36_91 VPWR VGND sg13g2_fill_2
XFILLER_43_960 VPWR VGND sg13g2_decap_8
XFILLER_21_109 VPWR VGND sg13g2_fill_2
XFILLER_30_621 VPWR VGND sg13g2_fill_2
Xinput11 uio_in[2] net11 VPWR VGND sg13g2_buf_1
X_3600_ _0447_ net1014 net946 VPWR VGND sg13g2_nand2_1
X_4580_ _1385_ _1376_ _1383_ VPWR VGND sg13g2_xnor2_1
X_3531_ _0368_ VPWR _0380_ VGND _0376_ _0378_ sg13g2_o21ai_1
X_3462_ _0301_ VPWR _0313_ VGND _0309_ _0311_ sg13g2_o21ai_1
X_6250_ net1068 VGND VPWR net134 mac1.sum_lvl2_ff\[51\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_5201_ _1979_ _1981_ _1982_ _1983_ VPWR VGND sg13g2_nor3_1
X_3393_ _2978_ _2964_ _2977_ VPWR VGND sg13g2_xnor2_1
X_6181_ net1081 VGND VPWR _0260_ DP_4.matrix\[72\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_5132_ VGND VPWR _1912_ _1913_ _1916_ _1878_ sg13g2_a21oi_1
XFILLER_28_0 VPWR VGND sg13g2_fill_2
X_5063_ _1848_ net858 net800 VPWR VGND sg13g2_nand2_1
X_4014_ _0845_ _0814_ _0843_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_938 VPWR VGND sg13g2_decap_8
XFILLER_16_28 VPWR VGND sg13g2_fill_2
X_5965_ net938 _0205_ VPWR VGND sg13g2_buf_1
X_4916_ _1710_ _1683_ _1706_ VPWR VGND sg13g2_nand2_1
X_5896_ _2466_ _2572_ net772 _2573_ VPWR VGND sg13g2_nand3_1
XFILLER_21_610 VPWR VGND sg13g2_fill_1
XFILLER_34_993 VPWR VGND sg13g2_decap_8
X_4847_ _1643_ _1640_ _1644_ VPWR VGND sg13g2_xor2_1
X_4778_ net845 net842 net888 net1029 _1577_ VPWR VGND sg13g2_and4_1
X_6517_ net1052 VGND VPWR DP_1.Q_range.data_plus_4\[6\] DP_1.Q_range.out_data\[5\]
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
X_3729_ VGND VPWR _0510_ _0540_ _0573_ _0542_ sg13g2_a21oi_1
X_6448_ net1053 VGND VPWR DP_1.I_range.data_plus_4\[6\] DP_1.I_range.out_data\[5\]
+ clknet_leaf_8_clk sg13g2_dfrbpq_1
X_6379_ net1105 VGND VPWR _0143_ mac2.products_ff\[14\] clknet_leaf_33_clk sg13g2_dfrbpq_1
XFILLER_29_710 VPWR VGND sg13g2_fill_1
XFILLER_29_743 VPWR VGND sg13g2_fill_2
XFILLER_29_754 VPWR VGND sg13g2_fill_1
XFILLER_32_908 VPWR VGND sg13g2_decap_8
XFILLER_19_1021 VPWR VGND sg13g2_decap_8
XFILLER_40_952 VPWR VGND sg13g2_decap_8
Xfanout1120 net1121 net1120 VPWR VGND sg13g2_buf_8
XFILLER_47_562 VPWR VGND sg13g2_fill_2
X_5750_ _2445_ _2444_ net783 net780 net279 VPWR VGND sg13g2_a22oi_1
XFILLER_22_429 VPWR VGND sg13g2_fill_2
X_5681_ _2375_ VPWR _2381_ VGND _2376_ _2380_ sg13g2_o21ai_1
X_4701_ _1499_ _1498_ _1468_ _1502_ VPWR VGND sg13g2_a21o_1
XFILLER_30_473 VPWR VGND sg13g2_fill_1
XFILLER_31_996 VPWR VGND sg13g2_decap_8
X_4632_ _1432_ _1406_ _1435_ VPWR VGND sg13g2_xor2_1
X_4563_ net847 net901 net843 net899 _1369_ VPWR VGND sg13g2_and4_1
X_6302_ net1050 VGND VPWR net100 mac1.sum_lvl3_ff\[21\] clknet_leaf_66_clk sg13g2_dfrbpq_1
X_3514_ _0363_ net1012 net950 VPWR VGND sg13g2_nand2_1
X_4494_ VGND VPWR _1260_ _1265_ _1306_ _1278_ sg13g2_a21oi_1
X_3445_ _0296_ net1020 net949 VPWR VGND sg13g2_nand2_1
X_6233_ net1114 VGND VPWR net190 mac1.sum_lvl2_ff\[31\] clknet_leaf_47_clk sg13g2_dfrbpq_2
X_3376_ _2962_ _2957_ _2960_ VPWR VGND sg13g2_xnor2_1
X_6164_ net1087 VGND VPWR _0245_ DP_4.matrix\[1\] clknet_leaf_27_clk sg13g2_dfrbpq_2
X_6095_ net1072 VGND VPWR _0199_ DP_2.matrix\[3\] clknet_leaf_57_clk sg13g2_dfrbpq_1
X_5115_ net813 net807 net851 net1024 _1899_ VPWR VGND sg13g2_and4_1
XFILLER_27_27 VPWR VGND sg13g2_fill_2
X_5046_ VGND VPWR _1829_ _1830_ _1832_ _1812_ sg13g2_a21oi_1
XFILLER_26_713 VPWR VGND sg13g2_decap_8
XFILLER_25_256 VPWR VGND sg13g2_fill_2
X_5948_ net1004 _0180_ VPWR VGND sg13g2_buf_1
XFILLER_40_204 VPWR VGND sg13g2_fill_2
XFILLER_22_941 VPWR VGND sg13g2_decap_8
X_5879_ net956 net771 _2562_ VPWR VGND sg13g2_nor2_1
XFILLER_1_834 VPWR VGND sg13g2_fill_1
XFILLER_44_521 VPWR VGND sg13g2_fill_2
XFILLER_44_510 VPWR VGND sg13g2_fill_2
XFILLER_44_565 VPWR VGND sg13g2_fill_1
XFILLER_32_716 VPWR VGND sg13g2_fill_1
XFILLER_16_289 VPWR VGND sg13g2_fill_1
XFILLER_13_930 VPWR VGND sg13g2_decap_8
XFILLER_12_495 VPWR VGND sg13g2_fill_1
XFILLER_40_793 VPWR VGND sg13g2_fill_2
X_3230_ _2819_ _2820_ _2821_ VPWR VGND sg13g2_nor2_1
X_3161_ net981 net979 net907 net905 _2753_ VPWR VGND sg13g2_and4_1
XFILLER_39_348 VPWR VGND sg13g2_fill_1
XFILLER_39_359 VPWR VGND sg13g2_fill_1
X_3092_ _2686_ net975 net913 VPWR VGND sg13g2_nand2_1
XFILLER_47_370 VPWR VGND sg13g2_fill_1
XFILLER_35_576 VPWR VGND sg13g2_fill_2
X_5802_ VGND VPWR _2493_ _2494_ _2496_ _2495_ sg13g2_a21oi_1
X_3994_ _0825_ _0815_ _0823_ VPWR VGND sg13g2_xnor2_1
X_5733_ net1007 DP_1.matrix\[42\] net788 _2429_ VPWR VGND sg13g2_mux2_1
X_5664_ _2367_ mac1.total_sum\[10\] mac2.total_sum\[10\] VPWR VGND sg13g2_nand2_1
X_5595_ _2309_ _2307_ _2308_ _2314_ VPWR VGND sg13g2_a21o_2
X_4615_ net850 net846 net895 net894 _1418_ VPWR VGND sg13g2_and4_1
X_4546_ _1342_ _1355_ _1356_ VPWR VGND sg13g2_nor2_1
Xhold400 _0022_ VPWR VGND net440 sg13g2_dlygate4sd3_1
Xhold411 mac2.sum_lvl2_ff\[4\] VPWR VGND net451 sg13g2_dlygate4sd3_1
Xhold444 mac2.sum_lvl3_ff\[3\] VPWR VGND net484 sg13g2_dlygate4sd3_1
Xhold433 mac2.sum_lvl3_ff\[22\] VPWR VGND net473 sg13g2_dlygate4sd3_1
Xhold422 _0005_ VPWR VGND net462 sg13g2_dlygate4sd3_1
X_4477_ _1289_ net1026 net819 net871 net818 VPWR VGND sg13g2_a22oi_1
Xhold455 DP_1.matrix\[38\] VPWR VGND net495 sg13g2_dlygate4sd3_1
Xhold466 _2124_ VPWR VGND net506 sg13g2_dlygate4sd3_1
Xhold477 mac2.sum_lvl2_ff\[6\] VPWR VGND net517 sg13g2_dlygate4sd3_1
Xhold488 _2278_ VPWR VGND net528 sg13g2_dlygate4sd3_1
Xfanout913 net914 net913 VPWR VGND sg13g2_buf_8
Xfanout924 net333 net924 VPWR VGND sg13g2_buf_1
X_3428_ _0280_ net1015 net954 VPWR VGND sg13g2_nand2_1
X_6216_ net1111 VGND VPWR net77 mac1.sum_lvl2_ff\[11\] clknet_leaf_46_clk sg13g2_dfrbpq_1
Xhold499 _2302_ VPWR VGND net539 sg13g2_dlygate4sd3_1
Xfanout902 net427 net902 VPWR VGND sg13g2_buf_8
X_6147_ net1096 VGND VPWR net116 mac1.sum_lvl1_ff\[8\] clknet_leaf_53_clk sg13g2_dfrbpq_1
Xfanout935 net936 net935 VPWR VGND sg13g2_buf_8
Xfanout957 net959 net957 VPWR VGND sg13g2_buf_2
Xfanout968 net315 net968 VPWR VGND sg13g2_buf_8
Xfanout946 net948 net946 VPWR VGND sg13g2_buf_8
X_3359_ _2945_ _2931_ _2946_ VPWR VGND sg13g2_xor2_1
Xfanout979 net980 net979 VPWR VGND sg13g2_buf_1
XFILLER_46_819 VPWR VGND sg13g2_fill_1
X_6078_ net1049 VGND VPWR _0065_ mac1.products_ff\[137\] clknet_leaf_67_clk sg13g2_dfrbpq_1
X_5029_ _1815_ net860 net802 VPWR VGND sg13g2_nand2_1
XFILLER_38_370 VPWR VGND sg13g2_fill_1
XFILLER_41_513 VPWR VGND sg13g2_fill_1
XFILLER_10_922 VPWR VGND sg13g2_fill_2
XFILLER_21_281 VPWR VGND sg13g2_fill_1
XFILLER_10_966 VPWR VGND sg13g2_decap_8
XFILLER_49_624 VPWR VGND sg13g2_fill_2
XFILLER_23_1006 VPWR VGND sg13g2_decap_8
XFILLER_48_167 VPWR VGND sg13g2_fill_1
XFILLER_29_370 VPWR VGND sg13g2_fill_1
XFILLER_45_896 VPWR VGND sg13g2_decap_8
XFILLER_9_786 VPWR VGND sg13g2_fill_1
X_4400_ _1215_ _1185_ _1214_ VPWR VGND sg13g2_nand2_1
X_5380_ mac1.sum_lvl2_ff\[30\] mac1.sum_lvl2_ff\[11\] _2146_ VPWR VGND sg13g2_nor2_1
XFILLER_5_981 VPWR VGND sg13g2_decap_8
X_4331_ _1147_ _1100_ _1146_ VPWR VGND sg13g2_xnor2_1
X_4262_ net827 net876 net829 _1080_ VPWR VGND net875 sg13g2_nand4_1
X_6001_ net818 _0257_ VPWR VGND sg13g2_buf_1
X_3213_ _2803_ _2752_ _2804_ VPWR VGND sg13g2_xor2_1
X_4193_ _1014_ _1005_ _1012_ VPWR VGND sg13g2_xnor2_1
X_3144_ _2737_ _2717_ _2735_ _2736_ VPWR VGND sg13g2_and3_1
X_3075_ _2668_ _2669_ _2651_ _2670_ VPWR VGND sg13g2_nand3_1
XFILLER_36_852 VPWR VGND sg13g2_decap_8
XFILLER_39_1024 VPWR VGND sg13g2_decap_4
X_3977_ _0809_ _0807_ _0808_ VPWR VGND sg13g2_nand2_1
X_5716_ net1013 net998 net788 _2412_ VPWR VGND sg13g2_mux2_1
X_5647_ _2349_ _2352_ _2353_ _2354_ VPWR VGND sg13g2_nor3_1
X_5578_ _2300_ mac2.sum_lvl3_ff\[27\] mac2.sum_lvl3_ff\[7\] VPWR VGND sg13g2_nand2_1
Xhold230 DP_4.matrix\[80\] VPWR VGND net270 sg13g2_dlygate4sd3_1
XFILLER_46_1006 VPWR VGND sg13g2_decap_8
X_4529_ _1339_ _1312_ _1335_ VPWR VGND sg13g2_nand2_1
Xhold241 DP_2.matrix\[43\] VPWR VGND net281 sg13g2_dlygate4sd3_1
Xhold252 DP_2.matrix\[7\] VPWR VGND net292 sg13g2_dlygate4sd3_1
Xhold285 _2585_ VPWR VGND net325 sg13g2_dlygate4sd3_1
Xhold263 DP_1.matrix\[75\] VPWR VGND net303 sg13g2_dlygate4sd3_1
Xhold274 DP_1.matrix\[80\] VPWR VGND net314 sg13g2_dlygate4sd3_1
Xhold296 mac2.sum_lvl3_ff\[30\] VPWR VGND net336 sg13g2_dlygate4sd3_1
Xfanout776 _2482_ net776 VPWR VGND sg13g2_buf_1
Xfanout798 net799 net798 VPWR VGND sg13g2_buf_8
Xfanout787 _2472_ net787 VPWR VGND sg13g2_buf_8
XFILLER_27_852 VPWR VGND sg13g2_decap_8
XFILLER_42_877 VPWR VGND sg13g2_decap_8
XFILLER_2_973 VPWR VGND sg13g2_decap_8
XFILLER_39_8 VPWR VGND sg13g2_fill_1
XFILLER_7_1011 VPWR VGND sg13g2_decap_8
XFILLER_1_494 VPWR VGND sg13g2_fill_1
XFILLER_36_126 VPWR VGND sg13g2_fill_1
Xinput9 uio_in[0] net9 VPWR VGND sg13g2_buf_1
XFILLER_33_800 VPWR VGND sg13g2_fill_1
X_4880_ _1674_ _1662_ _1676_ VPWR VGND sg13g2_xor2_1
X_3900_ _0715_ _0705_ _0713_ _0733_ VPWR VGND sg13g2_a21o_1
XFILLER_32_332 VPWR VGND sg13g2_fill_1
X_3831_ _0665_ _0645_ _0078_ VPWR VGND sg13g2_xor2_1
XFILLER_33_877 VPWR VGND sg13g2_decap_8
X_3762_ _0604_ net947 net1037 VPWR VGND sg13g2_nand2_1
XFILLER_32_387 VPWR VGND sg13g2_fill_1
XFILLER_9_550 VPWR VGND sg13g2_fill_1
X_5501_ _2240_ mac2.sum_lvl2_ff\[25\] net517 VPWR VGND sg13g2_xnor2_1
X_6481_ net1126 VGND VPWR net179 mac2.sum_lvl2_ff\[34\] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_3693_ _0537_ _0515_ _0538_ VPWR VGND sg13g2_nor2b_1
X_5432_ _2186_ net419 mac1.sum_lvl3_ff\[7\] VPWR VGND sg13g2_nand2_1
X_5363_ _2125_ _2128_ net530 _2133_ VPWR VGND sg13g2_or3_1
X_4314_ _1128_ _1127_ _1097_ _1131_ VPWR VGND sg13g2_a21o_1
X_5294_ _2047_ _2072_ _2073_ VPWR VGND sg13g2_nor2_1
X_4245_ _1061_ _1035_ _1064_ VPWR VGND sg13g2_xor2_1
X_4176_ net831 net885 net825 net882 _0998_ VPWR VGND sg13g2_and4_1
X_3127_ _2720_ net913 net973 VPWR VGND sg13g2_nand2_1
X_3058_ _2653_ net979 net911 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_62_clk clknet_4_2_0_clk clknet_leaf_62_clk VPWR VGND sg13g2_buf_8
XFILLER_13_1005 VPWR VGND sg13g2_decap_8
XFILLER_19_649 VPWR VGND sg13g2_decap_4
XFILLER_47_969 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_53_clk clknet_4_8_0_clk clknet_leaf_53_clk VPWR VGND sg13g2_buf_8
XFILLER_30_869 VPWR VGND sg13g2_decap_8
Xclkbuf_4_6_0_clk clknet_0_clk clknet_4_6_0_clk VPWR VGND sg13g2_buf_8
XFILLER_10_582 VPWR VGND sg13g2_fill_2
XFILLER_29_1023 VPWR VGND sg13g2_decap_4
X_4030_ _0859_ _0855_ _0860_ VPWR VGND sg13g2_xor2_1
XFILLER_38_947 VPWR VGND sg13g2_decap_8
X_5981_ net884 _0229_ VPWR VGND sg13g2_buf_1
X_4932_ _1724_ _1714_ _1726_ VPWR VGND sg13g2_xor2_1
XFILLER_18_693 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_44_clk clknet_4_9_0_clk clknet_leaf_44_clk VPWR VGND sg13g2_buf_8
XFILLER_36_1027 VPWR VGND sg13g2_fill_2
X_4863_ _1659_ net1028 net838 net889 DP_4.matrix\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_33_685 VPWR VGND sg13g2_fill_1
X_3814_ VPWR _0650_ _0649_ VGND sg13g2_inv_1
X_4794_ _1592_ _1553_ _0148_ VPWR VGND sg13g2_xor2_1
X_3745_ _0562_ _0587_ _0588_ VPWR VGND sg13g2_nor2_1
X_6464_ net1122 VGND VPWR net43 mac2.sum_lvl2_ff\[14\] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_5415_ _2173_ net361 mac1.sum_lvl3_ff\[3\] VPWR VGND sg13g2_nand2_1
X_3676_ _0521_ _0495_ _0519_ VPWR VGND sg13g2_xnor2_1
X_6395_ net1127 VGND VPWR _0132_ mac2.products_ff\[82\] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_5346_ _2117_ VPWR _2119_ VGND _2116_ _2118_ sg13g2_o21ai_1
XFILLER_43_1009 VPWR VGND sg13g2_decap_8
X_5277_ VGND VPWR _1994_ _2025_ _2057_ _2027_ sg13g2_a21oi_1
X_4228_ net830 net827 net878 net876 _1047_ VPWR VGND sg13g2_and4_1
XFILLER_29_925 VPWR VGND sg13g2_decap_8
X_4159_ _0971_ _0984_ _0985_ VPWR VGND sg13g2_nor2_1
XFILLER_37_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_35_clk clknet_4_15_0_clk clknet_leaf_35_clk VPWR VGND sg13g2_buf_8
XFILLER_24_663 VPWR VGND sg13g2_decap_4
XFILLER_3_578 VPWR VGND sg13g2_fill_1
XFILLER_4_1014 VPWR VGND sg13g2_decap_8
XFILLER_19_435 VPWR VGND sg13g2_fill_1
XFILLER_34_438 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_26_clk clknet_4_7_0_clk clknet_leaf_26_clk VPWR VGND sg13g2_buf_8
XFILLER_42_482 VPWR VGND sg13g2_fill_2
XFILLER_14_162 VPWR VGND sg13g2_fill_2
XFILLER_42_493 VPWR VGND sg13g2_decap_4
Xinput12 uio_in[3] net12 VPWR VGND sg13g2_buf_1
X_3530_ _0368_ _0376_ _0378_ _0379_ VPWR VGND sg13g2_or3_1
X_3461_ _0301_ _0309_ _0311_ _0312_ VPWR VGND sg13g2_or3_1
X_5200_ _1982_ net851 net803 net854 net801 VPWR VGND sg13g2_a22oi_1
X_6180_ net1106 VGND VPWR _0259_ DP_4.matrix\[43\] clknet_leaf_32_clk sg13g2_dfrbpq_2
X_3392_ _2977_ _2974_ _2976_ VPWR VGND sg13g2_xnor2_1
X_5131_ _1912_ _1913_ _1878_ _1915_ VPWR VGND sg13g2_nand3_1
X_5062_ _1847_ net863 net798 VPWR VGND sg13g2_nand2_1
X_4013_ _0844_ _0814_ _0843_ VPWR VGND sg13g2_nand2_1
XFILLER_26_917 VPWR VGND sg13g2_decap_8
X_5964_ net942 _0204_ VPWR VGND sg13g2_buf_1
Xclkbuf_leaf_17_clk clknet_4_4_0_clk clknet_leaf_17_clk VPWR VGND sg13g2_buf_8
XFILLER_34_972 VPWR VGND sg13g2_decap_8
X_4915_ _1684_ _1707_ _1709_ VPWR VGND sg13g2_and2_1
X_5895_ _2572_ _2441_ _2465_ VPWR VGND sg13g2_nand2b_1
X_4846_ _1643_ _1598_ _1641_ VPWR VGND sg13g2_xnor2_1
X_4777_ _1576_ net842 net1029 VPWR VGND sg13g2_nand2_1
X_6516_ net1052 VGND VPWR net7 DP_1.Q_range.out_data\[4\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_10_1008 VPWR VGND sg13g2_decap_8
X_3728_ VGND VPWR _0509_ _0540_ _0572_ _0542_ sg13g2_a21oi_1
X_6447_ net1052 VGND VPWR net3 DP_1.I_range.out_data\[4\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_3659_ _0505_ _0480_ _0504_ VPWR VGND sg13g2_nand2_1
X_6378_ net1105 VGND VPWR _0142_ mac2.products_ff\[13\] clknet_leaf_33_clk sg13g2_dfrbpq_1
X_5329_ _2106_ _2103_ _2105_ VPWR VGND sg13g2_xnor2_1
XFILLER_43_224 VPWR VGND sg13g2_fill_2
XFILLER_43_202 VPWR VGND sg13g2_fill_1
XFILLER_19_1000 VPWR VGND sg13g2_decap_8
XFILLER_40_931 VPWR VGND sg13g2_decap_8
XFILLER_7_114 VPWR VGND sg13g2_fill_2
XFILLER_12_688 VPWR VGND sg13g2_decap_8
Xfanout1110 net1112 net1110 VPWR VGND sg13g2_buf_8
XFILLER_26_1015 VPWR VGND sg13g2_decap_8
Xfanout1121 net1129 net1121 VPWR VGND sg13g2_buf_8
XFILLER_16_994 VPWR VGND sg13g2_decap_8
X_5680_ net21 _2377_ _2380_ VPWR VGND sg13g2_xnor2_1
X_4700_ VGND VPWR _1498_ _1499_ _1501_ _1468_ sg13g2_a21oi_1
XFILLER_31_975 VPWR VGND sg13g2_decap_8
X_4631_ VGND VPWR _1430_ _1431_ _1434_ _1406_ sg13g2_a21oi_1
X_4562_ _1368_ net903 net841 VPWR VGND sg13g2_nand2_1
X_4493_ _1303_ _1292_ _1305_ VPWR VGND sg13g2_xor2_1
X_6301_ net1049 VGND VPWR net107 mac1.sum_lvl3_ff\[20\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3513_ _0362_ net1016 net949 VPWR VGND sg13g2_nand2_1
X_3444_ _0286_ VPWR _0295_ VGND _0278_ _0287_ sg13g2_o21ai_1
X_6232_ net1115 VGND VPWR net241 mac1.sum_lvl2_ff\[30\] clknet_leaf_48_clk sg13g2_dfrbpq_2
Xclkbuf_leaf_6_clk clknet_4_1_0_clk clknet_leaf_6_clk VPWR VGND sg13g2_buf_8
X_3375_ _2961_ _2960_ _2957_ VPWR VGND sg13g2_nand2b_1
X_6163_ net1087 VGND VPWR _0244_ DP_4.matrix\[0\] clknet_leaf_27_clk sg13g2_dfrbpq_2
X_6094_ net1076 VGND VPWR net394 DP_2.matrix\[2\] clknet_leaf_61_clk sg13g2_dfrbpq_2
X_5114_ _1898_ net804 net854 VPWR VGND sg13g2_nand2_1
X_5045_ _1829_ _1830_ _1812_ _1831_ VPWR VGND sg13g2_nand3_1
XFILLER_26_758 VPWR VGND sg13g2_decap_4
XFILLER_41_706 VPWR VGND sg13g2_fill_2
X_5947_ net270 _0171_ VPWR VGND sg13g2_buf_1
XFILLER_22_920 VPWR VGND sg13g2_decap_8
X_5878_ _0196_ net960 _2395_ VPWR VGND sg13g2_xnor2_1
XFILLER_22_997 VPWR VGND sg13g2_decap_8
X_4829_ VGND VPWR _1626_ _1627_ _1592_ _1552_ sg13g2_a21oi_2
XFILLER_5_618 VPWR VGND sg13g2_fill_1
XFILLER_40_772 VPWR VGND sg13g2_fill_2
XFILLER_8_434 VPWR VGND sg13g2_fill_2
XFILLER_8_456 VPWR VGND sg13g2_fill_2
XFILLER_3_172 VPWR VGND sg13g2_fill_1
XFILLER_3_183 VPWR VGND sg13g2_fill_1
X_3160_ _2752_ net978 net905 VPWR VGND sg13g2_nand2_1
Xhold1 mac2.sum_lvl1_ff\[12\] VPWR VGND net41 sg13g2_dlygate4sd3_1
X_3091_ _2685_ net975 net911 VPWR VGND sg13g2_nand2_1
X_5801_ net901 _2493_ _2495_ VPWR VGND sg13g2_nor2_1
X_5732_ _2411_ _2424_ _2426_ _2428_ VPWR VGND sg13g2_nor3_1
X_3993_ _0815_ _0823_ _0824_ VPWR VGND sg13g2_nor2_1
X_5663_ net18 _2363_ _2366_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_783 VPWR VGND sg13g2_fill_1
X_5594_ VPWR _2313_ _2312_ VGND sg13g2_inv_1
X_4614_ _1417_ net841 net898 VPWR VGND sg13g2_nand2_1
X_4545_ _1353_ _1343_ _1355_ VPWR VGND sg13g2_xor2_1
XFILLER_8_990 VPWR VGND sg13g2_decap_8
Xhold401 DP_1.matrix\[1\] VPWR VGND net441 sg13g2_dlygate4sd3_1
Xhold423 mac2.sum_lvl3_ff\[6\] VPWR VGND net463 sg13g2_dlygate4sd3_1
Xhold445 _2288_ VPWR VGND net485 sg13g2_dlygate4sd3_1
Xhold434 _2285_ VPWR VGND net474 sg13g2_dlygate4sd3_1
Xhold412 _2235_ VPWR VGND net452 sg13g2_dlygate4sd3_1
X_4476_ _1274_ _1268_ _1276_ _1288_ VPWR VGND sg13g2_a21o_1
Xhold467 _0011_ VPWR VGND net507 sg13g2_dlygate4sd3_1
Xhold478 _2240_ VPWR VGND net518 sg13g2_dlygate4sd3_1
Xhold456 DP_4.matrix\[40\] VPWR VGND net496 sg13g2_dlygate4sd3_1
X_3427_ _2993_ VPWR _0279_ VGND _2991_ _2994_ sg13g2_o21ai_1
Xhold489 mac1.sum_lvl2_ff\[7\] VPWR VGND net529 sg13g2_dlygate4sd3_1
Xfanout914 DP_2.matrix\[75\] net914 VPWR VGND sg13g2_buf_1
Xfanout925 net926 net925 VPWR VGND sg13g2_buf_8
X_6215_ net1112 VGND VPWR net113 mac1.sum_lvl2_ff\[10\] clknet_leaf_46_clk sg13g2_dfrbpq_1
Xfanout903 net332 net903 VPWR VGND sg13g2_buf_8
X_6146_ net1122 VGND VPWR _0233_ DP_3.matrix\[41\] clknet_leaf_35_clk sg13g2_dfrbpq_2
Xfanout958 net959 net958 VPWR VGND sg13g2_buf_8
Xfanout936 net488 net936 VPWR VGND sg13g2_buf_8
X_3358_ _2943_ _2918_ _2945_ VPWR VGND sg13g2_xor2_1
Xfanout947 net948 net947 VPWR VGND sg13g2_buf_1
Xfanout969 net970 net969 VPWR VGND sg13g2_buf_8
XFILLER_38_49 VPWR VGND sg13g2_fill_2
X_3289_ _2877_ _2874_ _2878_ VPWR VGND sg13g2_xor2_1
X_6077_ net1110 VGND VPWR _0187_ DP_1.matrix\[43\] clknet_leaf_45_clk sg13g2_dfrbpq_2
XFILLER_26_500 VPWR VGND sg13g2_fill_2
X_5028_ _1814_ net860 net800 VPWR VGND sg13g2_nand2_1
XFILLER_26_533 VPWR VGND sg13g2_fill_2
XFILLER_26_544 VPWR VGND sg13g2_fill_1
XFILLER_41_547 VPWR VGND sg13g2_decap_8
XFILLER_41_569 VPWR VGND sg13g2_decap_8
XFILLER_28_71 VPWR VGND sg13g2_fill_1
XFILLER_45_875 VPWR VGND sg13g2_decap_8
XFILLER_17_577 VPWR VGND sg13g2_fill_1
XFILLER_44_81 VPWR VGND sg13g2_fill_1
XFILLER_9_732 VPWR VGND sg13g2_fill_1
XFILLER_8_220 VPWR VGND sg13g2_fill_2
XFILLER_12_260 VPWR VGND sg13g2_fill_2
XFILLER_5_960 VPWR VGND sg13g2_decap_8
X_4330_ _1146_ _1137_ _1144_ VPWR VGND sg13g2_xnor2_1
X_4261_ net829 net827 net876 net875 _1079_ VPWR VGND sg13g2_and4_1
X_3212_ _2803_ net975 net907 VPWR VGND sg13g2_nand2_1
X_6000_ net819 _0256_ VPWR VGND sg13g2_buf_1
X_4192_ _1013_ _1005_ _1012_ VPWR VGND sg13g2_nand2_1
X_3143_ _2724_ VPWR _2736_ VGND _2732_ _2734_ sg13g2_o21ai_1
X_3074_ _2657_ VPWR _2669_ VGND _2665_ _2667_ sg13g2_o21ai_1
XFILLER_36_831 VPWR VGND sg13g2_decap_8
XFILLER_39_1003 VPWR VGND sg13g2_decap_8
X_3976_ _0805_ _0804_ _0806_ _0808_ VPWR VGND sg13g2_a21o_1
X_5715_ _2411_ _2410_ net783 net780 net327 VPWR VGND sg13g2_a22oi_1
X_5646_ VPWR VGND _2347_ _2346_ _2345_ mac1.total_sum\[5\] _2353_ mac2.total_sum\[5\]
+ sg13g2_a221oi_1
X_5577_ _2298_ net465 _0060_ VPWR VGND sg13g2_nor2b_1
Xhold220 mac1.products_ff\[14\] VPWR VGND net260 sg13g2_dlygate4sd3_1
X_4528_ _1313_ _1336_ _1338_ VPWR VGND sg13g2_and2_1
Xhold231 DP_2.matrix\[80\] VPWR VGND net271 sg13g2_dlygate4sd3_1
Xhold253 DP_3.matrix\[73\] VPWR VGND net293 sg13g2_dlygate4sd3_1
Xhold242 DP_4.matrix\[72\] VPWR VGND net282 sg13g2_dlygate4sd3_1
Xhold286 DP_3.matrix\[40\] VPWR VGND net326 sg13g2_dlygate4sd3_1
X_4459_ VGND VPWR _1272_ _1270_ _1228_ sg13g2_or2_1
Xhold275 DP_1.matrix\[78\] VPWR VGND net315 sg13g2_dlygate4sd3_1
Xhold264 DP_1.matrix\[79\] VPWR VGND net304 sg13g2_dlygate4sd3_1
Xhold297 _2311_ VPWR VGND net337 sg13g2_dlygate4sd3_1
Xfanout799 net297 net799 VPWR VGND sg13g2_buf_8
X_6129_ net1072 VGND VPWR net186 mac1.sum_lvl1_ff\[2\] clknet_leaf_56_clk sg13g2_dfrbpq_1
Xfanout788 net789 net788 VPWR VGND sg13g2_buf_8
Xfanout777 net779 net777 VPWR VGND sg13g2_buf_8
XFILLER_27_831 VPWR VGND sg13g2_decap_8
XFILLER_42_856 VPWR VGND sg13g2_decap_8
XFILLER_14_84 VPWR VGND sg13g2_fill_1
XFILLER_2_952 VPWR VGND sg13g2_decap_8
XFILLER_49_400 VPWR VGND sg13g2_fill_2
XFILLER_18_842 VPWR VGND sg13g2_fill_1
XFILLER_33_856 VPWR VGND sg13g2_decap_8
X_3830_ VGND VPWR _0666_ _0665_ _0645_ sg13g2_or2_1
X_3761_ _0603_ net944 net1038 VPWR VGND sg13g2_nand2_1
X_5500_ mac2.sum_lvl2_ff\[25\] mac2.sum_lvl2_ff\[6\] _2239_ VPWR VGND sg13g2_and2_1
X_6480_ net1127 VGND VPWR net243 mac2.sum_lvl2_ff\[33\] clknet_leaf_37_clk sg13g2_dfrbpq_2
X_3692_ _0537_ _0516_ _0536_ VPWR VGND sg13g2_xnor2_1
X_5431_ _2184_ net503 _0028_ VPWR VGND sg13g2_nor2b_1
X_5362_ net530 VPWR _2132_ VGND _2125_ _2128_ sg13g2_o21ai_1
X_4313_ VGND VPWR _1127_ _1128_ _1130_ _1097_ sg13g2_a21oi_1
X_5293_ _2072_ _2032_ _2070_ VPWR VGND sg13g2_xnor2_1
X_4244_ VGND VPWR _1059_ _1060_ _1063_ _1035_ sg13g2_a21oi_1
X_4175_ _0997_ net886 net823 VPWR VGND sg13g2_nand2_1
X_3126_ _2719_ net973 net911 VPWR VGND sg13g2_nand2_1
X_3057_ _2652_ net984 net909 VPWR VGND sg13g2_nand2_1
X_3959_ _0791_ _0784_ _0789_ _0790_ VPWR VGND sg13g2_and3_1
XFILLER_13_1028 VPWR VGND sg13g2_fill_1
X_5629_ mac1.total_sum\[2\] mac2.total_sum\[2\] _2340_ VPWR VGND sg13g2_and2_1
XFILLER_2_237 VPWR VGND sg13g2_fill_2
XFILLER_47_948 VPWR VGND sg13g2_decap_8
XFILLER_46_469 VPWR VGND sg13g2_fill_2
XFILLER_30_815 VPWR VGND sg13g2_fill_2
XFILLER_29_1002 VPWR VGND sg13g2_decap_8
XFILLER_49_241 VPWR VGND sg13g2_fill_1
XFILLER_2_54 VPWR VGND sg13g2_fill_2
XFILLER_38_926 VPWR VGND sg13g2_decap_8
X_5980_ net886 _0228_ VPWR VGND sg13g2_buf_1
X_4931_ _1724_ _1714_ _1725_ VPWR VGND sg13g2_nor2b_1
XFILLER_46_992 VPWR VGND sg13g2_decap_8
X_4862_ _1644_ _1639_ _1646_ _1658_ VPWR VGND sg13g2_a21o_1
XFILLER_36_1006 VPWR VGND sg13g2_decap_8
X_3813_ _0646_ _0648_ _0649_ VPWR VGND sg13g2_nor2_1
XFILLER_20_347 VPWR VGND sg13g2_fill_1
X_4793_ _1590_ _1591_ _1592_ VPWR VGND sg13g2_nor2b_1
X_3744_ _0587_ _0547_ _0585_ VPWR VGND sg13g2_xnor2_1
X_6463_ net1123 VGND VPWR net42 mac2.sum_lvl2_ff\[13\] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_3675_ VGND VPWR _0520_ _0519_ _0495_ sg13g2_or2_1
X_5414_ VGND VPWR _2169_ _2171_ _2172_ _2170_ sg13g2_a21oi_1
X_6394_ net1126 VGND VPWR _0131_ mac2.products_ff\[81\] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_5345_ net371 _2116_ _0009_ VPWR VGND sg13g2_xor2_1
X_5276_ _2054_ _2053_ _2056_ VPWR VGND sg13g2_xor2_1
XFILLER_29_904 VPWR VGND sg13g2_decap_8
X_4227_ _1046_ net824 net881 VPWR VGND sg13g2_nand2_1
X_4158_ _0982_ _0972_ _0984_ VPWR VGND sg13g2_xor2_1
X_3109_ VGND VPWR _2700_ _2701_ _2703_ _2683_ sg13g2_a21oi_1
X_4089_ _0917_ net1036 net932 net988 net929 VPWR VGND sg13g2_a22oi_1
XFILLER_37_970 VPWR VGND sg13g2_decap_8
XFILLER_36_480 VPWR VGND sg13g2_decap_4
XFILLER_36_491 VPWR VGND sg13g2_fill_2
XFILLER_11_347 VPWR VGND sg13g2_fill_1
XFILLER_23_185 VPWR VGND sg13g2_fill_1
XFILLER_28_992 VPWR VGND sg13g2_decap_8
XFILLER_36_93 VPWR VGND sg13g2_fill_1
XFILLER_43_995 VPWR VGND sg13g2_decap_8
XFILLER_42_461 VPWR VGND sg13g2_decap_4
XFILLER_14_141 VPWR VGND sg13g2_fill_2
XFILLER_14_196 VPWR VGND sg13g2_decap_4
Xinput13 uio_in[4] net13 VPWR VGND sg13g2_buf_1
X_3460_ VGND VPWR _0307_ _0308_ _0311_ _0302_ sg13g2_a21oi_1
X_3391_ _2975_ _2958_ _2976_ VPWR VGND sg13g2_xor2_1
X_5130_ _1914_ _1878_ _1912_ _1913_ VPWR VGND sg13g2_and3_1
XFILLER_42_1010 VPWR VGND sg13g2_decap_8
XFILLER_28_2 VPWR VGND sg13g2_fill_1
X_5061_ _1828_ _1818_ _1826_ _1846_ VPWR VGND sg13g2_a21o_1
X_4012_ _0842_ _0825_ _0843_ VPWR VGND sg13g2_xor2_1
X_5963_ net966 _0195_ VPWR VGND sg13g2_buf_1
X_4914_ _0142_ _1707_ _1708_ VPWR VGND sg13g2_xnor2_1
XFILLER_34_951 VPWR VGND sg13g2_decap_8
X_5894_ _2571_ net948 _2395_ _0202_ VPWR VGND sg13g2_mux2_1
X_4845_ VGND VPWR _1642_ _1641_ _1598_ sg13g2_or2_1
XFILLER_21_656 VPWR VGND sg13g2_fill_2
X_4776_ _1529_ VPWR _1575_ VGND _1527_ _1530_ sg13g2_o21ai_1
X_6515_ net1052 VGND VPWR net6 DP_1.Q_range.out_data\[3\] clknet_leaf_4_clk sg13g2_dfrbpq_2
X_3727_ _0569_ _0568_ _0571_ VPWR VGND sg13g2_xor2_1
X_6446_ net1053 VGND VPWR net2 DP_1.I_range.out_data\[3\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3658_ _0503_ _0491_ _0504_ VPWR VGND sg13g2_xor2_1
X_6377_ net1105 VGND VPWR _0141_ mac2.products_ff\[12\] clknet_leaf_33_clk sg13g2_dfrbpq_1
X_3589_ _0437_ _0435_ _0436_ VPWR VGND sg13g2_nand2_1
X_5328_ _2104_ _2088_ _2105_ VPWR VGND sg13g2_xor2_1
X_5259_ net856 net854 net796 net793 _2039_ VPWR VGND sg13g2_and4_1
Xclkbuf_4_5_0_clk clknet_0_clk clknet_4_5_0_clk VPWR VGND sg13g2_buf_8
XFILLER_16_428 VPWR VGND sg13g2_fill_1
XFILLER_25_984 VPWR VGND sg13g2_decap_8
XFILLER_40_910 VPWR VGND sg13g2_decap_8
XFILLER_40_987 VPWR VGND sg13g2_decap_8
XFILLER_8_649 VPWR VGND sg13g2_fill_2
XFILLER_11_166 VPWR VGND sg13g2_fill_2
Xfanout1122 net1124 net1122 VPWR VGND sg13g2_buf_8
Xfanout1111 net1112 net1111 VPWR VGND sg13g2_buf_8
Xfanout1100 net1101 net1100 VPWR VGND sg13g2_buf_8
XFILLER_47_564 VPWR VGND sg13g2_fill_1
XFILLER_47_81 VPWR VGND sg13g2_fill_2
XFILLER_47_586 VPWR VGND sg13g2_fill_2
XFILLER_16_973 VPWR VGND sg13g2_decap_8
XFILLER_31_954 VPWR VGND sg13g2_decap_8
X_4630_ _1430_ _1431_ _1406_ _1433_ VPWR VGND sg13g2_nand3_1
X_6300_ net1057 VGND VPWR net257 mac2.sum_lvl1_ff\[87\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_4561_ _1366_ _1367_ _0085_ VPWR VGND sg13g2_nor2_1
X_4492_ VGND VPWR _1304_ _1303_ _1292_ sg13g2_or2_1
X_3512_ _0343_ _0333_ _0341_ _0361_ VPWR VGND sg13g2_a21o_1
X_3443_ _0293_ _0273_ _0073_ VPWR VGND sg13g2_xor2_1
X_6231_ net1115 VGND VPWR net209 mac1.sum_lvl2_ff\[29\] clknet_leaf_48_clk sg13g2_dfrbpq_2
X_6162_ net1116 VGND VPWR net213 mac1.sum_lvl1_ff\[13\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_3374_ _2959_ _2934_ _2960_ VPWR VGND sg13g2_xor2_1
X_5113_ _1857_ VPWR _1897_ VGND _1855_ _1858_ sg13g2_o21ai_1
X_6093_ net1064 VGND VPWR _0101_ mac1.products_ff\[142\] clknet_leaf_65_clk sg13g2_dfrbpq_1
X_5044_ _1828_ _1827_ _1818_ _1830_ VPWR VGND sg13g2_a21o_1
XFILLER_27_29 VPWR VGND sg13g2_fill_1
XFILLER_38_586 VPWR VGND sg13g2_decap_8
X_5946_ net1022 _0170_ VPWR VGND sg13g2_buf_1
X_5877_ _2561_ VPWR _0179_ VGND _2605_ net773 sg13g2_o21ai_1
XFILLER_21_420 VPWR VGND sg13g2_fill_1
XFILLER_22_976 VPWR VGND sg13g2_decap_8
X_4828_ VGND VPWR _1549_ _1591_ _1626_ _1590_ sg13g2_a21oi_1
XFILLER_21_475 VPWR VGND sg13g2_decap_4
X_4759_ _1523_ VPWR _1558_ VGND _1520_ _1524_ sg13g2_o21ai_1
XFILLER_49_1027 VPWR VGND sg13g2_fill_2
X_6429_ net1084 VGND VPWR net114 mac2.sum_lvl1_ff\[36\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_1_825 VPWR VGND sg13g2_fill_1
XFILLER_44_578 VPWR VGND sg13g2_fill_1
XFILLER_9_936 VPWR VGND sg13g2_decap_4
XFILLER_13_998 VPWR VGND sg13g2_decap_8
XFILLER_32_1020 VPWR VGND sg13g2_decap_8
Xhold2 mac2.sum_lvl1_ff\[13\] VPWR VGND net42 sg13g2_dlygate4sd3_1
X_3090_ _2684_ net982 net909 VPWR VGND sg13g2_nand2_1
XFILLER_0_891 VPWR VGND sg13g2_decap_8
XFILLER_48_884 VPWR VGND sg13g2_decap_8
X_3992_ _0823_ _0816_ _0822_ VPWR VGND sg13g2_xnor2_1
XFILLER_35_578 VPWR VGND sg13g2_fill_1
X_5800_ _2494_ net786 net867 net777 net885 VPWR VGND sg13g2_a22oi_1
X_5731_ _2424_ _2426_ _2427_ VPWR VGND sg13g2_nor2_1
XFILLER_15_291 VPWR VGND sg13g2_decap_8
X_5662_ _2366_ _2365_ _2364_ VPWR VGND sg13g2_nand2b_1
X_5593_ net444 net336 _2312_ VPWR VGND sg13g2_xor2_1
X_4613_ _1396_ VPWR _1416_ VGND _1394_ _1397_ sg13g2_o21ai_1
X_4544_ _1353_ _1343_ _1354_ VPWR VGND sg13g2_nor2b_1
Xhold402 _2981_ VPWR VGND net442 sg13g2_dlygate4sd3_1
XFILLER_7_490 VPWR VGND sg13g2_fill_2
Xhold435 _0056_ VPWR VGND net475 sg13g2_dlygate4sd3_1
Xhold424 _2296_ VPWR VGND net464 sg13g2_dlygate4sd3_1
Xhold413 _0042_ VPWR VGND net453 sg13g2_dlygate4sd3_1
Xhold457 DP_4.matrix\[39\] VPWR VGND net497 sg13g2_dlygate4sd3_1
Xhold468 mac1.sum_lvl2_ff\[6\] VPWR VGND net508 sg13g2_dlygate4sd3_1
X_6214_ net1110 VGND VPWR net246 mac1.sum_lvl2_ff\[9\] clknet_leaf_45_clk sg13g2_dfrbpq_1
Xhold446 _0057_ VPWR VGND net486 sg13g2_dlygate4sd3_1
X_4475_ _0129_ _1286_ _1287_ VPWR VGND sg13g2_xnor2_1
X_3426_ VPWR _0278_ _0277_ VGND sg13g2_inv_1
Xfanout915 net916 net915 VPWR VGND sg13g2_buf_8
Xhold479 _2243_ VPWR VGND net519 sg13g2_dlygate4sd3_1
Xfanout904 DP_3.matrix\[0\] net904 VPWR VGND sg13g2_buf_1
Xfanout937 net938 net937 VPWR VGND sg13g2_buf_2
Xfanout926 DP_2.matrix\[43\] net926 VPWR VGND sg13g2_buf_1
X_3357_ _2918_ _2943_ _2944_ VPWR VGND sg13g2_nor2_1
Xfanout948 net411 net948 VPWR VGND sg13g2_buf_2
X_6145_ net1106 VGND VPWR _0232_ DP_3.matrix\[40\] clknet_leaf_32_clk sg13g2_dfrbpq_2
Xfanout959 net523 net959 VPWR VGND sg13g2_buf_8
X_6076_ net1111 VGND VPWR _0186_ DP_1.matrix\[42\] clknet_leaf_45_clk sg13g2_dfrbpq_2
X_3288_ _2877_ _2851_ _2875_ VPWR VGND sg13g2_xnor2_1
X_5027_ _1813_ net866 net798 VPWR VGND sg13g2_nand2_1
XFILLER_39_884 VPWR VGND sg13g2_decap_8
XFILLER_14_707 VPWR VGND sg13g2_fill_1
XFILLER_16_1015 VPWR VGND sg13g2_decap_8
X_5929_ net837 net770 _2593_ VPWR VGND sg13g2_nor2_1
XFILLER_40_592 VPWR VGND sg13g2_decap_4
X_4260_ _1078_ net824 net879 VPWR VGND sg13g2_nand2_1
X_3211_ _2802_ net976 net905 VPWR VGND sg13g2_nand2_1
X_4191_ _1010_ _1011_ _1012_ VPWR VGND sg13g2_nor2b_1
X_3142_ _2724_ _2732_ _2734_ _2735_ VPWR VGND sg13g2_or3_1
XFILLER_39_158 VPWR VGND sg13g2_fill_2
X_3073_ _2657_ _2665_ _2667_ _2668_ VPWR VGND sg13g2_or3_1
XFILLER_36_887 VPWR VGND sg13g2_decap_8
X_3975_ _0805_ _0806_ _0804_ _0807_ VPWR VGND sg13g2_nand3_1
X_5714_ net1009 DP_1.matrix\[41\] net788 _2410_ VPWR VGND sg13g2_mux2_1
X_5645_ _2352_ mac1.total_sum\[6\] mac2.total_sum\[6\] VPWR VGND sg13g2_xnor2_1
X_5576_ net464 VPWR _2299_ VGND _2293_ _2297_ sg13g2_o21ai_1
Xhold210 mac1.products_ff\[146\] VPWR VGND net250 sg13g2_dlygate4sd3_1
X_4527_ _0131_ _1336_ _1337_ VPWR VGND sg13g2_xnor2_1
Xhold232 DP_2.matrix\[73\] VPWR VGND net272 sg13g2_dlygate4sd3_1
Xhold221 mac2.products_ff\[147\] VPWR VGND net261 sg13g2_dlygate4sd3_1
Xhold243 _0089_ VPWR VGND net283 sg13g2_dlygate4sd3_1
XFILLER_49_27 VPWR VGND sg13g2_fill_2
Xhold287 DP_1.matrix\[77\] VPWR VGND net327 sg13g2_dlygate4sd3_1
Xhold265 mac2.sum_lvl2_ff\[2\] VPWR VGND net305 sg13g2_dlygate4sd3_1
Xhold254 _1738_ VPWR VGND net294 sg13g2_dlygate4sd3_1
Xhold276 DP_4.matrix\[0\] VPWR VGND net316 sg13g2_dlygate4sd3_1
X_4458_ _1271_ net877 net816 VPWR VGND sg13g2_nand2_1
X_3409_ VGND VPWR _2990_ _2985_ _2983_ sg13g2_or2_1
Xhold298 _2318_ VPWR VGND net338 sg13g2_dlygate4sd3_1
Xfanout767 _2479_ net767 VPWR VGND sg13g2_buf_8
X_6128_ net1088 VGND VPWR _0221_ DP_3.matrix\[1\] clknet_leaf_28_clk sg13g2_dfrbpq_2
X_4389_ _1158_ VPWR _1204_ VGND _1156_ _1159_ sg13g2_o21ai_1
Xfanout778 net779 net778 VPWR VGND sg13g2_buf_8
Xfanout789 _2400_ net789 VPWR VGND sg13g2_buf_8
X_6059_ net1105 VGND VPWR _0170_ DP_4.matrix\[44\] clknet_leaf_34_clk sg13g2_dfrbpq_2
XFILLER_18_309 VPWR VGND sg13g2_decap_8
XFILLER_38_180 VPWR VGND sg13g2_fill_1
XFILLER_27_887 VPWR VGND sg13g2_decap_8
XFILLER_42_835 VPWR VGND sg13g2_decap_8
XFILLER_41_334 VPWR VGND sg13g2_fill_2
XFILLER_2_931 VPWR VGND sg13g2_decap_8
XFILLER_33_835 VPWR VGND sg13g2_decap_8
XFILLER_13_570 VPWR VGND sg13g2_decap_8
X_3760_ _0602_ DP_1.matrix\[6\] DP_2.matrix\[8\] VPWR VGND sg13g2_nand2_1
X_5430_ net502 VPWR _2185_ VGND _2179_ _2183_ sg13g2_o21ai_1
X_3691_ _0536_ _0525_ _0535_ VPWR VGND sg13g2_xnor2_1
X_5361_ net529 mac1.sum_lvl2_ff\[26\] _2131_ VPWR VGND sg13g2_xor2_1
X_5292_ _2032_ _2070_ _2071_ VPWR VGND sg13g2_nor2_1
X_4312_ _1127_ _1128_ _1097_ _1129_ VPWR VGND sg13g2_nand3_1
X_4243_ _1059_ _1060_ _1035_ _1062_ VPWR VGND sg13g2_nand3_1
X_4174_ _0995_ net401 _0080_ VPWR VGND sg13g2_nor2_1
X_3125_ _2718_ net979 net909 VPWR VGND sg13g2_nand2_1
X_3056_ _2642_ VPWR _2651_ VGND _2634_ _2643_ sg13g2_o21ai_1
XFILLER_24_857 VPWR VGND sg13g2_decap_4
X_3958_ _0785_ VPWR _0790_ VGND _0786_ _0788_ sg13g2_o21ai_1
X_3889_ _0722_ _0694_ _0723_ VPWR VGND sg13g2_nor2b_1
X_5628_ _2336_ VPWR _2339_ VGND _2335_ _2337_ sg13g2_o21ai_1
X_5559_ net474 _2283_ _0056_ VPWR VGND sg13g2_xor2_1
XFILLER_47_927 VPWR VGND sg13g2_decap_8
XFILLER_41_131 VPWR VGND sg13g2_fill_2
XFILLER_41_197 VPWR VGND sg13g2_fill_1
XFILLER_38_905 VPWR VGND sg13g2_decap_8
XFILLER_37_404 VPWR VGND sg13g2_decap_4
XFILLER_46_971 VPWR VGND sg13g2_decap_8
XFILLER_18_662 VPWR VGND sg13g2_fill_2
X_4930_ _1724_ _1699_ _1723_ VPWR VGND sg13g2_xnor2_1
X_4861_ _0140_ _1656_ _1657_ VPWR VGND sg13g2_xnor2_1
X_3812_ net1003 net1001 net933 net932 _0648_ VPWR VGND sg13g2_and4_1
XFILLER_32_175 VPWR VGND sg13g2_fill_1
X_4792_ _1591_ _1554_ _1589_ VPWR VGND sg13g2_nand2_1
X_3743_ _0547_ _0585_ _0586_ VPWR VGND sg13g2_nor2_1
X_6462_ net1122 VGND VPWR net41 mac2.sum_lvl2_ff\[12\] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_3674_ _0519_ net953 net1037 VPWR VGND sg13g2_nand2_1
X_6393_ net1126 VGND VPWR _0130_ mac2.products_ff\[80\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_5413_ net455 _2169_ _0024_ VPWR VGND sg13g2_xor2_1
X_5344_ _2118_ mac1.sum_lvl2_ff\[22\] net370 VPWR VGND sg13g2_xnor2_1
X_5275_ _2053_ _2054_ _2055_ VPWR VGND sg13g2_nor2_1
X_4226_ _1025_ VPWR _1045_ VGND _1023_ _1026_ sg13g2_o21ai_1
X_4157_ _0982_ _0972_ _0983_ VPWR VGND sg13g2_nor2b_1
X_3108_ _2700_ _2701_ _2683_ _2702_ VPWR VGND sg13g2_nand3_1
X_4088_ _0902_ _0897_ _0904_ _0916_ VPWR VGND sg13g2_a21o_1
X_3039_ _2621_ VPWR _2635_ VGND _2619_ _2622_ sg13g2_o21ai_1
XFILLER_7_319 VPWR VGND sg13g2_fill_1
XFILLER_11_75 VPWR VGND sg13g2_fill_2
XFILLER_47_713 VPWR VGND sg13g2_fill_2
XFILLER_46_223 VPWR VGND sg13g2_fill_1
XFILLER_28_971 VPWR VGND sg13g2_decap_8
XFILLER_43_974 VPWR VGND sg13g2_decap_8
XFILLER_42_484 VPWR VGND sg13g2_fill_1
Xinput14 uio_in[5] net14 VPWR VGND sg13g2_buf_1
XFILLER_11_871 VPWR VGND sg13g2_fill_2
XFILLER_7_853 VPWR VGND sg13g2_fill_2
XFILLER_6_363 VPWR VGND sg13g2_fill_2
X_3390_ _2975_ net965 net1030 VPWR VGND sg13g2_nand2_1
X_5060_ _1845_ _1840_ _1843_ VPWR VGND sg13g2_xnor2_1
X_4011_ _0842_ _0826_ _0840_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_735 VPWR VGND sg13g2_fill_2
X_5962_ net968 _0194_ VPWR VGND sg13g2_buf_1
XFILLER_19_993 VPWR VGND sg13g2_decap_8
XFILLER_46_790 VPWR VGND sg13g2_fill_2
X_4913_ VGND VPWR _1684_ _1687_ _1708_ _1683_ sg13g2_a21oi_1
XFILLER_18_481 VPWR VGND sg13g2_fill_1
XFILLER_34_930 VPWR VGND sg13g2_decap_8
X_5893_ _2571_ _2462_ _2464_ VPWR VGND sg13g2_xnor2_1
X_4844_ _1641_ net893 net834 VPWR VGND sg13g2_nand2_2
X_4775_ _1574_ _1569_ _1573_ VPWR VGND sg13g2_xnor2_1
X_6514_ net1053 VGND VPWR net5 DP_1.Q_range.out_data\[2\] clknet_leaf_9_clk sg13g2_dfrbpq_2
X_3726_ _0568_ _0569_ _0570_ VPWR VGND sg13g2_nor2_1
X_6445_ net1053 VGND VPWR net1 DP_1.I_range.out_data\[2\] clknet_leaf_9_clk sg13g2_dfrbpq_2
X_3657_ _0501_ _0492_ _0503_ VPWR VGND sg13g2_xor2_1
X_3588_ _0433_ _0432_ _0434_ _0436_ VPWR VGND sg13g2_a21o_1
X_6376_ net1104 VGND VPWR _0140_ mac2.products_ff\[11\] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_5327_ _2104_ net852 net1021 VPWR VGND sg13g2_nand2_1
X_5258_ _2038_ net854 net792 VPWR VGND sg13g2_nand2_1
X_5189_ VGND VPWR _1971_ _1969_ _1932_ sg13g2_or2_1
X_4209_ _1027_ _1028_ _1022_ _1029_ VPWR VGND sg13g2_nand3_1
XFILLER_17_908 VPWR VGND sg13g2_decap_8
XFILLER_44_749 VPWR VGND sg13g2_fill_2
XFILLER_44_738 VPWR VGND sg13g2_fill_1
XFILLER_25_963 VPWR VGND sg13g2_decap_8
XFILLER_8_628 VPWR VGND sg13g2_fill_1
XFILLER_12_679 VPWR VGND sg13g2_decap_4
XFILLER_40_966 VPWR VGND sg13g2_decap_8
XFILLER_7_116 VPWR VGND sg13g2_fill_1
Xfanout1112 net1118 net1112 VPWR VGND sg13g2_buf_8
Xfanout1101 net1107 net1101 VPWR VGND sg13g2_buf_8
Xfanout1123 net1124 net1123 VPWR VGND sg13g2_buf_2
XFILLER_47_510 VPWR VGND sg13g2_fill_2
XFILLER_19_267 VPWR VGND sg13g2_fill_2
XFILLER_16_952 VPWR VGND sg13g2_decap_8
XFILLER_15_473 VPWR VGND sg13g2_fill_2
XFILLER_31_933 VPWR VGND sg13g2_decap_8
X_4560_ _1367_ net843 net903 net901 net847 VPWR VGND sg13g2_a22oi_1
X_4491_ _1301_ _1293_ _1303_ VPWR VGND sg13g2_xor2_1
X_3511_ _0360_ _0355_ _0358_ VPWR VGND sg13g2_xnor2_1
XFILLER_6_182 VPWR VGND sg13g2_fill_2
X_3442_ VGND VPWR _0294_ _0293_ _0273_ sg13g2_or2_1
X_6230_ net1113 VGND VPWR net135 mac1.sum_lvl2_ff\[28\] clknet_leaf_49_clk sg13g2_dfrbpq_2
X_6161_ net1087 VGND VPWR _0243_ DP_3.matrix\[79\] clknet_leaf_24_clk sg13g2_dfrbpq_1
X_3373_ _2959_ net908 net1034 VPWR VGND sg13g2_nand2_1
X_5112_ _1896_ _1891_ _1895_ VPWR VGND sg13g2_xnor2_1
X_6092_ net1075 VGND VPWR _0197_ DP_2.matrix\[1\] clknet_leaf_61_clk sg13g2_dfrbpq_1
XFILLER_26_0 VPWR VGND sg13g2_fill_1
X_5043_ _1827_ _1828_ _1818_ _1829_ VPWR VGND sg13g2_nand3_1
X_5945_ net1024 _0168_ VPWR VGND sg13g2_buf_1
XFILLER_41_708 VPWR VGND sg13g2_fill_1
XFILLER_41_719 VPWR VGND sg13g2_fill_2
X_5876_ _2432_ _2560_ net773 _2561_ VPWR VGND sg13g2_nand3_1
XFILLER_22_955 VPWR VGND sg13g2_decap_8
X_4827_ _1625_ _1624_ _1623_ VPWR VGND sg13g2_nand2b_1
X_4758_ _1511_ _1514_ _1557_ VPWR VGND sg13g2_nor2_1
XFILLER_49_1006 VPWR VGND sg13g2_decap_8
X_3709_ _0553_ net1008 net945 VPWR VGND sg13g2_nand2_1
X_4689_ _1490_ _1483_ _1488_ _1489_ VPWR VGND sg13g2_and3_1
X_6428_ net1122 VGND VPWR net47 mac2.sum_lvl1_ff\[15\] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_6359_ net1044 VGND VPWR net350 mac1.total_sum\[10\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_29_554 VPWR VGND sg13g2_fill_1
XFILLER_1_1008 VPWR VGND sg13g2_decap_8
XFILLER_13_944 VPWR VGND sg13g2_decap_4
XFILLER_31_218 VPWR VGND sg13g2_fill_2
XFILLER_8_458 VPWR VGND sg13g2_fill_1
Xhold3 mac2.sum_lvl1_ff\[14\] VPWR VGND net43 sg13g2_dlygate4sd3_1
X_3991_ _0822_ _0817_ _0820_ VPWR VGND sg13g2_xnor2_1
X_5730_ _2426_ _2425_ net783 net780 net974 VPWR VGND sg13g2_a22oi_1
XFILLER_15_270 VPWR VGND sg13g2_decap_4
X_5661_ VGND VPWR _2365_ mac2.total_sum\[9\] mac1.total_sum\[9\] sg13g2_or2_1
X_5592_ _2311_ net336 mac2.sum_lvl3_ff\[10\] VPWR VGND sg13g2_nand2_1
Xclkbuf_4_4_0_clk clknet_0_clk clknet_4_4_0_clk VPWR VGND sg13g2_buf_8
X_4612_ _1413_ _1410_ _1415_ VPWR VGND sg13g2_xor2_1
X_4543_ _1353_ _1328_ _1352_ VPWR VGND sg13g2_xnor2_1
Xhold414 mac1.sum_lvl3_ff\[2\] VPWR VGND net454 sg13g2_dlygate4sd3_1
Xhold403 DP_1.I_range.out_data\[3\] VPWR VGND net443 sg13g2_dlygate4sd3_1
Xhold425 _2299_ VPWR VGND net465 sg13g2_dlygate4sd3_1
Xhold436 DP_3.matrix\[2\] VPWR VGND net476 sg13g2_dlygate4sd3_1
Xhold458 DP_1.matrix\[39\] VPWR VGND net498 sg13g2_dlygate4sd3_1
X_6213_ net1109 VGND VPWR net50 mac1.sum_lvl2_ff\[8\] clknet_leaf_52_clk sg13g2_dfrbpq_1
Xhold469 _2126_ VPWR VGND net509 sg13g2_dlygate4sd3_1
Xhold447 DP_1.matrix\[40\] VPWR VGND net487 sg13g2_dlygate4sd3_1
X_4474_ _1252_ _1257_ _1287_ VPWR VGND sg13g2_nor2_1
X_3425_ _0274_ _0276_ _0277_ VPWR VGND sg13g2_nor2_1
Xfanout916 net413 net916 VPWR VGND sg13g2_buf_1
Xfanout905 net906 net905 VPWR VGND sg13g2_buf_8
Xfanout938 net939 net938 VPWR VGND sg13g2_buf_1
X_6144_ net1096 VGND VPWR net88 mac1.sum_lvl1_ff\[7\] clknet_leaf_53_clk sg13g2_dfrbpq_1
Xfanout927 net928 net927 VPWR VGND sg13g2_buf_8
X_3356_ _2943_ _2904_ _2941_ VPWR VGND sg13g2_xnor2_1
Xfanout949 net472 net949 VPWR VGND sg13g2_buf_8
X_6075_ net1041 VGND VPWR _0064_ mac1.products_ff\[136\] clknet_leaf_67_clk sg13g2_dfrbpq_1
X_3287_ VGND VPWR _2876_ _2875_ _2851_ sg13g2_or2_1
X_5026_ _1795_ VPWR _1812_ VGND _1786_ _1796_ sg13g2_o21ai_1
XFILLER_39_863 VPWR VGND sg13g2_decap_8
XFILLER_41_527 VPWR VGND sg13g2_decap_8
X_5928_ VGND VPWR net769 _2592_ _0247_ _2591_ sg13g2_a21oi_1
X_5859_ net1018 net771 _2550_ VPWR VGND sg13g2_nor2_1
XFILLER_5_428 VPWR VGND sg13g2_fill_1
XFILLER_0_166 VPWR VGND sg13g2_fill_2
XFILLER_32_549 VPWR VGND sg13g2_fill_1
XFILLER_8_222 VPWR VGND sg13g2_fill_1
XFILLER_12_295 VPWR VGND sg13g2_fill_2
XFILLER_5_995 VPWR VGND sg13g2_decap_8
X_3210_ _2801_ net981 net1030 VPWR VGND sg13g2_nand2_1
X_4190_ _1006_ VPWR _1011_ VGND _1007_ _1009_ sg13g2_o21ai_1
X_3141_ VGND VPWR _2730_ _2731_ _2734_ _2725_ sg13g2_a21oi_1
XFILLER_48_671 VPWR VGND sg13g2_fill_1
X_3072_ VGND VPWR _2663_ _2664_ _2667_ _2658_ sg13g2_a21oi_1
XFILLER_47_181 VPWR VGND sg13g2_fill_1
XFILLER_36_866 VPWR VGND sg13g2_decap_8
X_3974_ _0758_ VPWR _0806_ VGND _0697_ _0759_ sg13g2_o21ai_1
X_5713_ _2409_ _2408_ net783 net780 net966 VPWR VGND sg13g2_a22oi_1
X_5644_ mac1.total_sum\[6\] mac2.total_sum\[6\] _2351_ VPWR VGND sg13g2_and2_1
Xhold211 mac1.products_ff\[73\] VPWR VGND net251 sg13g2_dlygate4sd3_1
X_5575_ _2293_ net464 _2297_ _2298_ VPWR VGND sg13g2_nor3_1
Xhold200 mac2.products_ff\[4\] VPWR VGND net240 sg13g2_dlygate4sd3_1
X_4526_ VGND VPWR _1313_ _1316_ _1337_ _1312_ sg13g2_a21oi_1
Xhold222 mac1.products_ff\[139\] VPWR VGND net262 sg13g2_dlygate4sd3_1
Xhold233 DP_1.matrix\[72\] VPWR VGND net273 sg13g2_dlygate4sd3_1
Xhold244 mac2.sum_lvl2_ff\[19\] VPWR VGND net284 sg13g2_dlygate4sd3_1
Xhold277 DP_3.matrix\[80\] VPWR VGND net317 sg13g2_dlygate4sd3_1
X_4457_ _1270_ net877 net815 VPWR VGND sg13g2_nand2_1
Xhold266 _2229_ VPWR VGND net306 sg13g2_dlygate4sd3_1
Xhold255 _0090_ VPWR VGND net295 sg13g2_dlygate4sd3_1
XFILLER_49_39 VPWR VGND sg13g2_fill_2
X_3408_ _2989_ net1019 net952 VPWR VGND sg13g2_nand2_1
Xhold299 _0050_ VPWR VGND net339 sg13g2_dlygate4sd3_1
Xhold288 mac2.sum_lvl3_ff\[14\] VPWR VGND net328 sg13g2_dlygate4sd3_1
X_6127_ net1081 VGND VPWR _0220_ DP_3.matrix\[0\] clknet_leaf_28_clk sg13g2_dfrbpq_2
X_4388_ _1203_ _1198_ _1202_ VPWR VGND sg13g2_xnor2_1
X_3339_ _2925_ _2924_ _2927_ VPWR VGND sg13g2_xor2_1
Xfanout768 net769 net768 VPWR VGND sg13g2_buf_2
Xfanout779 _2471_ net779 VPWR VGND sg13g2_buf_2
X_6058_ net1101 VGND VPWR _0169_ DP_4.matrix\[8\] clknet_leaf_27_clk sg13g2_dfrbpq_2
XFILLER_27_800 VPWR VGND sg13g2_decap_4
XFILLER_45_129 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_65_clk clknet_4_3_0_clk clknet_leaf_65_clk VPWR VGND sg13g2_buf_8
X_5009_ VGND VPWR _1792_ _1793_ _1796_ _1787_ sg13g2_a21oi_1
XFILLER_39_682 VPWR VGND sg13g2_fill_1
XFILLER_27_866 VPWR VGND sg13g2_decap_8
XFILLER_22_560 VPWR VGND sg13g2_fill_1
XFILLER_6_704 VPWR VGND sg13g2_fill_2
XFILLER_49_402 VPWR VGND sg13g2_fill_1
XFILLER_7_1025 VPWR VGND sg13g2_decap_4
XFILLER_2_987 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_56_clk clknet_4_8_0_clk clknet_leaf_56_clk VPWR VGND sg13g2_buf_8
XFILLER_29_170 VPWR VGND sg13g2_decap_4
XFILLER_33_814 VPWR VGND sg13g2_decap_8
XFILLER_45_696 VPWR VGND sg13g2_fill_1
XFILLER_44_162 VPWR VGND sg13g2_decap_4
XFILLER_44_184 VPWR VGND sg13g2_fill_1
X_3690_ _0535_ _0526_ _0533_ VPWR VGND sg13g2_xnor2_1
X_5360_ _2130_ mac1.sum_lvl2_ff\[26\] mac1.sum_lvl2_ff\[7\] VPWR VGND sg13g2_nand2_1
X_5291_ _2070_ _2061_ _2069_ VPWR VGND sg13g2_xnor2_1
X_4311_ _1103_ VPWR _1128_ VGND _1124_ _1126_ sg13g2_o21ai_1
X_4242_ _1059_ _1060_ _1061_ VPWR VGND sg13g2_and2_1
X_4173_ _0996_ net825 net886 net885 net831 VPWR VGND sg13g2_a22oi_1
X_3124_ _2699_ _2689_ _2697_ _2717_ VPWR VGND sg13g2_a21o_1
X_3055_ _2649_ _2629_ _0068_ VPWR VGND sg13g2_xor2_1
Xclkbuf_leaf_47_clk clknet_4_11_0_clk clknet_leaf_47_clk VPWR VGND sg13g2_buf_8
XFILLER_23_302 VPWR VGND sg13g2_fill_2
XFILLER_35_151 VPWR VGND sg13g2_fill_2
X_3957_ _0785_ _0786_ _0788_ _0789_ VPWR VGND sg13g2_or3_1
XFILLER_32_880 VPWR VGND sg13g2_decap_8
X_3888_ _0722_ _0698_ _0721_ VPWR VGND sg13g2_xnor2_1
XFILLER_13_1019 VPWR VGND sg13g2_decap_8
XFILLER_31_390 VPWR VGND sg13g2_fill_1
X_5627_ net26 _2335_ _2338_ VPWR VGND sg13g2_xnor2_1
X_5558_ mac2.sum_lvl3_ff\[2\] net473 _2285_ VPWR VGND sg13g2_xor2_1
X_4509_ _1320_ net870 net814 VPWR VGND sg13g2_nand2_1
X_5489_ _2231_ mac2.sum_lvl2_ff\[22\] net353 VPWR VGND sg13g2_nand2_1
XFILLER_47_906 VPWR VGND sg13g2_decap_8
XFILLER_46_449 VPWR VGND sg13g2_fill_1
XFILLER_14_346 VPWR VGND sg13g2_fill_2
XFILLER_15_858 VPWR VGND sg13g2_fill_2
XFILLER_30_817 VPWR VGND sg13g2_fill_1
XFILLER_10_563 VPWR VGND sg13g2_fill_2
XFILLER_6_534 VPWR VGND sg13g2_fill_2
XFILLER_41_73 VPWR VGND sg13g2_fill_1
XFILLER_46_950 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_29_clk clknet_4_12_0_clk clknet_leaf_29_clk VPWR VGND sg13g2_buf_8
XFILLER_45_482 VPWR VGND sg13g2_fill_2
X_4860_ _1623_ _1628_ _1657_ VPWR VGND sg13g2_nor2_1
X_3811_ _0647_ net1001 net932 VPWR VGND sg13g2_nand2_1
X_4791_ _1554_ _1589_ _1590_ VPWR VGND sg13g2_nor2_1
XFILLER_13_390 VPWR VGND sg13g2_fill_1
X_3742_ _0585_ _0576_ _0584_ VPWR VGND sg13g2_xnor2_1
X_3673_ _0518_ DP_2.matrix\[5\] net1008 VPWR VGND sg13g2_nand2_1
X_6461_ net1119 VGND VPWR net56 mac2.sum_lvl2_ff\[11\] clknet_leaf_42_clk sg13g2_dfrbpq_1
X_5412_ net454 mac1.sum_lvl3_ff\[22\] _2171_ VPWR VGND sg13g2_xor2_1
X_6392_ net1125 VGND VPWR _0129_ mac2.products_ff\[79\] clknet_leaf_41_clk sg13g2_dfrbpq_1
X_5343_ _2117_ mac1.sum_lvl2_ff\[22\] net370 VPWR VGND sg13g2_nand2_1
X_5274_ VGND VPWR _2001_ _2021_ _2054_ _2023_ sg13g2_a21oi_1
X_4225_ _1042_ _1039_ _1044_ VPWR VGND sg13g2_xor2_1
X_4156_ _0982_ _0957_ _0981_ VPWR VGND sg13g2_xnor2_1
XFILLER_29_939 VPWR VGND sg13g2_decap_8
X_3107_ _2699_ _2698_ _2689_ _2701_ VPWR VGND sg13g2_a21o_1
XFILLER_44_909 VPWR VGND sg13g2_decap_8
X_4087_ _0118_ _0914_ _0915_ VPWR VGND sg13g2_xnor2_1
X_3038_ VPWR _2634_ _2633_ VGND sg13g2_inv_1
XFILLER_24_611 VPWR VGND sg13g2_fill_1
XFILLER_24_644 VPWR VGND sg13g2_fill_2
XFILLER_36_493 VPWR VGND sg13g2_fill_1
XFILLER_12_828 VPWR VGND sg13g2_fill_2
XFILLER_24_688 VPWR VGND sg13g2_decap_8
X_4989_ _1775_ _1776_ _1777_ VPWR VGND sg13g2_nor2b_2
XFILLER_4_1028 VPWR VGND sg13g2_fill_1
XFILLER_28_950 VPWR VGND sg13g2_decap_8
XFILLER_35_909 VPWR VGND sg13g2_decap_8
XFILLER_34_419 VPWR VGND sg13g2_fill_2
XFILLER_43_953 VPWR VGND sg13g2_decap_8
XFILLER_14_143 VPWR VGND sg13g2_fill_1
Xinput15 uio_in[6] net15 VPWR VGND sg13g2_buf_1
XFILLER_6_331 VPWR VGND sg13g2_fill_1
X_4010_ _0841_ _0826_ _0840_ VPWR VGND sg13g2_nand2_1
XFILLER_37_246 VPWR VGND sg13g2_fill_1
X_5961_ net971 _0193_ VPWR VGND sg13g2_buf_1
XFILLER_19_972 VPWR VGND sg13g2_decap_8
X_4912_ _1705_ _1706_ _1707_ VPWR VGND sg13g2_and2_1
XFILLER_45_290 VPWR VGND sg13g2_fill_1
X_5892_ _2570_ net949 _2395_ _0201_ VPWR VGND sg13g2_mux2_1
XFILLER_34_986 VPWR VGND sg13g2_decap_8
X_4843_ _1640_ net898 net1023 VPWR VGND sg13g2_nand2_1
XFILLER_33_485 VPWR VGND sg13g2_fill_1
X_4774_ _1573_ _1521_ _1570_ VPWR VGND sg13g2_xnor2_1
XFILLER_21_658 VPWR VGND sg13g2_fill_1
XFILLER_21_669 VPWR VGND sg13g2_fill_1
X_3725_ VGND VPWR _0516_ _0536_ _0569_ _0538_ sg13g2_a21oi_1
X_6513_ net1054 VGND VPWR net345 mac2.total_sum\[15\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_6444_ net1126 VGND VPWR net151 mac2.sum_lvl1_ff\[51\] clknet_leaf_36_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_9_clk clknet_4_3_0_clk clknet_leaf_9_clk VPWR VGND sg13g2_buf_8
X_3656_ _0502_ _0492_ _0501_ VPWR VGND sg13g2_nand2b_1
X_3587_ _0433_ _0434_ _0432_ _0435_ VPWR VGND sg13g2_nand3_1
X_6375_ net1104 VGND VPWR _0139_ mac2.products_ff\[10\] clknet_leaf_43_clk sg13g2_dfrbpq_1
X_5326_ _2091_ VPWR _2103_ VGND _2063_ _2089_ sg13g2_o21ai_1
X_5257_ _2037_ net858 net1021 VPWR VGND sg13g2_nand2_1
X_4208_ _1023_ VPWR _1028_ VGND _1024_ _1026_ sg13g2_o21ai_1
X_5188_ _1970_ net858 net795 VPWR VGND sg13g2_nand2_1
XFILLER_28_202 VPWR VGND sg13g2_fill_1
X_4139_ VGND VPWR _0942_ _0945_ _0966_ _0941_ sg13g2_a21oi_1
XFILLER_25_942 VPWR VGND sg13g2_decap_8
XFILLER_19_1014 VPWR VGND sg13g2_decap_8
XFILLER_36_290 VPWR VGND sg13g2_fill_2
XFILLER_40_945 VPWR VGND sg13g2_decap_8
XFILLER_11_168 VPWR VGND sg13g2_fill_1
XFILLER_4_868 VPWR VGND sg13g2_fill_1
Xfanout1113 net1117 net1113 VPWR VGND sg13g2_buf_8
Xfanout1102 net1104 net1102 VPWR VGND sg13g2_buf_8
Xfanout1124 net1129 net1124 VPWR VGND sg13g2_buf_1
XFILLER_19_213 VPWR VGND sg13g2_fill_2
XFILLER_47_83 VPWR VGND sg13g2_fill_1
XFILLER_31_912 VPWR VGND sg13g2_decap_8
XFILLER_15_496 VPWR VGND sg13g2_decap_4
XFILLER_31_989 VPWR VGND sg13g2_decap_8
X_3510_ _0359_ _0355_ _0358_ VPWR VGND sg13g2_nand2_1
X_4490_ _1301_ _1293_ _1302_ VPWR VGND sg13g2_nor2b_1
XFILLER_10_190 VPWR VGND sg13g2_fill_2
XFILLER_7_684 VPWR VGND sg13g2_fill_1
X_3441_ _0291_ _0290_ _0293_ VPWR VGND sg13g2_xor2_1
X_6160_ net1081 VGND VPWR _0242_ DP_3.matrix\[78\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_3372_ _2958_ net906 net1034 VPWR VGND sg13g2_nand2_1
X_5111_ _1895_ _1848_ _1893_ VPWR VGND sg13g2_xnor2_1
X_6091_ net1073 VGND VPWR _0196_ DP_2.matrix\[0\] clknet_leaf_61_clk sg13g2_dfrbpq_2
X_5042_ _1825_ _1824_ _1819_ _1828_ VPWR VGND sg13g2_a21o_1
XFILLER_19_0 VPWR VGND sg13g2_fill_1
XFILLER_26_706 VPWR VGND sg13g2_decap_8
XFILLER_19_791 VPWR VGND sg13g2_fill_1
X_5944_ net1026 _0167_ VPWR VGND sg13g2_buf_1
X_5875_ _2560_ _2409_ _2431_ VPWR VGND sg13g2_nand2b_1
XFILLER_22_934 VPWR VGND sg13g2_decap_8
XFILLER_34_783 VPWR VGND sg13g2_fill_2
XFILLER_40_219 VPWR VGND sg13g2_fill_2
X_4826_ _1588_ _1622_ _1586_ _1624_ VPWR VGND sg13g2_nand3_1
X_4757_ _1539_ VPWR _1556_ VGND _1518_ _1540_ sg13g2_o21ai_1
X_3708_ _0552_ net1012 net1032 VPWR VGND sg13g2_nand2_1
X_4688_ _1484_ VPWR _1489_ VGND _1485_ _1487_ sg13g2_o21ai_1
X_6427_ net1105 VGND VPWR net125 mac2.sum_lvl1_ff\[14\] clknet_leaf_33_clk sg13g2_dfrbpq_1
X_3639_ _0485_ net1012 net946 VPWR VGND sg13g2_nand2_1
X_6358_ net1044 VGND VPWR net360 mac1.total_sum\[9\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_5309_ _2087_ net854 net1021 VPWR VGND sg13g2_nand2_1
X_6289_ net1080 VGND VPWR net65 mac2.sum_lvl1_ff\[76\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_44_536 VPWR VGND sg13g2_fill_2
XFILLER_13_923 VPWR VGND sg13g2_decap_8
XFILLER_9_905 VPWR VGND sg13g2_decap_4
XFILLER_33_74 VPWR VGND sg13g2_fill_2
XFILLER_40_786 VPWR VGND sg13g2_decap_8
Xhold4 mac2.sum_lvl2_ff\[42\] VPWR VGND net44 sg13g2_dlygate4sd3_1
X_3990_ _0821_ _0820_ _0817_ VPWR VGND sg13g2_nand2b_1
XFILLER_16_783 VPWR VGND sg13g2_fill_2
X_5660_ mac1.total_sum\[9\] mac2.total_sum\[9\] _2364_ VPWR VGND sg13g2_and2_1
XFILLER_31_797 VPWR VGND sg13g2_fill_2
X_4611_ _1414_ _1413_ _1410_ VPWR VGND sg13g2_nand2b_1
X_5591_ _0063_ _2307_ _2310_ VPWR VGND sg13g2_xnor2_1
X_4542_ _1350_ _1349_ _1352_ VPWR VGND sg13g2_xor2_1
XFILLER_7_492 VPWR VGND sg13g2_fill_1
Xhold415 _2171_ VPWR VGND net455 sg13g2_dlygate4sd3_1
Xhold426 _0060_ VPWR VGND net466 sg13g2_dlygate4sd3_1
Xhold404 mac2.sum_lvl3_ff\[10\] VPWR VGND net444 sg13g2_dlygate4sd3_1
X_4473_ _1284_ _1285_ _1286_ VPWR VGND sg13g2_nor2_1
Xhold459 DP_2.matrix\[39\] VPWR VGND net499 sg13g2_dlygate4sd3_1
Xhold448 DP_2.matrix\[38\] VPWR VGND net488 sg13g2_dlygate4sd3_1
X_6212_ net1109 VGND VPWR net92 mac1.sum_lvl2_ff\[7\] clknet_leaf_53_clk sg13g2_dfrbpq_1
X_3424_ net1019 net1017 net952 net951 _0276_ VPWR VGND sg13g2_and4_1
Xhold437 mac1.sum_lvl3_ff\[14\] VPWR VGND net477 sg13g2_dlygate4sd3_1
Xfanout906 net298 net906 VPWR VGND sg13g2_buf_8
Xfanout939 net431 net939 VPWR VGND sg13g2_buf_2
Xfanout917 net919 net917 VPWR VGND sg13g2_buf_8
Xfanout928 net412 net928 VPWR VGND sg13g2_buf_2
X_3355_ _2904_ _2941_ _2942_ VPWR VGND sg13g2_nor2_1
X_6143_ net1124 VGND VPWR _0231_ DP_3.matrix\[39\] clknet_leaf_35_clk sg13g2_dfrbpq_2
X_3286_ _2875_ net914 net1034 VPWR VGND sg13g2_nand2_1
X_6074_ net1111 VGND VPWR _0185_ DP_1.matrix\[41\] clknet_leaf_49_clk sg13g2_dfrbpq_2
X_5025_ _1809_ _1808_ _1811_ VPWR VGND sg13g2_xor2_1
XFILLER_39_842 VPWR VGND sg13g2_decap_8
XFILLER_38_341 VPWR VGND sg13g2_fill_1
X_5927_ _2533_ _2524_ _2592_ VPWR VGND sg13g2_xor2_1
X_5858_ _0172_ net1019 _2395_ VPWR VGND sg13g2_xnor2_1
X_4809_ VGND VPWR net846 net888 _1607_ _1576_ sg13g2_a21oi_1
XFILLER_10_959 VPWR VGND sg13g2_decap_8
X_5789_ _2483_ DP_3.matrix\[77\] net775 VPWR VGND sg13g2_nand2_1
XFILLER_28_30 VPWR VGND sg13g2_fill_2
XFILLER_44_300 VPWR VGND sg13g2_fill_1
XFILLER_17_514 VPWR VGND sg13g2_decap_4
XFILLER_45_889 VPWR VGND sg13g2_decap_8
XFILLER_17_569 VPWR VGND sg13g2_fill_1
XFILLER_9_768 VPWR VGND sg13g2_fill_2
XFILLER_5_974 VPWR VGND sg13g2_decap_8
X_3140_ _2730_ _2731_ _2725_ _2733_ VPWR VGND sg13g2_nand3_1
X_3071_ _2663_ _2664_ _2658_ _2666_ VPWR VGND sg13g2_nand3_1
XFILLER_36_845 VPWR VGND sg13g2_decap_8
XFILLER_39_1017 VPWR VGND sg13g2_decap_8
XFILLER_39_1028 VPWR VGND sg13g2_fill_1
X_3973_ _0731_ VPWR _0805_ VGND _0801_ _0803_ sg13g2_o21ai_1
X_5712_ VGND VPWR _2605_ net791 _2408_ _2407_ sg13g2_a21oi_1
X_5643_ net30 _2348_ _2350_ VPWR VGND sg13g2_xnor2_1
X_5574_ VPWR VGND _2291_ _2290_ _2289_ mac2.sum_lvl3_ff\[25\] _2297_ net396 sg13g2_a221oi_1
X_4525_ _1334_ _1335_ _1336_ VPWR VGND sg13g2_and2_1
Xhold201 mac1.sum_lvl1_ff\[47\] VPWR VGND net241 sg13g2_dlygate4sd3_1
Xhold223 mac1.sum_lvl2_ff\[42\] VPWR VGND net263 sg13g2_dlygate4sd3_1
Xhold212 mac2.sum_lvl1_ff\[41\] VPWR VGND net252 sg13g2_dlygate4sd3_1
Xhold234 DP_3.matrix\[76\] VPWR VGND net274 sg13g2_dlygate4sd3_1
Xhold278 DP_1.matrix\[76\] VPWR VGND net318 sg13g2_dlygate4sd3_1
Xhold256 DP_1.matrix\[73\] VPWR VGND net296 sg13g2_dlygate4sd3_1
Xhold267 _0040_ VPWR VGND net307 sg13g2_dlygate4sd3_1
Xhold245 _0039_ VPWR VGND net285 sg13g2_dlygate4sd3_1
X_4456_ _1269_ net881 net1022 VPWR VGND sg13g2_nand2_1
XFILLER_49_29 VPWR VGND sg13g2_fill_1
X_3407_ _2987_ _2980_ _0071_ VPWR VGND sg13g2_xor2_1
Xhold289 _2332_ VPWR VGND net329 sg13g2_dlygate4sd3_1
X_4387_ _1202_ _1150_ _1199_ VPWR VGND sg13g2_xnor2_1
X_6126_ net1070 VGND VPWR net182 mac1.sum_lvl1_ff\[1\] clknet_leaf_62_clk sg13g2_dfrbpq_1
X_3338_ _2924_ _2925_ _2926_ VPWR VGND sg13g2_nor2_1
Xfanout769 net770 net769 VPWR VGND sg13g2_buf_2
X_6057_ net1062 VGND VPWR _0168_ DP_3.matrix\[80\] clknet_leaf_24_clk sg13g2_dfrbpq_1
X_3269_ _2857_ _2848_ _2859_ VPWR VGND sg13g2_xor2_1
X_5008_ _1792_ _1793_ _1787_ _1795_ VPWR VGND sg13g2_nand3_1
XFILLER_41_336 VPWR VGND sg13g2_fill_1
XFILLER_30_31 VPWR VGND sg13g2_fill_2
XFILLER_2_900 VPWR VGND sg13g2_fill_1
XFILLER_2_966 VPWR VGND sg13g2_decap_8
XFILLER_7_1004 VPWR VGND sg13g2_decap_8
XFILLER_49_425 VPWR VGND sg13g2_fill_1
Xclkbuf_4_3_0_clk clknet_0_clk clknet_4_3_0_clk VPWR VGND sg13g2_buf_8
XFILLER_18_878 VPWR VGND sg13g2_decap_4
XFILLER_9_598 VPWR VGND sg13g2_decap_4
X_5290_ _2069_ _2033_ _2067_ VPWR VGND sg13g2_xnor2_1
X_4310_ _1103_ _1124_ _1126_ _1127_ VPWR VGND sg13g2_or3_1
X_4241_ _1058_ _1057_ _1019_ _1060_ VPWR VGND sg13g2_a21o_1
X_4172_ _0995_ net885 net825 _0079_ VPWR VGND sg13g2_and3_2
X_3123_ _2716_ _2711_ _2714_ VPWR VGND sg13g2_xnor2_1
XFILLER_49_992 VPWR VGND sg13g2_decap_8
X_3054_ VGND VPWR _2650_ _2649_ _2629_ sg13g2_or2_1
XFILLER_35_130 VPWR VGND sg13g2_decap_4
XFILLER_36_664 VPWR VGND sg13g2_fill_2
XFILLER_35_163 VPWR VGND sg13g2_fill_2
XFILLER_35_185 VPWR VGND sg13g2_fill_2
X_3956_ _0788_ net1035 net942 net986 net937 VPWR VGND sg13g2_a22oi_1
X_5626_ mac2.total_sum\[1\] mac1.total_sum\[1\] _2338_ VPWR VGND sg13g2_xor2_1
X_3887_ _0721_ _0718_ _0720_ VPWR VGND sg13g2_nand2_1
X_5557_ net473 mac2.sum_lvl3_ff\[2\] _2284_ VPWR VGND sg13g2_and2_1
X_4508_ _1319_ net877 net1022 VPWR VGND sg13g2_nand2_1
X_5488_ VGND VPWR _2227_ net306 _2230_ _2228_ sg13g2_a21oi_1
X_4439_ _1217_ _1251_ _1215_ _1253_ VPWR VGND sg13g2_nand3_1
X_6109_ net1108 VGND VPWR _0208_ DP_2.matrix\[40\] clknet_leaf_49_clk sg13g2_dfrbpq_2
XFILLER_18_108 VPWR VGND sg13g2_fill_2
XFILLER_23_870 VPWR VGND sg13g2_fill_1
XFILLER_41_133 VPWR VGND sg13g2_fill_1
XFILLER_29_1016 VPWR VGND sg13g2_decap_8
XFILLER_29_1027 VPWR VGND sg13g2_fill_2
XFILLER_17_130 VPWR VGND sg13g2_fill_2
XFILLER_45_461 VPWR VGND sg13g2_decap_4
XFILLER_18_664 VPWR VGND sg13g2_fill_1
X_3810_ _0646_ net932 net1003 net933 net1001 VPWR VGND sg13g2_a22oi_1
XFILLER_21_829 VPWR VGND sg13g2_decap_8
XFILLER_32_133 VPWR VGND sg13g2_fill_2
XFILLER_32_144 VPWR VGND sg13g2_fill_2
X_4790_ _1589_ _1555_ _1587_ VPWR VGND sg13g2_xnor2_1
X_3741_ _0584_ _0548_ _0582_ VPWR VGND sg13g2_xnor2_1
X_3672_ _0500_ _0493_ _0463_ _0517_ VPWR VGND sg13g2_a21o_2
X_6460_ net1119 VGND VPWR net52 mac2.sum_lvl2_ff\[10\] clknet_leaf_42_clk sg13g2_dfrbpq_1
X_5411_ mac1.sum_lvl3_ff\[22\] mac1.sum_lvl3_ff\[2\] _2170_ VPWR VGND sg13g2_and2_1
X_6391_ net1121 VGND VPWR _0128_ mac2.products_ff\[78\] clknet_leaf_41_clk sg13g2_dfrbpq_1
X_5342_ VGND VPWR _2113_ _2115_ _2116_ _2114_ sg13g2_a21oi_1
X_5273_ _2051_ _2030_ _2053_ VPWR VGND sg13g2_xor2_1
X_4224_ _1043_ _1042_ _1039_ VPWR VGND sg13g2_nand2b_1
X_4155_ _0979_ _0973_ _0981_ VPWR VGND sg13g2_xor2_1
XFILLER_29_918 VPWR VGND sg13g2_decap_8
X_3106_ _2698_ _2699_ _2689_ _2700_ VPWR VGND sg13g2_nand3_1
X_4086_ _0881_ _0886_ _0915_ VPWR VGND sg13g2_nor2_1
X_3037_ _2630_ _2632_ _2633_ VPWR VGND sg13g2_nor2_1
XFILLER_37_984 VPWR VGND sg13g2_decap_8
X_4988_ _1755_ VPWR _1776_ VGND _1746_ _1756_ sg13g2_o21ai_1
X_3939_ VGND VPWR _0771_ _0770_ _0769_ sg13g2_or2_1
X_5609_ _2319_ VPWR _2325_ VGND _2320_ _2324_ sg13g2_o21ai_1
XFILLER_4_1007 VPWR VGND sg13g2_decap_8
XFILLER_43_932 VPWR VGND sg13g2_decap_8
XFILLER_42_497 VPWR VGND sg13g2_fill_2
XFILLER_11_840 VPWR VGND sg13g2_fill_1
Xinput16 uio_in[7] net16 VPWR VGND sg13g2_buf_1
XFILLER_10_350 VPWR VGND sg13g2_fill_2
XFILLER_6_365 VPWR VGND sg13g2_fill_1
XFILLER_42_1024 VPWR VGND sg13g2_decap_4
X_5960_ net974 _0192_ VPWR VGND sg13g2_buf_1
X_4911_ _1678_ _1680_ _1704_ _1706_ VPWR VGND sg13g2_or3_1
X_5891_ _2570_ _2443_ _2461_ VPWR VGND sg13g2_xnor2_1
XFILLER_34_965 VPWR VGND sg13g2_decap_8
X_4842_ VGND VPWR _1639_ _1612_ _1610_ sg13g2_or2_1
X_4773_ _1521_ _1570_ _1572_ VPWR VGND sg13g2_and2_1
X_3724_ _0566_ _0545_ _0568_ VPWR VGND sg13g2_xor2_1
X_6512_ net1045 VGND VPWR net330 mac2.total_sum\[14\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_6443_ net1127 VGND VPWR net64 mac2.sum_lvl1_ff\[50\] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_3655_ _0501_ _0493_ _0500_ VPWR VGND sg13g2_xnor2_1
X_3586_ _0386_ VPWR _0434_ VGND _0325_ _0387_ sg13g2_o21ai_1
X_6374_ net1102 VGND VPWR _0148_ mac2.products_ff\[9\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_5325_ VGND VPWR _2071_ _2094_ _2102_ _2096_ sg13g2_a21oi_1
X_5256_ _2005_ VPWR _2036_ VGND _2003_ _2006_ sg13g2_o21ai_1
X_4207_ _1023_ _1024_ _1026_ _1027_ VPWR VGND sg13g2_or3_1
X_5187_ _1969_ net858 net793 VPWR VGND sg13g2_nand2_1
X_4138_ _0963_ _0964_ _0965_ VPWR VGND sg13g2_and2_1
XFILLER_28_247 VPWR VGND sg13g2_fill_1
X_4069_ _0898_ net997 net1031 VPWR VGND sg13g2_nand2_1
XFILLER_25_921 VPWR VGND sg13g2_decap_8
XFILLER_25_998 VPWR VGND sg13g2_decap_8
XFILLER_40_924 VPWR VGND sg13g2_decap_8
XFILLER_3_324 VPWR VGND sg13g2_fill_2
Xfanout1103 net1104 net1103 VPWR VGND sg13g2_buf_8
XFILLER_26_1008 VPWR VGND sg13g2_decap_8
Xfanout1114 net1115 net1114 VPWR VGND sg13g2_buf_8
Xfanout1125 net1128 net1125 VPWR VGND sg13g2_buf_8
XFILLER_19_236 VPWR VGND sg13g2_fill_1
XFILLER_15_442 VPWR VGND sg13g2_fill_2
XFILLER_16_987 VPWR VGND sg13g2_decap_8
XFILLER_15_475 VPWR VGND sg13g2_fill_1
XFILLER_31_968 VPWR VGND sg13g2_decap_8
X_3440_ _0290_ _0291_ _0292_ VPWR VGND sg13g2_nor2b_2
X_3371_ _2957_ net968 net1030 VPWR VGND sg13g2_nand2_1
X_6090_ net1041 VGND VPWR _0094_ mac1.products_ff\[141\] clknet_leaf_67_clk sg13g2_dfrbpq_1
X_5110_ VGND VPWR _1894_ _1892_ _1849_ sg13g2_or2_1
X_5041_ _1824_ _1825_ _1819_ _1827_ VPWR VGND sg13g2_nand3_1
X_5943_ net271 _0165_ VPWR VGND sg13g2_buf_1
X_5874_ _2559_ net1008 _2395_ _0178_ VPWR VGND sg13g2_mux2_1
X_4825_ VGND VPWR _1586_ _1588_ _1623_ _1622_ sg13g2_a21oi_1
X_4756_ _1516_ VPWR _1555_ VGND _1471_ _1517_ sg13g2_o21ai_1
X_3707_ _0520_ VPWR _0551_ VGND _0518_ _0521_ sg13g2_o21ai_1
X_4687_ _1484_ _1485_ _1487_ _1488_ VPWR VGND sg13g2_or3_1
X_6426_ net1105 VGND VPWR net75 mac2.sum_lvl1_ff\[13\] clknet_leaf_33_clk sg13g2_dfrbpq_1
X_3638_ _0484_ net1012 net945 VPWR VGND sg13g2_nand2_1
X_3569_ _0413_ _0414_ _0416_ _0417_ VPWR VGND sg13g2_or3_1
X_6357_ net1040 VGND VPWR net422 mac1.total_sum\[8\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_5308_ _2066_ VPWR _2086_ VGND _2038_ _2064_ sg13g2_o21ai_1
X_6288_ net1078 VGND VPWR net54 mac2.sum_lvl1_ff\[75\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_5239_ _2020_ _2011_ _2018_ VPWR VGND sg13g2_xnor2_1
XFILLER_29_501 VPWR VGND sg13g2_fill_1
XFILLER_13_913 VPWR VGND sg13g2_fill_2
XFILLER_33_31 VPWR VGND sg13g2_fill_2
XFILLER_33_86 VPWR VGND sg13g2_fill_2
Xhold5 mac2.sum_lvl1_ff\[8\] VPWR VGND net45 sg13g2_dlygate4sd3_1
XFILLER_48_898 VPWR VGND sg13g2_decap_8
XFILLER_15_283 VPWR VGND sg13g2_fill_2
X_4610_ _1412_ _1389_ _1413_ VPWR VGND sg13g2_xor2_1
X_5590_ _2310_ _2309_ _2308_ VPWR VGND sg13g2_nand2b_1
XFILLER_30_297 VPWR VGND sg13g2_fill_1
X_4541_ _1351_ _1349_ _1350_ VPWR VGND sg13g2_nand2_1
XFILLER_8_983 VPWR VGND sg13g2_decap_8
Xhold416 _0024_ VPWR VGND net456 sg13g2_dlygate4sd3_1
Xhold405 _0049_ VPWR VGND net445 sg13g2_dlygate4sd3_1
Xhold427 mac2.sum_lvl3_ff\[13\] VPWR VGND net467 sg13g2_dlygate4sd3_1
X_4472_ VGND VPWR _1248_ _1250_ _1285_ _1282_ sg13g2_a21oi_1
X_3423_ _0275_ net1017 net950 VPWR VGND sg13g2_nand2_1
X_6211_ net1096 VGND VPWR net76 mac1.sum_lvl2_ff\[6\] clknet_leaf_53_clk sg13g2_dfrbpq_1
Xhold438 _2218_ VPWR VGND net478 sg13g2_dlygate4sd3_1
Xhold449 DP_3.matrix\[72\] VPWR VGND net489 sg13g2_dlygate4sd3_1
Xfanout907 net908 net907 VPWR VGND sg13g2_buf_8
X_6142_ net1106 VGND VPWR _0230_ DP_3.matrix\[38\] clknet_leaf_32_clk sg13g2_dfrbpq_2
Xfanout929 net930 net929 VPWR VGND sg13g2_buf_8
Xfanout918 net919 net918 VPWR VGND sg13g2_buf_2
X_3354_ _2941_ _2932_ _2940_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_0 VPWR VGND sg13g2_fill_1
X_6073_ net1108 VGND VPWR _0184_ DP_1.matrix\[40\] clknet_leaf_49_clk sg13g2_dfrbpq_1
X_3285_ _2874_ net909 net968 VPWR VGND sg13g2_nand2_1
X_5024_ _1810_ _1808_ _1809_ VPWR VGND sg13g2_nand2b_1
XFILLER_0_1010 VPWR VGND sg13g2_decap_8
XFILLER_39_898 VPWR VGND sg13g2_decap_8
X_5926_ net839 net769 _2591_ VPWR VGND sg13g2_nor2_1
X_5857_ _2516_ _2518_ _2549_ _0169_ VPWR VGND sg13g2_mux2_1
X_4808_ _1580_ VPWR _1606_ VGND _1574_ _1581_ sg13g2_o21ai_1
X_5788_ _2469_ net785 _2482_ VPWR VGND sg13g2_nor2_1
XFILLER_6_909 VPWR VGND sg13g2_decap_4
X_4739_ _1536_ _1537_ _1519_ _1539_ VPWR VGND sg13g2_nand3_1
X_6409_ net1056 VGND VPWR _0152_ mac2.products_ff\[148\] clknet_leaf_21_clk sg13g2_dfrbpq_1
XFILLER_0_168 VPWR VGND sg13g2_fill_1
XFILLER_17_548 VPWR VGND sg13g2_fill_2
XFILLER_25_570 VPWR VGND sg13g2_fill_2
XFILLER_44_74 VPWR VGND sg13g2_decap_8
XFILLER_25_581 VPWR VGND sg13g2_fill_1
XFILLER_8_235 VPWR VGND sg13g2_fill_2
XFILLER_5_953 VPWR VGND sg13g2_decap_8
X_3070_ _2665_ _2658_ _2663_ _2664_ VPWR VGND sg13g2_and3_1
X_3972_ _0731_ _0801_ _0803_ _0804_ VPWR VGND sg13g2_or3_1
X_5711_ DP_1.matrix\[43\] net791 _2407_ VPWR VGND sg13g2_nor2_1
X_5642_ mac2.total_sum\[5\] mac1.total_sum\[5\] _2350_ VPWR VGND sg13g2_xor2_1
X_5573_ _2296_ mac2.sum_lvl3_ff\[26\] net463 VPWR VGND sg13g2_xnor2_1
X_4524_ _1307_ _1309_ _1333_ _1335_ VPWR VGND sg13g2_or3_1
Xhold202 mac2.sum_lvl1_ff\[72\] VPWR VGND net242 sg13g2_dlygate4sd3_1
Xhold235 DP_3.matrix\[79\] VPWR VGND net275 sg13g2_dlygate4sd3_1
Xhold213 mac2.products_ff\[148\] VPWR VGND net253 sg13g2_dlygate4sd3_1
Xhold224 mac2.sum_lvl1_ff\[86\] VPWR VGND net264 sg13g2_dlygate4sd3_1
Xhold257 DP_4.matrix\[77\] VPWR VGND net297 sg13g2_dlygate4sd3_1
X_4455_ VGND VPWR _1268_ _1241_ _1239_ sg13g2_or2_1
Xhold246 mac1.sum_lvl2_ff\[0\] VPWR VGND net286 sg13g2_dlygate4sd3_1
Xhold268 DP_4.matrix\[74\] VPWR VGND net308 sg13g2_dlygate4sd3_1
X_3406_ _2988_ _2980_ _2987_ VPWR VGND sg13g2_nand2_1
X_4386_ _1150_ _1199_ _1201_ VPWR VGND sg13g2_and2_1
Xhold279 DP_4.matrix\[38\] VPWR VGND net319 sg13g2_dlygate4sd3_1
X_6125_ net1073 VGND VPWR _0219_ DP_2.matrix\[79\] clknet_leaf_59_clk sg13g2_dfrbpq_1
X_3337_ VGND VPWR _2872_ _2893_ _2925_ _2895_ sg13g2_a21oi_1
X_6056_ net1124 VGND VPWR _0167_ DP_3.matrix\[44\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_3268_ _2858_ _2848_ _2857_ VPWR VGND sg13g2_nand2b_1
XFILLER_22_1011 VPWR VGND sg13g2_decap_8
X_3199_ _2789_ _2790_ _2788_ _2791_ VPWR VGND sg13g2_nand3_1
X_5007_ _1794_ _1787_ _1792_ _1793_ VPWR VGND sg13g2_and3_1
XFILLER_42_849 VPWR VGND sg13g2_decap_8
X_5909_ _2581_ _2501_ _2503_ VPWR VGND sg13g2_xnor2_1
XFILLER_2_945 VPWR VGND sg13g2_decap_8
XFILLER_39_63 VPWR VGND sg13g2_fill_1
XFILLER_33_849 VPWR VGND sg13g2_decap_8
XFILLER_41_893 VPWR VGND sg13g2_decap_8
XFILLER_4_260 VPWR VGND sg13g2_fill_2
X_4240_ _1057_ _1058_ _1019_ _1059_ VPWR VGND sg13g2_nand3_1
XFILLER_45_1022 VPWR VGND sg13g2_decap_8
X_4171_ net886 net831 _0079_ VPWR VGND sg13g2_and2_1
X_3122_ _2715_ _2711_ _2714_ VPWR VGND sg13g2_nand2_1
XFILLER_49_971 VPWR VGND sg13g2_decap_8
X_3053_ _2647_ _2646_ _2649_ VPWR VGND sg13g2_xor2_1
X_3955_ net937 net986 net941 _0787_ VPWR VGND net1035 sg13g2_nand4_1
X_5625_ mac1.total_sum\[1\] mac2.total_sum\[1\] _2337_ VPWR VGND sg13g2_nor2_1
X_3886_ _0717_ _0716_ _0699_ _0720_ VPWR VGND sg13g2_a21o_1
X_5556_ _2280_ VPWR _2283_ VGND _2279_ _2281_ sg13g2_o21ai_1
X_4507_ _1299_ VPWR _1318_ VGND _1270_ _1297_ sg13g2_o21ai_1
X_5487_ net306 _2227_ _0040_ VPWR VGND sg13g2_xor2_1
X_4438_ VGND VPWR _1215_ _1217_ _1252_ _1251_ sg13g2_a21oi_1
X_4369_ _1145_ VPWR _1184_ VGND _1100_ _1146_ sg13g2_o21ai_1
X_6108_ net1046 VGND VPWR _0096_ mac1.products_ff\[147\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_46_429 VPWR VGND sg13g2_fill_1
X_6039_ net1096 VGND VPWR _0123_ mac1.products_ff\[74\] clknet_leaf_51_clk sg13g2_dfrbpq_1
XFILLER_42_657 VPWR VGND sg13g2_fill_2
XFILLER_30_808 VPWR VGND sg13g2_decap_8
XFILLER_10_510 VPWR VGND sg13g2_decap_4
XFILLER_10_565 VPWR VGND sg13g2_fill_1
XFILLER_10_554 VPWR VGND sg13g2_fill_2
XFILLER_6_536 VPWR VGND sg13g2_fill_1
XFILLER_38_919 VPWR VGND sg13g2_decap_8
XFILLER_46_985 VPWR VGND sg13g2_decap_8
XFILLER_14_893 VPWR VGND sg13g2_fill_1
X_3740_ _0548_ _0582_ _0583_ VPWR VGND sg13g2_nor2b_1
XFILLER_32_189 VPWR VGND sg13g2_fill_2
XFILLER_12_1010 VPWR VGND sg13g2_decap_8
X_3671_ _0502_ VPWR _0516_ VGND _0491_ _0503_ sg13g2_o21ai_1
X_5410_ _2166_ VPWR _2169_ VGND _2165_ _2167_ sg13g2_o21ai_1
X_6390_ net1119 VGND VPWR _0137_ mac2.products_ff\[77\] clknet_leaf_42_clk sg13g2_dfrbpq_1
X_5341_ net381 _2113_ _0008_ VPWR VGND sg13g2_xor2_1
X_5272_ _2051_ _2030_ _2052_ VPWR VGND sg13g2_nor2b_1
X_4223_ _1041_ _1018_ _1042_ VPWR VGND sg13g2_xor2_1
X_4154_ _0980_ _0973_ _0979_ VPWR VGND sg13g2_nand2_1
X_3105_ _2696_ _2695_ _2690_ _2699_ VPWR VGND sg13g2_a21o_1
X_4085_ _0912_ _0913_ _0914_ VPWR VGND sg13g2_nor2_1
XFILLER_49_790 VPWR VGND sg13g2_fill_2
X_3036_ net984 net981 net913 net911 _2632_ VPWR VGND sg13g2_and4_1
XFILLER_24_602 VPWR VGND sg13g2_decap_8
XFILLER_37_963 VPWR VGND sg13g2_decap_8
XFILLER_23_112 VPWR VGND sg13g2_fill_1
XFILLER_11_307 VPWR VGND sg13g2_fill_1
X_4987_ _1775_ _1763_ _1774_ VPWR VGND sg13g2_xnor2_1
X_3938_ _0770_ net925 DP_1.matrix\[37\] net927 net999 VPWR VGND sg13g2_a22oi_1
X_3869_ _0702_ _0669_ _0703_ VPWR VGND sg13g2_xor2_1
XFILLER_20_874 VPWR VGND sg13g2_decap_4
Xclkbuf_4_2_0_clk clknet_0_clk clknet_4_2_0_clk VPWR VGND sg13g2_buf_8
X_5608_ _0051_ net311 _2324_ VPWR VGND sg13g2_xnor2_1
X_5539_ VGND VPWR _2271_ mac2.sum_lvl2_ff\[13\] mac2.sum_lvl2_ff\[32\] sg13g2_or2_1
XFILLER_43_911 VPWR VGND sg13g2_decap_8
XFILLER_28_985 VPWR VGND sg13g2_decap_8
XFILLER_15_635 VPWR VGND sg13g2_fill_2
XFILLER_43_988 VPWR VGND sg13g2_decap_8
XFILLER_42_465 VPWR VGND sg13g2_fill_2
XFILLER_14_189 VPWR VGND sg13g2_decap_8
XFILLER_35_1021 VPWR VGND sg13g2_decap_8
XFILLER_7_878 VPWR VGND sg13g2_fill_2
XFILLER_42_1003 VPWR VGND sg13g2_decap_8
XFILLER_19_930 VPWR VGND sg13g2_fill_1
XFILLER_37_259 VPWR VGND sg13g2_fill_2
X_4910_ _1704_ VPWR _1705_ VGND _1678_ _1680_ sg13g2_o21ai_1
X_5890_ VGND VPWR net772 _2569_ _0200_ _2568_ sg13g2_a21oi_1
XFILLER_34_944 VPWR VGND sg13g2_decap_8
X_4841_ _1600_ VPWR _1638_ VGND _1597_ _1601_ sg13g2_o21ai_1
X_4772_ VGND VPWR _1571_ _1570_ _1521_ sg13g2_or2_1
X_3723_ _0566_ _0545_ _0567_ VPWR VGND sg13g2_nor2b_1
X_6511_ net1045 VGND VPWR net470 mac2.total_sum\[13\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_6442_ net1126 VGND VPWR net222 mac2.sum_lvl1_ff\[49\] clknet_leaf_37_clk sg13g2_dfrbpq_1
XFILLER_9_193 VPWR VGND sg13g2_fill_1
X_3654_ _0498_ _0499_ _0500_ VPWR VGND sg13g2_nor2b_1
X_3585_ _0359_ VPWR _0433_ VGND _0429_ _0431_ sg13g2_o21ai_1
X_6373_ net1102 VGND VPWR _0147_ mac2.products_ff\[8\] clknet_leaf_43_clk sg13g2_dfrbpq_1
X_5324_ _2098_ VPWR _2101_ VGND _2083_ _2100_ sg13g2_o21ai_1
X_5255_ _2015_ VPWR _2035_ VGND _2013_ _2016_ sg13g2_o21ai_1
X_4206_ _1026_ net878 net830 net880 net827 VPWR VGND sg13g2_a22oi_1
X_5186_ _1968_ net863 net1021 VPWR VGND sg13g2_nand2_1
X_4137_ _0936_ _0938_ _0962_ _0964_ VPWR VGND sg13g2_or3_1
X_4068_ VGND VPWR _0897_ _0870_ _0868_ sg13g2_or2_1
XFILLER_25_911 VPWR VGND sg13g2_fill_1
X_3019_ _2615_ _2608_ _0066_ VPWR VGND sg13g2_xor2_1
XFILLER_25_977 VPWR VGND sg13g2_decap_8
XFILLER_40_903 VPWR VGND sg13g2_decap_8
Xfanout1104 net1107 net1104 VPWR VGND sg13g2_buf_8
Xfanout1126 net1127 net1126 VPWR VGND sg13g2_buf_8
Xfanout1115 net1116 net1115 VPWR VGND sg13g2_buf_8
XFILLER_47_502 VPWR VGND sg13g2_fill_2
XFILLER_47_546 VPWR VGND sg13g2_fill_2
XFILLER_34_218 VPWR VGND sg13g2_fill_2
XFILLER_16_966 VPWR VGND sg13g2_decap_8
XFILLER_43_796 VPWR VGND sg13g2_decap_4
XFILLER_42_251 VPWR VGND sg13g2_fill_2
XFILLER_31_947 VPWR VGND sg13g2_decap_8
XFILLER_7_642 VPWR VGND sg13g2_fill_2
XFILLER_10_192 VPWR VGND sg13g2_fill_1
XFILLER_7_653 VPWR VGND sg13g2_decap_4
XFILLER_6_152 VPWR VGND sg13g2_fill_1
X_3370_ _2940_ _2932_ _2939_ _2956_ VPWR VGND sg13g2_a21o_1
X_5040_ _1826_ _1819_ _1824_ _1825_ VPWR VGND sg13g2_and3_1
XFILLER_38_557 VPWR VGND sg13g2_decap_4
X_5942_ net1031 _0164_ VPWR VGND sg13g2_buf_1
X_5873_ _2559_ _2428_ _2430_ VPWR VGND sg13g2_xnor2_1
XFILLER_22_969 VPWR VGND sg13g2_decap_8
X_4824_ _1620_ _1593_ _1622_ VPWR VGND sg13g2_xor2_1
XFILLER_21_479 VPWR VGND sg13g2_fill_1
X_4755_ _1544_ VPWR _1554_ VGND _1473_ _1545_ sg13g2_o21ai_1
X_3706_ _0530_ VPWR _0550_ VGND _0528_ _0531_ sg13g2_o21ai_1
X_4686_ _1487_ net890 net849 net891 net845 VPWR VGND sg13g2_a22oi_1
X_6425_ net1105 VGND VPWR net62 mac2.sum_lvl1_ff\[12\] clknet_leaf_33_clk sg13g2_dfrbpq_1
X_3637_ _0483_ net1016 net1032 VPWR VGND sg13g2_nand2_1
X_6356_ net1040 VGND VPWR _0029_ mac1.total_sum\[7\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3568_ _0416_ net1037 net961 net1006 net957 VPWR VGND sg13g2_a22oi_1
X_5307_ _2069_ _2061_ _2068_ _2085_ VPWR VGND sg13g2_a21o_1
X_3499_ _0349_ _0346_ _0348_ VPWR VGND sg13g2_nand2_1
X_6287_ net1078 VGND VPWR net164 mac2.sum_lvl1_ff\[74\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_5238_ _2018_ _2011_ _2019_ VPWR VGND sg13g2_nor2b_1
X_5169_ _1952_ _1946_ _1950_ VPWR VGND sg13g2_xnor2_1
XFILLER_25_752 VPWR VGND sg13g2_fill_2
XFILLER_40_711 VPWR VGND sg13g2_fill_2
XFILLER_12_424 VPWR VGND sg13g2_fill_2
XFILLER_32_1013 VPWR VGND sg13g2_decap_8
XFILLER_33_76 VPWR VGND sg13g2_fill_1
XFILLER_0_884 VPWR VGND sg13g2_decap_8
Xhold6 mac1.sum_lvl2_ff\[50\] VPWR VGND net46 sg13g2_dlygate4sd3_1
XFILLER_48_877 VPWR VGND sg13g2_decap_8
XFILLER_16_763 VPWR VGND sg13g2_fill_2
XFILLER_16_774 VPWR VGND sg13g2_fill_1
X_4540_ _1323_ VPWR _1350_ VGND _1296_ _1321_ sg13g2_o21ai_1
XFILLER_11_490 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_10_clk clknet_4_3_0_clk clknet_leaf_10_clk VPWR VGND sg13g2_buf_8
XFILLER_7_461 VPWR VGND sg13g2_fill_1
Xhold406 DP_1.matrix\[6\] VPWR VGND net446 sg13g2_dlygate4sd3_1
Xhold417 mac2.sum_lvl3_ff\[4\] VPWR VGND net457 sg13g2_dlygate4sd3_1
X_4471_ VPWR _1284_ _1283_ VGND sg13g2_inv_1
X_3422_ _0274_ net951 net1019 net952 net1017 VPWR VGND sg13g2_a22oi_1
X_6210_ net1097 VGND VPWR net140 mac1.sum_lvl2_ff\[5\] clknet_leaf_54_clk sg13g2_dfrbpq_1
Xhold439 _0021_ VPWR VGND net479 sg13g2_dlygate4sd3_1
Xhold428 _2327_ VPWR VGND net468 sg13g2_dlygate4sd3_1
X_6141_ net1096 VGND VPWR net144 mac1.sum_lvl1_ff\[6\] clknet_leaf_53_clk sg13g2_dfrbpq_1
Xfanout919 net920 net919 VPWR VGND sg13g2_buf_8
Xfanout908 net300 net908 VPWR VGND sg13g2_buf_8
X_3353_ _2940_ _2905_ _2938_ VPWR VGND sg13g2_xnor2_1
X_6072_ net1118 VGND VPWR _0183_ DP_1.matrix\[39\] clknet_leaf_52_clk sg13g2_dfrbpq_1
X_3284_ _2856_ _2849_ _2819_ _2873_ VPWR VGND sg13g2_a21o_2
XFILLER_24_0 VPWR VGND sg13g2_fill_2
X_5023_ _1809_ net868 net795 VPWR VGND sg13g2_nand2_1
XFILLER_39_877 VPWR VGND sg13g2_decap_8
XFILLER_22_711 VPWR VGND sg13g2_fill_1
X_5925_ VGND VPWR net769 _2590_ _0246_ _2589_ sg13g2_a21oi_1
X_5856_ _2549_ net770 _2548_ VPWR VGND sg13g2_nand2_1
XFILLER_16_1008 VPWR VGND sg13g2_decap_8
X_4807_ _1603_ _1595_ _1605_ VPWR VGND sg13g2_xor2_1
X_5787_ _2480_ VPWR _2481_ VGND _2475_ net767 sg13g2_o21ai_1
XFILLER_22_799 VPWR VGND sg13g2_fill_2
X_2999_ VPWR _2603_ DP_3.I_range.out_data\[5\] VGND sg13g2_inv_1
X_4738_ _1538_ _1519_ _1536_ _1537_ VPWR VGND sg13g2_and3_1
X_4669_ _1470_ net832 net904 net834 net902 VPWR VGND sg13g2_a22oi_1
X_6408_ net1052 VGND VPWR _0151_ mac2.products_ff\[147\] clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_1_615 VPWR VGND sg13g2_fill_1
X_6339_ net1077 VGND VPWR net122 mac2.sum_lvl3_ff\[26\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_12_276 VPWR VGND sg13g2_fill_2
XFILLER_40_585 VPWR VGND sg13g2_decap_8
XFILLER_40_596 VPWR VGND sg13g2_fill_1
XFILLER_5_910 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_59_clk clknet_4_9_0_clk clknet_leaf_59_clk VPWR VGND sg13g2_buf_8
XFILLER_47_151 VPWR VGND sg13g2_fill_1
X_3971_ VGND VPWR _0799_ _0800_ _0803_ _0765_ sg13g2_a21oi_1
X_5710_ _2395_ net1037 _2404_ _2406_ VPWR VGND sg13g2_a21o_1
X_5641_ mac1.total_sum\[5\] mac2.total_sum\[5\] _2349_ VPWR VGND sg13g2_nor2_1
X_5572_ mac2.sum_lvl3_ff\[26\] net463 _2295_ VPWR VGND sg13g2_and2_1
X_4523_ _1333_ VPWR _1334_ VGND _1307_ _1309_ sg13g2_o21ai_1
Xhold203 mac2.sum_lvl1_ff\[50\] VPWR VGND net243 sg13g2_dlygate4sd3_1
Xhold225 mac1.sum_lvl3_ff\[0\] VPWR VGND net265 sg13g2_dlygate4sd3_1
Xhold214 mac1.sum_lvl1_ff\[86\] VPWR VGND net254 sg13g2_dlygate4sd3_1
Xhold236 DP_4.matrix\[76\] VPWR VGND net276 sg13g2_dlygate4sd3_1
Xhold269 DP_1.matrix\[74\] VPWR VGND net309 sg13g2_dlygate4sd3_1
Xhold247 _0000_ VPWR VGND net287 sg13g2_dlygate4sd3_1
Xhold258 DP_2.matrix\[79\] VPWR VGND net298 sg13g2_dlygate4sd3_1
X_4454_ _1229_ VPWR _1267_ VGND _1226_ _1230_ sg13g2_o21ai_1
X_3405_ _2985_ _2986_ _2987_ VPWR VGND sg13g2_nor2b_1
X_4385_ VGND VPWR _1200_ _1199_ _1150_ sg13g2_or2_1
X_6124_ net1073 VGND VPWR _0218_ DP_2.matrix\[78\] clknet_leaf_61_clk sg13g2_dfrbpq_1
X_3336_ _2922_ _2902_ _2924_ VPWR VGND sg13g2_xor2_1
X_6055_ net1101 VGND VPWR _0166_ DP_3.matrix\[8\] clknet_leaf_26_clk sg13g2_dfrbpq_1
X_3267_ _2857_ _2849_ _2856_ VPWR VGND sg13g2_xnor2_1
X_5006_ _1788_ VPWR _1793_ VGND _1789_ _1791_ sg13g2_o21ai_1
X_3198_ _2742_ VPWR _2790_ VGND _2681_ _2743_ sg13g2_o21ai_1
XFILLER_42_828 VPWR VGND sg13g2_decap_8
X_5908_ net895 net769 _2580_ VPWR VGND sg13g2_nor2_1
X_5839_ _2532_ _2531_ net777 net775 net805 VPWR VGND sg13g2_a22oi_1
XFILLER_5_239 VPWR VGND sg13g2_fill_1
XFILLER_30_33 VPWR VGND sg13g2_fill_1
XFILLER_2_924 VPWR VGND sg13g2_decap_8
XFILLER_39_97 VPWR VGND sg13g2_fill_2
XFILLER_29_184 VPWR VGND sg13g2_fill_1
XFILLER_33_828 VPWR VGND sg13g2_decap_8
XFILLER_40_371 VPWR VGND sg13g2_fill_2
XFILLER_41_872 VPWR VGND sg13g2_decap_8
XFILLER_45_1001 VPWR VGND sg13g2_decap_8
X_4170_ _0122_ _0987_ _0994_ VPWR VGND sg13g2_xnor2_1
X_3121_ _2712_ _2713_ _2714_ VPWR VGND sg13g2_nor2b_1
XFILLER_49_950 VPWR VGND sg13g2_decap_8
X_3052_ _2646_ _2647_ _2648_ VPWR VGND sg13g2_nor2b_2
XFILLER_36_600 VPWR VGND sg13g2_fill_2
XFILLER_35_121 VPWR VGND sg13g2_fill_1
XFILLER_36_666 VPWR VGND sg13g2_fill_1
XFILLER_35_187 VPWR VGND sg13g2_fill_1
XFILLER_36_699 VPWR VGND sg13g2_decap_4
X_3954_ DP_2.matrix\[36\] net937 net986 net1035 _0786_ VPWR VGND sg13g2_and4_1
X_3885_ VGND VPWR _0716_ _0717_ _0719_ _0699_ sg13g2_a21oi_1
XFILLER_32_894 VPWR VGND sg13g2_decap_8
X_5624_ _2336_ mac1.total_sum\[1\] mac2.total_sum\[1\] VPWR VGND sg13g2_nand2_1
X_5555_ _0055_ _2279_ _2282_ VPWR VGND sg13g2_xnor2_1
X_4506_ _1300_ _1294_ _1302_ _1317_ VPWR VGND sg13g2_a21o_1
X_5486_ net305 mac2.sum_lvl2_ff\[21\] _2229_ VPWR VGND sg13g2_xor2_1
X_4437_ _1249_ _1222_ _1251_ VPWR VGND sg13g2_xor2_1
X_6107_ net1098 VGND VPWR _0207_ DP_2.matrix\[39\] clknet_leaf_52_clk sg13g2_dfrbpq_1
X_4368_ _1173_ VPWR _1183_ VGND _1102_ _1174_ sg13g2_o21ai_1
X_3319_ _2887_ VPWR _2907_ VGND _2884_ _2888_ sg13g2_o21ai_1
X_4299_ _1116_ net871 net829 net874 net826 VPWR VGND sg13g2_a22oi_1
X_6038_ net1096 VGND VPWR _0116_ mac1.products_ff\[73\] clknet_leaf_51_clk sg13g2_dfrbpq_1
XFILLER_26_121 VPWR VGND sg13g2_decap_4
XFILLER_41_124 VPWR VGND sg13g2_fill_2
XFILLER_41_157 VPWR VGND sg13g2_decap_8
XFILLER_41_87 VPWR VGND sg13g2_fill_2
XFILLER_37_408 VPWR VGND sg13g2_fill_2
XFILLER_17_110 VPWR VGND sg13g2_fill_1
XFILLER_18_633 VPWR VGND sg13g2_fill_1
XFILLER_46_964 VPWR VGND sg13g2_decap_8
XFILLER_18_655 VPWR VGND sg13g2_decap_8
XFILLER_17_198 VPWR VGND sg13g2_fill_1
XFILLER_9_353 VPWR VGND sg13g2_fill_2
X_3670_ _0488_ _0482_ _0490_ _0515_ VPWR VGND sg13g2_a21o_1
X_5340_ net380 mac1.sum_lvl2_ff\[21\] _2115_ VPWR VGND sg13g2_xor2_1
X_5271_ _2049_ _2048_ _2051_ VPWR VGND sg13g2_xor2_1
X_4222_ _1041_ net883 net821 VPWR VGND sg13g2_nand2_1
X_4153_ _0979_ _0974_ _0977_ VPWR VGND sg13g2_xnor2_1
X_3104_ _2695_ _2696_ _2690_ _2698_ VPWR VGND sg13g2_nand3_1
X_4084_ VGND VPWR _0877_ _0879_ _0913_ _0910_ sg13g2_a21oi_1
X_3035_ _2631_ net982 net911 VPWR VGND sg13g2_nand2_1
XFILLER_37_942 VPWR VGND sg13g2_decap_8
XFILLER_23_102 VPWR VGND sg13g2_fill_2
X_4986_ _1774_ _1771_ _1773_ VPWR VGND sg13g2_nand2_1
X_3937_ net1001 net999 net927 net925 _0769_ VPWR VGND sg13g2_and4_1
X_3868_ _0702_ net998 net933 VPWR VGND sg13g2_nand2_1
XFILLER_20_853 VPWR VGND sg13g2_fill_2
X_3799_ net943 net940 net1000 net998 _0636_ VPWR VGND sg13g2_and4_1
X_5607_ VPWR VGND _2323_ _2322_ _2314_ mac2.sum_lvl3_ff\[31\] _2324_ mac2.sum_lvl3_ff\[11\]
+ sg13g2_a221oi_1
X_5538_ mac2.sum_lvl2_ff\[32\] mac2.sum_lvl2_ff\[13\] _2270_ VPWR VGND sg13g2_and2_1
XFILLER_3_507 VPWR VGND sg13g2_fill_2
X_5469_ _2216_ mac1.sum_lvl3_ff\[34\] mac1.sum_lvl3_ff\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_28_964 VPWR VGND sg13g2_decap_8
XFILLER_43_967 VPWR VGND sg13g2_decap_8
XFILLER_35_1000 VPWR VGND sg13g2_decap_8
XFILLER_10_352 VPWR VGND sg13g2_fill_1
XFILLER_7_868 VPWR VGND sg13g2_fill_1
XFILLER_19_986 VPWR VGND sg13g2_decap_8
XFILLER_46_783 VPWR VGND sg13g2_fill_2
XFILLER_34_923 VPWR VGND sg13g2_decap_8
X_4840_ _1637_ _1631_ _1636_ VPWR VGND sg13g2_xnor2_1
XFILLER_33_444 VPWR VGND sg13g2_fill_2
XFILLER_21_606 VPWR VGND sg13g2_decap_4
X_4771_ _1570_ net839 net891 VPWR VGND sg13g2_nand2_1
XFILLER_21_639 VPWR VGND sg13g2_fill_2
X_6510_ net1045 VGND VPWR net312 mac2.total_sum\[12\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_3722_ _0564_ _0563_ _0566_ VPWR VGND sg13g2_xor2_1
X_6441_ net1126 VGND VPWR net244 mac2.sum_lvl1_ff\[48\] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_3653_ _0494_ VPWR _0499_ VGND _0496_ _0497_ sg13g2_o21ai_1
X_6372_ net1102 VGND VPWR _0146_ mac2.products_ff\[7\] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_5323_ _0154_ _2083_ _2099_ VPWR VGND sg13g2_xnor2_1
X_3584_ _0359_ _0429_ _0431_ _0432_ VPWR VGND sg13g2_or3_1
X_5254_ _2034_ _2033_ _2031_ VPWR VGND sg13g2_nand2b_1
X_4205_ net827 net880 net830 _1025_ VPWR VGND net878 sg13g2_nand4_1
X_5185_ _1942_ VPWR _1967_ VGND _1940_ _1943_ sg13g2_o21ai_1
X_4136_ _0962_ VPWR _0963_ VGND _0936_ _0938_ sg13g2_o21ai_1
X_4067_ _0858_ VPWR _0896_ VGND _0855_ _0859_ sg13g2_o21ai_1
X_3018_ _2616_ _2608_ _2615_ VPWR VGND sg13g2_nand2_1
XFILLER_25_956 VPWR VGND sg13g2_decap_8
XFILLER_12_606 VPWR VGND sg13g2_decap_4
XFILLER_19_1028 VPWR VGND sg13g2_fill_1
X_4969_ _1758_ _1757_ _1745_ VPWR VGND sg13g2_nand2b_1
XFILLER_40_959 VPWR VGND sg13g2_decap_8
XFILLER_3_326 VPWR VGND sg13g2_fill_1
Xfanout1105 net1106 net1105 VPWR VGND sg13g2_buf_8
Xfanout1116 net1117 net1116 VPWR VGND sg13g2_buf_8
Xfanout1127 net1128 net1127 VPWR VGND sg13g2_buf_8
XFILLER_47_536 VPWR VGND sg13g2_fill_2
XFILLER_47_97 VPWR VGND sg13g2_fill_2
XFILLER_16_945 VPWR VGND sg13g2_decap_8
XFILLER_31_926 VPWR VGND sg13g2_decap_8
XFILLER_30_469 VPWR VGND sg13g2_decap_4
XFILLER_7_632 VPWR VGND sg13g2_fill_1
Xclkbuf_4_1_0_clk clknet_0_clk clknet_4_1_0_clk VPWR VGND sg13g2_buf_8
X_5941_ net1033 _0162_ VPWR VGND sg13g2_buf_1
X_5872_ _2558_ net1010 _2395_ _0177_ VPWR VGND sg13g2_mux2_1
XFILLER_22_948 VPWR VGND sg13g2_decap_8
X_4823_ _1621_ _1620_ _1593_ VPWR VGND sg13g2_nand2b_1
X_4754_ _1549_ VPWR _1553_ VGND _1506_ _1551_ sg13g2_o21ai_1
X_3705_ _0549_ _0548_ _0546_ VPWR VGND sg13g2_nand2b_1
XFILLER_30_981 VPWR VGND sg13g2_decap_8
X_4685_ net845 net891 net849 _1486_ VPWR VGND net890 sg13g2_nand4_1
X_3636_ _0457_ VPWR _0482_ VGND _0455_ _0458_ sg13g2_o21ai_1
X_6424_ net1120 VGND VPWR net97 mac2.sum_lvl1_ff\[11\] clknet_leaf_41_clk sg13g2_dfrbpq_1
X_6355_ net1040 VGND VPWR net504 mac1.total_sum\[6\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3567_ net957 net1006 net961 _0415_ VPWR VGND net1037 sg13g2_nand4_1
X_5306_ VGND VPWR _2060_ _2074_ _2084_ _2073_ sg13g2_a21oi_1
X_6286_ net1079 VGND VPWR net71 mac2.sum_lvl1_ff\[73\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_5237_ _2018_ _2012_ _2017_ VPWR VGND sg13g2_xnor2_1
X_3498_ _0345_ _0344_ _0327_ _0348_ VPWR VGND sg13g2_a21o_1
X_5168_ _1951_ _1946_ _1950_ VPWR VGND sg13g2_nand2_1
XFILLER_29_536 VPWR VGND sg13g2_fill_1
X_4119_ _0929_ _0922_ _0931_ _0946_ VPWR VGND sg13g2_a21o_1
X_5099_ _1883_ net792 net866 net795 net863 VPWR VGND sg13g2_a22oi_1
XFILLER_44_517 VPWR VGND sg13g2_decap_4
XFILLER_16_219 VPWR VGND sg13g2_fill_1
XFILLER_25_720 VPWR VGND sg13g2_decap_4
XFILLER_13_937 VPWR VGND sg13g2_decap_8
XFILLER_33_33 VPWR VGND sg13g2_fill_1
XFILLER_40_756 VPWR VGND sg13g2_decap_4
XFILLER_21_992 VPWR VGND sg13g2_decap_8
XFILLER_3_156 VPWR VGND sg13g2_fill_1
Xhold7 mac2.products_ff\[15\] VPWR VGND net47 sg13g2_dlygate4sd3_1
XFILLER_15_263 VPWR VGND sg13g2_decap_8
XFILLER_15_274 VPWR VGND sg13g2_fill_1
XFILLER_15_285 VPWR VGND sg13g2_fill_1
XFILLER_31_778 VPWR VGND sg13g2_fill_1
Xhold407 DP_1.matrix\[7\] VPWR VGND net447 sg13g2_dlygate4sd3_1
Xhold418 _2291_ VPWR VGND net458 sg13g2_dlygate4sd3_1
X_4470_ _1250_ _1282_ _1248_ _1283_ VPWR VGND sg13g2_nand3_1
XFILLER_48_1010 VPWR VGND sg13g2_decap_8
X_3421_ _0072_ _2988_ _0272_ VPWR VGND sg13g2_xnor2_1
Xhold429 _2328_ VPWR VGND net469 sg13g2_dlygate4sd3_1
X_3352_ _2905_ _2938_ _2939_ VPWR VGND sg13g2_nor2b_1
X_6140_ net1122 VGND VPWR _0229_ DP_3.matrix\[37\] clknet_leaf_32_clk sg13g2_dfrbpq_1
Xfanout909 net910 net909 VPWR VGND sg13g2_buf_8
X_6071_ net1108 VGND VPWR _0182_ DP_1.matrix\[38\] clknet_leaf_52_clk sg13g2_dfrbpq_1
X_3283_ _2858_ VPWR _2872_ VGND _2847_ _2859_ sg13g2_o21ai_1
X_5022_ _1785_ VPWR _1808_ VGND _1760_ _1783_ sg13g2_o21ai_1
XFILLER_17_0 VPWR VGND sg13g2_fill_1
XFILLER_39_856 VPWR VGND sg13g2_decap_8
X_5924_ _2532_ _2530_ _2590_ VPWR VGND sg13g2_xor2_1
X_5855_ _2548_ _2545_ _2547_ VPWR VGND sg13g2_nand2b_1
X_4806_ _1603_ _1595_ _1604_ VPWR VGND sg13g2_nor2b_1
X_5786_ _2480_ net1028 net767 VPWR VGND sg13g2_nand2_1
X_2998_ VPWR _2602_ DP_1.Q_range.out_data\[5\] VGND sg13g2_inv_1
X_4737_ _1525_ VPWR _1537_ VGND _1533_ _1535_ sg13g2_o21ai_1
X_4668_ _1446_ VPWR _1469_ VGND _1411_ _1444_ sg13g2_o21ai_1
X_3619_ _0466_ _0461_ _0465_ VPWR VGND sg13g2_nand2_1
X_6407_ net1054 VGND VPWR _0150_ mac2.products_ff\[146\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_4599_ _1403_ _1400_ _1402_ VPWR VGND sg13g2_nand2_1
X_6338_ net1077 VGND VPWR net94 mac2.sum_lvl3_ff\[25\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_6269_ net1041 VGND VPWR net155 mac1.sum_lvl1_ff\[72\] clknet_leaf_67_clk sg13g2_dfrbpq_1
XFILLER_13_712 VPWR VGND sg13g2_fill_2
XFILLER_44_98 VPWR VGND sg13g2_fill_2
XFILLER_5_988 VPWR VGND sg13g2_decap_8
XFILLER_36_859 VPWR VGND sg13g2_decap_8
X_3970_ _0799_ _0800_ _0765_ _0802_ VPWR VGND sg13g2_nand3_1
XFILLER_44_881 VPWR VGND sg13g2_decap_8
X_5640_ VGND VPWR _2345_ _2347_ _2348_ _2346_ sg13g2_a21oi_1
XFILLER_31_575 VPWR VGND sg13g2_fill_1
X_5571_ _0059_ _2292_ net397 VPWR VGND sg13g2_xnor2_1
X_4522_ _1331_ _1317_ _1333_ VPWR VGND sg13g2_xor2_1
Xhold204 mac2.products_ff\[80\] VPWR VGND net244 sg13g2_dlygate4sd3_1
Xhold226 _0016_ VPWR VGND net266 sg13g2_dlygate4sd3_1
Xhold215 mac2.sum_lvl1_ff\[84\] VPWR VGND net255 sg13g2_dlygate4sd3_1
X_4453_ _1266_ _1260_ _1265_ VPWR VGND sg13g2_xnor2_1
Xhold259 DP_3.matrix\[43\] VPWR VGND net299 sg13g2_dlygate4sd3_1
Xhold237 DP_3.matrix\[77\] VPWR VGND net277 sg13g2_dlygate4sd3_1
X_3404_ _2982_ VPWR _2986_ VGND _2983_ _2984_ sg13g2_o21ai_1
Xhold248 mac1.sum_lvl3_ff\[20\] VPWR VGND net288 sg13g2_dlygate4sd3_1
X_4384_ _1199_ net821 net873 VPWR VGND sg13g2_nand2_1
X_6123_ net1067 VGND VPWR net210 mac1.sum_lvl1_ff\[0\] clknet_leaf_63_clk sg13g2_dfrbpq_1
X_3335_ _2922_ _2902_ _2923_ VPWR VGND sg13g2_nor2b_1
X_3266_ _2854_ _2855_ _2856_ VPWR VGND sg13g2_nor2b_1
X_6054_ net1068 VGND VPWR _0165_ DP_2.matrix\[80\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_5005_ _1788_ _1789_ _1791_ _1792_ VPWR VGND sg13g2_or3_1
X_3197_ _2715_ VPWR _2789_ VGND _2785_ _2787_ sg13g2_o21ai_1
XFILLER_27_804 VPWR VGND sg13g2_fill_1
XFILLER_27_859 VPWR VGND sg13g2_decap_8
XFILLER_35_881 VPWR VGND sg13g2_decap_8
X_5907_ VGND VPWR net768 _2579_ _0223_ _2578_ sg13g2_a21oi_1
X_5838_ net823 net841 net786 _2531_ VPWR VGND sg13g2_mux2_1
X_5769_ _2464_ _2463_ net784 net781 net908 VPWR VGND sg13g2_a22oi_1
XFILLER_49_439 VPWR VGND sg13g2_fill_1
XFILLER_7_1018 VPWR VGND sg13g2_decap_8
XFILLER_17_303 VPWR VGND sg13g2_fill_1
XFILLER_44_100 VPWR VGND sg13g2_fill_1
XFILLER_18_848 VPWR VGND sg13g2_fill_1
XFILLER_29_174 VPWR VGND sg13g2_fill_1
XFILLER_45_667 VPWR VGND sg13g2_fill_2
XFILLER_44_155 VPWR VGND sg13g2_decap_8
XFILLER_44_144 VPWR VGND sg13g2_fill_1
XFILLER_41_851 VPWR VGND sg13g2_decap_8
XFILLER_1_980 VPWR VGND sg13g2_decap_8
X_3120_ net982 net907 net985 _2713_ VPWR VGND net905 sg13g2_nand4_1
X_3051_ _2626_ VPWR _2647_ VGND _2617_ _2627_ sg13g2_o21ai_1
XFILLER_35_111 VPWR VGND sg13g2_fill_2
X_3953_ _0785_ net935 net989 VPWR VGND sg13g2_nand2_1
XFILLER_16_391 VPWR VGND sg13g2_fill_1
X_3884_ _0716_ _0717_ _0699_ _0718_ VPWR VGND sg13g2_nand3_1
XFILLER_32_873 VPWR VGND sg13g2_decap_8
X_5623_ _2335_ mac1.total_sum\[0\] mac2.total_sum\[0\] VPWR VGND sg13g2_nand2_1
X_5554_ mac2.sum_lvl3_ff\[1\] mac2.sum_lvl3_ff\[21\] _2282_ VPWR VGND sg13g2_xor2_1
X_4505_ _1316_ _1313_ _0130_ VPWR VGND sg13g2_xor2_1
X_5485_ mac2.sum_lvl2_ff\[21\] net305 _2228_ VPWR VGND sg13g2_and2_1
X_4436_ _1250_ _1249_ _1222_ VPWR VGND sg13g2_nand2b_1
X_4367_ _1178_ VPWR _1182_ VGND _1135_ _1180_ sg13g2_o21ai_1
X_6106_ net1109 VGND VPWR _0206_ DP_2.matrix\[38\] clknet_leaf_52_clk sg13g2_dfrbpq_1
X_3318_ _2906_ _2905_ _2903_ VPWR VGND sg13g2_nand2b_1
X_4298_ net826 net874 net830 _1115_ VPWR VGND net871 sg13g2_nand4_1
X_6037_ net1097 VGND VPWR _0078_ mac1.products_ff\[72\] clknet_leaf_54_clk sg13g2_dfrbpq_1
X_3249_ _2839_ net978 net1030 VPWR VGND sg13g2_nand2_1
XFILLER_27_689 VPWR VGND sg13g2_decap_4
XFILLER_42_659 VPWR VGND sg13g2_fill_1
XFILLER_41_169 VPWR VGND sg13g2_fill_1
XFILLER_10_556 VPWR VGND sg13g2_fill_1
XFILLER_2_700 VPWR VGND sg13g2_fill_1
XFILLER_46_943 VPWR VGND sg13g2_decap_8
XFILLER_17_144 VPWR VGND sg13g2_fill_2
XFILLER_17_188 VPWR VGND sg13g2_fill_1
XFILLER_14_884 VPWR VGND sg13g2_fill_1
XFILLER_41_681 VPWR VGND sg13g2_fill_1
X_5270_ _2049_ _2048_ _2050_ VPWR VGND sg13g2_nor2b_1
XFILLER_5_593 VPWR VGND sg13g2_fill_2
X_4221_ _1040_ net883 net819 VPWR VGND sg13g2_nand2_1
X_4152_ _0978_ _0977_ _0974_ VPWR VGND sg13g2_nand2b_1
X_3103_ _2697_ _2690_ _2695_ _2696_ VPWR VGND sg13g2_and3_1
X_4083_ VPWR _0912_ _0911_ VGND sg13g2_inv_1
X_3034_ _2630_ net911 net984 net913 net981 VPWR VGND sg13g2_a22oi_1
XFILLER_37_921 VPWR VGND sg13g2_decap_8
XFILLER_36_453 VPWR VGND sg13g2_decap_4
XFILLER_37_998 VPWR VGND sg13g2_decap_8
X_4985_ _1770_ _1769_ _1764_ _1773_ VPWR VGND sg13g2_a21o_1
X_3936_ _0768_ net999 net925 VPWR VGND sg13g2_nand2_1
X_3867_ _0701_ net998 net931 VPWR VGND sg13g2_nand2_1
X_3798_ _0635_ net1002 net936 VPWR VGND sg13g2_nand2_1
XFILLER_20_898 VPWR VGND sg13g2_fill_1
X_5606_ _2313_ _2317_ _2323_ VPWR VGND sg13g2_nor2_1
X_5537_ _2263_ VPWR _2269_ VGND _2264_ _2268_ sg13g2_o21ai_1
X_5468_ _0020_ _2213_ net368 VPWR VGND sg13g2_xnor2_1
X_5399_ net460 mac1.sum_lvl2_ff\[33\] _2162_ VPWR VGND sg13g2_xor2_1
X_4419_ _1232_ _1224_ _1233_ VPWR VGND sg13g2_nor2b_1
XFILLER_28_943 VPWR VGND sg13g2_decap_8
XFILLER_43_946 VPWR VGND sg13g2_decap_8
XFILLER_42_423 VPWR VGND sg13g2_fill_2
XFILLER_19_965 VPWR VGND sg13g2_decap_8
XFILLER_34_902 VPWR VGND sg13g2_decap_8
XFILLER_34_979 VPWR VGND sg13g2_decap_8
X_4770_ _1569_ net896 net836 VPWR VGND sg13g2_nand2_1
X_3721_ _0564_ _0563_ _0565_ VPWR VGND sg13g2_nor2b_1
X_3652_ _0494_ _0496_ _0497_ _0498_ VPWR VGND sg13g2_nor3_1
X_6440_ net1125 VGND VPWR net223 mac2.sum_lvl1_ff\[47\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_3583_ VGND VPWR _0427_ _0428_ _0431_ _0393_ sg13g2_a21oi_1
X_6371_ net1100 VGND VPWR _0145_ mac2.products_ff\[6\] clknet_leaf_29_clk sg13g2_dfrbpq_1
X_5322_ VPWR _2100_ _2099_ VGND sg13g2_inv_1
XFILLER_6_880 VPWR VGND sg13g2_fill_2
X_5253_ VGND VPWR _2033_ _2032_ _1980_ sg13g2_or2_1
X_4204_ net830 net828 net880 net878 _1024_ VPWR VGND sg13g2_and4_1
X_5184_ _1934_ VPWR _1966_ VGND _1881_ _1932_ sg13g2_o21ai_1
X_4135_ _0960_ _0946_ _0962_ VPWR VGND sg13g2_xor2_1
XFILLER_3_1010 VPWR VGND sg13g2_decap_8
X_4066_ _0895_ _0889_ _0894_ VPWR VGND sg13g2_xnor2_1
X_3017_ _2613_ _2614_ _2615_ VPWR VGND sg13g2_nor2b_1
XFILLER_25_935 VPWR VGND sg13g2_decap_8
XFILLER_19_1007 VPWR VGND sg13g2_decap_8
XFILLER_24_423 VPWR VGND sg13g2_fill_2
X_4968_ _1756_ _1746_ _1757_ VPWR VGND sg13g2_xor2_1
XFILLER_40_938 VPWR VGND sg13g2_decap_8
X_4899_ _1694_ _1693_ _1690_ VPWR VGND sg13g2_nand2b_1
X_3919_ _0740_ VPWR _0752_ VGND _0748_ _0750_ sg13g2_o21ai_1
Xfanout1117 net1118 net1117 VPWR VGND sg13g2_buf_8
Xfanout1128 net1129 net1128 VPWR VGND sg13g2_buf_8
Xfanout1106 net1107 net1106 VPWR VGND sg13g2_buf_8
XFILLER_47_504 VPWR VGND sg13g2_fill_1
XFILLER_47_43 VPWR VGND sg13g2_fill_1
XFILLER_47_548 VPWR VGND sg13g2_fill_1
XFILLER_16_913 VPWR VGND sg13g2_fill_1
XFILLER_31_905 VPWR VGND sg13g2_decap_8
XFILLER_42_253 VPWR VGND sg13g2_fill_1
XFILLER_42_297 VPWR VGND sg13g2_fill_1
XFILLER_8_48 VPWR VGND sg13g2_fill_2
XFILLER_7_600 VPWR VGND sg13g2_fill_2
XFILLER_11_673 VPWR VGND sg13g2_fill_1
XFILLER_7_644 VPWR VGND sg13g2_fill_1
XFILLER_3_861 VPWR VGND sg13g2_fill_2
XFILLER_3_894 VPWR VGND sg13g2_fill_2
XFILLER_38_537 VPWR VGND sg13g2_decap_8
X_5940_ net1036 _0161_ VPWR VGND sg13g2_buf_1
X_5871_ _2558_ _2411_ _2427_ VPWR VGND sg13g2_xnor2_1
XFILLER_22_927 VPWR VGND sg13g2_decap_8
XFILLER_15_990 VPWR VGND sg13g2_decap_8
X_4822_ _1618_ _1594_ _1620_ VPWR VGND sg13g2_xor2_1
XFILLER_30_960 VPWR VGND sg13g2_decap_8
X_4753_ _1551_ _1506_ _0147_ VPWR VGND sg13g2_xor2_1
X_3704_ VGND VPWR _0548_ _0547_ _0495_ sg13g2_or2_1
X_6423_ net1119 VGND VPWR net48 mac2.sum_lvl1_ff\[10\] clknet_leaf_41_clk sg13g2_dfrbpq_1
X_4684_ net849 net845 net892 net890 _1485_ VPWR VGND sg13g2_and4_1
X_3635_ _0449_ VPWR _0481_ VGND _0396_ _0447_ sg13g2_o21ai_1
X_6354_ net1040 VGND VPWR net322 mac1.total_sum\[5\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_3566_ net961 net957 net1006 net1037 _0414_ VPWR VGND sg13g2_and4_1
X_5305_ _2083_ _2082_ _2077_ _2081_ _2059_ VPWR VGND sg13g2_a22oi_1
X_3497_ VGND VPWR _0344_ _0345_ _0347_ _0327_ sg13g2_a21oi_1
X_6285_ net1079 VGND VPWR net74 mac2.sum_lvl1_ff\[72\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_5236_ _2016_ _2013_ _2017_ VPWR VGND sg13g2_xor2_1
X_5167_ _1948_ _1949_ _1950_ VPWR VGND sg13g2_nor2_1
X_4118_ _0945_ _0942_ _0119_ VPWR VGND sg13g2_xor2_1
X_5098_ net866 net863 net795 net792 _1882_ VPWR VGND sg13g2_and4_1
X_4049_ _0879_ _0878_ _0851_ VPWR VGND sg13g2_nand2b_1
XFILLER_8_408 VPWR VGND sg13g2_fill_1
XFILLER_40_779 VPWR VGND sg13g2_fill_2
XFILLER_21_971 VPWR VGND sg13g2_decap_8
XFILLER_20_470 VPWR VGND sg13g2_fill_2
Xhold8 mac2.products_ff\[10\] VPWR VGND net48 sg13g2_dlygate4sd3_1
XFILLER_15_231 VPWR VGND sg13g2_fill_2
XFILLER_16_765 VPWR VGND sg13g2_fill_1
XFILLER_12_982 VPWR VGND sg13g2_decap_8
XFILLER_8_997 VPWR VGND sg13g2_decap_8
Xhold408 DP_1.matrix\[5\] VPWR VGND net448 sg13g2_dlygate4sd3_1
X_3420_ _0273_ _0272_ _2988_ VPWR VGND sg13g2_nand2b_1
Xhold419 _0058_ VPWR VGND net459 sg13g2_dlygate4sd3_1
X_3351_ _2938_ _2933_ _2936_ VPWR VGND sg13g2_xnor2_1
X_6070_ net1108 VGND VPWR _0181_ DP_1.matrix\[37\] clknet_leaf_51_clk sg13g2_dfrbpq_1
X_3282_ _2844_ _2838_ _2846_ _2871_ VPWR VGND sg13g2_a21o_1
XFILLER_24_2 VPWR VGND sg13g2_fill_1
X_5021_ _1807_ _1799_ _1801_ VPWR VGND sg13g2_nand2_1
XFILLER_39_835 VPWR VGND sg13g2_decap_8
XFILLER_0_1024 VPWR VGND sg13g2_decap_4
X_5923_ net841 net769 _2589_ VPWR VGND sg13g2_nor2_1
X_5854_ _2547_ _2546_ net778 net776 net794 VPWR VGND sg13g2_a22oi_1
X_4805_ _1603_ _1596_ _1602_ VPWR VGND sg13g2_xnor2_1
XFILLER_22_768 VPWR VGND sg13g2_fill_2
X_2997_ VPWR _2601_ DP_1.I_range.out_data\[5\] VGND sg13g2_inv_1
X_5785_ _2476_ _2477_ _2468_ _2479_ VPWR VGND sg13g2_nand3_1
X_4736_ _1525_ _1533_ _1535_ _1536_ VPWR VGND sg13g2_or3_1
X_4667_ _1460_ VPWR _1468_ VGND _1440_ _1461_ sg13g2_o21ai_1
X_3618_ _0463_ _0464_ _0465_ VPWR VGND sg13g2_nor2_1
X_6406_ net1060 VGND VPWR _0159_ mac2.products_ff\[145\] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_6337_ net1078 VGND VPWR net44 mac2.sum_lvl3_ff\[24\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_4598_ _1399_ _1398_ _1393_ _1402_ VPWR VGND sg13g2_a21o_1
XFILLER_1_639 VPWR VGND sg13g2_fill_1
X_3549_ net1017 net1016 net946 net944 _0397_ VPWR VGND sg13g2_and4_1
X_6268_ net1057 VGND VPWR net235 mac2.sum_lvl2_ff\[53\] clknet_leaf_23_clk sg13g2_dfrbpq_1
XFILLER_0_149 VPWR VGND sg13g2_fill_1
X_6199_ net1115 VGND VPWR net206 mac1.sum_lvl1_ff\[46\] clknet_leaf_48_clk sg13g2_dfrbpq_1
X_5219_ _1973_ _1967_ _1975_ _2000_ VPWR VGND sg13g2_a21o_1
XFILLER_45_838 VPWR VGND sg13g2_fill_1
XFILLER_17_518 VPWR VGND sg13g2_fill_2
XFILLER_25_595 VPWR VGND sg13g2_decap_8
XFILLER_8_249 VPWR VGND sg13g2_fill_1
XFILLER_5_967 VPWR VGND sg13g2_decap_8
Xclkbuf_4_0_0_clk clknet_0_clk clknet_4_0_0_clk VPWR VGND sg13g2_buf_8
XFILLER_4_444 VPWR VGND sg13g2_fill_1
XFILLER_48_610 VPWR VGND sg13g2_fill_1
XFILLER_29_890 VPWR VGND sg13g2_decap_8
XFILLER_35_326 VPWR VGND sg13g2_fill_1
XFILLER_36_838 VPWR VGND sg13g2_decap_8
XFILLER_16_573 VPWR VGND sg13g2_fill_1
X_5570_ net396 mac2.sum_lvl3_ff\[25\] _2294_ VPWR VGND sg13g2_xor2_1
X_4521_ _1332_ _1317_ _1331_ VPWR VGND sg13g2_nand2_1
X_4452_ _1264_ _1261_ _1265_ VPWR VGND sg13g2_xor2_1
Xhold216 mac1.sum_lvl1_ff\[74\] VPWR VGND net256 sg13g2_dlygate4sd3_1
Xhold205 mac2.products_ff\[9\] VPWR VGND net245 sg13g2_dlygate4sd3_1
X_3403_ _2982_ _2983_ _2984_ _2985_ VPWR VGND sg13g2_nor3_1
Xhold249 _0023_ VPWR VGND net289 sg13g2_dlygate4sd3_1
Xhold238 DP_1.matrix\[43\] VPWR VGND net278 sg13g2_dlygate4sd3_1
Xhold227 mac2.sum_lvl2_ff\[0\] VPWR VGND net267 sg13g2_dlygate4sd3_1
X_4383_ _1198_ net879 DP_4.matrix\[41\] VPWR VGND sg13g2_nand2_1
X_6122_ net1073 VGND VPWR _0217_ DP_2.matrix\[77\] clknet_leaf_60_clk sg13g2_dfrbpq_1
X_3334_ _2920_ _2919_ _2922_ VPWR VGND sg13g2_xor2_1
X_3265_ _2850_ VPWR _2855_ VGND _2852_ _2853_ sg13g2_o21ai_1
X_6053_ net1111 VGND VPWR _0164_ DP_2.matrix\[44\] clknet_leaf_46_clk sg13g2_dfrbpq_2
XFILLER_22_1025 VPWR VGND sg13g2_decap_4
X_5004_ _1791_ net857 net811 net859 net808 VPWR VGND sg13g2_a22oi_1
X_3196_ _2715_ _2785_ _2787_ _2788_ VPWR VGND sg13g2_or3_1
XFILLER_38_153 VPWR VGND sg13g2_fill_2
XFILLER_26_326 VPWR VGND sg13g2_fill_1
XFILLER_27_838 VPWR VGND sg13g2_fill_1
XFILLER_35_860 VPWR VGND sg13g2_decap_8
X_5906_ _2500_ _2488_ _2579_ VPWR VGND sg13g2_xor2_1
X_5837_ _2526_ _2529_ _2530_ VPWR VGND sg13g2_nor2_1
X_5768_ net948 DP_2.matrix\[42\] net788 _2463_ VPWR VGND sg13g2_mux2_1
X_4719_ _1491_ VPWR _1519_ VGND _1482_ _1492_ sg13g2_o21ai_1
X_5699_ DP_1.Q_range.out_data\[2\] DP_1.I_range.out_data\[6\] _2391_ _2394_ _2395_
+ VPWR VGND sg13g2_or4_1
XFILLER_2_959 VPWR VGND sg13g2_decap_8
XFILLER_44_134 VPWR VGND sg13g2_fill_1
XFILLER_26_871 VPWR VGND sg13g2_decap_8
XFILLER_38_1010 VPWR VGND sg13g2_decap_8
XFILLER_41_830 VPWR VGND sg13g2_decap_8
XFILLER_40_373 VPWR VGND sg13g2_fill_1
X_3050_ _2646_ _2634_ _2645_ VPWR VGND sg13g2_xnor2_1
XFILLER_49_985 VPWR VGND sg13g2_decap_8
XFILLER_36_602 VPWR VGND sg13g2_fill_1
X_3952_ _0744_ VPWR _0784_ VGND _0742_ _0745_ sg13g2_o21ai_1
XFILLER_32_852 VPWR VGND sg13g2_decap_8
X_3883_ _0715_ _0714_ _0705_ _0717_ VPWR VGND sg13g2_a21o_1
XFILLER_31_340 VPWR VGND sg13g2_fill_2
X_5622_ net290 mac2.sum_lvl3_ff\[20\] _0048_ VPWR VGND sg13g2_xor2_1
X_5553_ mac2.sum_lvl3_ff\[21\] mac2.sum_lvl3_ff\[1\] _2281_ VPWR VGND sg13g2_nor2_1
X_4504_ VGND VPWR _1315_ _1316_ _1314_ _1256_ sg13g2_a21oi_2
X_5484_ _2224_ VPWR _2227_ VGND _2223_ _2225_ sg13g2_o21ai_1
X_4435_ _1247_ _1223_ _1249_ VPWR VGND sg13g2_xor2_1
X_4366_ _1180_ _1135_ _0136_ VPWR VGND sg13g2_xor2_1
X_3317_ VGND VPWR _2905_ _2904_ _2851_ sg13g2_or2_1
X_6105_ net1044 VGND VPWR _0095_ mac1.products_ff\[146\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_4297_ DP_4.matrix\[36\] net826 net874 net872 _1114_ VPWR VGND sg13g2_and4_1
X_6036_ net1092 VGND VPWR _0077_ mac1.products_ff\[71\] clknet_leaf_56_clk sg13g2_dfrbpq_1
X_3248_ _2813_ VPWR _2838_ VGND _2811_ _2814_ sg13g2_o21ai_1
X_3179_ net919 net964 net922 _2771_ VPWR VGND net1033 sg13g2_nand4_1
XFILLER_35_690 VPWR VGND sg13g2_fill_2
XFILLER_22_373 VPWR VGND sg13g2_fill_2
XFILLER_29_1009 VPWR VGND sg13g2_decap_8
XFILLER_46_922 VPWR VGND sg13g2_decap_8
XFILLER_18_624 VPWR VGND sg13g2_fill_1
XFILLER_45_432 VPWR VGND sg13g2_fill_2
XFILLER_46_999 VPWR VGND sg13g2_decap_8
XFILLER_45_465 VPWR VGND sg13g2_fill_1
XFILLER_32_159 VPWR VGND sg13g2_fill_2
XFILLER_12_1024 VPWR VGND sg13g2_decap_4
XFILLER_5_583 VPWR VGND sg13g2_fill_2
X_4220_ _1039_ net886 net818 VPWR VGND sg13g2_nand2_1
X_4151_ _0976_ _0949_ _0977_ VPWR VGND sg13g2_xor2_1
X_3102_ _2691_ VPWR _2696_ VGND _2692_ _2694_ sg13g2_o21ai_1
X_4082_ _0879_ _0910_ _0877_ _0911_ VPWR VGND sg13g2_nand3_1
XFILLER_37_900 VPWR VGND sg13g2_decap_8
X_3033_ _0067_ _2616_ _2628_ VPWR VGND sg13g2_xnor2_1
XFILLER_37_977 VPWR VGND sg13g2_decap_8
X_4984_ VGND VPWR _1769_ _1770_ _1772_ _1764_ sg13g2_a21oi_1
X_3935_ _0767_ net1004 net1031 VPWR VGND sg13g2_nand2_1
X_3866_ _0700_ net1001 net930 VPWR VGND sg13g2_nand2_1
X_5605_ _2311_ _2316_ _2322_ VPWR VGND sg13g2_nor2_1
X_3797_ VGND VPWR _0634_ _0629_ _0627_ sg13g2_or2_1
X_5536_ _0035_ _2265_ _2268_ VPWR VGND sg13g2_xnor2_1
X_5467_ _2215_ mac1.sum_lvl3_ff\[33\] net367 VPWR VGND sg13g2_xnor2_1
X_4418_ _1232_ _1225_ _1231_ VPWR VGND sg13g2_xnor2_1
X_5398_ mac1.sum_lvl2_ff\[33\] mac1.sum_lvl2_ff\[14\] _2161_ VPWR VGND sg13g2_nor2_1
XFILLER_28_1020 VPWR VGND sg13g2_decap_8
X_4349_ _1154_ _1162_ _1164_ _1165_ VPWR VGND sg13g2_or3_1
XFILLER_46_207 VPWR VGND sg13g2_fill_2
X_6019_ net1072 VGND VPWR _0071_ mac1.products_ff\[2\] clknet_leaf_56_clk sg13g2_dfrbpq_1
XFILLER_28_922 VPWR VGND sg13g2_decap_8
XFILLER_43_925 VPWR VGND sg13g2_decap_8
XFILLER_28_999 VPWR VGND sg13g2_decap_8
XFILLER_10_310 VPWR VGND sg13g2_fill_1
XFILLER_23_693 VPWR VGND sg13g2_decap_4
XFILLER_11_899 VPWR VGND sg13g2_decap_4
XFILLER_7_0 VPWR VGND sg13g2_fill_2
XFILLER_42_1017 VPWR VGND sg13g2_decap_8
XFILLER_42_1028 VPWR VGND sg13g2_fill_1
Xfanout890 net324 net890 VPWR VGND sg13g2_buf_8
XFILLER_18_454 VPWR VGND sg13g2_fill_1
XFILLER_33_424 VPWR VGND sg13g2_fill_1
XFILLER_34_958 VPWR VGND sg13g2_decap_8
X_3720_ VGND VPWR _0524_ _0535_ _0564_ _0523_ sg13g2_a21oi_1
Xclkbuf_leaf_40_clk clknet_4_14_0_clk clknet_leaf_40_clk VPWR VGND sg13g2_buf_8
X_3651_ _0497_ net1005 net953 net1008 net950 VPWR VGND sg13g2_a22oi_1
X_3582_ _0427_ _0428_ _0393_ _0430_ VPWR VGND sg13g2_nand3_1
X_6370_ net1099 VGND VPWR _0138_ mac2.products_ff\[5\] clknet_leaf_29_clk sg13g2_dfrbpq_1
X_5321_ _2097_ _2084_ _2099_ VPWR VGND sg13g2_xor2_1
XFILLER_6_892 VPWR VGND sg13g2_fill_1
X_5252_ _2032_ net799 net1024 VPWR VGND sg13g2_nand2_2
X_4203_ _1023_ net882 net823 VPWR VGND sg13g2_nand2_1
X_5183_ _1954_ VPWR _1965_ VGND _1938_ _1955_ sg13g2_o21ai_1
X_4134_ _0961_ _0946_ _0960_ VPWR VGND sg13g2_nand2_1
XFILLER_29_708 VPWR VGND sg13g2_fill_2
X_4065_ _0893_ _0890_ _0894_ VPWR VGND sg13g2_xor2_1
X_3016_ _2610_ VPWR _2614_ VGND _2611_ _2612_ sg13g2_o21ai_1
XFILLER_36_262 VPWR VGND sg13g2_fill_1
XFILLER_40_917 VPWR VGND sg13g2_decap_8
X_4967_ _1756_ _1747_ _1754_ VPWR VGND sg13g2_xnor2_1
X_4898_ _1692_ _1666_ _1693_ VPWR VGND sg13g2_xor2_1
X_3918_ _0740_ _0748_ _0750_ _0751_ VPWR VGND sg13g2_or3_1
Xclkbuf_leaf_31_clk clknet_4_13_0_clk clknet_leaf_31_clk VPWR VGND sg13g2_buf_8
X_3849_ _0673_ _0681_ _0683_ _0684_ VPWR VGND sg13g2_or3_1
X_5519_ _0047_ _2251_ _2254_ VPWR VGND sg13g2_xnor2_1
X_6499_ net1039 VGND VPWR net450 mac2.total_sum\[1\] clknet_leaf_3_clk sg13g2_dfrbpq_1
Xfanout1118 net1129 net1118 VPWR VGND sg13g2_buf_8
Xfanout1129 rst_n net1129 VPWR VGND sg13g2_buf_8
Xfanout1107 rst_n net1107 VPWR VGND sg13g2_buf_8
XFILLER_8_27 VPWR VGND sg13g2_fill_2
XFILLER_11_641 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_22_clk clknet_4_5_0_clk clknet_leaf_22_clk VPWR VGND sg13g2_buf_8
X_5870_ VGND VPWR net772 _2557_ _0176_ _2556_ sg13g2_a21oi_1
X_4821_ _1619_ _1594_ _1618_ VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_13_clk clknet_4_6_0_clk clknet_leaf_13_clk VPWR VGND sg13g2_buf_8
X_4752_ _1504_ _1505_ _1549_ _1550_ _1552_ VPWR VGND sg13g2_and4_1
X_3703_ _0547_ net949 net1038 VPWR VGND sg13g2_nand2_1
X_4683_ _1484_ net841 net893 VPWR VGND sg13g2_nand2_1
X_3634_ _0469_ VPWR _0480_ VGND _0453_ _0470_ sg13g2_o21ai_1
X_6422_ net1103 VGND VPWR net245 mac2.sum_lvl1_ff\[9\] clknet_leaf_43_clk sg13g2_dfrbpq_1
X_6353_ net1039 VGND VPWR net408 mac1.total_sum\[4\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_3565_ _0413_ net955 net1007 VPWR VGND sg13g2_nand2_1
X_5304_ _2076_ VPWR _2082_ VGND _2053_ _2054_ sg13g2_o21ai_1
X_3496_ _0344_ _0345_ _0327_ _0346_ VPWR VGND sg13g2_nand3_1
X_6284_ net1073 VGND VPWR net211 mac1.sum_lvl1_ff\[87\] clknet_leaf_59_clk sg13g2_dfrbpq_1
X_5235_ _2016_ _1969_ _2014_ VPWR VGND sg13g2_xnor2_1
XFILLER_25_1012 VPWR VGND sg13g2_decap_8
X_5166_ _1949_ net1025 net806 net851 net804 VPWR VGND sg13g2_a22oi_1
X_4117_ VGND VPWR _0944_ _0945_ _0943_ _0885_ sg13g2_a21oi_2
X_5097_ _1881_ net863 net792 VPWR VGND sg13g2_nand2_1
X_4048_ _0876_ _0852_ _0878_ VPWR VGND sg13g2_xor2_1
XFILLER_37_560 VPWR VGND sg13g2_decap_4
XFILLER_13_906 VPWR VGND sg13g2_decap_8
X_5999_ net821 _0255_ VPWR VGND sg13g2_buf_1
XFILLER_21_950 VPWR VGND sg13g2_decap_8
XFILLER_32_1027 VPWR VGND sg13g2_fill_2
XFILLER_0_898 VPWR VGND sg13g2_decap_8
Xhold9 mac2.sum_lvl1_ff\[36\] VPWR VGND net49 sg13g2_dlygate4sd3_1
XFILLER_15_254 VPWR VGND sg13g2_fill_1
XFILLER_8_976 VPWR VGND sg13g2_decap_8
Xhold409 mac2.sum_lvl3_ff\[20\] VPWR VGND net449 sg13g2_dlygate4sd3_1
X_3350_ _2937_ _2936_ _2933_ VPWR VGND sg13g2_nand2b_1
X_3281_ _2869_ _2867_ _0095_ VPWR VGND sg13g2_xor2_1
X_5020_ _0149_ _1779_ _1806_ VPWR VGND sg13g2_xnor2_1
Xclkbuf_leaf_2_clk clknet_4_0_0_clk clknet_leaf_2_clk VPWR VGND sg13g2_buf_8
XFILLER_0_1003 VPWR VGND sg13g2_decap_8
X_5922_ VGND VPWR net768 _2588_ _0245_ _2587_ sg13g2_a21oi_1
X_5853_ DP_4.matrix\[43\] net832 _2472_ _2546_ VPWR VGND sg13g2_mux2_1
X_4804_ _1601_ _1597_ _1602_ VPWR VGND sg13g2_xor2_1
X_5784_ _2478_ _2468_ _2476_ _2477_ VPWR VGND sg13g2_and3_2
X_2996_ VPWR _2600_ DP_1.Q_range.out_data\[3\] VGND sg13g2_inv_1
XFILLER_21_279 VPWR VGND sg13g2_fill_2
X_4735_ VGND VPWR _1531_ _1532_ _1535_ _1526_ sg13g2_a21oi_1
X_4666_ _1467_ _1466_ _0145_ VPWR VGND sg13g2_xor2_1
X_3617_ _0464_ net1038 net958 net1005 net955 VPWR VGND sg13g2_a22oi_1
X_6405_ net1060 VGND VPWR _0158_ mac2.products_ff\[144\] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_4597_ VGND VPWR _1398_ _1399_ _1401_ _1393_ sg13g2_a21oi_1
X_3548_ _0396_ net1016 net944 VPWR VGND sg13g2_nand2_1
X_6336_ net1083 VGND VPWR net137 mac2.sum_lvl3_ff\[23\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_3479_ _0329_ net1014 net950 VPWR VGND sg13g2_nand2_1
X_6267_ net1058 VGND VPWR net264 mac2.sum_lvl2_ff\[52\] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_6198_ net1113 VGND VPWR net219 mac1.sum_lvl1_ff\[45\] clknet_leaf_49_clk sg13g2_dfrbpq_1
X_5218_ _1998_ _1996_ _0150_ VPWR VGND sg13g2_xor2_1
X_5149_ _1932_ net860 net795 VPWR VGND sg13g2_nand2_1
XFILLER_38_891 VPWR VGND sg13g2_decap_8
XFILLER_44_34 VPWR VGND sg13g2_fill_2
XFILLER_13_714 VPWR VGND sg13g2_fill_1
XFILLER_12_235 VPWR VGND sg13g2_fill_2
XFILLER_12_246 VPWR VGND sg13g2_fill_2
XFILLER_5_946 VPWR VGND sg13g2_decap_8
XFILLER_48_699 VPWR VGND sg13g2_fill_1
XFILLER_15_1011 VPWR VGND sg13g2_decap_8
XFILLER_8_740 VPWR VGND sg13g2_fill_2
X_4520_ _1331_ _1304_ _1329_ VPWR VGND sg13g2_xnor2_1
XFILLER_7_250 VPWR VGND sg13g2_fill_1
Xhold217 mac2.products_ff\[151\] VPWR VGND net257 sg13g2_dlygate4sd3_1
X_4451_ _1264_ _1238_ _1262_ VPWR VGND sg13g2_xnor2_1
Xhold206 mac1.sum_lvl1_ff\[9\] VPWR VGND net246 sg13g2_dlygate4sd3_1
Xhold239 DP_2.matrix\[75\] VPWR VGND net279 sg13g2_dlygate4sd3_1
X_3402_ _2984_ net1015 net960 net956 net1018 VPWR VGND sg13g2_a22oi_1
Xhold228 _0032_ VPWR VGND net268 sg13g2_dlygate4sd3_1
X_6121_ net1067 VGND VPWR _0216_ DP_2.matrix\[76\] clknet_leaf_60_clk sg13g2_dfrbpq_1
X_4382_ _1163_ VPWR _1197_ VGND _1154_ _1164_ sg13g2_o21ai_1
X_3333_ _2920_ _2919_ _2921_ VPWR VGND sg13g2_nor2b_1
X_3264_ _2850_ _2852_ _2853_ _2854_ VPWR VGND sg13g2_nor3_1
X_6052_ net1093 VGND VPWR _0163_ DP_2.matrix\[8\] clknet_leaf_58_clk sg13g2_dfrbpq_2
XFILLER_22_1004 VPWR VGND sg13g2_decap_8
X_5003_ net808 net858 net811 _1790_ VPWR VGND net857 sg13g2_nand4_1
X_3195_ VGND VPWR _2783_ _2784_ _2787_ _2749_ sg13g2_a21oi_1
X_5905_ net897 net768 _2578_ VPWR VGND sg13g2_nor2_1
XFILLER_22_577 VPWR VGND sg13g2_fill_2
X_5836_ _2527_ _2493_ _2528_ _2529_ VPWR VGND sg13g2_a21o_1
X_5767_ _2443_ _2461_ _2462_ VPWR VGND sg13g2_nor2b_1
XFILLER_5_209 VPWR VGND sg13g2_fill_1
X_5698_ DP_1.I_range.out_data\[3\] _2600_ DP_1.I_range.out_data\[2\] _2601_ _2394_
+ VPWR VGND sg13g2_or4_1
X_4718_ _1518_ _1471_ _1517_ VPWR VGND sg13g2_xnor2_1
X_4649_ net845 net893 net849 _1451_ VPWR VGND net892 sg13g2_nand4_1
XFILLER_2_905 VPWR VGND sg13g2_decap_4
XFILLER_2_938 VPWR VGND sg13g2_decap_8
X_6319_ net1065 VGND VPWR net382 mac1.sum_lvl3_ff\[2\] clknet_leaf_64_clk sg13g2_dfrbpq_1
XFILLER_44_124 VPWR VGND sg13g2_fill_2
XFILLER_26_850 VPWR VGND sg13g2_decap_8
XFILLER_13_577 VPWR VGND sg13g2_decap_4
XFILLER_40_352 VPWR VGND sg13g2_fill_2
XFILLER_41_886 VPWR VGND sg13g2_decap_8
XFILLER_45_1015 VPWR VGND sg13g2_decap_8
XFILLER_49_964 VPWR VGND sg13g2_decap_8
XFILLER_35_113 VPWR VGND sg13g2_fill_1
X_3951_ _0783_ _0778_ _0782_ VPWR VGND sg13g2_xnor2_1
XFILLER_32_831 VPWR VGND sg13g2_decap_8
X_3882_ _0714_ _0715_ _0705_ _0716_ VPWR VGND sg13g2_nand3_1
X_5621_ _0054_ _2333_ net344 VPWR VGND sg13g2_xnor2_1
X_5552_ _2280_ mac2.sum_lvl3_ff\[21\] mac2.sum_lvl3_ff\[1\] VPWR VGND sg13g2_nand2_1
X_4503_ VGND VPWR _1253_ _1283_ _1315_ _1285_ sg13g2_a21oi_1
X_5483_ _0039_ _2223_ _2226_ VPWR VGND sg13g2_xnor2_1
X_4434_ _1248_ _1223_ _1247_ VPWR VGND sg13g2_nand2_1
X_4365_ _1133_ _1134_ _1178_ _1179_ _1181_ VPWR VGND sg13g2_and4_1
X_6104_ net1113 VGND VPWR _0205_ DP_2.matrix\[37\] clknet_leaf_49_clk sg13g2_dfrbpq_2
X_3316_ _2904_ net909 net1034 VPWR VGND sg13g2_nand2_1
XFILLER_6_1020 VPWR VGND sg13g2_decap_8
X_6035_ net1072 VGND VPWR _0076_ mac1.products_ff\[70\] clknet_leaf_62_clk sg13g2_dfrbpq_1
X_4296_ _1113_ net824 net877 VPWR VGND sg13g2_nand2_1
X_3247_ _2805_ VPWR _2837_ VGND _2752_ _2803_ sg13g2_o21ai_1
X_3178_ net922 net919 net964 net1033 _2770_ VPWR VGND sg13g2_and4_1
XFILLER_27_647 VPWR VGND sg13g2_fill_2
XFILLER_14_319 VPWR VGND sg13g2_decap_4
XFILLER_25_69 VPWR VGND sg13g2_fill_2
X_5819_ _2513_ _2510_ _2512_ VPWR VGND sg13g2_nand2b_1
XFILLER_10_514 VPWR VGND sg13g2_fill_1
XFILLER_9_4 VPWR VGND sg13g2_fill_1
XFILLER_2_757 VPWR VGND sg13g2_fill_2
XFILLER_1_256 VPWR VGND sg13g2_fill_1
XFILLER_1_289 VPWR VGND sg13g2_fill_1
XFILLER_46_901 VPWR VGND sg13g2_decap_8
XFILLER_18_603 VPWR VGND sg13g2_fill_1
XFILLER_46_978 VPWR VGND sg13g2_decap_8
XFILLER_17_146 VPWR VGND sg13g2_fill_1
XFILLER_45_488 VPWR VGND sg13g2_fill_1
XFILLER_12_1003 VPWR VGND sg13g2_decap_8
XFILLER_40_182 VPWR VGND sg13g2_fill_2
X_4150_ _0976_ net928 net1036 VPWR VGND sg13g2_nand2_1
X_3101_ _2691_ _2692_ _2694_ _2695_ VPWR VGND sg13g2_or3_1
X_4081_ _0908_ _0887_ _0910_ VPWR VGND sg13g2_xor2_1
X_3032_ _2629_ _2628_ _2616_ VPWR VGND sg13g2_nand2b_1
XFILLER_37_956 VPWR VGND sg13g2_decap_8
X_4983_ _1769_ _1770_ _1764_ _1771_ VPWR VGND sg13g2_nand3_1
X_3934_ _0737_ VPWR _0766_ VGND _0734_ _0738_ sg13g2_o21ai_1
X_3865_ _0682_ VPWR _0699_ VGND _0673_ _0683_ sg13g2_o21ai_1
X_5604_ net310 mac2.sum_lvl3_ff\[32\] _2321_ VPWR VGND sg13g2_xor2_1
X_3796_ _0633_ net1003 net934 VPWR VGND sg13g2_nand2_1
XFILLER_20_878 VPWR VGND sg13g2_fill_2
X_5535_ VPWR VGND _2267_ _2266_ _2258_ mac2.sum_lvl2_ff\[30\] _2268_ mac2.sum_lvl2_ff\[11\]
+ sg13g2_a221oi_1
X_5466_ _2214_ mac1.sum_lvl3_ff\[33\] mac1.sum_lvl3_ff\[13\] VPWR VGND sg13g2_nand2_1
X_4417_ _1230_ _1226_ _1231_ VPWR VGND sg13g2_xor2_1
X_5397_ _2160_ mac1.sum_lvl2_ff\[33\] mac1.sum_lvl2_ff\[14\] VPWR VGND sg13g2_nand2_1
X_4348_ VGND VPWR _1160_ _1161_ _1164_ _1155_ sg13g2_a21oi_1
XFILLER_28_901 VPWR VGND sg13g2_decap_8
X_4279_ _1096_ _1095_ _0134_ VPWR VGND sg13g2_xor2_1
X_6018_ net1070 VGND VPWR _0070_ mac1.products_ff\[1\] clknet_leaf_61_clk sg13g2_dfrbpq_1
XFILLER_43_904 VPWR VGND sg13g2_decap_8
XFILLER_15_617 VPWR VGND sg13g2_fill_2
XFILLER_28_978 VPWR VGND sg13g2_decap_8
XFILLER_42_414 VPWR VGND sg13g2_fill_1
XFILLER_42_425 VPWR VGND sg13g2_fill_1
XFILLER_11_823 VPWR VGND sg13g2_fill_2
XFILLER_35_1014 VPWR VGND sg13g2_decap_8
XFILLER_2_587 VPWR VGND sg13g2_decap_4
Xfanout891 net892 net891 VPWR VGND sg13g2_buf_8
XFILLER_18_400 VPWR VGND sg13g2_decap_4
Xfanout880 net334 net880 VPWR VGND sg13g2_buf_8
XFILLER_34_937 VPWR VGND sg13g2_decap_8
X_3650_ net953 net950 net1008 net1005 _0496_ VPWR VGND sg13g2_and4_1
X_3581_ _0429_ _0393_ _0427_ _0428_ VPWR VGND sg13g2_and3_1
X_5320_ VGND VPWR _2098_ _2097_ _2084_ sg13g2_or2_1
X_5251_ _2031_ net1024 net801 net852 net798 VPWR VGND sg13g2_a22oi_1
X_4202_ _1008_ VPWR _1022_ VGND _1006_ _1009_ sg13g2_o21ai_1
X_5182_ VGND VPWR _1929_ _1935_ _1964_ _1937_ sg13g2_a21oi_1
X_4133_ _0960_ _0933_ _0958_ VPWR VGND sg13g2_xnor2_1
X_4064_ _0893_ _0867_ _0891_ VPWR VGND sg13g2_xnor2_1
X_3015_ _2610_ _2611_ _2612_ _2613_ VPWR VGND sg13g2_nor3_1
XFILLER_37_720 VPWR VGND sg13g2_fill_1
XFILLER_37_764 VPWR VGND sg13g2_fill_2
X_4966_ _1755_ _1747_ _1754_ VPWR VGND sg13g2_nand2_1
X_4897_ _1692_ net835 net889 VPWR VGND sg13g2_nand2_1
X_3917_ VGND VPWR _0746_ _0747_ _0750_ _0741_ sg13g2_a21oi_1
X_3848_ VGND VPWR _0679_ _0680_ _0683_ _0674_ sg13g2_a21oi_1
XFILLER_20_675 VPWR VGND sg13g2_decap_4
X_3779_ _0619_ _0603_ _0620_ VPWR VGND sg13g2_xor2_1
X_5518_ _2254_ _2253_ _2252_ VPWR VGND sg13g2_nand2b_1
X_6498_ net1039 VGND VPWR net291 mac2.total_sum\[0\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_5449_ mac1.sum_lvl3_ff\[10\] net348 _2200_ VPWR VGND sg13g2_xor2_1
Xfanout1108 net1109 net1108 VPWR VGND sg13g2_buf_8
Xfanout1119 net1120 net1119 VPWR VGND sg13g2_buf_8
XFILLER_16_959 VPWR VGND sg13g2_decap_8
XFILLER_7_602 VPWR VGND sg13g2_fill_1
XFILLER_7_657 VPWR VGND sg13g2_fill_1
XFILLER_3_896 VPWR VGND sg13g2_fill_1
XFILLER_2_362 VPWR VGND sg13g2_fill_2
XFILLER_18_252 VPWR VGND sg13g2_fill_1
XFILLER_18_274 VPWR VGND sg13g2_fill_2
X_4820_ _1617_ _1605_ _1618_ VPWR VGND sg13g2_xor2_1
XFILLER_34_778 VPWR VGND sg13g2_fill_1
X_4751_ _1551_ _1549_ _1550_ VPWR VGND sg13g2_nand2_1
X_3702_ _0546_ net1037 net951 DP_1.matrix\[7\] DP_2.matrix\[5\] VPWR VGND sg13g2_a22oi_1
X_4682_ _1451_ VPWR _1483_ VGND _1449_ _1452_ sg13g2_o21ai_1
X_3633_ VGND VPWR _0444_ _0450_ _0479_ _0452_ sg13g2_a21oi_1
X_6421_ net1103 VGND VPWR net104 mac2.sum_lvl1_ff\[8\] clknet_leaf_43_clk sg13g2_dfrbpq_1
XFILLER_30_995 VPWR VGND sg13g2_decap_8
X_6352_ net1039 VGND VPWR net363 mac1.total_sum\[3\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3564_ _0372_ VPWR _0412_ VGND _0370_ _0373_ sg13g2_o21ai_1
X_5303_ VPWR _2081_ _2080_ VGND sg13g2_inv_1
X_3495_ _0343_ _0342_ _0333_ _0345_ VPWR VGND sg13g2_a21o_1
X_6283_ net1074 VGND VPWR net103 mac1.sum_lvl1_ff\[86\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_5234_ VGND VPWR _2015_ _2014_ _1969_ sg13g2_or2_1
X_5165_ net807 net804 net851 net1025 _1948_ VPWR VGND sg13g2_and4_1
X_4116_ VGND VPWR _0882_ _0911_ _0944_ _0913_ sg13g2_a21oi_1
X_5096_ _1880_ net868 net1021 VPWR VGND sg13g2_nand2_1
X_4047_ _0877_ _0852_ _0876_ VPWR VGND sg13g2_nand2_1
X_5998_ net823 _0254_ VPWR VGND sg13g2_buf_1
XFILLER_12_439 VPWR VGND sg13g2_fill_1
X_4949_ _1739_ net869 net805 VPWR VGND sg13g2_nand2_1
XFILLER_32_1006 VPWR VGND sg13g2_decap_8
XFILLER_47_336 VPWR VGND sg13g2_fill_2
XFILLER_47_314 VPWR VGND sg13g2_fill_2
XFILLER_35_509 VPWR VGND sg13g2_decap_8
XFILLER_43_542 VPWR VGND sg13g2_fill_2
XFILLER_15_233 VPWR VGND sg13g2_fill_1
XFILLER_7_498 VPWR VGND sg13g2_fill_2
XFILLER_48_1024 VPWR VGND sg13g2_decap_4
X_3280_ _2867_ _2869_ _2870_ VPWR VGND sg13g2_nor2_1
XFILLER_47_892 VPWR VGND sg13g2_decap_8
X_5921_ _2588_ _2526_ _2529_ VPWR VGND sg13g2_xnor2_1
XFILLER_19_594 VPWR VGND sg13g2_fill_2
XFILLER_34_520 VPWR VGND sg13g2_fill_1
X_5852_ _2540_ _2544_ _2545_ VPWR VGND sg13g2_nor2b_1
X_4803_ _1601_ _1560_ _1599_ VPWR VGND sg13g2_xnor2_1
X_5783_ DP_3.I_range.out_data\[6\] DP_3.I_range.out_data\[2\] _2603_ DP_3.I_range.out_data\[4\]
+ _2477_ VPWR VGND sg13g2_nor4_1
X_4734_ _1531_ _1532_ _1526_ _1534_ VPWR VGND sg13g2_nand3_1
X_4665_ _1433_ VPWR _1467_ VGND _1408_ _1434_ sg13g2_o21ai_1
X_3616_ net957 net955 net1005 net1038 _0463_ VPWR VGND sg13g2_and4_1
X_6404_ net1060 VGND VPWR _0157_ mac2.products_ff\[143\] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_4596_ _1398_ _1399_ _1393_ _1400_ VPWR VGND sg13g2_nand3_1
X_3547_ _0395_ net1020 net1032 VPWR VGND sg13g2_nand2_1
X_6335_ net1083 VGND VPWR net214 mac2.sum_lvl3_ff\[22\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_3478_ _0328_ net1017 net949 VPWR VGND sg13g2_nand2_1
X_6266_ net1059 VGND VPWR net194 mac2.sum_lvl2_ff\[51\] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_6197_ net1117 VGND VPWR net224 mac1.sum_lvl1_ff\[44\] clknet_leaf_50_clk sg13g2_dfrbpq_1
X_5217_ _1996_ _1998_ _1999_ VPWR VGND sg13g2_nor2_1
X_5148_ _1931_ net860 net793 VPWR VGND sg13g2_nand2_1
XFILLER_28_69 VPWR VGND sg13g2_fill_2
X_5079_ _1853_ _1861_ _1863_ _1864_ VPWR VGND sg13g2_or3_1
XFILLER_38_870 VPWR VGND sg13g2_decap_8
XFILLER_8_207 VPWR VGND sg13g2_fill_1
XFILLER_40_578 VPWR VGND sg13g2_decap_8
XFILLER_47_199 VPWR VGND sg13g2_fill_1
XFILLER_44_895 VPWR VGND sg13g2_decap_8
XFILLER_16_586 VPWR VGND sg13g2_fill_2
X_4450_ VGND VPWR _1263_ _1262_ _1238_ sg13g2_or2_1
Xhold207 mac2.sum_lvl2_ff\[46\] VPWR VGND net247 sg13g2_dlygate4sd3_1
X_3401_ net960 net1018 net956 net1015 _2983_ VPWR VGND sg13g2_and4_1
Xhold229 DP_2.matrix\[76\] VPWR VGND net269 sg13g2_dlygate4sd3_1
Xhold218 mac1.products_ff\[83\] VPWR VGND net258 sg13g2_dlygate4sd3_1
X_4381_ _1196_ _1186_ _1194_ VPWR VGND sg13g2_xnor2_1
X_3332_ VGND VPWR _2880_ _2892_ _2920_ _2879_ sg13g2_a21oi_1
X_6120_ net1074 VGND VPWR _0100_ mac1.products_ff\[151\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_3263_ _2853_ net965 net914 net968 net912 VPWR VGND sg13g2_a22oi_1
X_6051_ net1068 VGND VPWR _0162_ DP_1.matrix\[80\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_3194_ _2783_ _2784_ _2749_ _2786_ VPWR VGND sg13g2_nand3_1
XFILLER_38_111 VPWR VGND sg13g2_fill_2
X_5002_ net811 net808 net858 net857 _1789_ VPWR VGND sg13g2_and4_1
XFILLER_39_623 VPWR VGND sg13g2_fill_2
XFILLER_38_155 VPWR VGND sg13g2_fill_1
XFILLER_39_678 VPWR VGND sg13g2_decap_4
X_5904_ VGND VPWR net768 _2577_ _0222_ _2576_ sg13g2_a21oi_1
XFILLER_41_309 VPWR VGND sg13g2_fill_2
XFILLER_35_895 VPWR VGND sg13g2_decap_8
X_5835_ net843 _2493_ _2528_ VPWR VGND sg13g2_nor2_1
XFILLER_10_718 VPWR VGND sg13g2_fill_1
X_5766_ _2456_ _2460_ _2461_ VPWR VGND sg13g2_nor2b_1
X_5697_ net443 _2600_ _2391_ _2392_ _2393_ VPWR VGND sg13g2_nor4_1
X_4717_ _1517_ _1508_ _1515_ VPWR VGND sg13g2_xnor2_1
X_4648_ net849 net846 net894 net892 _1450_ VPWR VGND sg13g2_and4_1
XFILLER_2_917 VPWR VGND sg13g2_decap_8
X_4579_ _1384_ _1376_ _1383_ VPWR VGND sg13g2_nand2_1
X_6318_ net1064 VGND VPWR net357 mac1.sum_lvl3_ff\[1\] clknet_leaf_64_clk sg13g2_dfrbpq_2
X_6249_ net1051 VGND VPWR net180 mac1.sum_lvl2_ff\[50\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_26_840 VPWR VGND sg13g2_fill_1
XFILLER_13_556 VPWR VGND sg13g2_fill_2
XFILLER_41_865 VPWR VGND sg13g2_decap_8
XFILLER_5_799 VPWR VGND sg13g2_fill_2
XFILLER_49_943 VPWR VGND sg13g2_decap_8
XFILLER_1_994 VPWR VGND sg13g2_decap_8
Xhold90 mac1.sum_lvl1_ff\[2\] VPWR VGND net130 sg13g2_dlygate4sd3_1
X_3950_ _0782_ _0735_ _0780_ VPWR VGND sg13g2_xnor2_1
XFILLER_16_361 VPWR VGND sg13g2_fill_1
X_3881_ _0712_ _0711_ _0706_ _0715_ VPWR VGND sg13g2_a21o_1
XFILLER_31_342 VPWR VGND sg13g2_fill_1
X_5620_ _2334_ mac2.sum_lvl3_ff\[35\] net343 VPWR VGND sg13g2_xnor2_1
XFILLER_32_887 VPWR VGND sg13g2_decap_8
X_5551_ _2279_ net449 net290 VPWR VGND sg13g2_nand2_1
XFILLER_8_560 VPWR VGND sg13g2_fill_2
X_4502_ VGND VPWR _1252_ _1283_ _1314_ _1285_ sg13g2_a21oi_1
X_5482_ mac2.sum_lvl2_ff\[1\] mac2.sum_lvl2_ff\[20\] _2226_ VPWR VGND sg13g2_xor2_1
X_4433_ _1246_ _1234_ _1247_ VPWR VGND sg13g2_xor2_1
X_4364_ _1180_ _1178_ _1179_ VPWR VGND sg13g2_nand2_1
X_6103_ net1113 VGND VPWR _0204_ DP_2.matrix\[36\] clknet_leaf_49_clk sg13g2_dfrbpq_2
X_3315_ _2903_ net1033 net912 net966 net910 VPWR VGND sg13g2_a22oi_1
X_4295_ _1080_ VPWR _1112_ VGND _1078_ _1081_ sg13g2_o21ai_1
X_6034_ net1070 VGND VPWR net433 mac1.products_ff\[69\] clknet_leaf_62_clk sg13g2_dfrbpq_1
X_3246_ _2825_ VPWR _2836_ VGND _2809_ _2826_ sg13g2_o21ai_1
X_3177_ _2769_ net915 net967 VPWR VGND sg13g2_nand2_1
XFILLER_39_464 VPWR VGND sg13g2_fill_1
XFILLER_26_114 VPWR VGND sg13g2_decap_8
XFILLER_23_832 VPWR VGND sg13g2_decap_8
XFILLER_41_117 VPWR VGND sg13g2_decap_8
X_5818_ _2512_ _2511_ net778 net776 net275 VPWR VGND sg13g2_a22oi_1
X_5749_ net952 net934 net788 _2444_ VPWR VGND sg13g2_mux2_1
XFILLER_45_401 VPWR VGND sg13g2_fill_2
XFILLER_46_957 VPWR VGND sg13g2_decap_8
XFILLER_45_445 VPWR VGND sg13g2_fill_2
XFILLER_33_629 VPWR VGND sg13g2_fill_1
XFILLER_9_324 VPWR VGND sg13g2_fill_2
XFILLER_41_695 VPWR VGND sg13g2_fill_2
XFILLER_5_585 VPWR VGND sg13g2_fill_1
X_3100_ _2694_ net967 net921 net969 net918 VPWR VGND sg13g2_a22oi_1
XFILLER_49_740 VPWR VGND sg13g2_fill_2
X_4080_ _0908_ _0887_ _0909_ VPWR VGND sg13g2_nor2b_1
X_3031_ _2627_ _2617_ _2628_ VPWR VGND sg13g2_xor2_1
XFILLER_37_935 VPWR VGND sg13g2_decap_8
XFILLER_24_629 VPWR VGND sg13g2_fill_1
X_4982_ _1765_ VPWR _1770_ VGND _1766_ _1768_ sg13g2_o21ai_1
X_3933_ _0754_ VPWR _0765_ VGND _0732_ _0755_ sg13g2_o21ai_1
X_3864_ _0696_ _0695_ _0698_ VPWR VGND sg13g2_xor2_1
X_5603_ mac2.sum_lvl3_ff\[32\] net310 _2320_ VPWR VGND sg13g2_nor2_1
X_3795_ _0631_ _0624_ _0076_ VPWR VGND sg13g2_xor2_1
X_5534_ _2257_ _2261_ _2267_ VPWR VGND sg13g2_nor2_1
X_5465_ _2213_ _2206_ _2211_ VPWR VGND sg13g2_nand2_1
X_4416_ _1230_ _1189_ _1228_ VPWR VGND sg13g2_xnor2_1
X_5396_ VGND VPWR _2155_ _2157_ _2159_ _2156_ sg13g2_a21oi_1
X_4347_ _1160_ _1161_ _1155_ _1163_ VPWR VGND sg13g2_nand3_1
X_4278_ _1062_ VPWR _1096_ VGND _1037_ _1063_ sg13g2_o21ai_1
XFILLER_46_209 VPWR VGND sg13g2_fill_1
X_3229_ _2820_ net1033 net918 net964 net915 VPWR VGND sg13g2_a22oi_1
X_6017_ net1066 VGND VPWR _0069_ mac1.products_ff\[0\] clknet_leaf_63_clk sg13g2_dfrbpq_1
XFILLER_28_957 VPWR VGND sg13g2_decap_8
XFILLER_36_36 VPWR VGND sg13g2_fill_2
XFILLER_7_2 VPWR VGND sg13g2_fill_1
Xhold390 _0063_ VPWR VGND net430 sg13g2_dlygate4sd3_1
Xfanout870 net871 net870 VPWR VGND sg13g2_buf_8
Xfanout892 net428 net892 VPWR VGND sg13g2_buf_8
Xfanout881 DP_3.matrix\[39\] net881 VPWR VGND sg13g2_buf_8
XFILLER_18_445 VPWR VGND sg13g2_fill_1
XFILLER_19_979 VPWR VGND sg13g2_decap_8
XFILLER_34_916 VPWR VGND sg13g2_decap_8
XFILLER_42_982 VPWR VGND sg13g2_decap_8
XFILLER_14_684 VPWR VGND sg13g2_decap_4
XFILLER_41_470 VPWR VGND sg13g2_fill_1
XFILLER_41_492 VPWR VGND sg13g2_fill_2
XFILLER_9_154 VPWR VGND sg13g2_fill_2
X_3580_ _0404_ VPWR _0428_ VGND _0424_ _0426_ sg13g2_o21ai_1
X_5250_ _2017_ _2012_ _2019_ _2030_ VPWR VGND sg13g2_a21o_1
X_4201_ VPWR _1021_ _1020_ VGND sg13g2_inv_1
X_5181_ _1963_ _1924_ _0159_ VPWR VGND sg13g2_xor2_1
X_4132_ _0959_ _0958_ _0933_ VPWR VGND sg13g2_nand2b_1
X_4063_ VGND VPWR _0892_ _0891_ _0867_ sg13g2_or2_1
XFILLER_3_1024 VPWR VGND sg13g2_decap_4
X_3014_ _2612_ net978 net923 net917 net981 VPWR VGND sg13g2_a22oi_1
XFILLER_25_949 VPWR VGND sg13g2_decap_8
X_4965_ _1752_ _1753_ _1754_ VPWR VGND sg13g2_nor2b_1
X_3916_ _0746_ _0747_ _0741_ _0749_ VPWR VGND sg13g2_nand3_1
XFILLER_33_982 VPWR VGND sg13g2_decap_8
X_4896_ _1691_ net889 net833 VPWR VGND sg13g2_nand2_1
X_3847_ _0679_ _0680_ _0674_ _0682_ VPWR VGND sg13g2_nand3_1
X_3778_ _0619_ net1005 DP_2.matrix\[8\] VPWR VGND sg13g2_nand2_1
X_5517_ VGND VPWR _2253_ net545 mac2.sum_lvl2_ff\[28\] sg13g2_or2_1
X_6497_ net1059 VGND VPWR _0038_ mac2.sum_lvl3_ff\[15\] clknet_leaf_24_clk sg13g2_dfrbpq_1
X_5448_ _2199_ net348 net364 VPWR VGND sg13g2_nand2_1
Xfanout1109 net1118 net1109 VPWR VGND sg13g2_buf_8
X_5379_ _0001_ _2143_ _2144_ VPWR VGND sg13g2_xnor2_1
XFILLER_16_938 VPWR VGND sg13g2_decap_8
XFILLER_31_919 VPWR VGND sg13g2_decap_8
XFILLER_24_982 VPWR VGND sg13g2_decap_8
XFILLER_8_29 VPWR VGND sg13g2_fill_1
XFILLER_33_234 VPWR VGND sg13g2_fill_1
XFILLER_18_1010 VPWR VGND sg13g2_decap_8
XFILLER_14_481 VPWR VGND sg13g2_fill_1
X_4750_ _1547_ _1546_ _1548_ _1550_ VPWR VGND sg13g2_a21o_1
X_3701_ _0532_ _0527_ _0534_ _0545_ VPWR VGND sg13g2_a21o_1
XFILLER_30_974 VPWR VGND sg13g2_decap_8
X_4681_ _1482_ _1476_ _1481_ VPWR VGND sg13g2_xnor2_1
X_3632_ _0478_ _0439_ _0115_ VPWR VGND sg13g2_xor2_1
X_6420_ net1104 VGND VPWR net234 mac2.sum_lvl1_ff\[7\] clknet_leaf_43_clk sg13g2_dfrbpq_1
X_6351_ net1039 VGND VPWR net456 mac1.total_sum\[2\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_5302_ _2080_ _2056_ _2078_ VPWR VGND sg13g2_nand2_1
X_3563_ _0411_ _0406_ _0410_ VPWR VGND sg13g2_xnor2_1
X_3494_ _0342_ _0343_ _0333_ _0344_ VPWR VGND sg13g2_nand3_1
X_6282_ net1068 VGND VPWR net212 mac1.sum_lvl1_ff\[85\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_5233_ _2014_ net856 net795 VPWR VGND sg13g2_nand2_1
X_5164_ _1947_ net804 net1025 VPWR VGND sg13g2_nand2_1
X_4115_ VGND VPWR _0881_ _0911_ _0943_ _0913_ sg13g2_a21oi_1
XFILLER_29_529 VPWR VGND sg13g2_decap_8
X_5095_ _1850_ VPWR _1879_ VGND _1847_ _1851_ sg13g2_o21ai_1
X_4046_ _0875_ _0863_ _0876_ VPWR VGND sg13g2_xor2_1
XFILLER_25_724 VPWR VGND sg13g2_fill_1
X_5997_ net826 _0253_ VPWR VGND sg13g2_buf_1
X_4948_ _1737_ net294 _0090_ VPWR VGND sg13g2_nor2_1
XFILLER_40_749 VPWR VGND sg13g2_decap_8
X_4879_ VGND VPWR _1675_ _1674_ _1662_ sg13g2_or2_1
XFILLER_21_985 VPWR VGND sg13g2_decap_8
XFILLER_0_856 VPWR VGND sg13g2_fill_1
XFILLER_12_941 VPWR VGND sg13g2_decap_4
XFILLER_8_934 VPWR VGND sg13g2_fill_2
XFILLER_12_996 VPWR VGND sg13g2_decap_8
XFILLER_7_455 VPWR VGND sg13g2_fill_1
XFILLER_23_92 VPWR VGND sg13g2_fill_2
XFILLER_48_1003 VPWR VGND sg13g2_decap_8
XFILLER_38_304 VPWR VGND sg13g2_fill_2
XFILLER_39_805 VPWR VGND sg13g2_fill_2
XFILLER_39_849 VPWR VGND sg13g2_decap_8
X_5920_ net843 net768 _2587_ VPWR VGND sg13g2_nor2_1
X_5851_ _2541_ VPWR _2544_ VGND _2542_ _2543_ sg13g2_o21ai_1
XFILLER_34_576 VPWR VGND sg13g2_fill_2
X_4802_ VGND VPWR _1600_ _1598_ _1561_ sg13g2_or2_1
X_5782_ DP_3.Q_range.out_data\[2\] _2604_ DP_3.Q_range.out_data\[4\] DP_3.Q_range.out_data\[6\]
+ _2476_ VPWR VGND sg13g2_nor4_1
X_4733_ _1533_ _1526_ _1531_ _1532_ VPWR VGND sg13g2_and3_1
X_6403_ net1061 VGND VPWR _0156_ mac2.products_ff\[142\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_4664_ _1466_ _1436_ _1464_ VPWR VGND sg13g2_xnor2_1
X_3615_ _0462_ net955 net1038 VPWR VGND sg13g2_nand2_1
X_4595_ _1394_ VPWR _1399_ VGND _1395_ _1397_ sg13g2_o21ai_1
X_3546_ _0365_ VPWR _0394_ VGND _0362_ _0366_ sg13g2_o21ai_1
X_6334_ net1083 VGND VPWR net230 mac2.sum_lvl3_ff\[21\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_6265_ net1055 VGND VPWR net255 mac2.sum_lvl2_ff\[50\] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_3477_ _0310_ VPWR _0327_ VGND _0301_ _0311_ sg13g2_o21ai_1
X_5216_ VGND VPWR _1997_ _1998_ _1963_ _1923_ sg13g2_a21oi_2
X_6196_ net1108 VGND VPWR net221 mac1.sum_lvl1_ff\[43\] clknet_leaf_51_clk sg13g2_dfrbpq_1
X_5147_ _1930_ net866 net1021 VPWR VGND sg13g2_nand2_1
XFILLER_28_59 VPWR VGND sg13g2_fill_1
X_5078_ VGND VPWR _1859_ _1860_ _1863_ _1854_ sg13g2_a21oi_1
X_4029_ _0859_ _0818_ _0857_ VPWR VGND sg13g2_xnor2_1
XFILLER_12_237 VPWR VGND sg13g2_fill_1
XFILLER_16_510 VPWR VGND sg13g2_fill_1
XFILLER_16_521 VPWR VGND sg13g2_decap_8
XFILLER_44_874 VPWR VGND sg13g2_decap_8
XFILLER_8_742 VPWR VGND sg13g2_fill_1
XFILLER_11_292 VPWR VGND sg13g2_fill_2
Xhold208 mac1.products_ff\[72\] VPWR VGND net248 sg13g2_dlygate4sd3_1
Xhold219 mac1.sum_lvl1_ff\[73\] VPWR VGND net259 sg13g2_dlygate4sd3_1
X_3400_ _2982_ net1019 net954 VPWR VGND sg13g2_nand2_1
X_4380_ _1186_ _1194_ _1195_ VPWR VGND sg13g2_nor2_1
X_3331_ _2917_ _2906_ _2919_ VPWR VGND sg13g2_xor2_1
X_3262_ net914 net911 net968 net965 _2852_ VPWR VGND sg13g2_and4_1
X_6050_ net1111 VGND VPWR _0161_ DP_1.matrix\[44\] clknet_leaf_46_clk sg13g2_dfrbpq_2
X_3193_ _2785_ _2749_ _2783_ _2784_ VPWR VGND sg13g2_and3_1
X_5001_ _1788_ net804 net861 VPWR VGND sg13g2_nand2_1
XFILLER_38_178 VPWR VGND sg13g2_fill_2
XFILLER_35_874 VPWR VGND sg13g2_decap_8
X_5903_ _2499_ _2497_ _2577_ VPWR VGND sg13g2_xor2_1
X_5834_ _2527_ net786 net810 net777 net825 VPWR VGND sg13g2_a22oi_1
X_5765_ _2457_ VPWR _2460_ VGND _2458_ _2459_ sg13g2_o21ai_1
XFILLER_22_579 VPWR VGND sg13g2_fill_1
X_5696_ DP_1.I_range.out_data\[2\] DP_1.Q_range.out_data\[2\] DP_1.I_range.out_data\[6\]
+ _2601_ _2392_ VPWR VGND sg13g2_or4_1
X_4716_ _1516_ _1508_ _1515_ VPWR VGND sg13g2_nand2_1
X_4647_ _1449_ net841 net896 VPWR VGND sg13g2_nand2_1
X_6317_ net1049 VGND VPWR net287 mac1.sum_lvl3_ff\[0\] clknet_leaf_67_clk sg13g2_dfrbpq_1
X_4578_ _1381_ _1382_ _1383_ VPWR VGND sg13g2_nor2b_1
X_3529_ VGND VPWR _0374_ _0375_ _0378_ _0369_ sg13g2_a21oi_1
X_6248_ net1046 VGND VPWR net167 mac1.sum_lvl2_ff\[49\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_6179_ net1123 VGND VPWR _0258_ DP_4.matrix\[42\] clknet_leaf_34_clk sg13g2_dfrbpq_1
XFILLER_26_896 VPWR VGND sg13g2_decap_8
XFILLER_38_1024 VPWR VGND sg13g2_decap_4
XFILLER_41_844 VPWR VGND sg13g2_decap_8
XFILLER_4_211 VPWR VGND sg13g2_fill_1
XFILLER_49_922 VPWR VGND sg13g2_decap_8
XFILLER_1_973 VPWR VGND sg13g2_decap_8
XFILLER_48_443 VPWR VGND sg13g2_fill_2
XFILLER_29_80 VPWR VGND sg13g2_fill_2
XFILLER_49_999 VPWR VGND sg13g2_decap_8
Xhold80 mac1.sum_lvl1_ff\[3\] VPWR VGND net120 sg13g2_dlygate4sd3_1
XFILLER_29_91 VPWR VGND sg13g2_fill_2
Xhold91 mac2.sum_lvl2_ff\[38\] VPWR VGND net131 sg13g2_dlygate4sd3_1
X_3880_ _0711_ _0712_ _0706_ _0714_ VPWR VGND sg13g2_nand3_1
XFILLER_32_866 VPWR VGND sg13g2_decap_8
X_5550_ net267 mac2.sum_lvl2_ff\[19\] _0032_ VPWR VGND sg13g2_xor2_1
X_4501_ _1311_ _1310_ _1313_ VPWR VGND sg13g2_xor2_1
X_5481_ mac2.sum_lvl2_ff\[20\] mac2.sum_lvl2_ff\[1\] _2225_ VPWR VGND sg13g2_nor2_1
X_4432_ _1244_ _1235_ _1246_ VPWR VGND sg13g2_xor2_1
X_4363_ _1176_ _1175_ _1177_ _1179_ VPWR VGND sg13g2_a21o_1
X_3314_ _2889_ _2883_ _2891_ _2902_ VPWR VGND sg13g2_a21o_1
X_6102_ net1047 VGND VPWR _0104_ mac1.products_ff\[145\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_4294_ _1111_ _1105_ _1110_ VPWR VGND sg13g2_xnor2_1
X_6033_ net1066 VGND VPWR _0074_ mac1.products_ff\[68\] clknet_leaf_63_clk sg13g2_dfrbpq_1
X_3245_ VGND VPWR _2800_ _2806_ _2835_ _2808_ sg13g2_a21oi_1
X_3176_ _2728_ VPWR _2768_ VGND _2726_ _2729_ sg13g2_o21ai_1
XFILLER_39_498 VPWR VGND sg13g2_fill_2
XFILLER_25_27 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_61_clk clknet_4_8_0_clk clknet_leaf_61_clk VPWR VGND sg13g2_buf_8
X_5817_ net872 net890 net787 _2511_ VPWR VGND sg13g2_mux2_1
X_5748_ _2443_ _2442_ net784 net780 net910 VPWR VGND sg13g2_a22oi_1
X_5679_ VPWR VGND _2379_ _2378_ _2370_ mac1.total_sum\[11\] _2380_ mac2.total_sum\[11\]
+ sg13g2_a221oi_1
XFILLER_2_759 VPWR VGND sg13g2_fill_1
XFILLER_46_936 VPWR VGND sg13g2_decap_8
XFILLER_26_660 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_52_clk clknet_4_10_0_clk clknet_leaf_52_clk VPWR VGND sg13g2_buf_8
XFILLER_14_899 VPWR VGND sg13g2_fill_1
XFILLER_40_184 VPWR VGND sg13g2_fill_1
XFILLER_31_81 VPWR VGND sg13g2_fill_1
XFILLER_0_280 VPWR VGND sg13g2_decap_8
X_3030_ _2627_ _2618_ _2625_ VPWR VGND sg13g2_xnor2_1
XFILLER_37_914 VPWR VGND sg13g2_decap_8
XFILLER_45_980 VPWR VGND sg13g2_decap_8
X_4981_ _1765_ _1766_ _1768_ _1769_ VPWR VGND sg13g2_or3_1
X_3932_ _0763_ _0762_ _0124_ VPWR VGND sg13g2_xor2_1
Xclkbuf_leaf_43_clk clknet_4_13_0_clk clknet_leaf_43_clk VPWR VGND sg13g2_buf_8
X_3863_ _0697_ _0695_ _0696_ VPWR VGND sg13g2_nand2b_1
XFILLER_20_836 VPWR VGND sg13g2_decap_4
X_5602_ _2319_ mac2.sum_lvl3_ff\[32\] net310 VPWR VGND sg13g2_nand2_1
X_3794_ _0632_ _0624_ _0631_ VPWR VGND sg13g2_nand2_2
X_5533_ _2255_ _2260_ _2266_ VPWR VGND sg13g2_nor2_1
X_5464_ _2211_ _2212_ _0019_ VPWR VGND sg13g2_and2_1
X_5395_ _0004_ _2155_ _2158_ VPWR VGND sg13g2_xnor2_1
X_4415_ VGND VPWR _1229_ _1227_ _1190_ sg13g2_or2_1
X_4346_ _1162_ _1155_ _1160_ _1161_ VPWR VGND sg13g2_and3_1
X_4277_ _1095_ _1065_ _1093_ VPWR VGND sg13g2_xnor2_1
X_3228_ net918 net915 net964 net1033 _2819_ VPWR VGND sg13g2_and4_1
X_6016_ net1056 VGND VPWR net12 DP_3.Q_range.out_data\[6\] clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_39_240 VPWR VGND sg13g2_fill_1
X_3159_ _2751_ net985 net1030 VPWR VGND sg13g2_nand2_1
XFILLER_28_936 VPWR VGND sg13g2_decap_8
XFILLER_43_939 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_34_clk clknet_4_15_0_clk clknet_leaf_34_clk VPWR VGND sg13g2_buf_8
XFILLER_11_825 VPWR VGND sg13g2_fill_1
XFILLER_10_302 VPWR VGND sg13g2_fill_2
Xhold380 _2186_ VPWR VGND net420 sg13g2_dlygate4sd3_1
Xhold391 DP_2.matrix\[37\] VPWR VGND net431 sg13g2_dlygate4sd3_1
Xfanout860 net862 net860 VPWR VGND sg13g2_buf_8
Xfanout871 net872 net871 VPWR VGND sg13g2_buf_8
Xfanout893 net894 net893 VPWR VGND sg13g2_buf_8
Xfanout882 net331 net882 VPWR VGND sg13g2_buf_8
XFILLER_19_958 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_25_clk clknet_4_7_0_clk clknet_leaf_25_clk VPWR VGND sg13g2_buf_8
XFILLER_42_961 VPWR VGND sg13g2_decap_8
XFILLER_14_663 VPWR VGND sg13g2_fill_1
XFILLER_13_195 VPWR VGND sg13g2_decap_8
XFILLER_10_880 VPWR VGND sg13g2_fill_1
X_4200_ _1017_ _1019_ _1020_ VPWR VGND sg13g2_nor2_1
X_5180_ _1961_ _1962_ _1963_ VPWR VGND sg13g2_nor2b_1
X_4131_ _0956_ _0918_ _0958_ VPWR VGND sg13g2_xor2_1
XFILLER_3_1003 VPWR VGND sg13g2_decap_8
X_4062_ _0891_ net934 net1035 VPWR VGND sg13g2_nand2_1
X_3013_ net923 net981 net917 net978 _2611_ VPWR VGND sg13g2_and4_1
XFILLER_25_928 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_16_clk clknet_4_6_0_clk clknet_leaf_16_clk VPWR VGND sg13g2_buf_8
X_4964_ _1748_ VPWR _1753_ VGND _1749_ _1751_ sg13g2_o21ai_1
X_3915_ _0748_ _0741_ _0746_ _0747_ VPWR VGND sg13g2_and3_1
XFILLER_33_961 VPWR VGND sg13g2_decap_8
X_4895_ _1690_ net893 net1023 VPWR VGND sg13g2_nand2_1
X_3846_ _0681_ _0674_ _0679_ _0680_ VPWR VGND sg13g2_and3_1
X_3777_ _0606_ VPWR _0618_ VGND _0578_ _0604_ sg13g2_o21ai_1
X_6496_ net1059 VGND VPWR _0037_ mac2.sum_lvl3_ff\[14\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_5516_ mac2.sum_lvl2_ff\[28\] mac2.sum_lvl2_ff\[9\] _2252_ VPWR VGND sg13g2_and2_1
X_5447_ _2198_ _2195_ _2197_ VPWR VGND sg13g2_nand2_1
X_5378_ _2145_ _2142_ _2144_ VPWR VGND sg13g2_nand2_1
X_4329_ _1145_ _1137_ _1144_ VPWR VGND sg13g2_nand2_1
XFILLER_28_700 VPWR VGND sg13g2_fill_2
XFILLER_28_788 VPWR VGND sg13g2_fill_2
XFILLER_24_961 VPWR VGND sg13g2_decap_8
XFILLER_30_408 VPWR VGND sg13g2_fill_2
XFILLER_12_61 VPWR VGND sg13g2_fill_2
XFILLER_3_810 VPWR VGND sg13g2_fill_2
XFILLER_18_276 VPWR VGND sg13g2_fill_1
XFILLER_15_983 VPWR VGND sg13g2_decap_8
X_3700_ _0107_ _0543_ _0544_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_953 VPWR VGND sg13g2_decap_8
X_4680_ _1481_ _1443_ _1478_ VPWR VGND sg13g2_xnor2_1
X_3631_ _0476_ _0477_ _0478_ VPWR VGND sg13g2_nor2b_1
X_6350_ net1040 VGND VPWR net289 mac1.total_sum\[1\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3562_ _0410_ _0363_ _0408_ VPWR VGND sg13g2_xnor2_1
X_5301_ _0153_ _2078_ _2079_ VPWR VGND sg13g2_xnor2_1
X_3493_ _0340_ _0339_ _0334_ _0343_ VPWR VGND sg13g2_a21o_1
X_6281_ net1051 VGND VPWR net238 mac1.sum_lvl1_ff\[84\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_5232_ _2013_ net860 net1021 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_5_clk clknet_4_1_0_clk clknet_leaf_5_clk VPWR VGND sg13g2_buf_8
X_5163_ _1900_ VPWR _1946_ VGND _1898_ _1901_ sg13g2_o21ai_1
X_4114_ _0940_ _0939_ _0942_ VPWR VGND sg13g2_xor2_1
XFILLER_25_1026 VPWR VGND sg13g2_fill_2
X_5094_ _1867_ VPWR _1878_ VGND _1845_ _1868_ sg13g2_o21ai_1
X_4045_ _0873_ _0864_ _0875_ VPWR VGND sg13g2_xor2_1
X_5996_ net829 _0252_ VPWR VGND sg13g2_buf_1
X_4947_ _1738_ net809 net869 net293 net812 VPWR VGND sg13g2_a22oi_1
X_4878_ _1672_ _1663_ _1674_ VPWR VGND sg13g2_xor2_1
XFILLER_21_964 VPWR VGND sg13g2_decap_8
X_3829_ _0663_ _0662_ _0665_ VPWR VGND sg13g2_xor2_1
X_6479_ net1127 VGND VPWR net123 mac2.sum_lvl2_ff\[32\] clknet_leaf_37_clk sg13g2_dfrbpq_1
XFILLER_0_846 VPWR VGND sg13g2_fill_1
XFILLER_47_316 VPWR VGND sg13g2_fill_1
XFILLER_15_202 VPWR VGND sg13g2_fill_2
XFILLER_8_924 VPWR VGND sg13g2_fill_2
XFILLER_12_975 VPWR VGND sg13g2_decap_8
XFILLER_23_60 VPWR VGND sg13g2_fill_1
XFILLER_39_828 VPWR VGND sg13g2_decap_8
XFILLER_0_1017 VPWR VGND sg13g2_decap_8
XFILLER_46_382 VPWR VGND sg13g2_fill_2
XFILLER_46_371 VPWR VGND sg13g2_fill_1
XFILLER_0_1028 VPWR VGND sg13g2_fill_1
X_5850_ net778 VPWR _2543_ VGND net835 _2473_ sg13g2_o21ai_1
X_4801_ _1599_ net896 net835 VPWR VGND sg13g2_nand2_1
X_5781_ VGND VPWR _2607_ net785 _2475_ _2474_ sg13g2_a21oi_1
XFILLER_22_739 VPWR VGND sg13g2_fill_2
X_4732_ _1527_ VPWR _1532_ VGND _1528_ _1530_ sg13g2_o21ai_1
X_4663_ _1464_ _1436_ _1465_ VPWR VGND sg13g2_nor2b_1
X_3614_ _0415_ VPWR _0461_ VGND _0413_ _0416_ sg13g2_o21ai_1
X_6402_ net1062 VGND VPWR _0149_ mac2.products_ff\[141\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_4594_ _1394_ _1395_ _1397_ _1398_ VPWR VGND sg13g2_or3_1
X_3545_ _0382_ VPWR _0393_ VGND _0360_ _0383_ sg13g2_o21ai_1
XFILLER_7_990 VPWR VGND sg13g2_decap_8
X_6333_ net1083 VGND VPWR net131 mac2.sum_lvl3_ff\[20\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_3476_ _0324_ _0323_ _0326_ VPWR VGND sg13g2_xor2_1
X_6264_ net1054 VGND VPWR net115 mac2.sum_lvl2_ff\[49\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_5215_ VGND VPWR _1920_ _1962_ _1997_ _1961_ sg13g2_a21oi_1
X_6195_ net1109 VGND VPWR net91 mac1.sum_lvl1_ff\[42\] clknet_leaf_51_clk sg13g2_dfrbpq_1
Xclkbuf_4_15_0_clk clknet_0_clk clknet_4_15_0_clk VPWR VGND sg13g2_buf_8
X_5146_ _1894_ VPWR _1929_ VGND _1891_ _1895_ sg13g2_o21ai_1
X_5077_ _1859_ _1860_ _1854_ _1862_ VPWR VGND sg13g2_nand3_1
X_4028_ VGND VPWR _0858_ _0856_ _0819_ sg13g2_or2_1
XFILLER_25_522 VPWR VGND sg13g2_fill_2
X_5979_ net906 _0219_ VPWR VGND sg13g2_buf_1
XFILLER_29_883 VPWR VGND sg13g2_decap_8
XFILLER_43_352 VPWR VGND sg13g2_fill_2
XFILLER_16_588 VPWR VGND sg13g2_fill_1
XFILLER_31_525 VPWR VGND sg13g2_decap_4
XFILLER_15_1025 VPWR VGND sg13g2_decap_4
Xhold209 mac1.sum_lvl1_ff\[76\] VPWR VGND net249 sg13g2_dlygate4sd3_1
X_3330_ VGND VPWR _2918_ _2917_ _2906_ sg13g2_or2_1
XFILLER_4_993 VPWR VGND sg13g2_decap_8
X_3261_ _2851_ net912 net965 VPWR VGND sg13g2_nand2_1
X_5000_ _1767_ VPWR _1787_ VGND _1765_ _1768_ sg13g2_o21ai_1
X_3192_ _2760_ VPWR _2784_ VGND _2780_ _2782_ sg13g2_o21ai_1
XFILLER_39_625 VPWR VGND sg13g2_fill_1
XFILLER_22_1018 VPWR VGND sg13g2_decap_8
XFILLER_35_853 VPWR VGND sg13g2_decap_8
X_5902_ net899 net768 _2576_ VPWR VGND sg13g2_nor2_1
XFILLER_34_385 VPWR VGND sg13g2_fill_2
X_5833_ _2526_ _2525_ net777 net775 net282 VPWR VGND sg13g2_a22oi_1
XFILLER_22_536 VPWR VGND sg13g2_fill_2
X_5764_ net783 VPWR _2459_ VGND net951 net788 sg13g2_o21ai_1
X_5695_ DP_1.I_range.out_data\[4\] _2602_ DP_1.Q_range.out_data\[4\] DP_1.Q_range.out_data\[6\]
+ _2391_ VPWR VGND sg13g2_or4_1
XFILLER_30_591 VPWR VGND sg13g2_fill_2
X_4715_ _1513_ _1509_ _1515_ VPWR VGND sg13g2_xor2_1
X_4646_ _1419_ VPWR _1448_ VGND _1417_ _1420_ sg13g2_o21ai_1
X_4577_ _1377_ VPWR _1382_ VGND _1378_ _1380_ sg13g2_o21ai_1
X_6316_ net1093 VGND VPWR net185 mac1.sum_lvl3_ff\[35\] clknet_leaf_59_clk sg13g2_dfrbpq_1
X_3528_ _0374_ _0375_ _0369_ _0377_ VPWR VGND sg13g2_nand3_1
X_3459_ _0307_ _0308_ _0302_ _0310_ VPWR VGND sg13g2_nand3_1
X_6247_ net1046 VGND VPWR net205 mac1.sum_lvl2_ff\[48\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_6178_ net1106 VGND VPWR _0257_ DP_4.matrix\[41\] clknet_leaf_32_clk sg13g2_dfrbpq_2
X_5129_ _1889_ VPWR _1913_ VGND _1909_ _1911_ sg13g2_o21ai_1
XFILLER_45_639 VPWR VGND sg13g2_fill_1
XFILLER_44_149 VPWR VGND sg13g2_fill_2
XFILLER_26_864 VPWR VGND sg13g2_decap_8
XFILLER_38_1003 VPWR VGND sg13g2_decap_8
XFILLER_41_823 VPWR VGND sg13g2_decap_8
XFILLER_13_558 VPWR VGND sg13g2_fill_1
XFILLER_9_529 VPWR VGND sg13g2_fill_2
XFILLER_20_50 VPWR VGND sg13g2_fill_1
XFILLER_49_901 VPWR VGND sg13g2_decap_8
XFILLER_1_952 VPWR VGND sg13g2_decap_8
XFILLER_49_978 VPWR VGND sg13g2_decap_8
XFILLER_48_466 VPWR VGND sg13g2_fill_2
Xhold70 mac2.sum_lvl2_ff\[49\] VPWR VGND net110 sg13g2_dlygate4sd3_1
Xhold92 mac2.sum_lvl1_ff\[79\] VPWR VGND net132 sg13g2_dlygate4sd3_1
Xhold81 mac2.sum_lvl1_ff\[46\] VPWR VGND net121 sg13g2_dlygate4sd3_1
XFILLER_45_80 VPWR VGND sg13g2_fill_1
XFILLER_16_374 VPWR VGND sg13g2_fill_2
XFILLER_32_845 VPWR VGND sg13g2_decap_8
XFILLER_31_388 VPWR VGND sg13g2_fill_2
X_4500_ _1310_ _1311_ _1312_ VPWR VGND sg13g2_nor2_1
XFILLER_8_562 VPWR VGND sg13g2_fill_1
X_5480_ _2224_ mac2.sum_lvl2_ff\[20\] mac2.sum_lvl2_ff\[1\] VPWR VGND sg13g2_nand2_1
X_4431_ _1245_ _1235_ _1244_ VPWR VGND sg13g2_nand2b_1
X_4362_ _1176_ _1177_ _1175_ _1178_ VPWR VGND sg13g2_nand3_1
X_3313_ _0096_ _2900_ _2901_ VPWR VGND sg13g2_xnor2_1
X_6101_ net1094 VGND VPWR _0203_ DP_2.matrix\[7\] clknet_leaf_58_clk sg13g2_dfrbpq_2
X_4293_ _1110_ _1072_ _1107_ VPWR VGND sg13g2_xnor2_1
X_3244_ _2834_ _2795_ _0104_ VPWR VGND sg13g2_xor2_1
X_6032_ net1125 VGND VPWR _0111_ mac1.products_ff\[15\] clknet_leaf_42_clk sg13g2_dfrbpq_1
XFILLER_20_0 VPWR VGND sg13g2_fill_2
X_3175_ _2767_ _2762_ _2766_ VPWR VGND sg13g2_xnor2_1
Xfanout1090 net1091 net1090 VPWR VGND sg13g2_buf_8
XFILLER_39_488 VPWR VGND sg13g2_decap_4
XFILLER_35_661 VPWR VGND sg13g2_fill_2
X_5816_ _2505_ _2509_ _2510_ VPWR VGND sg13g2_nor2b_1
X_5747_ net949 net930 net788 _2442_ VPWR VGND sg13g2_mux2_1
X_5678_ _2369_ _2373_ _2379_ VPWR VGND sg13g2_nor2_1
X_4629_ _1430_ _1431_ _1432_ VPWR VGND sg13g2_and2_1
XFILLER_46_915 VPWR VGND sg13g2_decap_8
XFILLER_45_403 VPWR VGND sg13g2_fill_1
XFILLER_17_116 VPWR VGND sg13g2_fill_2
XFILLER_40_152 VPWR VGND sg13g2_decap_4
XFILLER_9_337 VPWR VGND sg13g2_fill_1
XFILLER_9_326 VPWR VGND sg13g2_fill_1
XFILLER_12_1017 VPWR VGND sg13g2_decap_8
XFILLER_12_1028 VPWR VGND sg13g2_fill_1
XFILLER_5_565 VPWR VGND sg13g2_fill_1
XFILLER_49_775 VPWR VGND sg13g2_fill_2
XFILLER_48_230 VPWR VGND sg13g2_fill_1
XFILLER_17_650 VPWR VGND sg13g2_fill_1
XFILLER_24_609 VPWR VGND sg13g2_fill_2
XFILLER_36_447 VPWR VGND sg13g2_fill_1
X_4980_ _1768_ net859 net811 net861 net808 VPWR VGND sg13g2_a22oi_1
XFILLER_44_491 VPWR VGND sg13g2_decap_8
X_3931_ _0764_ _0762_ _0763_ VPWR VGND sg13g2_nand2_1
XFILLER_32_620 VPWR VGND sg13g2_fill_2
X_3862_ _0696_ net1004 net927 VPWR VGND sg13g2_nand2_1
XFILLER_20_826 VPWR VGND sg13g2_fill_2
X_5601_ _0050_ _2317_ net338 VPWR VGND sg13g2_xnor2_1
X_5532_ mac2.sum_lvl2_ff\[12\] mac2.sum_lvl2_ff\[31\] _2265_ VPWR VGND sg13g2_xor2_1
X_3793_ _0629_ _0630_ _0631_ VPWR VGND sg13g2_nor2b_2
X_5463_ _2207_ _2208_ _2210_ _2212_ VPWR VGND sg13g2_or3_1
X_5394_ _2158_ _2157_ _2156_ VPWR VGND sg13g2_nand2b_1
X_4414_ _1228_ net879 net816 VPWR VGND sg13g2_nand2_1
XFILLER_28_1013 VPWR VGND sg13g2_decap_8
X_4345_ _1156_ VPWR _1161_ VGND _1157_ _1159_ sg13g2_o21ai_1
X_4276_ _1093_ _1065_ _1094_ VPWR VGND sg13g2_nor2b_1
X_3227_ _2818_ net916 net1033 VPWR VGND sg13g2_nand2_1
XFILLER_28_915 VPWR VGND sg13g2_decap_8
X_6015_ net1056 VGND VPWR DP_3.Q_range.data_plus_4\[6\] DP_3.Q_range.out_data\[5\]
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
X_3158_ _2721_ VPWR _2750_ VGND _2718_ _2722_ sg13g2_o21ai_1
XFILLER_43_918 VPWR VGND sg13g2_decap_8
X_3089_ _2666_ VPWR _2683_ VGND _2657_ _2667_ sg13g2_o21ai_1
XFILLER_36_992 VPWR VGND sg13g2_decap_8
XFILLER_35_1028 VPWR VGND sg13g2_fill_1
XFILLER_23_686 VPWR VGND sg13g2_decap_8
XFILLER_23_697 VPWR VGND sg13g2_fill_1
XFILLER_11_859 VPWR VGND sg13g2_fill_2
XFILLER_6_329 VPWR VGND sg13g2_fill_2
Xhold381 _2193_ VPWR VGND net421 sg13g2_dlygate4sd3_1
XFILLER_2_557 VPWR VGND sg13g2_fill_2
Xhold370 DP_4.matrix\[2\] VPWR VGND net410 sg13g2_dlygate4sd3_1
Xhold392 _0625_ VPWR VGND net432 sg13g2_dlygate4sd3_1
Xfanout850 DP_4.matrix\[0\] net850 VPWR VGND sg13g2_buf_1
Xfanout861 net862 net861 VPWR VGND sg13g2_buf_1
Xfanout872 net299 net872 VPWR VGND sg13g2_buf_8
Xfanout894 net416 net894 VPWR VGND sg13g2_buf_8
Xfanout883 DP_3.matrix\[38\] net883 VPWR VGND sg13g2_buf_8
XFILLER_45_288 VPWR VGND sg13g2_fill_2
XFILLER_42_940 VPWR VGND sg13g2_decap_8
XFILLER_26_82 VPWR VGND sg13g2_fill_1
XFILLER_27_992 VPWR VGND sg13g2_decap_8
X_4130_ _0918_ _0956_ _0957_ VPWR VGND sg13g2_nor2_1
XFILLER_49_550 VPWR VGND sg13g2_fill_1
X_4061_ _0890_ net929 net989 VPWR VGND sg13g2_nand2_1
XFILLER_49_572 VPWR VGND sg13g2_fill_2
X_3012_ _2610_ net984 net915 VPWR VGND sg13g2_nand2_1
XFILLER_25_907 VPWR VGND sg13g2_decap_4
XFILLER_33_940 VPWR VGND sg13g2_decap_8
X_4963_ _1748_ _1749_ _1751_ _1752_ VPWR VGND sg13g2_nor3_1
X_3914_ _0742_ VPWR _0747_ VGND _0743_ _0745_ sg13g2_o21ai_1
XFILLER_32_450 VPWR VGND sg13g2_fill_2
X_4894_ _1668_ VPWR _1689_ VGND _1665_ _1669_ sg13g2_o21ai_1
XFILLER_32_483 VPWR VGND sg13g2_fill_2
X_3845_ _0675_ VPWR _0680_ VGND _0676_ _0678_ sg13g2_o21ai_1
X_3776_ VGND VPWR _0586_ _0609_ _0617_ _0611_ sg13g2_a21oi_1
X_5515_ net490 mac2.sum_lvl2_ff\[27\] _2249_ _2251_ VPWR VGND sg13g2_a21o_1
X_6495_ net1059 VGND VPWR _0036_ mac2.sum_lvl3_ff\[13\] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_5446_ _0031_ _2194_ net359 VPWR VGND sg13g2_xnor2_1
X_5377_ _2139_ _2137_ _2138_ _2144_ VPWR VGND sg13g2_a21o_2
X_4328_ _1142_ _1138_ _1144_ VPWR VGND sg13g2_xor2_1
X_4259_ _1048_ VPWR _1077_ VGND _1046_ _1049_ sg13g2_o21ai_1
XFILLER_43_726 VPWR VGND sg13g2_fill_2
XFILLER_15_428 VPWR VGND sg13g2_fill_1
XFILLER_24_940 VPWR VGND sg13g2_decap_8
XFILLER_11_667 VPWR VGND sg13g2_fill_1
XFILLER_46_520 VPWR VGND sg13g2_fill_2
XFILLER_15_962 VPWR VGND sg13g2_decap_8
XFILLER_30_932 VPWR VGND sg13g2_decap_8
X_3630_ _0477_ _0440_ _0475_ VPWR VGND sg13g2_nand2_1
X_3561_ VGND VPWR _0409_ _0407_ _0364_ sg13g2_or2_1
X_5300_ VGND VPWR _2056_ _2059_ _2079_ _2055_ sg13g2_a21oi_1
X_3492_ _0339_ _0340_ _0334_ _0342_ VPWR VGND sg13g2_nand3_1
X_6280_ net1046 VGND VPWR net166 mac1.sum_lvl1_ff\[83\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_5231_ VGND VPWR _2012_ _1983_ _1981_ sg13g2_or2_1
XFILLER_25_1005 VPWR VGND sg13g2_decap_8
X_5162_ _1945_ _1940_ _1944_ VPWR VGND sg13g2_xnor2_1
X_4113_ _0939_ _0940_ _0941_ VPWR VGND sg13g2_nor2_1
X_5093_ _1876_ _1875_ _0157_ VPWR VGND sg13g2_xor2_1
X_4044_ _0874_ _0864_ _0873_ VPWR VGND sg13g2_nand2b_1
XFILLER_37_553 VPWR VGND sg13g2_decap_8
X_5995_ net275 _0243_ VPWR VGND sg13g2_buf_1
XFILLER_24_247 VPWR VGND sg13g2_fill_2
X_4946_ _1737_ net867 net810 _0089_ VPWR VGND sg13g2_and3_2
X_4877_ _1672_ _1663_ _1673_ VPWR VGND sg13g2_nor2b_1
XFILLER_20_442 VPWR VGND sg13g2_fill_1
XFILLER_21_943 VPWR VGND sg13g2_decap_8
X_3828_ _0662_ _0663_ _0664_ VPWR VGND sg13g2_nor2b_2
XFILLER_3_107 VPWR VGND sg13g2_fill_2
X_3759_ _0581_ VPWR _0601_ VGND _0553_ _0579_ sg13g2_o21ai_1
X_6478_ net1126 VGND VPWR net108 mac2.sum_lvl2_ff\[31\] clknet_leaf_36_clk sg13g2_dfrbpq_2
X_5429_ _2179_ net502 _2183_ _2184_ VPWR VGND sg13g2_nor3_1
XFILLER_31_707 VPWR VGND sg13g2_fill_2
XFILLER_30_228 VPWR VGND sg13g2_decap_4
XFILLER_8_914 VPWR VGND sg13g2_fill_2
XFILLER_8_969 VPWR VGND sg13g2_decap_8
XFILLER_23_83 VPWR VGND sg13g2_fill_1
X_4800_ _1598_ net896 net833 VPWR VGND sg13g2_nand2_1
XFILLER_34_578 VPWR VGND sg13g2_fill_1
X_5780_ net778 VPWR _2474_ VGND net1028 net785 sg13g2_o21ai_1
X_4731_ _1527_ _1528_ _1530_ _1531_ VPWR VGND sg13g2_or3_1
XFILLER_30_773 VPWR VGND sg13g2_decap_4
X_4662_ _1464_ _1440_ _1463_ VPWR VGND sg13g2_xnor2_1
X_3613_ _0460_ _0455_ _0459_ VPWR VGND sg13g2_xnor2_1
X_6401_ net1077 VGND VPWR _0093_ mac2.products_ff\[140\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_4593_ _1397_ net895 net848 net897 net844 VPWR VGND sg13g2_a22oi_1
X_3544_ _0391_ _0390_ _0113_ VPWR VGND sg13g2_xor2_1
X_6332_ net1094 VGND VPWR net392 mac1.sum_lvl3_ff\[15\] clknet_leaf_58_clk sg13g2_dfrbpq_1
X_3475_ _0325_ _0323_ _0324_ VPWR VGND sg13g2_nand2b_1
X_6263_ net1055 VGND VPWR net112 mac2.sum_lvl2_ff\[48\] clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_9_1021 VPWR VGND sg13g2_decap_8
X_5214_ _1996_ _1995_ _1994_ VPWR VGND sg13g2_nand2b_1
X_6194_ net1096 VGND VPWR net251 mac1.sum_lvl1_ff\[41\] clknet_leaf_54_clk sg13g2_dfrbpq_1
X_5145_ _1882_ _1885_ _1928_ VPWR VGND sg13g2_nor2_1
X_5076_ _1861_ _1854_ _1859_ _1860_ VPWR VGND sg13g2_and3_1
XFILLER_44_309 VPWR VGND sg13g2_fill_1
X_4027_ _0857_ net994 net927 VPWR VGND sg13g2_nand2_1
XFILLER_38_884 VPWR VGND sg13g2_decap_8
X_5978_ net908 _0218_ VPWR VGND sg13g2_buf_1
X_4929_ _1721_ _1715_ _1723_ VPWR VGND sg13g2_xor2_1
XFILLER_21_762 VPWR VGND sg13g2_fill_1
XFILLER_29_862 VPWR VGND sg13g2_decap_8
XFILLER_28_372 VPWR VGND sg13g2_fill_2
XFILLER_43_375 VPWR VGND sg13g2_fill_1
XFILLER_15_1004 VPWR VGND sg13g2_decap_8
XFILLER_11_294 VPWR VGND sg13g2_fill_1
XFILLER_4_972 VPWR VGND sg13g2_decap_8
X_3260_ _2850_ net970 net909 VPWR VGND sg13g2_nand2_1
X_3191_ _2760_ _2780_ _2782_ _2783_ VPWR VGND sg13g2_or3_1
XFILLER_38_125 VPWR VGND sg13g2_fill_2
XFILLER_35_832 VPWR VGND sg13g2_decap_8
X_5901_ VGND VPWR net768 _2575_ _0221_ _2574_ sg13g2_a21oi_1
X_5832_ net831 net847 net786 _2525_ VPWR VGND sg13g2_mux2_1
X_5763_ DP_2.matrix\[40\] net791 _2458_ VPWR VGND sg13g2_nor2_1
X_4714_ _1509_ _1513_ _1514_ VPWR VGND sg13g2_nor2_1
X_5694_ mac2.total_sum\[0\] mac1.total_sum\[0\] net25 VPWR VGND sg13g2_xor2_1
X_4645_ _1447_ _1442_ _1445_ VPWR VGND sg13g2_xnor2_1
X_4576_ _1377_ _1378_ _1380_ _1381_ VPWR VGND sg13g2_nor3_1
X_3527_ _0376_ _0369_ _0374_ _0375_ VPWR VGND sg13g2_and3_1
X_6315_ net1074 VGND VPWR net81 mac1.sum_lvl3_ff\[34\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_3458_ _0309_ _0302_ _0307_ _0308_ VPWR VGND sg13g2_and3_1
X_6246_ net1047 VGND VPWR net83 mac1.sum_lvl2_ff\[47\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_6177_ net1122 VGND VPWR _0256_ DP_4.matrix\[40\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_3389_ _2961_ VPWR _2974_ VGND _2934_ _2959_ sg13g2_o21ai_1
X_5128_ _1889_ _1909_ _1911_ _1912_ VPWR VGND sg13g2_or3_1
X_5059_ _1844_ _1840_ _1843_ VPWR VGND sg13g2_nand2_1
XFILLER_25_397 VPWR VGND sg13g2_fill_2
XFILLER_40_345 VPWR VGND sg13g2_fill_2
XFILLER_41_879 VPWR VGND sg13g2_decap_8
XFILLER_5_714 VPWR VGND sg13g2_fill_1
XFILLER_4_246 VPWR VGND sg13g2_fill_2
XFILLER_45_1008 VPWR VGND sg13g2_decap_8
XFILLER_1_931 VPWR VGND sg13g2_decap_8
XFILLER_48_401 VPWR VGND sg13g2_fill_1
XFILLER_49_957 VPWR VGND sg13g2_decap_8
Xhold60 mac1.sum_lvl2_ff\[39\] VPWR VGND net100 sg13g2_dlygate4sd3_1
Xhold82 mac2.sum_lvl2_ff\[44\] VPWR VGND net122 sg13g2_dlygate4sd3_1
Xhold71 mac2.products_ff\[5\] VPWR VGND net111 sg13g2_dlygate4sd3_1
XFILLER_17_810 VPWR VGND sg13g2_fill_2
Xhold93 mac1.sum_lvl1_ff\[14\] VPWR VGND net133 sg13g2_dlygate4sd3_1
XFILLER_43_161 VPWR VGND sg13g2_decap_8
XFILLER_31_301 VPWR VGND sg13g2_fill_1
XFILLER_32_824 VPWR VGND sg13g2_decap_8
Xclkbuf_4_14_0_clk clknet_0_clk clknet_4_14_0_clk VPWR VGND sg13g2_buf_8
X_4430_ _1244_ _1236_ _1243_ VPWR VGND sg13g2_xnor2_1
X_6100_ net1093 VGND VPWR _0202_ DP_2.matrix\[6\] clknet_leaf_59_clk sg13g2_dfrbpq_1
X_4361_ _1129_ VPWR _1177_ VGND _1068_ _1130_ sg13g2_o21ai_1
X_3312_ _2865_ _2870_ _2901_ VPWR VGND sg13g2_nor2_1
X_4292_ _1072_ _1107_ _1109_ VPWR VGND sg13g2_and2_1
X_3243_ _2832_ _2833_ _2834_ VPWR VGND sg13g2_nor2b_1
X_6031_ net1111 VGND VPWR _0110_ mac1.products_ff\[14\] clknet_leaf_44_clk sg13g2_dfrbpq_1
XFILLER_6_1013 VPWR VGND sg13g2_decap_8
X_3174_ _2766_ _2719_ _2764_ VPWR VGND sg13g2_xnor2_1
Xfanout1091 rst_n net1091 VPWR VGND sg13g2_buf_8
Xfanout1080 net1090 net1080 VPWR VGND sg13g2_buf_8
XFILLER_25_29 VPWR VGND sg13g2_fill_1
X_5815_ _2506_ VPWR _2509_ VGND _2507_ _2508_ sg13g2_o21ai_1
XFILLER_23_868 VPWR VGND sg13g2_fill_2
X_5746_ _2441_ _2440_ net783 net780 net906 VPWR VGND sg13g2_a22oi_1
X_5677_ _2367_ _2372_ _2378_ VPWR VGND sg13g2_nor2_1
X_4628_ _1429_ _1428_ _1390_ _1431_ VPWR VGND sg13g2_a21o_1
X_4559_ _1366_ net901 net843 _0084_ VPWR VGND sg13g2_and3_2
X_6229_ net1113 VGND VPWR net159 mac1.sum_lvl2_ff\[27\] clknet_leaf_50_clk sg13g2_dfrbpq_2
XFILLER_45_426 VPWR VGND sg13g2_fill_1
Xheichips25_template_40 VPWR VGND uio_oe[7] sg13g2_tiehi
XFILLER_22_890 VPWR VGND sg13g2_fill_2
XFILLER_5_555 VPWR VGND sg13g2_fill_2
XFILLER_36_415 VPWR VGND sg13g2_decap_4
XFILLER_37_949 VPWR VGND sg13g2_decap_8
XFILLER_36_437 VPWR VGND sg13g2_fill_2
X_3930_ _0725_ _0724_ _0723_ _0763_ VPWR VGND sg13g2_a21o_2
XFILLER_44_470 VPWR VGND sg13g2_fill_2
X_3861_ _0672_ VPWR _0695_ VGND _0647_ _0670_ sg13g2_o21ai_1
XFILLER_20_816 VPWR VGND sg13g2_fill_2
XFILLER_32_676 VPWR VGND sg13g2_decap_8
X_3792_ _0626_ VPWR _0630_ VGND _0627_ _0628_ sg13g2_o21ai_1
X_5600_ _2318_ net337 _2315_ VPWR VGND sg13g2_nand2_1
X_5531_ mac2.sum_lvl2_ff\[31\] mac2.sum_lvl2_ff\[12\] _2264_ VPWR VGND sg13g2_nor2_1
XFILLER_8_393 VPWR VGND sg13g2_fill_1
X_5462_ _2207_ VPWR _2211_ VGND _2208_ _2210_ sg13g2_o21ai_1
X_5393_ VGND VPWR _2157_ mac1.sum_lvl2_ff\[13\] mac1.sum_lvl2_ff\[32\] sg13g2_or2_1
X_4413_ _1227_ net879 net815 VPWR VGND sg13g2_nand2_1
X_4344_ _1156_ _1157_ _1159_ _1160_ VPWR VGND sg13g2_or3_1
X_4275_ _1093_ _1069_ _1092_ VPWR VGND sg13g2_xnor2_1
X_6014_ net1056 VGND VPWR net11 DP_3.Q_range.out_data\[4\] clknet_leaf_22_clk sg13g2_dfrbpq_1
X_3226_ _2771_ VPWR _2817_ VGND _2769_ _2772_ sg13g2_o21ai_1
X_3157_ _2738_ VPWR _2749_ VGND _2716_ _2739_ sg13g2_o21ai_1
X_3088_ _2680_ _2679_ _2682_ VPWR VGND sg13g2_xor2_1
XFILLER_36_971 VPWR VGND sg13g2_decap_8
XFILLER_35_481 VPWR VGND sg13g2_fill_1
XFILLER_35_1007 VPWR VGND sg13g2_decap_8
XFILLER_7_809 VPWR VGND sg13g2_fill_1
X_5729_ net1011 net996 net788 _2425_ VPWR VGND sg13g2_mux2_1
Xhold371 DP_2.matrix\[6\] VPWR VGND net411 sg13g2_dlygate4sd3_1
Xhold360 DP_4.matrix\[37\] VPWR VGND net400 sg13g2_dlygate4sd3_1
Xhold393 _0075_ VPWR VGND net433 sg13g2_dlygate4sd3_1
Xhold382 _0030_ VPWR VGND net422 sg13g2_dlygate4sd3_1
Xfanout851 net853 net851 VPWR VGND sg13g2_buf_2
Xfanout840 DP_4.matrix\[3\] net840 VPWR VGND sg13g2_buf_1
Xfanout862 net351 net862 VPWR VGND sg13g2_buf_1
XFILLER_19_905 VPWR VGND sg13g2_decap_8
Xfanout884 net885 net884 VPWR VGND sg13g2_buf_8
Xfanout873 net874 net873 VPWR VGND sg13g2_buf_8
XFILLER_18_404 VPWR VGND sg13g2_fill_2
Xfanout895 net385 net895 VPWR VGND sg13g2_buf_8
XFILLER_46_746 VPWR VGND sg13g2_fill_1
XFILLER_27_971 VPWR VGND sg13g2_decap_8
XFILLER_26_72 VPWR VGND sg13g2_fill_2
XFILLER_42_996 VPWR VGND sg13g2_decap_8
X_4060_ _0872_ _0865_ _0835_ _0889_ VPWR VGND sg13g2_a21o_1
X_3011_ _2608_ _2609_ _0065_ VPWR VGND sg13g2_nor2_1
XFILLER_18_982 VPWR VGND sg13g2_decap_8
XFILLER_36_256 VPWR VGND sg13g2_fill_1
X_4962_ _1751_ net860 net812 net864 net809 VPWR VGND sg13g2_a22oi_1
X_4893_ _1671_ _1664_ _1673_ _1688_ VPWR VGND sg13g2_a21o_1
X_3913_ _0742_ _0743_ _0745_ _0746_ VPWR VGND sg13g2_or3_1
X_3844_ _0675_ _0676_ _0678_ _0679_ VPWR VGND sg13g2_or3_1
XFILLER_33_996 VPWR VGND sg13g2_decap_8
XFILLER_20_679 VPWR VGND sg13g2_fill_1
X_3775_ _0613_ VPWR _0616_ VGND _0598_ _0615_ sg13g2_o21ai_1
X_5514_ net492 _2250_ _0046_ VPWR VGND sg13g2_nor2b_2
X_6494_ net1054 VGND VPWR _0035_ mac2.sum_lvl3_ff\[12\] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_5445_ _2196_ VPWR _2197_ VGND _2190_ _2192_ sg13g2_o21ai_1
X_5376_ VPWR _2143_ _2142_ VGND sg13g2_inv_1
X_4327_ _1138_ _1142_ _1143_ VPWR VGND sg13g2_nor2_1
X_4258_ _1076_ _1071_ _1074_ VPWR VGND sg13g2_xnor2_1
X_3209_ _2765_ VPWR _2800_ VGND _2762_ _2766_ sg13g2_o21ai_1
XFILLER_28_702 VPWR VGND sg13g2_fill_1
X_4189_ _1006_ _1007_ _1009_ _1010_ VPWR VGND sg13g2_nor3_1
XFILLER_24_996 VPWR VGND sg13g2_decap_8
Xhold190 mac2.sum_lvl2_ff\[39\] VPWR VGND net230 sg13g2_dlygate4sd3_1
XFILLER_46_543 VPWR VGND sg13g2_fill_1
XFILLER_15_941 VPWR VGND sg13g2_fill_1
XFILLER_18_1024 VPWR VGND sg13g2_decap_4
XFILLER_30_911 VPWR VGND sg13g2_decap_8
XFILLER_30_988 VPWR VGND sg13g2_decap_8
X_3560_ _0408_ net952 net1010 VPWR VGND sg13g2_nand2_1
X_3491_ _0341_ _0334_ _0339_ _0340_ VPWR VGND sg13g2_and3_1
X_5230_ _1971_ VPWR _2011_ VGND _1968_ _1972_ sg13g2_o21ai_1
X_5161_ _1944_ _1892_ _1941_ VPWR VGND sg13g2_xnor2_1
X_4112_ VGND VPWR _0888_ _0907_ _0940_ _0909_ sg13g2_a21oi_1
XFILLER_25_1028 VPWR VGND sg13g2_fill_1
X_5092_ _1877_ _1875_ _1876_ VPWR VGND sg13g2_nand2_1
X_4043_ _0873_ _0865_ _0872_ VPWR VGND sg13g2_xnor2_1
X_5994_ net280 _0242_ VPWR VGND sg13g2_buf_1
X_4945_ net869 net282 _0089_ VPWR VGND sg13g2_and2_1
X_4876_ _1672_ _1664_ _1671_ VPWR VGND sg13g2_xnor2_1
X_3827_ _0642_ VPWR _0663_ VGND _0633_ _0643_ sg13g2_o21ai_1
XFILLER_21_999 VPWR VGND sg13g2_decap_8
X_3758_ _0584_ _0576_ _0583_ _0600_ VPWR VGND sg13g2_a21o_1
X_3689_ _0533_ _0526_ _0534_ VPWR VGND sg13g2_nor2b_1
X_6477_ net1125 VGND VPWR net82 mac2.sum_lvl2_ff\[30\] clknet_leaf_39_clk sg13g2_dfrbpq_2
X_5428_ VPWR VGND _2177_ _2176_ _2175_ mac1.sum_lvl3_ff\[25\] _2183_ net320 sg13g2_a221oi_1
X_5359_ _2128_ net510 _0012_ VPWR VGND sg13g2_nor2b_2
XFILLER_43_524 VPWR VGND sg13g2_fill_2
XFILLER_24_760 VPWR VGND sg13g2_fill_1
XFILLER_23_292 VPWR VGND sg13g2_fill_1
XFILLER_48_1017 VPWR VGND sg13g2_decap_8
XFILLER_48_1028 VPWR VGND sg13g2_fill_1
XFILLER_2_141 VPWR VGND sg13g2_fill_2
XFILLER_47_885 VPWR VGND sg13g2_decap_8
XFILLER_46_384 VPWR VGND sg13g2_fill_1
X_4730_ _1530_ net1028 net849 net888 net845 VPWR VGND sg13g2_a22oi_1
XFILLER_9_75 VPWR VGND sg13g2_fill_2
X_4661_ _1463_ _1460_ _1462_ VPWR VGND sg13g2_nand2_1
X_3612_ _0459_ _0407_ _0456_ VPWR VGND sg13g2_xnor2_1
X_6400_ net1077 VGND VPWR _0092_ mac2.products_ff\[139\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_31_1010 VPWR VGND sg13g2_decap_8
X_6331_ net1075 VGND VPWR net462 mac1.sum_lvl3_ff\[14\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_4592_ net844 net897 net848 _1396_ VPWR VGND net895 sg13g2_nand4_1
X_3543_ _0392_ _0390_ _0391_ VPWR VGND sg13g2_nand2_1
X_3474_ _0324_ net1020 net946 VPWR VGND sg13g2_nand2_1
X_6262_ net1060 VGND VPWR net154 mac2.sum_lvl2_ff\[47\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_6193_ net1097 VGND VPWR net248 mac1.sum_lvl1_ff\[40\] clknet_leaf_54_clk sg13g2_dfrbpq_1
XFILLER_9_1000 VPWR VGND sg13g2_decap_8
X_5213_ _1959_ _1993_ _1957_ _1995_ VPWR VGND sg13g2_nand3_1
X_5144_ _1910_ VPWR _1927_ VGND _1889_ _1911_ sg13g2_o21ai_1
XFILLER_29_307 VPWR VGND sg13g2_fill_2
X_5075_ _1855_ VPWR _1860_ VGND _1856_ _1858_ sg13g2_o21ai_1
X_4026_ _0856_ net994 net925 VPWR VGND sg13g2_nand2_1
XFILLER_38_863 VPWR VGND sg13g2_decap_8
XFILLER_25_524 VPWR VGND sg13g2_fill_1
XFILLER_37_384 VPWR VGND sg13g2_fill_2
X_5977_ net910 _0217_ VPWR VGND sg13g2_buf_1
X_4928_ _1722_ _1715_ _1721_ VPWR VGND sg13g2_nand2_1
X_4859_ _1654_ _1655_ _1656_ VPWR VGND sg13g2_nor2_1
XFILLER_0_623 VPWR VGND sg13g2_fill_2
XFILLER_48_638 VPWR VGND sg13g2_fill_1
XFILLER_44_888 VPWR VGND sg13g2_decap_8
XFILLER_4_951 VPWR VGND sg13g2_decap_8
X_3190_ VGND VPWR _2778_ _2779_ _2782_ _2761_ sg13g2_a21oi_1
XFILLER_19_351 VPWR VGND sg13g2_fill_1
XFILLER_35_811 VPWR VGND sg13g2_decap_8
X_5900_ _2575_ _2492_ _2496_ VPWR VGND sg13g2_xnor2_1
XFILLER_35_888 VPWR VGND sg13g2_decap_8
X_5831_ _2524_ _2523_ net779 net776 net374 VPWR VGND sg13g2_a22oi_1
X_5762_ _2457_ net269 net781 VPWR VGND sg13g2_nand2_1
XFILLER_34_387 VPWR VGND sg13g2_fill_1
X_4713_ VGND VPWR _1513_ _1512_ _1511_ sg13g2_or2_1
X_5693_ net24 _2389_ _2390_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_593 VPWR VGND sg13g2_fill_1
X_4644_ _1446_ _1445_ _1442_ VPWR VGND sg13g2_nand2b_1
X_4575_ _1380_ net897 net848 net899 net843 VPWR VGND sg13g2_a22oi_1
X_3526_ _0370_ VPWR _0375_ VGND _0371_ _0373_ sg13g2_o21ai_1
X_6314_ net1069 VGND VPWR net99 mac1.sum_lvl3_ff\[33\] clknet_leaf_10_clk sg13g2_dfrbpq_2
X_6245_ net1042 VGND VPWR net177 mac1.sum_lvl2_ff\[46\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3457_ _0303_ VPWR _0308_ VGND _0304_ _0306_ sg13g2_o21ai_1
X_6176_ net1106 VGND VPWR _0255_ DP_4.matrix\[39\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_3388_ VGND VPWR _2942_ _2965_ _2973_ _2967_ sg13g2_a21oi_1
X_5127_ VGND VPWR _1907_ _1908_ _1911_ _1890_ sg13g2_a21oi_1
X_5058_ _1841_ _1842_ _1843_ VPWR VGND sg13g2_nor2b_1
X_4009_ _0839_ _0832_ _0840_ VPWR VGND sg13g2_xor2_1
Xclkbuf_leaf_64_clk clknet_4_2_0_clk clknet_leaf_64_clk VPWR VGND sg13g2_buf_8
XFILLER_13_505 VPWR VGND sg13g2_fill_1
XFILLER_13_516 VPWR VGND sg13g2_fill_2
XFILLER_40_302 VPWR VGND sg13g2_fill_1
XFILLER_41_858 VPWR VGND sg13g2_decap_8
XFILLER_21_582 VPWR VGND sg13g2_fill_2
XFILLER_1_910 VPWR VGND sg13g2_decap_8
XFILLER_1_987 VPWR VGND sg13g2_decap_8
XFILLER_49_936 VPWR VGND sg13g2_decap_8
Xhold50 mac1.sum_lvl2_ff\[46\] VPWR VGND net90 sg13g2_dlygate4sd3_1
Xhold83 mac2.sum_lvl1_ff\[49\] VPWR VGND net123 sg13g2_dlygate4sd3_1
XFILLER_21_1020 VPWR VGND sg13g2_decap_8
Xhold72 mac2.sum_lvl1_ff\[82\] VPWR VGND net112 sg13g2_dlygate4sd3_1
Xhold61 mac2.sum_lvl1_ff\[1\] VPWR VGND net101 sg13g2_dlygate4sd3_1
XFILLER_17_822 VPWR VGND sg13g2_fill_2
Xhold94 mac1.sum_lvl1_ff\[85\] VPWR VGND net134 sg13g2_dlygate4sd3_1
XFILLER_29_682 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_55_clk clknet_4_8_0_clk clknet_leaf_55_clk VPWR VGND sg13g2_buf_8
XFILLER_17_888 VPWR VGND sg13g2_fill_2
XFILLER_8_520 VPWR VGND sg13g2_fill_1
XFILLER_12_582 VPWR VGND sg13g2_decap_8
XFILLER_6_43 VPWR VGND sg13g2_fill_2
X_4360_ _1102_ VPWR _1176_ VGND _1172_ _1174_ sg13g2_o21ai_1
X_3311_ _2898_ _2899_ _2900_ VPWR VGND sg13g2_nor2_1
X_4291_ VGND VPWR _1108_ _1106_ _1073_ sg13g2_or2_1
X_3242_ _2833_ _2796_ _2831_ VPWR VGND sg13g2_nand2_1
X_6030_ net1111 VGND VPWR _0109_ mac1.products_ff\[13\] clknet_leaf_44_clk sg13g2_dfrbpq_1
XFILLER_39_402 VPWR VGND sg13g2_fill_2
X_3173_ VGND VPWR _2765_ _2763_ _2720_ sg13g2_or2_1
Xfanout1081 net1090 net1081 VPWR VGND sg13g2_buf_8
Xfanout1070 net1072 net1070 VPWR VGND sg13g2_buf_8
Xfanout1092 net1095 net1092 VPWR VGND sg13g2_buf_8
XFILLER_39_446 VPWR VGND sg13g2_fill_1
XFILLER_19_170 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_46_clk clknet_4_11_0_clk clknet_leaf_46_clk VPWR VGND sg13g2_buf_8
XFILLER_35_663 VPWR VGND sg13g2_fill_1
X_5814_ net778 VPWR _2508_ VGND net892 net785 sg13g2_o21ai_1
X_5745_ VGND VPWR _2606_ net791 _2440_ _2439_ sg13g2_a21oi_1
XFILLER_31_891 VPWR VGND sg13g2_decap_8
X_5676_ mac2.total_sum\[12\] mac1.total_sum\[12\] _2377_ VPWR VGND sg13g2_xor2_1
X_4627_ _1428_ _1429_ _1390_ _1430_ VPWR VGND sg13g2_nand3_1
X_4558_ net903 net847 _0084_ VPWR VGND sg13g2_and2_1
X_4489_ _1301_ _1294_ _1300_ VPWR VGND sg13g2_xnor2_1
XFILLER_1_228 VPWR VGND sg13g2_fill_1
X_3509_ _0356_ _0357_ _0358_ VPWR VGND sg13g2_nor2b_1
X_6228_ net1108 VGND VPWR net184 mac1.sum_lvl2_ff\[26\] clknet_leaf_50_clk sg13g2_dfrbpq_2
X_6159_ net1111 VGND VPWR net175 mac1.sum_lvl1_ff\[12\] clknet_leaf_46_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_37_clk clknet_4_15_0_clk clknet_leaf_37_clk VPWR VGND sg13g2_buf_8
XFILLER_13_324 VPWR VGND sg13g2_decap_8
XFILLER_41_633 VPWR VGND sg13g2_fill_1
XFILLER_13_335 VPWR VGND sg13g2_fill_1
XFILLER_5_523 VPWR VGND sg13g2_fill_2
XFILLER_5_512 VPWR VGND sg13g2_fill_2
XFILLER_49_777 VPWR VGND sg13g2_fill_1
XFILLER_37_928 VPWR VGND sg13g2_decap_8
XFILLER_17_641 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_28_clk clknet_4_7_0_clk clknet_leaf_28_clk VPWR VGND sg13g2_buf_8
XFILLER_45_994 VPWR VGND sg13g2_decap_8
XFILLER_16_162 VPWR VGND sg13g2_fill_2
XFILLER_17_685 VPWR VGND sg13g2_decap_8
X_3860_ _0694_ _0686_ _0688_ VPWR VGND sg13g2_nand2_1
X_3791_ _0626_ _0627_ _0628_ _0629_ VPWR VGND sg13g2_nor3_1
X_5530_ _2263_ mac2.sum_lvl2_ff\[31\] mac2.sum_lvl2_ff\[12\] VPWR VGND sg13g2_nand2_1
X_5461_ VGND VPWR _2195_ _2197_ _2210_ _2209_ sg13g2_a21oi_1
X_4412_ _1226_ net883 net1022 VPWR VGND sg13g2_nand2_1
X_5392_ mac1.sum_lvl2_ff\[32\] mac1.sum_lvl2_ff\[13\] _2156_ VPWR VGND sg13g2_and2_1
X_4343_ _1159_ net1026 net829 net871 net828 VPWR VGND sg13g2_a22oi_1
X_4274_ _1092_ _1089_ _1091_ VPWR VGND sg13g2_nand2_1
X_3225_ _2816_ _2811_ _2815_ VPWR VGND sg13g2_xnor2_1
X_6013_ net1056 VGND VPWR net10 DP_3.Q_range.out_data\[3\] clknet_leaf_22_clk sg13g2_dfrbpq_1
X_3156_ _2747_ _2746_ _0102_ VPWR VGND sg13g2_xor2_1
X_3087_ _2681_ _2679_ _2680_ VPWR VGND sg13g2_nand2b_1
Xclkbuf_leaf_19_clk clknet_4_4_0_clk clknet_leaf_19_clk VPWR VGND sg13g2_buf_8
XFILLER_36_950 VPWR VGND sg13g2_decap_8
X_5728_ VGND VPWR _2424_ _2423_ _2413_ sg13g2_or2_1
X_3989_ _0819_ _0768_ _0820_ VPWR VGND sg13g2_xor2_1
XFILLER_22_187 VPWR VGND sg13g2_fill_2
X_5659_ mac2.total_sum\[8\] mac1.total_sum\[8\] _2361_ _2363_ VPWR VGND sg13g2_a21o_1
Xhold350 mac1.sum_lvl2_ff\[15\] VPWR VGND net390 sg13g2_dlygate4sd3_1
Xhold361 _0996_ VPWR VGND net401 sg13g2_dlygate4sd3_1
XFILLER_2_559 VPWR VGND sg13g2_fill_1
Xhold372 DP_2.matrix\[42\] VPWR VGND net412 sg13g2_dlygate4sd3_1
Xhold394 mac1.sum_lvl2_ff\[9\] VPWR VGND net434 sg13g2_dlygate4sd3_1
Xhold383 mac2.sum_lvl3_ff\[8\] VPWR VGND net423 sg13g2_dlygate4sd3_1
Xfanout852 net853 net852 VPWR VGND sg13g2_buf_1
Xfanout830 net373 net830 VPWR VGND sg13g2_buf_8
Xfanout841 net410 net841 VPWR VGND sg13g2_buf_8
Xclkbuf_4_13_0_clk clknet_0_clk clknet_4_13_0_clk VPWR VGND sg13g2_buf_8
Xfanout885 net516 net885 VPWR VGND sg13g2_buf_8
Xfanout863 net865 net863 VPWR VGND sg13g2_buf_8
Xfanout874 net875 net874 VPWR VGND sg13g2_buf_1
XFILLER_19_928 VPWR VGND sg13g2_fill_2
Xfanout896 DP_3.matrix\[4\] net896 VPWR VGND sg13g2_buf_2
XFILLER_34_909 VPWR VGND sg13g2_decap_8
XFILLER_27_950 VPWR VGND sg13g2_decap_8
XFILLER_42_975 VPWR VGND sg13g2_decap_8
XFILLER_14_655 VPWR VGND sg13g2_fill_2
XFILLER_14_677 VPWR VGND sg13g2_decap_8
XFILLER_14_688 VPWR VGND sg13g2_fill_1
XFILLER_41_463 VPWR VGND sg13g2_fill_1
XFILLER_42_61 VPWR VGND sg13g2_fill_1
XFILLER_10_894 VPWR VGND sg13g2_decap_4
XFILLER_5_375 VPWR VGND sg13g2_fill_2
XFILLER_49_541 VPWR VGND sg13g2_decap_8
XFILLER_49_574 VPWR VGND sg13g2_fill_1
X_3010_ _2609_ net917 net984 net981 net923 VPWR VGND sg13g2_a22oi_1
XFILLER_3_1017 VPWR VGND sg13g2_decap_8
XFILLER_3_1028 VPWR VGND sg13g2_fill_1
XFILLER_18_961 VPWR VGND sg13g2_decap_8
X_4961_ net809 net864 net812 _1750_ VPWR VGND net860 sg13g2_nand4_1
X_4892_ _1687_ _1684_ _0141_ VPWR VGND sg13g2_xor2_1
X_3912_ _0745_ net987 net941 net989 net938 VPWR VGND sg13g2_a22oi_1
X_3843_ _0678_ net993 net942 net994 net939 VPWR VGND sg13g2_a22oi_1
XFILLER_33_975 VPWR VGND sg13g2_decap_8
X_3774_ _0110_ _0598_ _0614_ VPWR VGND sg13g2_xnor2_1
X_5513_ _2246_ net491 _2244_ _2250_ VPWR VGND sg13g2_nand3_1
X_6493_ net1054 VGND VPWR _0034_ mac2.sum_lvl3_ff\[11\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_5444_ mac1.sum_lvl3_ff\[9\] net358 _2196_ VPWR VGND sg13g2_xor2_1
Xclkbuf_leaf_8_clk clknet_4_4_0_clk clknet_leaf_8_clk VPWR VGND sg13g2_buf_8
X_5375_ mac1.sum_lvl2_ff\[10\] mac1.sum_lvl2_ff\[29\] _2142_ VPWR VGND sg13g2_xor2_1
X_4326_ VGND VPWR _1142_ _1141_ _1140_ sg13g2_or2_1
X_4257_ _1075_ _1074_ _1071_ VPWR VGND sg13g2_nand2b_1
XFILLER_41_1012 VPWR VGND sg13g2_decap_8
X_3208_ _2753_ _2756_ _2799_ VPWR VGND sg13g2_nor2_1
X_4188_ _1009_ net880 net831 net882 net825 VPWR VGND sg13g2_a22oi_1
X_3139_ _2732_ _2725_ _2730_ _2731_ VPWR VGND sg13g2_and3_1
XFILLER_24_975 VPWR VGND sg13g2_decap_8
XFILLER_10_113 VPWR VGND sg13g2_fill_2
XFILLER_23_485 VPWR VGND sg13g2_fill_2
Xhold180 mac2.sum_lvl1_ff\[15\] VPWR VGND net220 sg13g2_dlygate4sd3_1
XFILLER_3_857 VPWR VGND sg13g2_decap_4
Xhold191 mac1.products_ff\[15\] VPWR VGND net231 sg13g2_dlygate4sd3_1
XFILLER_46_588 VPWR VGND sg13g2_fill_2
XFILLER_34_728 VPWR VGND sg13g2_fill_1
XFILLER_18_1003 VPWR VGND sg13g2_decap_8
XFILLER_42_783 VPWR VGND sg13g2_fill_2
XFILLER_15_997 VPWR VGND sg13g2_decap_8
XFILLER_30_967 VPWR VGND sg13g2_decap_8
X_3490_ _0335_ VPWR _0340_ VGND _0336_ _0338_ sg13g2_o21ai_1
X_5160_ _1892_ _1941_ _1943_ VPWR VGND sg13g2_and2_1
X_4111_ _0937_ _0916_ _0939_ VPWR VGND sg13g2_xor2_1
X_5091_ _1838_ _1837_ _1836_ _1876_ VPWR VGND sg13g2_a21o_2
X_4042_ _0870_ _0871_ _0872_ VPWR VGND sg13g2_nor2b_1
XFILLER_49_382 VPWR VGND sg13g2_fill_2
XFILLER_37_544 VPWR VGND sg13g2_fill_1
X_5993_ net277 _0241_ VPWR VGND sg13g2_buf_1
X_4944_ _0144_ _1729_ _1736_ VPWR VGND sg13g2_xnor2_1
XFILLER_24_249 VPWR VGND sg13g2_fill_1
X_4875_ _1671_ _1665_ _1670_ VPWR VGND sg13g2_xnor2_1
X_3826_ _0662_ _0650_ _0661_ VPWR VGND sg13g2_xnor2_1
XFILLER_21_978 VPWR VGND sg13g2_decap_8
X_3757_ VGND VPWR _0575_ _0589_ _0599_ _0588_ sg13g2_a21oi_1
X_3688_ _0533_ _0527_ _0532_ VPWR VGND sg13g2_xnor2_1
X_6476_ net1125 VGND VPWR net121 mac2.sum_lvl2_ff\[29\] clknet_leaf_39_clk sg13g2_dfrbpq_2
X_5427_ _2182_ mac1.sum_lvl3_ff\[26\] net501 VPWR VGND sg13g2_xnor2_1
X_5358_ net509 VPWR _2129_ VGND _2123_ _2127_ sg13g2_o21ai_1
X_4309_ VGND VPWR _1122_ _1123_ _1126_ _1104_ sg13g2_a21oi_1
X_5289_ _2033_ _2067_ _2068_ VPWR VGND sg13g2_nor2b_1
XFILLER_16_717 VPWR VGND sg13g2_fill_1
XFILLER_31_709 VPWR VGND sg13g2_fill_1
XFILLER_12_934 VPWR VGND sg13g2_decap_8
XFILLER_12_945 VPWR VGND sg13g2_fill_2
XFILLER_8_916 VPWR VGND sg13g2_fill_1
XFILLER_12_989 VPWR VGND sg13g2_decap_8
XFILLER_7_448 VPWR VGND sg13g2_fill_1
XFILLER_11_488 VPWR VGND sg13g2_fill_2
XFILLER_3_643 VPWR VGND sg13g2_fill_2
XFILLER_9_87 VPWR VGND sg13g2_fill_2
X_4660_ _1459_ _1458_ _1441_ _1462_ VPWR VGND sg13g2_a21o_1
X_3611_ _0407_ _0456_ _0458_ VPWR VGND sg13g2_and2_1
X_6330_ net1068 VGND VPWR _0004_ mac1.sum_lvl3_ff\[13\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_4591_ net848 net844 net897 net895 _1395_ VPWR VGND sg13g2_and4_1
X_3542_ _0353_ _0352_ _0351_ _0391_ VPWR VGND sg13g2_a21o_2
X_3473_ _0300_ VPWR _0323_ VGND _0275_ _0298_ sg13g2_o21ai_1
X_6261_ net1061 VGND VPWR net117 mac2.sum_lvl2_ff\[46\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_6192_ net1095 VGND VPWR net228 mac1.sum_lvl1_ff\[39\] clknet_leaf_55_clk sg13g2_dfrbpq_1
X_5212_ VGND VPWR _1957_ _1959_ _1994_ _1993_ sg13g2_a21oi_1
X_5143_ _1887_ VPWR _1926_ VGND _1842_ _1888_ sg13g2_o21ai_1
X_5074_ _1855_ _1856_ _1858_ _1859_ VPWR VGND sg13g2_or3_1
X_4025_ _0855_ net999 net1031 VPWR VGND sg13g2_nand2_1
XFILLER_38_842 VPWR VGND sg13g2_decap_8
X_5976_ net269 _0216_ VPWR VGND sg13g2_buf_1
X_4927_ _1721_ _1716_ _1719_ VPWR VGND sg13g2_xnor2_1
X_4858_ VGND VPWR _1619_ _1621_ _1655_ _1652_ sg13g2_a21oi_1
X_3809_ _0077_ _0632_ _0644_ VPWR VGND sg13g2_xnor2_1
X_4789_ _1588_ _1555_ _1587_ VPWR VGND sg13g2_nand2b_1
X_6459_ net1103 VGND VPWR net189 mac2.sum_lvl2_ff\[9\] clknet_leaf_43_clk sg13g2_dfrbpq_1
XFILLER_29_897 VPWR VGND sg13g2_decap_8
XFILLER_44_867 VPWR VGND sg13g2_decap_8
XFILLER_38_127 VPWR VGND sg13g2_fill_1
XFILLER_19_396 VPWR VGND sg13g2_fill_1
XFILLER_34_322 VPWR VGND sg13g2_fill_1
XFILLER_35_867 VPWR VGND sg13g2_decap_8
X_5830_ net822 net839 net787 _2523_ VPWR VGND sg13g2_mux2_1
X_5761_ VGND VPWR _2456_ _2455_ _2445_ sg13g2_or2_1
X_4712_ _1512_ net832 net902 net834 net900 VPWR VGND sg13g2_a22oi_1
X_5692_ _2390_ mac1.total_sum\[15\] mac2.total_sum\[15\] VPWR VGND sg13g2_xnor2_1
X_4643_ _1444_ _1411_ _1445_ VPWR VGND sg13g2_xor2_1
X_4574_ net844 net899 net847 _1379_ VPWR VGND net897 sg13g2_nand4_1
X_3525_ _0370_ _0371_ _0373_ _0374_ VPWR VGND sg13g2_or3_1
X_6313_ net1068 VGND VPWR net46 mac1.sum_lvl3_ff\[32\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_6244_ net1041 VGND VPWR net165 mac1.sum_lvl2_ff\[45\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3456_ _0303_ _0304_ _0306_ _0307_ VPWR VGND sg13g2_or3_1
X_3387_ _2969_ VPWR _2972_ VGND _2954_ _2971_ sg13g2_o21ai_1
X_6175_ net1122 VGND VPWR _0254_ DP_4.matrix\[38\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_5126_ _1907_ _1908_ _1890_ _1910_ VPWR VGND sg13g2_nand3_1
X_5057_ net866 net795 net868 _1842_ VPWR VGND net792 sg13g2_nand4_1
X_4008_ _0839_ _0833_ _0837_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_878 VPWR VGND sg13g2_fill_2
XFILLER_26_889 VPWR VGND sg13g2_decap_8
XFILLER_38_1017 VPWR VGND sg13g2_decap_8
XFILLER_38_1028 VPWR VGND sg13g2_fill_1
X_5959_ net977 _0191_ VPWR VGND sg13g2_buf_1
XFILLER_25_399 VPWR VGND sg13g2_fill_1
XFILLER_41_837 VPWR VGND sg13g2_decap_8
XFILLER_49_915 VPWR VGND sg13g2_decap_8
XFILLER_1_966 VPWR VGND sg13g2_decap_8
Xhold40 mac1.products_ff\[5\] VPWR VGND net80 sg13g2_dlygate4sd3_1
XFILLER_29_40 VPWR VGND sg13g2_fill_2
Xhold51 mac1.products_ff\[74\] VPWR VGND net91 sg13g2_dlygate4sd3_1
Xhold73 mac1.sum_lvl1_ff\[10\] VPWR VGND net113 sg13g2_dlygate4sd3_1
Xhold62 mac1.sum_lvl1_ff\[51\] VPWR VGND net102 sg13g2_dlygate4sd3_1
Xhold95 mac1.sum_lvl1_ff\[45\] VPWR VGND net135 sg13g2_dlygate4sd3_1
Xhold84 mac2.sum_lvl1_ff\[75\] VPWR VGND net124 sg13g2_dlygate4sd3_1
XFILLER_35_119 VPWR VGND sg13g2_fill_2
XFILLER_44_620 VPWR VGND sg13g2_fill_2
XFILLER_32_859 VPWR VGND sg13g2_decap_8
XFILLER_6_88 VPWR VGND sg13g2_fill_2
XFILLER_6_77 VPWR VGND sg13g2_fill_2
X_3310_ VGND VPWR _2861_ _2863_ _2899_ _2896_ sg13g2_a21oi_1
X_4290_ _1107_ net821 net879 VPWR VGND sg13g2_nand2_1
X_3241_ _2796_ _2831_ _2832_ VPWR VGND sg13g2_nor2_1
X_3172_ _2764_ net913 net970 VPWR VGND sg13g2_nand2_1
Xfanout1071 net1072 net1071 VPWR VGND sg13g2_buf_1
Xfanout1060 net1061 net1060 VPWR VGND sg13g2_buf_8
Xfanout1082 net1090 net1082 VPWR VGND sg13g2_buf_1
Xfanout1093 net1094 net1093 VPWR VGND sg13g2_buf_8
XFILLER_23_804 VPWR VGND sg13g2_fill_1
X_5813_ net875 _2472_ _2507_ VPWR VGND sg13g2_nor2_1
X_5744_ DP_2.matrix\[43\] net790 _2439_ VPWR VGND sg13g2_nor2_1
XFILLER_31_870 VPWR VGND sg13g2_decap_8
X_5675_ mac1.total_sum\[12\] mac2.total_sum\[12\] _2376_ VPWR VGND sg13g2_nor2_1
X_4626_ _1427_ _1426_ _1409_ _1429_ VPWR VGND sg13g2_a21o_1
X_4557_ _0133_ _1358_ _1365_ VPWR VGND sg13g2_xnor2_1
X_4488_ _1300_ _1295_ _1298_ VPWR VGND sg13g2_xnor2_1
X_3508_ net1017 net946 net1020 _0357_ VPWR VGND net944 sg13g2_nand4_1
XFILLER_44_1021 VPWR VGND sg13g2_decap_8
X_3439_ _0270_ VPWR _0291_ VGND _2989_ _0271_ sg13g2_o21ai_1
X_6227_ net1109 VGND VPWR net178 mac1.sum_lvl2_ff\[25\] clknet_leaf_51_clk sg13g2_dfrbpq_1
X_6158_ net1081 VGND VPWR _0241_ DP_3.matrix\[77\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_5109_ _1893_ net802 net856 VPWR VGND sg13g2_nand2_1
XFILLER_46_929 VPWR VGND sg13g2_decap_8
XFILLER_17_108 VPWR VGND sg13g2_fill_2
X_6089_ net1073 VGND VPWR _0195_ DP_1.matrix\[79\] clknet_leaf_59_clk sg13g2_dfrbpq_1
XFILLER_26_664 VPWR VGND sg13g2_decap_4
XFILLER_40_199 VPWR VGND sg13g2_fill_1
Xoutput30 net30 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_37_907 VPWR VGND sg13g2_decap_8
XFILLER_45_973 VPWR VGND sg13g2_decap_8
XFILLER_44_472 VPWR VGND sg13g2_fill_1
XFILLER_44_461 VPWR VGND sg13g2_decap_4
XFILLER_17_675 VPWR VGND sg13g2_fill_1
XFILLER_32_656 VPWR VGND sg13g2_fill_2
X_3790_ _0628_ net1000 net943 net940 net1002 VPWR VGND sg13g2_a22oi_1
XFILLER_13_870 VPWR VGND sg13g2_fill_1
X_5460_ _2203_ _2200_ _2209_ VPWR VGND _2202_ sg13g2_nand3b_1
X_4411_ _1200_ VPWR _1225_ VGND _1198_ _1201_ sg13g2_o21ai_1
X_5391_ _2149_ VPWR _2155_ VGND _2150_ _2154_ sg13g2_o21ai_1
X_4342_ net826 net871 net829 _1158_ VPWR VGND net1026 sg13g2_nand4_1
XFILLER_28_1027 VPWR VGND sg13g2_fill_2
X_4273_ _1088_ _1087_ _1070_ _1091_ VPWR VGND sg13g2_a21o_1
X_3224_ _2815_ _2763_ _2812_ VPWR VGND sg13g2_xnor2_1
X_6012_ net1056 VGND VPWR net9 DP_3.Q_range.out_data\[2\] clknet_leaf_22_clk sg13g2_dfrbpq_2
.ends

