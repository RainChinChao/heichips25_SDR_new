module heichips25_template (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \DP_1.matrix[0] ;
 wire \DP_1.matrix[112] ;
 wire \DP_1.matrix[113] ;
 wire \DP_1.matrix[128] ;
 wire \DP_1.matrix[129] ;
 wire \DP_1.matrix[16] ;
 wire \DP_1.matrix[17] ;
 wire \DP_1.matrix[1] ;
 wire \DP_1.matrix[32] ;
 wire \DP_1.matrix[33] ;
 wire \DP_1.matrix[48] ;
 wire \DP_1.matrix[49] ;
 wire \DP_1.matrix[64] ;
 wire \DP_1.matrix[65] ;
 wire \DP_1.matrix[80] ;
 wire \DP_1.matrix[81] ;
 wire \DP_1.matrix[96] ;
 wire \DP_1.matrix[97] ;
 wire \DP_2.matrix[0] ;
 wire \DP_2.matrix[112] ;
 wire \DP_2.matrix[113] ;
 wire \DP_2.matrix[128] ;
 wire \DP_2.matrix[129] ;
 wire \DP_2.matrix[16] ;
 wire \DP_2.matrix[17] ;
 wire \DP_2.matrix[1] ;
 wire \DP_2.matrix[32] ;
 wire \DP_2.matrix[33] ;
 wire \DP_2.matrix[48] ;
 wire \DP_2.matrix[49] ;
 wire \DP_2.matrix[64] ;
 wire \DP_2.matrix[65] ;
 wire \DP_2.matrix[80] ;
 wire \DP_2.matrix[81] ;
 wire \DP_2.matrix[96] ;
 wire \DP_2.matrix[97] ;
 wire \DP_3.matrix[0] ;
 wire \DP_3.matrix[112] ;
 wire \DP_3.matrix[113] ;
 wire \DP_3.matrix[128] ;
 wire \DP_3.matrix[129] ;
 wire \DP_3.matrix[16] ;
 wire \DP_3.matrix[17] ;
 wire \DP_3.matrix[1] ;
 wire \DP_3.matrix[32] ;
 wire \DP_3.matrix[33] ;
 wire \DP_3.matrix[48] ;
 wire \DP_3.matrix[49] ;
 wire \DP_3.matrix[64] ;
 wire \DP_3.matrix[65] ;
 wire \DP_3.matrix[80] ;
 wire \DP_3.matrix[81] ;
 wire \DP_3.matrix[96] ;
 wire \DP_3.matrix[97] ;
 wire \DP_4.matrix[0] ;
 wire \DP_4.matrix[112] ;
 wire \DP_4.matrix[113] ;
 wire \DP_4.matrix[128] ;
 wire \DP_4.matrix[129] ;
 wire \DP_4.matrix[16] ;
 wire \DP_4.matrix[17] ;
 wire \DP_4.matrix[1] ;
 wire \DP_4.matrix[32] ;
 wire \DP_4.matrix[33] ;
 wire \DP_4.matrix[48] ;
 wire \DP_4.matrix[49] ;
 wire \DP_4.matrix[64] ;
 wire \DP_4.matrix[65] ;
 wire \DP_4.matrix[80] ;
 wire \DP_4.matrix[81] ;
 wire \DP_4.matrix[96] ;
 wire \DP_4.matrix[97] ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire \mac1.products_ff[0] ;
 wire \mac1.products_ff[112] ;
 wire \mac1.products_ff[113] ;
 wire \mac1.products_ff[128] ;
 wire \mac1.products_ff[129] ;
 wire \mac1.products_ff[16] ;
 wire \mac1.products_ff[17] ;
 wire \mac1.products_ff[1] ;
 wire \mac1.products_ff[32] ;
 wire \mac1.products_ff[33] ;
 wire \mac1.products_ff[48] ;
 wire \mac1.products_ff[49] ;
 wire \mac1.products_ff[64] ;
 wire \mac1.products_ff[65] ;
 wire \mac1.products_ff[80] ;
 wire \mac1.products_ff[81] ;
 wire \mac1.products_ff[96] ;
 wire \mac1.products_ff[97] ;
 wire \mac1.sum_lvl1_ff[0] ;
 wire \mac1.sum_lvl1_ff[16] ;
 wire \mac1.sum_lvl1_ff[17] ;
 wire \mac1.sum_lvl1_ff[1] ;
 wire \mac1.sum_lvl1_ff[24] ;
 wire \mac1.sum_lvl1_ff[25] ;
 wire \mac1.sum_lvl1_ff[32] ;
 wire \mac1.sum_lvl1_ff[33] ;
 wire \mac1.sum_lvl1_ff[8] ;
 wire \mac1.sum_lvl1_ff[9] ;
 wire \mac1.sum_lvl2_ff[0] ;
 wire \mac1.sum_lvl2_ff[1] ;
 wire \mac1.sum_lvl2_ff[4] ;
 wire \mac1.sum_lvl2_ff[5] ;
 wire \mac1.sum_lvl2_ff[8] ;
 wire \mac1.sum_lvl2_ff[9] ;
 wire \mac1.sum_lvl3_ff[0] ;
 wire \mac1.sum_lvl3_ff[1] ;
 wire \mac1.sum_lvl3_ff[2] ;
 wire \mac1.sum_lvl3_ff[3] ;
 wire \mac1.total_sum[0] ;
 wire \mac1.total_sum[1] ;
 wire \mac1.total_sum[2] ;
 wire \mac2.products_ff[0] ;
 wire \mac2.products_ff[112] ;
 wire \mac2.products_ff[113] ;
 wire \mac2.products_ff[128] ;
 wire \mac2.products_ff[129] ;
 wire \mac2.products_ff[16] ;
 wire \mac2.products_ff[17] ;
 wire \mac2.products_ff[1] ;
 wire \mac2.products_ff[32] ;
 wire \mac2.products_ff[33] ;
 wire \mac2.products_ff[48] ;
 wire \mac2.products_ff[49] ;
 wire \mac2.products_ff[64] ;
 wire \mac2.products_ff[65] ;
 wire \mac2.products_ff[80] ;
 wire \mac2.products_ff[81] ;
 wire \mac2.products_ff[96] ;
 wire \mac2.products_ff[97] ;
 wire \mac2.sum_lvl1_ff[0] ;
 wire \mac2.sum_lvl1_ff[16] ;
 wire \mac2.sum_lvl1_ff[17] ;
 wire \mac2.sum_lvl1_ff[1] ;
 wire \mac2.sum_lvl1_ff[24] ;
 wire \mac2.sum_lvl1_ff[25] ;
 wire \mac2.sum_lvl1_ff[32] ;
 wire \mac2.sum_lvl1_ff[33] ;
 wire \mac2.sum_lvl1_ff[8] ;
 wire \mac2.sum_lvl1_ff[9] ;
 wire \mac2.sum_lvl2_ff[0] ;
 wire \mac2.sum_lvl2_ff[1] ;
 wire \mac2.sum_lvl2_ff[4] ;
 wire \mac2.sum_lvl2_ff[5] ;
 wire \mac2.sum_lvl2_ff[8] ;
 wire \mac2.sum_lvl2_ff[9] ;
 wire \mac2.sum_lvl3_ff[0] ;
 wire \mac2.sum_lvl3_ff[1] ;
 wire \mac2.sum_lvl3_ff[2] ;
 wire \mac2.sum_lvl3_ff[3] ;
 wire \mac2.total_sum[0] ;
 wire \mac2.total_sum[1] ;
 wire \mac2.total_sum[2] ;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire clknet_0_clk;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net5;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;

 sg13g2_and2_1 _222_ (.A(net155),
    .B(net125),
    .X(_034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _223_ (.A(net124),
    .B(net142),
    .X(_036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _224_ (.A(net144),
    .B(net138),
    .X(_038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _225_ (.A(net136),
    .B(net137),
    .X(_040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _226_ (.A(net154),
    .B(net156),
    .X(_042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _227_ (.A(net143),
    .B(net146),
    .X(_044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _228_ (.A(net151),
    .B(net140),
    .X(_046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _229_ (.A(net162),
    .B(net158),
    .X(_048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _230_ (.A(net131),
    .B(net157),
    .X(_050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _231_ (.A(net164),
    .B(net132),
    .X(_052_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _232_ (.A(net160),
    .B(net123),
    .X(_054_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _233_ (.A(net128),
    .B(net135),
    .X(_056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _234_ (.A(net119),
    .B(net150),
    .X(_058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _235_ (.A(net134),
    .B(net141),
    .X(_060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _236_ (.A(net159),
    .B(net120),
    .X(_062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _237_ (.A(net145),
    .B(net149),
    .X(_064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _238_ (.A(net139),
    .B(net163),
    .X(_066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _239_ (.A(net133),
    .B(net161),
    .X(_068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _240_ (.Y(_142_),
    .A(\mac1.total_sum[0] ),
    .B(\mac2.total_sum[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _241_ (.Y(_143_),
    .A(\mac1.total_sum[1] ),
    .B(\mac2.total_sum[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _242_ (.A(\mac1.total_sum[1] ),
    .B(\mac2.total_sum[1] ),
    .Y(_144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _243_ (.B(\mac2.total_sum[1] ),
    .A(\mac1.total_sum[1] ),
    .X(_145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _244_ (.Y(net2),
    .A(_142_),
    .B(_145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _245_ (.B1(_143_),
    .VDD(VPWR),
    .Y(_146_),
    .VSS(VGND),
    .A1(_142_),
    .A2(_144_));
 sg13g2_and2_1 _246_ (.A(\mac1.total_sum[2] ),
    .B(\mac2.total_sum[2] ),
    .X(_147_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _247_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_148_),
    .B(\mac2.total_sum[2] ),
    .A(\mac1.total_sum[2] ));
 sg13g2_nand2b_1 _248_ (.Y(_149_),
    .B(_148_),
    .A_N(_147_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _249_ (.Y(net3),
    .A(_146_),
    .B(_149_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _250_ (.B(\mac2.total_sum[0] ),
    .A(\mac1.total_sum[0] ),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _251_ (.Y(_150_),
    .A(net178),
    .B(net126),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _252_ (.B(\mac1.products_ff[17] ),
    .A(\mac1.products_ff[1] ),
    .X(_151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _253_ (.Y(_001_),
    .A(_150_),
    .B(_151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _254_ (.B(net126),
    .A(\mac1.products_ff[0] ),
    .X(_000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _255_ (.Y(_152_),
    .A(net203),
    .B(net115),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _256_ (.B(\mac1.sum_lvl2_ff[1] ),
    .A(\mac1.sum_lvl2_ff[5] ),
    .X(_153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _257_ (.Y(_013_),
    .A(_152_),
    .B(_153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _258_ (.B(net115),
    .A(\mac1.sum_lvl2_ff[4] ),
    .X(_012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _259_ (.Y(_154_),
    .A(net173),
    .B(net102),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _260_ (.B(\mac1.sum_lvl1_ff[17] ),
    .A(\mac1.sum_lvl1_ff[25] ),
    .X(_155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _261_ (.Y(_011_),
    .A(_154_),
    .B(_155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _262_ (.B(net102),
    .A(\mac1.sum_lvl1_ff[24] ),
    .X(_010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _263_ (.Y(_156_),
    .A(net191),
    .B(net129),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _264_ (.B(\mac1.sum_lvl1_ff[1] ),
    .A(\mac1.sum_lvl1_ff[9] ),
    .X(_157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _265_ (.Y(_009_),
    .A(_156_),
    .B(_157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _266_ (.B(net129),
    .A(\mac1.sum_lvl1_ff[8] ),
    .X(_008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _267_ (.Y(_158_),
    .A(\mac1.products_ff[112] ),
    .B(net37),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _268_ (.B(net193),
    .A(\mac1.products_ff[113] ),
    .X(_159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _269_ (.Y(_007_),
    .A(_158_),
    .B(net194),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _270_ (.B(net37),
    .A(\mac1.products_ff[112] ),
    .X(_006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _271_ (.Y(_160_),
    .A(\mac1.products_ff[80] ),
    .B(net97),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _272_ (.B(net188),
    .A(\mac1.products_ff[81] ),
    .X(_161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _273_ (.Y(_005_),
    .A(_160_),
    .B(net189),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _274_ (.B(net97),
    .A(\mac1.products_ff[80] ),
    .X(_004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _275_ (.Y(_162_),
    .A(net182),
    .B(net109),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _276_ (.B(\mac1.products_ff[49] ),
    .A(\mac1.products_ff[33] ),
    .X(_163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _277_ (.Y(_003_),
    .A(_162_),
    .B(_163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _278_ (.B(net109),
    .A(\mac1.products_ff[32] ),
    .X(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _279_ (.Y(_164_),
    .A(net201),
    .B(net147),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _280_ (.B(\mac2.products_ff[1] ),
    .A(\mac2.products_ff[17] ),
    .X(_165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _281_ (.Y(_018_),
    .A(_164_),
    .B(_165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _282_ (.B(net147),
    .A(\mac2.products_ff[16] ),
    .X(_017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _283_ (.Y(_166_),
    .A(net205),
    .B(net165),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _284_ (.Y(_167_),
    .A(net167),
    .B(\mac1.sum_lvl3_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _285_ (.A(net167),
    .B(\mac1.sum_lvl3_ff[1] ),
    .Y(_168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _286_ (.B(\mac1.sum_lvl3_ff[1] ),
    .A(net167),
    .X(_169_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _287_ (.Y(_016_),
    .A(_166_),
    .B(_169_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _288_ (.B(net165),
    .A(\mac1.sum_lvl3_ff[2] ),
    .X(_015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _289_ (.Y(_170_),
    .A(net196),
    .B(net152),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _290_ (.B(\mac2.sum_lvl2_ff[1] ),
    .A(\mac2.sum_lvl2_ff[5] ),
    .X(_171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _291_ (.Y(_030_),
    .A(_170_),
    .B(_171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _292_ (.B(net152),
    .A(\mac2.sum_lvl2_ff[4] ),
    .X(_029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _293_ (.Y(_172_),
    .A(net186),
    .B(net105),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _294_ (.B(\mac2.sum_lvl1_ff[17] ),
    .A(\mac2.sum_lvl1_ff[25] ),
    .X(_173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _295_ (.Y(_028_),
    .A(_172_),
    .B(_173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _296_ (.B(net105),
    .A(\mac2.sum_lvl1_ff[24] ),
    .X(_027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _297_ (.Y(_174_),
    .A(net121),
    .B(\mac2.sum_lvl1_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _298_ (.B(net198),
    .A(\mac2.sum_lvl1_ff[9] ),
    .X(_175_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _299_ (.Y(_026_),
    .A(_174_),
    .B(net199),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _300_ (.B(\mac2.sum_lvl1_ff[0] ),
    .A(net121),
    .X(_025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _301_ (.Y(_176_),
    .A(net180),
    .B(net113),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _302_ (.B(\mac2.products_ff[113] ),
    .A(\mac2.products_ff[97] ),
    .X(_177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _303_ (.Y(_024_),
    .A(_176_),
    .B(_177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _304_ (.B(net113),
    .A(\mac2.products_ff[96] ),
    .X(_023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _305_ (.Y(_178_),
    .A(net111),
    .B(\mac2.products_ff[80] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _306_ (.B(net175),
    .A(\mac2.products_ff[65] ),
    .X(_179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _307_ (.Y(_022_),
    .A(_178_),
    .B(net176),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _308_ (.B(\mac2.products_ff[80] ),
    .A(net111),
    .X(_021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _309_ (.Y(_180_),
    .A(net184),
    .B(net117),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _310_ (.B(\mac2.products_ff[33] ),
    .A(\mac2.products_ff[49] ),
    .X(_181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _311_ (.Y(_020_),
    .A(_180_),
    .B(_181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _312_ (.B(net117),
    .A(\mac2.products_ff[48] ),
    .X(_019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _313_ (.Y(_182_),
    .A(net207),
    .B(net107),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _314_ (.Y(_183_),
    .A(net170),
    .B(\mac2.sum_lvl3_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _315_ (.A(net170),
    .B(\mac2.sum_lvl3_ff[3] ),
    .Y(_184_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _316_ (.B(\mac2.sum_lvl3_ff[3] ),
    .A(net170),
    .X(_185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _317_ (.Y(_033_),
    .A(_182_),
    .B(_185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _318_ (.B(net107),
    .A(\mac2.sum_lvl3_ff[0] ),
    .X(_032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _319_ (.Y(_186_),
    .A(net155),
    .B(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _320_ (.Y(_187_),
    .A(net125),
    .B(net41),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _321_ (.B(_187_),
    .A(_186_),
    .X(_035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _322_ (.Y(_188_),
    .A(net124),
    .B(net87),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _323_ (.Y(_189_),
    .A(net142),
    .B(net83),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _324_ (.B(_189_),
    .A(_188_),
    .X(_037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _325_ (.A2(_148_),
    .A1(_146_),
    .B1(_147_),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _326_ (.Y(_190_),
    .A(net144),
    .B(net52),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _327_ (.Y(_191_),
    .A(net138),
    .B(net50),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _328_ (.B(_191_),
    .A(_190_),
    .X(_039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _329_ (.Y(_192_),
    .A(net136),
    .B(net85),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _330_ (.Y(_193_),
    .A(net137),
    .B(net94),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _331_ (.B(_193_),
    .A(_192_),
    .X(_041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _332_ (.Y(_194_),
    .A(net46),
    .B(net156),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _333_ (.Y(_195_),
    .A(net154),
    .B(net55),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _334_ (.B(_195_),
    .A(_194_),
    .X(_043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _335_ (.Y(_196_),
    .A(net143),
    .B(net45),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _336_ (.Y(_197_),
    .A(net146),
    .B(net51),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _337_ (.B(_197_),
    .A(_196_),
    .X(_045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _338_ (.Y(_198_),
    .A(net48),
    .B(net140),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _339_ (.Y(_199_),
    .A(net151),
    .B(net95),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _340_ (.B(_199_),
    .A(_198_),
    .X(_047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _341_ (.Y(_200_),
    .A(net89),
    .B(net158),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _342_ (.Y(_201_),
    .A(net162),
    .B(net84),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _343_ (.B(_201_),
    .A(_200_),
    .X(_049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _344_ (.Y(_202_),
    .A(net101),
    .B(net157),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _345_ (.Y(_203_),
    .A(net131),
    .B(net91),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _346_ (.B(_203_),
    .A(_202_),
    .X(_051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _347_ (.Y(_204_),
    .A(net86),
    .B(net132),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _348_ (.Y(_205_),
    .A(net164),
    .B(net100),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _349_ (.B(_205_),
    .A(_204_),
    .X(_053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _350_ (.Y(_206_),
    .A(net92),
    .B(net123),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _351_ (.Y(_207_),
    .A(net160),
    .B(net53),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _352_ (.B(_207_),
    .A(_206_),
    .X(_055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _353_ (.Y(_208_),
    .A(net40),
    .B(net135),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _354_ (.Y(_209_),
    .A(net128),
    .B(net49),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _355_ (.B(_209_),
    .A(_208_),
    .X(_057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _356_ (.B1(net168),
    .VDD(VPWR),
    .Y(_014_),
    .VSS(VGND),
    .A1(_166_),
    .A2(_168_));
 sg13g2_nand2_1 _357_ (.Y(_210_),
    .A(net104),
    .B(net150),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _358_ (.Y(_211_),
    .A(net119),
    .B(net96),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _359_ (.B(_211_),
    .A(_210_),
    .X(_059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _360_ (.Y(_212_),
    .A(net134),
    .B(net93),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _361_ (.Y(_213_),
    .A(net141),
    .B(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _362_ (.B(_213_),
    .A(_212_),
    .X(_061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _363_ (.Y(_214_),
    .A(net47),
    .B(net120),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _364_ (.Y(_215_),
    .A(net159),
    .B(net88),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _365_ (.B(_215_),
    .A(_214_),
    .X(_063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _366_ (.Y(_216_),
    .A(net145),
    .B(net42),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _367_ (.Y(_217_),
    .A(net149),
    .B(net90),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _368_ (.B(_217_),
    .A(_216_),
    .X(_065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _369_ (.Y(_218_),
    .A(net139),
    .B(net99),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _370_ (.Y(_219_),
    .A(net163),
    .B(net54),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _371_ (.B(_219_),
    .A(_218_),
    .X(_067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _372_ (.Y(_220_),
    .A(net133),
    .B(net82),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _373_ (.Y(_221_),
    .A(net161),
    .B(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _374_ (.B(_221_),
    .A(_220_),
    .X(_069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _375_ (.B1(net171),
    .VDD(VPWR),
    .Y(_031_),
    .VSS(VGND),
    .A1(_182_),
    .A2(_184_));
 sg13g2_buf_1 _376_ (.A(net154),
    .X(_070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _377_ (.A(net46),
    .X(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _378_ (.A(net128),
    .X(_072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _379_ (.A(net40),
    .X(_073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _380_ (.A(net160),
    .X(_074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _381_ (.A(net92),
    .X(_075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _382_ (.A(net164),
    .X(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _383_ (.A(net86),
    .X(_077_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _384_ (.A(net131),
    .X(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _385_ (.A(net101),
    .X(_079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _386_ (.A(net162),
    .X(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _387_ (.A(net89),
    .X(_081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _388_ (.A(net151),
    .X(_082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _389_ (.A(net48),
    .X(_083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _390_ (.A(net159),
    .X(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _391_ (.A(net47),
    .X(_085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _392_ (.A(net119),
    .X(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _393_ (.A(net104),
    .X(_087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _394_ (.A(net156),
    .X(_088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _395_ (.A(net55),
    .X(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _396_ (.A(net135),
    .X(_090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _397_ (.A(net49),
    .X(_091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _398_ (.A(net123),
    .X(_092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _399_ (.A(net53),
    .X(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _400_ (.A(net132),
    .X(_094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _401_ (.A(net100),
    .X(_095_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _402_ (.A(net157),
    .X(_096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _403_ (.A(net91),
    .X(_097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _404_ (.A(net158),
    .X(_098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _405_ (.A(net84),
    .X(_099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _406_ (.A(net140),
    .X(_100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _407_ (.A(net95),
    .X(_101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _408_ (.A(net120),
    .X(_102_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _409_ (.A(net88),
    .X(_103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _410_ (.A(net150),
    .X(_104_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _411_ (.A(net96),
    .X(_105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _412_ (.A(net146),
    .X(_106_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _413_ (.A(net45),
    .X(_107_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _414_ (.A(net161),
    .X(_108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _415_ (.A(net82),
    .X(_109_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _416_ (.A(net163),
    .X(_110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _417_ (.A(net99),
    .X(_111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _418_ (.A(net149),
    .X(_112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _419_ (.A(net42),
    .X(_113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _420_ (.A(net141),
    .X(_114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _421_ (.A(net93),
    .X(_115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _422_ (.A(net138),
    .X(_116_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _423_ (.A(net52),
    .X(_117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _424_ (.A(net137),
    .X(_118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _425_ (.A(net85),
    .X(_119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _426_ (.A(net125),
    .X(_120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _427_ (.A(net43),
    .X(_121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _428_ (.A(net142),
    .X(_122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _429_ (.A(net87),
    .X(_123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _430_ (.A(net143),
    .X(_124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _431_ (.A(net51),
    .X(_125_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _432_ (.A(net133),
    .X(_126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _433_ (.A(net39),
    .X(_127_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _434_ (.A(net139),
    .X(_128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _435_ (.A(net54),
    .X(_129_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _436_ (.A(net145),
    .X(_130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _437_ (.A(net90),
    .X(_131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _438_ (.A(net134),
    .X(_132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _439_ (.A(net44),
    .X(_133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _440_ (.A(net144),
    .X(_134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _441_ (.A(net50),
    .X(_135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _442_ (.A(net136),
    .X(_136_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _443_ (.A(net94),
    .X(_137_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _444_ (.A(net155),
    .X(_138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _445_ (.A(net41),
    .X(_139_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _446_ (.A(net124),
    .X(_140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _447_ (.A(net83),
    .X(_141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbpq_1 _448_ (.RESET_B(net72),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_070_),
    .Q(\DP_1.matrix[0] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _449_ (.RESET_B(net72),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_071_),
    .Q(\DP_1.matrix[1] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _450_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_072_),
    .Q(\DP_1.matrix[16] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _451_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_073_),
    .Q(\DP_1.matrix[17] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _452_ (.RESET_B(net69),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_074_),
    .Q(\DP_1.matrix[32] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _453_ (.RESET_B(net69),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_075_),
    .Q(\DP_1.matrix[33] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _454_ (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_076_),
    .Q(\DP_1.matrix[48] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _455_ (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_077_),
    .Q(\DP_1.matrix[49] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _456_ (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_078_),
    .Q(\DP_1.matrix[64] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _457_ (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_079_),
    .Q(\DP_1.matrix[65] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _458_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_080_),
    .Q(\DP_1.matrix[80] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _459_ (.RESET_B(net80),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_081_),
    .Q(\DP_1.matrix[81] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _460_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_082_),
    .Q(\DP_1.matrix[96] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _461_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_083_),
    .Q(\DP_1.matrix[97] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _462_ (.RESET_B(net62),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_084_),
    .Q(\DP_1.matrix[112] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _463_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_085_),
    .Q(\DP_1.matrix[113] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _464_ (.RESET_B(net56),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_086_),
    .Q(\DP_1.matrix[128] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _465_ (.RESET_B(net56),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_087_),
    .Q(\DP_1.matrix[129] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _466_ (.RESET_B(net72),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_088_),
    .Q(\DP_2.matrix[0] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _467_ (.RESET_B(net72),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_089_),
    .Q(\DP_2.matrix[1] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _468_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_090_),
    .Q(\DP_2.matrix[16] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _469_ (.RESET_B(net74),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_091_),
    .Q(\DP_2.matrix[17] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _470_ (.RESET_B(net69),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_092_),
    .Q(\DP_2.matrix[32] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _471_ (.RESET_B(net69),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_093_),
    .Q(\DP_2.matrix[33] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _472_ (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_094_),
    .Q(\DP_2.matrix[48] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _473_ (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_095_),
    .Q(\DP_2.matrix[49] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _474_ (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_096_),
    .Q(\DP_2.matrix[64] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _475_ (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_097_),
    .Q(\DP_2.matrix[65] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _476_ (.RESET_B(net78),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_098_),
    .Q(\DP_2.matrix[80] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _477_ (.RESET_B(net78),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_099_),
    .Q(\DP_2.matrix[81] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _478_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_100_),
    .Q(\DP_2.matrix[96] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _479_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_101_),
    .Q(\DP_2.matrix[97] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _480_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_102_),
    .Q(\DP_2.matrix[112] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _481_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_103_),
    .Q(\DP_2.matrix[113] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _482_ (.RESET_B(net59),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_104_),
    .Q(\DP_2.matrix[128] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _483_ (.RESET_B(net59),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_105_),
    .Q(\DP_2.matrix[129] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _484_ (.RESET_B(net78),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_106_),
    .Q(\DP_3.matrix[0] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _485_ (.RESET_B(net78),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_107_),
    .Q(\DP_3.matrix[1] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _486_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_108_),
    .Q(\DP_3.matrix[16] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _487_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_109_),
    .Q(\DP_3.matrix[17] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _488_ (.RESET_B(net76),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_110_),
    .Q(\DP_3.matrix[32] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _489_ (.RESET_B(net76),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_111_),
    .Q(\DP_3.matrix[33] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _490_ (.RESET_B(net66),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_112_),
    .Q(\DP_3.matrix[48] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _491_ (.RESET_B(net66),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_113_),
    .Q(\DP_3.matrix[49] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _492_ (.RESET_B(net68),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_114_),
    .Q(\DP_3.matrix[64] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _493_ (.RESET_B(net63),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_115_),
    .Q(\DP_3.matrix[65] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _494_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_116_),
    .Q(\DP_3.matrix[80] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _495_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_117_),
    .Q(\DP_3.matrix[81] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _496_ (.RESET_B(net63),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_118_),
    .Q(\DP_3.matrix[96] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _497_ (.RESET_B(net63),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_119_),
    .Q(\DP_3.matrix[97] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _498_ (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_120_),
    .Q(\DP_3.matrix[112] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _499_ (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_121_),
    .Q(\DP_3.matrix[113] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _500_ (.RESET_B(net57),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_122_),
    .Q(\DP_3.matrix[128] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _501_ (.RESET_B(net57),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_123_),
    .Q(\DP_3.matrix[129] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _502_ (.RESET_B(net78),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_124_),
    .Q(\DP_4.matrix[0] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _503_ (.RESET_B(net78),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_125_),
    .Q(\DP_4.matrix[1] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _504_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_126_),
    .Q(\DP_4.matrix[16] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _505_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_127_),
    .Q(\DP_4.matrix[17] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _506_ (.RESET_B(net76),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_128_),
    .Q(\DP_4.matrix[32] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _507_ (.RESET_B(net76),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_129_),
    .Q(\DP_4.matrix[33] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _508_ (.RESET_B(net66),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_130_),
    .Q(\DP_4.matrix[48] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _509_ (.RESET_B(net66),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_131_),
    .Q(\DP_4.matrix[49] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _510_ (.RESET_B(net68),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_132_),
    .Q(\DP_4.matrix[64] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _511_ (.RESET_B(net63),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_133_),
    .Q(\DP_4.matrix[65] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _512_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_134_),
    .Q(\DP_4.matrix[80] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _513_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_135_),
    .Q(\DP_4.matrix[81] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _514_ (.RESET_B(net63),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_136_),
    .Q(\DP_4.matrix[96] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _515_ (.RESET_B(net63),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_137_),
    .Q(\DP_4.matrix[97] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _516_ (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_138_),
    .Q(\DP_4.matrix[112] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _517_ (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_139_),
    .Q(\DP_4.matrix[113] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _518_ (.RESET_B(net57),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_140_),
    .Q(\DP_4.matrix[128] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _519_ (.RESET_B(net57),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_141_),
    .Q(\DP_4.matrix[129] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _520_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_048_),
    .Q(\mac1.products_ff[80] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _521_ (.RESET_B(net78),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_049_),
    .Q(\mac1.products_ff[81] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _522_ (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_050_),
    .Q(\mac1.products_ff[64] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _523_ (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_051_),
    .Q(\mac1.products_ff[65] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _524_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net127),
    .Q(\mac1.sum_lvl1_ff[0] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _525_ (.RESET_B(net72),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net179),
    .Q(\mac1.sum_lvl1_ff[1] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _526_ (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net110),
    .Q(\mac1.sum_lvl1_ff[8] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _527_ (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net183),
    .Q(\mac1.sum_lvl1_ff[9] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _528_ (.RESET_B(net59),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_058_),
    .Q(\mac1.products_ff[128] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _529_ (.RESET_B(net61),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_059_),
    .Q(\mac1.products_ff[129] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _530_ (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net98),
    .Q(\mac1.sum_lvl1_ff[16] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _531_ (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net190),
    .Q(\mac1.sum_lvl1_ff[17] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _532_ (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_052_),
    .Q(\mac1.products_ff[48] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _533_ (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_053_),
    .Q(\mac1.products_ff[49] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _534_ (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net38),
    .Q(\mac1.sum_lvl1_ff[24] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _535_ (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net195),
    .Q(\mac1.sum_lvl1_ff[25] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _536_ (.RESET_B(net61),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net35),
    .Q(\mac1.sum_lvl1_ff[32] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _537_ (.RESET_B(net61),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net27),
    .Q(\mac1.sum_lvl1_ff[33] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _538_ (.RESET_B(net62),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_062_),
    .Q(\mac1.products_ff[112] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _539_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_063_),
    .Q(\mac1.products_ff[113] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _540_ (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_054_),
    .Q(\mac1.products_ff[32] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _541_ (.RESET_B(net69),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_055_),
    .Q(\mac1.products_ff[33] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _542_ (.RESET_B(net69),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net130),
    .Q(\mac1.sum_lvl2_ff[0] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _543_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net192),
    .Q(\mac1.sum_lvl2_ff[1] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _544_ (.RESET_B(net74),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_056_),
    .Q(\mac1.products_ff[16] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _545_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_057_),
    .Q(\mac1.products_ff[17] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _546_ (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net103),
    .Q(\mac1.sum_lvl2_ff[4] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _547_ (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net174),
    .Q(\mac1.sum_lvl2_ff[5] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _548_ (.RESET_B(net61),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net34),
    .Q(\mac1.sum_lvl2_ff[8] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _549_ (.RESET_B(net61),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net26),
    .Q(\mac1.sum_lvl2_ff[9] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _550_ (.RESET_B(net72),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_042_),
    .Q(\mac1.products_ff[0] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _551_ (.RESET_B(net72),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_043_),
    .Q(\mac1.products_ff[1] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _552_ (.RESET_B(net75),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_046_),
    .Q(\mac1.products_ff[96] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _553_ (.RESET_B(net75),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_047_),
    .Q(\mac1.products_ff[97] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _554_ (.RESET_B(net56),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net166),
    .Q(\mac1.total_sum[0] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _555_ (.RESET_B(net56),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net206),
    .Q(\mac1.total_sum[1] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _556_ (.RESET_B(net56),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net169),
    .Q(\mac1.total_sum[2] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _557_ (.RESET_B(net69),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net116),
    .Q(\mac1.sum_lvl3_ff[0] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _558_ (.RESET_B(net69),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net204),
    .Q(\mac1.sum_lvl3_ff[1] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _559_ (.RESET_B(net61),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net31),
    .Q(\mac1.sum_lvl3_ff[2] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _560_ (.RESET_B(net61),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net29),
    .Q(\mac1.sum_lvl3_ff[3] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _561_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_038_),
    .Q(\mac2.products_ff[80] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _562_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_039_),
    .Q(\mac2.products_ff[81] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _563_ (.RESET_B(net63),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_060_),
    .Q(\mac2.products_ff[64] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _564_ (.RESET_B(net68),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_061_),
    .Q(\mac2.products_ff[65] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_2 _565_ (.RESET_B(net78),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net148),
    .Q(\mac2.sum_lvl1_ff[0] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _566_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net202),
    .Q(\mac2.sum_lvl1_ff[1] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _567_ (.RESET_B(net81),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net118),
    .Q(\mac2.sum_lvl1_ff[8] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _568_ (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net185),
    .Q(\mac2.sum_lvl1_ff[9] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _569_ (.RESET_B(net57),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_036_),
    .Q(\mac2.products_ff[128] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _570_ (.RESET_B(net57),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_037_),
    .Q(\mac2.products_ff[129] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _571_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net112),
    .Q(\mac2.sum_lvl1_ff[16] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _572_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net177),
    .Q(\mac2.sum_lvl1_ff[17] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _573_ (.RESET_B(net76),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_064_),
    .Q(\mac2.products_ff[48] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _574_ (.RESET_B(net76),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_065_),
    .Q(\mac2.products_ff[49] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _575_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net114),
    .Q(\mac2.sum_lvl1_ff[24] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _576_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net181),
    .Q(\mac2.sum_lvl1_ff[25] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _577_ (.RESET_B(net57),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net28),
    .Q(\mac2.sum_lvl1_ff[32] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _578_ (.RESET_B(net58),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net32),
    .Q(\mac2.sum_lvl1_ff[33] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _579_ (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_034_),
    .Q(\mac2.products_ff[112] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _580_ (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_035_),
    .Q(\mac2.products_ff[113] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _581_ (.RESET_B(net76),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_066_),
    .Q(\mac2.products_ff[32] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _582_ (.RESET_B(net76),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_067_),
    .Q(\mac2.products_ff[33] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _583_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net122),
    .Q(\mac2.sum_lvl2_ff[0] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _584_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net200),
    .Q(\mac2.sum_lvl2_ff[1] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _585_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_068_),
    .Q(\mac2.products_ff[16] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _586_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_069_),
    .Q(\mac2.products_ff[17] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _587_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net106),
    .Q(\mac2.sum_lvl2_ff[4] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _588_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net187),
    .Q(\mac2.sum_lvl2_ff[5] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _589_ (.RESET_B(net57),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net30),
    .Q(\mac2.sum_lvl2_ff[8] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _590_ (.RESET_B(net58),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net25),
    .Q(\mac2.sum_lvl2_ff[9] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _591_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_044_),
    .Q(\mac2.products_ff[0] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _592_ (.RESET_B(net80),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_045_),
    .Q(\mac2.products_ff[1] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _593_ (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_040_),
    .Q(\mac2.products_ff[96] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _594_ (.RESET_B(net63),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_041_),
    .Q(\mac2.products_ff[97] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _595_ (.RESET_B(net56),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net108),
    .Q(\mac2.total_sum[0] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _596_ (.RESET_B(net56),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net208),
    .Q(\mac2.total_sum[1] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _597_ (.RESET_B(net56),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net172),
    .Q(\mac2.total_sum[2] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _598_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net153),
    .Q(\mac2.sum_lvl3_ff[0] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_2 _599_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net197),
    .Q(\mac2.sum_lvl3_ff[1] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _600_ (.RESET_B(net58),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net36),
    .Q(\mac2.sum_lvl3_ff[2] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _601_ (.RESET_B(net58),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net33),
    .Q(\mac2.sum_lvl3_ff[3] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_tiehi heichips25_template_18 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net18));
 sg13g2_tiehi heichips25_template_19 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net19));
 sg13g2_tiehi heichips25_template_20 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net20));
 sg13g2_tiehi heichips25_template_21 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net21));
 sg13g2_tiehi heichips25_template_22 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net22));
 sg13g2_tiehi heichips25_template_23 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net23));
 sg13g2_tiehi heichips25_template_24 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net24));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_template_6 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net6));
 sg13g2_tielo heichips25_template_7 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net7));
 sg13g2_tielo heichips25_template_8 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net8));
 sg13g2_tielo heichips25_template_9 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net9));
 sg13g2_tielo heichips25_template_10 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net10));
 sg13g2_tielo heichips25_template_11 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net11));
 sg13g2_tielo heichips25_template_12 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net12));
 sg13g2_tielo heichips25_template_13 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net13));
 sg13g2_tielo heichips25_template_14 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net14));
 sg13g2_tielo heichips25_template_15 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net15));
 sg13g2_tielo heichips25_template_16 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net16));
 sg13g2_tiehi heichips25_template_17 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net17));
 sg13g2_buf_8 fanout56 (.A(net59),
    .X(net56),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout57 (.A(net59),
    .X(net57),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout58 (.A(net59),
    .X(net58),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout59 (.A(net62),
    .X(net59),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout60 (.A(net61),
    .X(net60),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout61 (.A(net62),
    .X(net61),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout62 (.A(rst_n),
    .X(net62),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout63 (.A(net64),
    .X(net63),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout64 (.A(net68),
    .X(net64),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout65 (.A(net68),
    .X(net65),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout66 (.A(net68),
    .X(net66),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout67 (.A(net68),
    .X(net67),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout68 (.A(rst_n),
    .X(net68),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout69 (.A(net70),
    .X(net69),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout70 (.A(net75),
    .X(net70),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout71 (.A(net74),
    .X(net71),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout72 (.A(net74),
    .X(net72),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout73 (.A(net74),
    .X(net73),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout74 (.A(net75),
    .X(net74),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout75 (.A(net81),
    .X(net75),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout76 (.A(net77),
    .X(net76),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout77 (.A(net81),
    .X(net77),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout78 (.A(net80),
    .X(net78),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout79 (.A(net80),
    .X(net79),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout80 (.A(net81),
    .X(net80),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout81 (.A(rst_n),
    .X(net81),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output1 (.A(net1),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uo_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_template_5 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net5));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload0 (.VDD(VPWR),
    .A(clknet_5_7__leaf_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload1 (.VDD(VPWR),
    .A(clknet_5_11__leaf_clk),
    .VSS(VGND));
 sg13g2_buf_1 clkload2 (.A(clknet_5_12__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload3 (.VDD(VPWR),
    .A(clknet_5_15__leaf_clk),
    .VSS(VGND));
 sg13g2_buf_1 clkload4 (.A(clknet_5_17__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 clkload5 (.A(clknet_5_19__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload6 (.VDD(VPWR),
    .A(clknet_5_23__leaf_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload7 (.VDD(VPWR),
    .A(clknet_5_27__leaf_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload8 (.VDD(VPWR),
    .A(clknet_5_31__leaf_clk),
    .VSS(VGND));
 sg13g2_dlygate4sd3_1 hold1 (.A(\mac2.sum_lvl1_ff[33] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold2 (.A(\mac1.sum_lvl1_ff[33] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold3 (.A(\mac1.products_ff[129] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold4 (.A(\mac2.products_ff[128] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold5 (.A(\mac1.sum_lvl2_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold6 (.A(\mac2.sum_lvl1_ff[32] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold7 (.A(\mac1.sum_lvl2_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold8 (.A(\mac2.products_ff[129] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold9 (.A(\mac2.sum_lvl2_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold10 (.A(\mac1.sum_lvl1_ff[32] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold11 (.A(\mac1.products_ff[128] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold12 (.A(\mac2.sum_lvl2_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold13 (.A(\mac1.products_ff[96] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold14 (.A(_006_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold15 (.A(\DP_4.matrix[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold16 (.A(\DP_1.matrix[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold17 (.A(\DP_4.matrix[113] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold18 (.A(\DP_3.matrix[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold19 (.A(\DP_3.matrix[113] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold20 (.A(\DP_4.matrix[65] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold21 (.A(\DP_3.matrix[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold22 (.A(\DP_1.matrix[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold23 (.A(\DP_1.matrix[113] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold24 (.A(\DP_1.matrix[97] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold25 (.A(\DP_2.matrix[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold26 (.A(\DP_4.matrix[81] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold27 (.A(\DP_4.matrix[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold28 (.A(\DP_3.matrix[81] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold29 (.A(\DP_2.matrix[33] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold30 (.A(\DP_4.matrix[33] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold31 (.A(\DP_2.matrix[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold32 (.A(\DP_3.matrix[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold33 (.A(\DP_4.matrix[129] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold34 (.A(\DP_2.matrix[81] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold35 (.A(\DP_3.matrix[97] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold36 (.A(\DP_1.matrix[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold37 (.A(\DP_3.matrix[129] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold38 (.A(\DP_2.matrix[113] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold39 (.A(\DP_1.matrix[81] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold40 (.A(\DP_4.matrix[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold41 (.A(\DP_2.matrix[65] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold42 (.A(\DP_1.matrix[33] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold43 (.A(\DP_3.matrix[65] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold44 (.A(\DP_4.matrix[97] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold45 (.A(\DP_2.matrix[97] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold46 (.A(\DP_2.matrix[129] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold47 (.A(\mac1.products_ff[64] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold48 (.A(_004_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold49 (.A(\DP_3.matrix[33] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold50 (.A(\DP_2.matrix[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold51 (.A(\DP_1.matrix[65] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold52 (.A(\mac1.sum_lvl1_ff[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold53 (.A(_010_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold54 (.A(\DP_1.matrix[129] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold55 (.A(\mac2.sum_lvl1_ff[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold56 (.A(_027_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold57 (.A(\mac2.sum_lvl3_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold58 (.A(_032_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold59 (.A(\mac1.products_ff[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold60 (.A(_002_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold61 (.A(\mac2.products_ff[64] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold62 (.A(_021_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold63 (.A(\mac2.products_ff[112] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold64 (.A(_023_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold65 (.A(\mac1.sum_lvl2_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold66 (.A(_012_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold67 (.A(\mac2.products_ff[32] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold68 (.A(_019_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold69 (.A(\DP_1.matrix[128] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold70 (.A(\DP_2.matrix[112] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold71 (.A(\mac2.sum_lvl1_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold72 (.A(_025_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold73 (.A(\DP_2.matrix[32] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold74 (.A(\DP_4.matrix[128] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold75 (.A(\DP_3.matrix[112] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold76 (.A(\mac1.products_ff[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold77 (.A(_000_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold78 (.A(\DP_1.matrix[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold79 (.A(\mac1.sum_lvl1_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold80 (.A(_008_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold81 (.A(\DP_1.matrix[64] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold82 (.A(\DP_2.matrix[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold83 (.A(\DP_4.matrix[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold84 (.A(\DP_4.matrix[64] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold85 (.A(\DP_2.matrix[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold86 (.A(\DP_4.matrix[96] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold87 (.A(\DP_3.matrix[96] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold88 (.A(\DP_3.matrix[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold89 (.A(\DP_4.matrix[32] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold90 (.A(\DP_2.matrix[96] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold91 (.A(\DP_3.matrix[64] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold92 (.A(\DP_3.matrix[128] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold93 (.A(\DP_4.matrix[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold94 (.A(\DP_4.matrix[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold95 (.A(\DP_4.matrix[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold96 (.A(\DP_3.matrix[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold97 (.A(\mac2.products_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold98 (.A(_017_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold99 (.A(\DP_3.matrix[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold100 (.A(\DP_2.matrix[128] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold101 (.A(\DP_1.matrix[96] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold102 (.A(\mac2.sum_lvl2_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold103 (.A(_029_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold104 (.A(\DP_1.matrix[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold105 (.A(\DP_4.matrix[112] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold106 (.A(\DP_2.matrix[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold107 (.A(\DP_2.matrix[64] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold108 (.A(\DP_2.matrix[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold109 (.A(\DP_1.matrix[112] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold110 (.A(\DP_1.matrix[32] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold111 (.A(\DP_3.matrix[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold112 (.A(\DP_1.matrix[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold113 (.A(\DP_3.matrix[32] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold114 (.A(\DP_1.matrix[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold115 (.A(\mac1.sum_lvl3_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold116 (.A(_015_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold117 (.A(\mac1.sum_lvl3_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold118 (.A(_167_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold119 (.A(_014_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold120 (.A(\mac2.sum_lvl3_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold121 (.A(_183_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold122 (.A(_031_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold123 (.A(\mac1.sum_lvl1_ff[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold124 (.A(_011_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold125 (.A(\mac2.products_ff[81] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold126 (.A(_179_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold127 (.A(_022_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold128 (.A(\mac1.products_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold129 (.A(_001_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold130 (.A(\mac2.products_ff[96] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold131 (.A(_024_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold132 (.A(\mac1.products_ff[32] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold133 (.A(_003_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold134 (.A(\mac2.products_ff[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold135 (.A(_020_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold136 (.A(\mac2.sum_lvl1_ff[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold137 (.A(_028_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold138 (.A(\mac1.products_ff[65] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold139 (.A(_161_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold140 (.A(_005_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold141 (.A(\mac1.sum_lvl1_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold142 (.A(_009_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold143 (.A(\mac1.products_ff[97] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold144 (.A(_159_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold145 (.A(_007_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold146 (.A(\mac2.sum_lvl2_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold147 (.A(_030_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold148 (.A(\mac2.sum_lvl1_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold149 (.A(_175_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold150 (.A(_026_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold151 (.A(\mac2.products_ff[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold152 (.A(_018_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold153 (.A(\mac1.sum_lvl2_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold154 (.A(_013_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold155 (.A(\mac1.sum_lvl3_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold156 (.A(_016_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold157 (.A(\mac2.sum_lvl3_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold158 (.A(_033_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net208));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_6 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_1028 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net17;
 assign uio_oe[1] = net18;
 assign uio_oe[2] = net19;
 assign uio_oe[3] = net20;
 assign uio_oe[4] = net21;
 assign uio_oe[5] = net22;
 assign uio_oe[6] = net23;
 assign uio_oe[7] = net24;
 assign uio_out[0] = net5;
 assign uio_out[1] = net6;
 assign uio_out[2] = net7;
 assign uio_out[3] = net8;
 assign uio_out[4] = net9;
 assign uio_out[5] = net10;
 assign uio_out[6] = net11;
 assign uio_out[7] = net12;
 assign uo_out[4] = net13;
 assign uo_out[5] = net14;
 assign uo_out[6] = net15;
 assign uo_out[7] = net16;
endmodule
