module heichips25_template (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \DP_1.matrix[0] ;
 wire \DP_1.matrix[112] ;
 wire \DP_1.matrix[113] ;
 wire \DP_1.matrix[128] ;
 wire \DP_1.matrix[129] ;
 wire \DP_1.matrix[16] ;
 wire \DP_1.matrix[17] ;
 wire \DP_1.matrix[1] ;
 wire \DP_1.matrix[32] ;
 wire \DP_1.matrix[33] ;
 wire \DP_1.matrix[48] ;
 wire \DP_1.matrix[49] ;
 wire \DP_1.matrix[64] ;
 wire \DP_1.matrix[65] ;
 wire \DP_1.matrix[80] ;
 wire \DP_1.matrix[81] ;
 wire \DP_1.matrix[96] ;
 wire \DP_1.matrix[97] ;
 wire \DP_2.matrix[0] ;
 wire \DP_2.matrix[112] ;
 wire \DP_2.matrix[113] ;
 wire \DP_2.matrix[128] ;
 wire \DP_2.matrix[129] ;
 wire \DP_2.matrix[16] ;
 wire \DP_2.matrix[17] ;
 wire \DP_2.matrix[1] ;
 wire \DP_2.matrix[32] ;
 wire \DP_2.matrix[33] ;
 wire \DP_2.matrix[48] ;
 wire \DP_2.matrix[49] ;
 wire \DP_2.matrix[64] ;
 wire \DP_2.matrix[65] ;
 wire \DP_2.matrix[80] ;
 wire \DP_2.matrix[81] ;
 wire \DP_2.matrix[96] ;
 wire \DP_2.matrix[97] ;
 wire \DP_3.matrix[0] ;
 wire \DP_3.matrix[112] ;
 wire \DP_3.matrix[113] ;
 wire \DP_3.matrix[128] ;
 wire \DP_3.matrix[129] ;
 wire \DP_3.matrix[16] ;
 wire \DP_3.matrix[17] ;
 wire \DP_3.matrix[1] ;
 wire \DP_3.matrix[32] ;
 wire \DP_3.matrix[33] ;
 wire \DP_3.matrix[48] ;
 wire \DP_3.matrix[49] ;
 wire \DP_3.matrix[64] ;
 wire \DP_3.matrix[65] ;
 wire \DP_3.matrix[80] ;
 wire \DP_3.matrix[81] ;
 wire \DP_3.matrix[96] ;
 wire \DP_3.matrix[97] ;
 wire \DP_4.matrix[0] ;
 wire \DP_4.matrix[112] ;
 wire \DP_4.matrix[113] ;
 wire \DP_4.matrix[128] ;
 wire \DP_4.matrix[129] ;
 wire \DP_4.matrix[16] ;
 wire \DP_4.matrix[17] ;
 wire \DP_4.matrix[1] ;
 wire \DP_4.matrix[32] ;
 wire \DP_4.matrix[33] ;
 wire \DP_4.matrix[48] ;
 wire \DP_4.matrix[49] ;
 wire \DP_4.matrix[64] ;
 wire \DP_4.matrix[65] ;
 wire \DP_4.matrix[80] ;
 wire \DP_4.matrix[81] ;
 wire \DP_4.matrix[96] ;
 wire \DP_4.matrix[97] ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire \mac1.products_ff[0] ;
 wire \mac1.products_ff[112] ;
 wire \mac1.products_ff[113] ;
 wire \mac1.products_ff[128] ;
 wire \mac1.products_ff[129] ;
 wire \mac1.products_ff[16] ;
 wire \mac1.products_ff[17] ;
 wire \mac1.products_ff[1] ;
 wire \mac1.products_ff[32] ;
 wire \mac1.products_ff[33] ;
 wire \mac1.products_ff[48] ;
 wire \mac1.products_ff[49] ;
 wire \mac1.products_ff[64] ;
 wire \mac1.products_ff[65] ;
 wire \mac1.products_ff[80] ;
 wire \mac1.products_ff[81] ;
 wire \mac1.products_ff[96] ;
 wire \mac1.products_ff[97] ;
 wire \mac1.sum_lvl1_ff[0] ;
 wire \mac1.sum_lvl1_ff[16] ;
 wire \mac1.sum_lvl1_ff[17] ;
 wire \mac1.sum_lvl1_ff[1] ;
 wire \mac1.sum_lvl1_ff[24] ;
 wire \mac1.sum_lvl1_ff[25] ;
 wire \mac1.sum_lvl1_ff[32] ;
 wire \mac1.sum_lvl1_ff[33] ;
 wire \mac1.sum_lvl1_ff[8] ;
 wire \mac1.sum_lvl1_ff[9] ;
 wire \mac1.sum_lvl2_ff[0] ;
 wire \mac1.sum_lvl2_ff[1] ;
 wire \mac1.sum_lvl2_ff[4] ;
 wire \mac1.sum_lvl2_ff[5] ;
 wire \mac1.sum_lvl2_ff[8] ;
 wire \mac1.sum_lvl2_ff[9] ;
 wire \mac1.sum_lvl3_ff[0] ;
 wire \mac1.sum_lvl3_ff[1] ;
 wire \mac1.sum_lvl3_ff[2] ;
 wire \mac1.sum_lvl3_ff[3] ;
 wire \mac1.total_sum[0] ;
 wire \mac1.total_sum[1] ;
 wire \mac1.total_sum[2] ;
 wire \mac2.products_ff[0] ;
 wire \mac2.products_ff[112] ;
 wire \mac2.products_ff[113] ;
 wire \mac2.products_ff[128] ;
 wire \mac2.products_ff[129] ;
 wire \mac2.products_ff[16] ;
 wire \mac2.products_ff[17] ;
 wire \mac2.products_ff[1] ;
 wire \mac2.products_ff[32] ;
 wire \mac2.products_ff[33] ;
 wire \mac2.products_ff[48] ;
 wire \mac2.products_ff[49] ;
 wire \mac2.products_ff[64] ;
 wire \mac2.products_ff[65] ;
 wire \mac2.products_ff[80] ;
 wire \mac2.products_ff[81] ;
 wire \mac2.products_ff[96] ;
 wire \mac2.products_ff[97] ;
 wire \mac2.sum_lvl1_ff[0] ;
 wire \mac2.sum_lvl1_ff[16] ;
 wire \mac2.sum_lvl1_ff[17] ;
 wire \mac2.sum_lvl1_ff[1] ;
 wire \mac2.sum_lvl1_ff[24] ;
 wire \mac2.sum_lvl1_ff[25] ;
 wire \mac2.sum_lvl1_ff[32] ;
 wire \mac2.sum_lvl1_ff[33] ;
 wire \mac2.sum_lvl1_ff[8] ;
 wire \mac2.sum_lvl1_ff[9] ;
 wire \mac2.sum_lvl2_ff[0] ;
 wire \mac2.sum_lvl2_ff[1] ;
 wire \mac2.sum_lvl2_ff[4] ;
 wire \mac2.sum_lvl2_ff[5] ;
 wire \mac2.sum_lvl2_ff[8] ;
 wire \mac2.sum_lvl2_ff[9] ;
 wire \mac2.sum_lvl3_ff[0] ;
 wire \mac2.sum_lvl3_ff[1] ;
 wire \mac2.sum_lvl3_ff[2] ;
 wire \mac2.sum_lvl3_ff[3] ;
 wire \mac2.total_sum[0] ;
 wire \mac2.total_sum[1] ;
 wire \mac2.total_sum[2] ;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire clknet_0_clk;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net5;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;

 sg13g2_and2_1 _222_ (.A(net155),
    .B(net125),
    .X(_034_));
 sg13g2_and2_1 _223_ (.A(net124),
    .B(net142),
    .X(_036_));
 sg13g2_and2_1 _224_ (.A(net144),
    .B(net138),
    .X(_038_));
 sg13g2_and2_1 _225_ (.A(net136),
    .B(net137),
    .X(_040_));
 sg13g2_and2_1 _226_ (.A(net154),
    .B(net156),
    .X(_042_));
 sg13g2_and2_1 _227_ (.A(net143),
    .B(net146),
    .X(_044_));
 sg13g2_and2_1 _228_ (.A(net151),
    .B(net140),
    .X(_046_));
 sg13g2_and2_1 _229_ (.A(net162),
    .B(net158),
    .X(_048_));
 sg13g2_and2_1 _230_ (.A(net131),
    .B(net157),
    .X(_050_));
 sg13g2_and2_1 _231_ (.A(net164),
    .B(net132),
    .X(_052_));
 sg13g2_and2_1 _232_ (.A(net160),
    .B(net123),
    .X(_054_));
 sg13g2_and2_1 _233_ (.A(net128),
    .B(net135),
    .X(_056_));
 sg13g2_and2_1 _234_ (.A(net119),
    .B(net150),
    .X(_058_));
 sg13g2_and2_1 _235_ (.A(net134),
    .B(net141),
    .X(_060_));
 sg13g2_and2_1 _236_ (.A(net159),
    .B(net120),
    .X(_062_));
 sg13g2_and2_1 _237_ (.A(net145),
    .B(net149),
    .X(_064_));
 sg13g2_and2_1 _238_ (.A(net139),
    .B(net163),
    .X(_066_));
 sg13g2_and2_1 _239_ (.A(net133),
    .B(net161),
    .X(_068_));
 sg13g2_nand2_1 _240_ (.Y(_142_),
    .A(\mac1.total_sum[0] ),
    .B(\mac2.total_sum[0] ));
 sg13g2_nand2_1 _241_ (.Y(_143_),
    .A(\mac1.total_sum[1] ),
    .B(\mac2.total_sum[1] ));
 sg13g2_nor2_1 _242_ (.A(\mac1.total_sum[1] ),
    .B(\mac2.total_sum[1] ),
    .Y(_144_));
 sg13g2_xor2_1 _243_ (.B(\mac2.total_sum[1] ),
    .A(\mac1.total_sum[1] ),
    .X(_145_));
 sg13g2_xnor2_1 _244_ (.Y(net2),
    .A(_142_),
    .B(_145_));
 sg13g2_o21ai_1 _245_ (.B1(_143_),
    .Y(_146_),
    .A1(_142_),
    .A2(_144_));
 sg13g2_and2_1 _246_ (.A(\mac1.total_sum[2] ),
    .B(\mac2.total_sum[2] ),
    .X(_147_));
 sg13g2_or2_1 _247_ (.X(_148_),
    .B(\mac2.total_sum[2] ),
    .A(\mac1.total_sum[2] ));
 sg13g2_nand2b_1 _248_ (.Y(_149_),
    .B(_148_),
    .A_N(_147_));
 sg13g2_xnor2_1 _249_ (.Y(net3),
    .A(_146_),
    .B(_149_));
 sg13g2_xor2_1 _250_ (.B(\mac2.total_sum[0] ),
    .A(\mac1.total_sum[0] ),
    .X(net1));
 sg13g2_nand2_1 _251_ (.Y(_150_),
    .A(net178),
    .B(net126));
 sg13g2_xor2_1 _252_ (.B(\mac1.products_ff[17] ),
    .A(\mac1.products_ff[1] ),
    .X(_151_));
 sg13g2_xnor2_1 _253_ (.Y(_001_),
    .A(_150_),
    .B(_151_));
 sg13g2_xor2_1 _254_ (.B(net126),
    .A(\mac1.products_ff[0] ),
    .X(_000_));
 sg13g2_nand2_1 _255_ (.Y(_152_),
    .A(net203),
    .B(net115));
 sg13g2_xor2_1 _256_ (.B(\mac1.sum_lvl2_ff[1] ),
    .A(\mac1.sum_lvl2_ff[5] ),
    .X(_153_));
 sg13g2_xnor2_1 _257_ (.Y(_013_),
    .A(_152_),
    .B(_153_));
 sg13g2_xor2_1 _258_ (.B(net115),
    .A(\mac1.sum_lvl2_ff[4] ),
    .X(_012_));
 sg13g2_nand2_1 _259_ (.Y(_154_),
    .A(net173),
    .B(net102));
 sg13g2_xor2_1 _260_ (.B(\mac1.sum_lvl1_ff[17] ),
    .A(\mac1.sum_lvl1_ff[25] ),
    .X(_155_));
 sg13g2_xnor2_1 _261_ (.Y(_011_),
    .A(_154_),
    .B(_155_));
 sg13g2_xor2_1 _262_ (.B(net102),
    .A(\mac1.sum_lvl1_ff[24] ),
    .X(_010_));
 sg13g2_nand2_1 _263_ (.Y(_156_),
    .A(net191),
    .B(net129));
 sg13g2_xor2_1 _264_ (.B(\mac1.sum_lvl1_ff[1] ),
    .A(\mac1.sum_lvl1_ff[9] ),
    .X(_157_));
 sg13g2_xnor2_1 _265_ (.Y(_009_),
    .A(_156_),
    .B(_157_));
 sg13g2_xor2_1 _266_ (.B(net129),
    .A(\mac1.sum_lvl1_ff[8] ),
    .X(_008_));
 sg13g2_nand2_1 _267_ (.Y(_158_),
    .A(\mac1.products_ff[112] ),
    .B(net37));
 sg13g2_xor2_1 _268_ (.B(net193),
    .A(\mac1.products_ff[113] ),
    .X(_159_));
 sg13g2_xnor2_1 _269_ (.Y(_007_),
    .A(_158_),
    .B(net194));
 sg13g2_xor2_1 _270_ (.B(net37),
    .A(\mac1.products_ff[112] ),
    .X(_006_));
 sg13g2_nand2_1 _271_ (.Y(_160_),
    .A(\mac1.products_ff[80] ),
    .B(net97));
 sg13g2_xor2_1 _272_ (.B(net188),
    .A(\mac1.products_ff[81] ),
    .X(_161_));
 sg13g2_xnor2_1 _273_ (.Y(_005_),
    .A(_160_),
    .B(net189));
 sg13g2_xor2_1 _274_ (.B(net97),
    .A(\mac1.products_ff[80] ),
    .X(_004_));
 sg13g2_nand2_1 _275_ (.Y(_162_),
    .A(net182),
    .B(net109));
 sg13g2_xor2_1 _276_ (.B(\mac1.products_ff[49] ),
    .A(\mac1.products_ff[33] ),
    .X(_163_));
 sg13g2_xnor2_1 _277_ (.Y(_003_),
    .A(_162_),
    .B(_163_));
 sg13g2_xor2_1 _278_ (.B(net109),
    .A(\mac1.products_ff[32] ),
    .X(_002_));
 sg13g2_nand2_1 _279_ (.Y(_164_),
    .A(net201),
    .B(net147));
 sg13g2_xor2_1 _280_ (.B(\mac2.products_ff[1] ),
    .A(\mac2.products_ff[17] ),
    .X(_165_));
 sg13g2_xnor2_1 _281_ (.Y(_018_),
    .A(_164_),
    .B(_165_));
 sg13g2_xor2_1 _282_ (.B(net147),
    .A(\mac2.products_ff[16] ),
    .X(_017_));
 sg13g2_nand2_1 _283_ (.Y(_166_),
    .A(net205),
    .B(net165));
 sg13g2_nand2_1 _284_ (.Y(_167_),
    .A(net167),
    .B(\mac1.sum_lvl3_ff[1] ));
 sg13g2_nor2_1 _285_ (.A(net167),
    .B(\mac1.sum_lvl3_ff[1] ),
    .Y(_168_));
 sg13g2_xor2_1 _286_ (.B(\mac1.sum_lvl3_ff[1] ),
    .A(net167),
    .X(_169_));
 sg13g2_xnor2_1 _287_ (.Y(_016_),
    .A(_166_),
    .B(_169_));
 sg13g2_xor2_1 _288_ (.B(net165),
    .A(\mac1.sum_lvl3_ff[2] ),
    .X(_015_));
 sg13g2_nand2_1 _289_ (.Y(_170_),
    .A(net196),
    .B(net152));
 sg13g2_xor2_1 _290_ (.B(\mac2.sum_lvl2_ff[1] ),
    .A(\mac2.sum_lvl2_ff[5] ),
    .X(_171_));
 sg13g2_xnor2_1 _291_ (.Y(_030_),
    .A(_170_),
    .B(_171_));
 sg13g2_xor2_1 _292_ (.B(net152),
    .A(\mac2.sum_lvl2_ff[4] ),
    .X(_029_));
 sg13g2_nand2_1 _293_ (.Y(_172_),
    .A(net186),
    .B(net105));
 sg13g2_xor2_1 _294_ (.B(\mac2.sum_lvl1_ff[17] ),
    .A(\mac2.sum_lvl1_ff[25] ),
    .X(_173_));
 sg13g2_xnor2_1 _295_ (.Y(_028_),
    .A(_172_),
    .B(_173_));
 sg13g2_xor2_1 _296_ (.B(net105),
    .A(\mac2.sum_lvl1_ff[24] ),
    .X(_027_));
 sg13g2_nand2_1 _297_ (.Y(_174_),
    .A(net121),
    .B(\mac2.sum_lvl1_ff[0] ));
 sg13g2_xor2_1 _298_ (.B(net198),
    .A(\mac2.sum_lvl1_ff[9] ),
    .X(_175_));
 sg13g2_xnor2_1 _299_ (.Y(_026_),
    .A(_174_),
    .B(net199));
 sg13g2_xor2_1 _300_ (.B(\mac2.sum_lvl1_ff[0] ),
    .A(net121),
    .X(_025_));
 sg13g2_nand2_1 _301_ (.Y(_176_),
    .A(net180),
    .B(net113));
 sg13g2_xor2_1 _302_ (.B(\mac2.products_ff[113] ),
    .A(\mac2.products_ff[97] ),
    .X(_177_));
 sg13g2_xnor2_1 _303_ (.Y(_024_),
    .A(_176_),
    .B(_177_));
 sg13g2_xor2_1 _304_ (.B(net113),
    .A(\mac2.products_ff[96] ),
    .X(_023_));
 sg13g2_nand2_1 _305_ (.Y(_178_),
    .A(net111),
    .B(\mac2.products_ff[80] ));
 sg13g2_xor2_1 _306_ (.B(net175),
    .A(\mac2.products_ff[65] ),
    .X(_179_));
 sg13g2_xnor2_1 _307_ (.Y(_022_),
    .A(_178_),
    .B(net176));
 sg13g2_xor2_1 _308_ (.B(\mac2.products_ff[80] ),
    .A(net111),
    .X(_021_));
 sg13g2_nand2_1 _309_ (.Y(_180_),
    .A(net184),
    .B(net117));
 sg13g2_xor2_1 _310_ (.B(\mac2.products_ff[33] ),
    .A(\mac2.products_ff[49] ),
    .X(_181_));
 sg13g2_xnor2_1 _311_ (.Y(_020_),
    .A(_180_),
    .B(_181_));
 sg13g2_xor2_1 _312_ (.B(net117),
    .A(\mac2.products_ff[48] ),
    .X(_019_));
 sg13g2_nand2_1 _313_ (.Y(_182_),
    .A(net207),
    .B(net107));
 sg13g2_nand2_1 _314_ (.Y(_183_),
    .A(net170),
    .B(\mac2.sum_lvl3_ff[3] ));
 sg13g2_nor2_1 _315_ (.A(net170),
    .B(\mac2.sum_lvl3_ff[3] ),
    .Y(_184_));
 sg13g2_xor2_1 _316_ (.B(\mac2.sum_lvl3_ff[3] ),
    .A(net170),
    .X(_185_));
 sg13g2_xnor2_1 _317_ (.Y(_033_),
    .A(_182_),
    .B(_185_));
 sg13g2_xor2_1 _318_ (.B(net107),
    .A(\mac2.sum_lvl3_ff[0] ),
    .X(_032_));
 sg13g2_nand2_1 _319_ (.Y(_186_),
    .A(net155),
    .B(net43));
 sg13g2_nand2_1 _320_ (.Y(_187_),
    .A(net125),
    .B(net41));
 sg13g2_xor2_1 _321_ (.B(_187_),
    .A(_186_),
    .X(_035_));
 sg13g2_nand2_1 _322_ (.Y(_188_),
    .A(net124),
    .B(net87));
 sg13g2_nand2_1 _323_ (.Y(_189_),
    .A(net142),
    .B(net83));
 sg13g2_xor2_1 _324_ (.B(_189_),
    .A(_188_),
    .X(_037_));
 sg13g2_a21o_2 _325_ (.A2(_148_),
    .A1(_146_),
    .B1(_147_),
    .X(net4));
 sg13g2_nand2_1 _326_ (.Y(_190_),
    .A(net144),
    .B(net52));
 sg13g2_nand2_1 _327_ (.Y(_191_),
    .A(net138),
    .B(net50));
 sg13g2_xor2_1 _328_ (.B(_191_),
    .A(_190_),
    .X(_039_));
 sg13g2_nand2_1 _329_ (.Y(_192_),
    .A(net136),
    .B(net85));
 sg13g2_nand2_1 _330_ (.Y(_193_),
    .A(net137),
    .B(net94));
 sg13g2_xor2_1 _331_ (.B(_193_),
    .A(_192_),
    .X(_041_));
 sg13g2_nand2_1 _332_ (.Y(_194_),
    .A(net46),
    .B(net156));
 sg13g2_nand2_1 _333_ (.Y(_195_),
    .A(net154),
    .B(net55));
 sg13g2_xor2_1 _334_ (.B(_195_),
    .A(_194_),
    .X(_043_));
 sg13g2_nand2_1 _335_ (.Y(_196_),
    .A(net143),
    .B(net45));
 sg13g2_nand2_1 _336_ (.Y(_197_),
    .A(net146),
    .B(net51));
 sg13g2_xor2_1 _337_ (.B(_197_),
    .A(_196_),
    .X(_045_));
 sg13g2_nand2_1 _338_ (.Y(_198_),
    .A(net48),
    .B(net140));
 sg13g2_nand2_1 _339_ (.Y(_199_),
    .A(net151),
    .B(net95));
 sg13g2_xor2_1 _340_ (.B(_199_),
    .A(_198_),
    .X(_047_));
 sg13g2_nand2_1 _341_ (.Y(_200_),
    .A(net89),
    .B(net158));
 sg13g2_nand2_1 _342_ (.Y(_201_),
    .A(net162),
    .B(net84));
 sg13g2_xor2_1 _343_ (.B(_201_),
    .A(_200_),
    .X(_049_));
 sg13g2_nand2_1 _344_ (.Y(_202_),
    .A(net101),
    .B(net157));
 sg13g2_nand2_1 _345_ (.Y(_203_),
    .A(net131),
    .B(net91));
 sg13g2_xor2_1 _346_ (.B(_203_),
    .A(_202_),
    .X(_051_));
 sg13g2_nand2_1 _347_ (.Y(_204_),
    .A(net86),
    .B(net132));
 sg13g2_nand2_1 _348_ (.Y(_205_),
    .A(net164),
    .B(net100));
 sg13g2_xor2_1 _349_ (.B(_205_),
    .A(_204_),
    .X(_053_));
 sg13g2_nand2_1 _350_ (.Y(_206_),
    .A(net92),
    .B(net123));
 sg13g2_nand2_1 _351_ (.Y(_207_),
    .A(net160),
    .B(net53));
 sg13g2_xor2_1 _352_ (.B(_207_),
    .A(_206_),
    .X(_055_));
 sg13g2_nand2_1 _353_ (.Y(_208_),
    .A(net40),
    .B(net135));
 sg13g2_nand2_1 _354_ (.Y(_209_),
    .A(net128),
    .B(net49));
 sg13g2_xor2_1 _355_ (.B(_209_),
    .A(_208_),
    .X(_057_));
 sg13g2_o21ai_1 _356_ (.B1(net168),
    .Y(_014_),
    .A1(_166_),
    .A2(_168_));
 sg13g2_nand2_1 _357_ (.Y(_210_),
    .A(net104),
    .B(net150));
 sg13g2_nand2_1 _358_ (.Y(_211_),
    .A(net119),
    .B(net96));
 sg13g2_xor2_1 _359_ (.B(_211_),
    .A(_210_),
    .X(_059_));
 sg13g2_nand2_1 _360_ (.Y(_212_),
    .A(net134),
    .B(net93));
 sg13g2_nand2_1 _361_ (.Y(_213_),
    .A(net141),
    .B(net44));
 sg13g2_xor2_1 _362_ (.B(_213_),
    .A(_212_),
    .X(_061_));
 sg13g2_nand2_1 _363_ (.Y(_214_),
    .A(net47),
    .B(net120));
 sg13g2_nand2_1 _364_ (.Y(_215_),
    .A(net159),
    .B(net88));
 sg13g2_xor2_1 _365_ (.B(_215_),
    .A(_214_),
    .X(_063_));
 sg13g2_nand2_1 _366_ (.Y(_216_),
    .A(net145),
    .B(net42));
 sg13g2_nand2_1 _367_ (.Y(_217_),
    .A(net149),
    .B(net90));
 sg13g2_xor2_1 _368_ (.B(_217_),
    .A(_216_),
    .X(_065_));
 sg13g2_nand2_1 _369_ (.Y(_218_),
    .A(net139),
    .B(net99));
 sg13g2_nand2_1 _370_ (.Y(_219_),
    .A(net163),
    .B(net54));
 sg13g2_xor2_1 _371_ (.B(_219_),
    .A(_218_),
    .X(_067_));
 sg13g2_nand2_1 _372_ (.Y(_220_),
    .A(net133),
    .B(net82));
 sg13g2_nand2_1 _373_ (.Y(_221_),
    .A(net161),
    .B(net39));
 sg13g2_xor2_1 _374_ (.B(_221_),
    .A(_220_),
    .X(_069_));
 sg13g2_o21ai_1 _375_ (.B1(net171),
    .Y(_031_),
    .A1(_182_),
    .A2(_184_));
 sg13g2_buf_1 _376_ (.A(net154),
    .X(_070_));
 sg13g2_buf_1 _377_ (.A(net46),
    .X(_071_));
 sg13g2_buf_1 _378_ (.A(net128),
    .X(_072_));
 sg13g2_buf_1 _379_ (.A(net40),
    .X(_073_));
 sg13g2_buf_1 _380_ (.A(net160),
    .X(_074_));
 sg13g2_buf_1 _381_ (.A(net92),
    .X(_075_));
 sg13g2_buf_1 _382_ (.A(net164),
    .X(_076_));
 sg13g2_buf_1 _383_ (.A(net86),
    .X(_077_));
 sg13g2_buf_1 _384_ (.A(net131),
    .X(_078_));
 sg13g2_buf_1 _385_ (.A(net101),
    .X(_079_));
 sg13g2_buf_1 _386_ (.A(net162),
    .X(_080_));
 sg13g2_buf_1 _387_ (.A(net89),
    .X(_081_));
 sg13g2_buf_1 _388_ (.A(net151),
    .X(_082_));
 sg13g2_buf_1 _389_ (.A(net48),
    .X(_083_));
 sg13g2_buf_1 _390_ (.A(net159),
    .X(_084_));
 sg13g2_buf_1 _391_ (.A(net47),
    .X(_085_));
 sg13g2_buf_1 _392_ (.A(net119),
    .X(_086_));
 sg13g2_buf_1 _393_ (.A(net104),
    .X(_087_));
 sg13g2_buf_1 _394_ (.A(net156),
    .X(_088_));
 sg13g2_buf_1 _395_ (.A(net55),
    .X(_089_));
 sg13g2_buf_1 _396_ (.A(net135),
    .X(_090_));
 sg13g2_buf_1 _397_ (.A(net49),
    .X(_091_));
 sg13g2_buf_1 _398_ (.A(net123),
    .X(_092_));
 sg13g2_buf_1 _399_ (.A(net53),
    .X(_093_));
 sg13g2_buf_1 _400_ (.A(net132),
    .X(_094_));
 sg13g2_buf_1 _401_ (.A(net100),
    .X(_095_));
 sg13g2_buf_1 _402_ (.A(net157),
    .X(_096_));
 sg13g2_buf_1 _403_ (.A(net91),
    .X(_097_));
 sg13g2_buf_1 _404_ (.A(net158),
    .X(_098_));
 sg13g2_buf_1 _405_ (.A(net84),
    .X(_099_));
 sg13g2_buf_1 _406_ (.A(net140),
    .X(_100_));
 sg13g2_buf_1 _407_ (.A(net95),
    .X(_101_));
 sg13g2_buf_1 _408_ (.A(net120),
    .X(_102_));
 sg13g2_buf_1 _409_ (.A(net88),
    .X(_103_));
 sg13g2_buf_1 _410_ (.A(net150),
    .X(_104_));
 sg13g2_buf_1 _411_ (.A(net96),
    .X(_105_));
 sg13g2_buf_1 _412_ (.A(net146),
    .X(_106_));
 sg13g2_buf_1 _413_ (.A(net45),
    .X(_107_));
 sg13g2_buf_1 _414_ (.A(net161),
    .X(_108_));
 sg13g2_buf_1 _415_ (.A(net82),
    .X(_109_));
 sg13g2_buf_1 _416_ (.A(net163),
    .X(_110_));
 sg13g2_buf_1 _417_ (.A(net99),
    .X(_111_));
 sg13g2_buf_1 _418_ (.A(net149),
    .X(_112_));
 sg13g2_buf_1 _419_ (.A(net42),
    .X(_113_));
 sg13g2_buf_1 _420_ (.A(net141),
    .X(_114_));
 sg13g2_buf_1 _421_ (.A(net93),
    .X(_115_));
 sg13g2_buf_1 _422_ (.A(net138),
    .X(_116_));
 sg13g2_buf_1 _423_ (.A(net52),
    .X(_117_));
 sg13g2_buf_1 _424_ (.A(net137),
    .X(_118_));
 sg13g2_buf_1 _425_ (.A(net85),
    .X(_119_));
 sg13g2_buf_1 _426_ (.A(net125),
    .X(_120_));
 sg13g2_buf_1 _427_ (.A(net43),
    .X(_121_));
 sg13g2_buf_1 _428_ (.A(net142),
    .X(_122_));
 sg13g2_buf_1 _429_ (.A(net87),
    .X(_123_));
 sg13g2_buf_1 _430_ (.A(net143),
    .X(_124_));
 sg13g2_buf_1 _431_ (.A(net51),
    .X(_125_));
 sg13g2_buf_1 _432_ (.A(net133),
    .X(_126_));
 sg13g2_buf_1 _433_ (.A(net39),
    .X(_127_));
 sg13g2_buf_1 _434_ (.A(net139),
    .X(_128_));
 sg13g2_buf_1 _435_ (.A(net54),
    .X(_129_));
 sg13g2_buf_1 _436_ (.A(net145),
    .X(_130_));
 sg13g2_buf_1 _437_ (.A(net90),
    .X(_131_));
 sg13g2_buf_1 _438_ (.A(net134),
    .X(_132_));
 sg13g2_buf_1 _439_ (.A(net44),
    .X(_133_));
 sg13g2_buf_1 _440_ (.A(net144),
    .X(_134_));
 sg13g2_buf_1 _441_ (.A(net50),
    .X(_135_));
 sg13g2_buf_1 _442_ (.A(net136),
    .X(_136_));
 sg13g2_buf_1 _443_ (.A(net94),
    .X(_137_));
 sg13g2_buf_1 _444_ (.A(net155),
    .X(_138_));
 sg13g2_buf_1 _445_ (.A(net41),
    .X(_139_));
 sg13g2_buf_1 _446_ (.A(net124),
    .X(_140_));
 sg13g2_buf_1 _447_ (.A(net83),
    .X(_141_));
 sg13g2_dfrbpq_1 _448_ (.RESET_B(net72),
    .D(_070_),
    .Q(\DP_1.matrix[0] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _449_ (.RESET_B(net72),
    .D(_071_),
    .Q(\DP_1.matrix[1] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _450_ (.RESET_B(net73),
    .D(_072_),
    .Q(\DP_1.matrix[16] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _451_ (.RESET_B(net73),
    .D(_073_),
    .Q(\DP_1.matrix[17] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _452_ (.RESET_B(net69),
    .D(_074_),
    .Q(\DP_1.matrix[32] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _453_ (.RESET_B(net69),
    .D(_075_),
    .Q(\DP_1.matrix[33] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _454_ (.RESET_B(net71),
    .D(_076_),
    .Q(\DP_1.matrix[48] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _455_ (.RESET_B(net71),
    .D(_077_),
    .Q(\DP_1.matrix[49] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _456_ (.RESET_B(net77),
    .D(_078_),
    .Q(\DP_1.matrix[64] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _457_ (.RESET_B(net77),
    .D(_079_),
    .Q(\DP_1.matrix[65] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _458_ (.RESET_B(net73),
    .D(_080_),
    .Q(\DP_1.matrix[80] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _459_ (.RESET_B(net80),
    .D(_081_),
    .Q(\DP_1.matrix[81] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _460_ (.RESET_B(net60),
    .D(_082_),
    .Q(\DP_1.matrix[96] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _461_ (.RESET_B(net67),
    .D(_083_),
    .Q(\DP_1.matrix[97] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _462_ (.RESET_B(net62),
    .D(_084_),
    .Q(\DP_1.matrix[112] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _463_ (.RESET_B(net60),
    .D(_085_),
    .Q(\DP_1.matrix[113] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _464_ (.RESET_B(net56),
    .D(_086_),
    .Q(\DP_1.matrix[128] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _465_ (.RESET_B(net56),
    .D(_087_),
    .Q(\DP_1.matrix[129] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _466_ (.RESET_B(net72),
    .D(_088_),
    .Q(\DP_2.matrix[0] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _467_ (.RESET_B(net72),
    .D(_089_),
    .Q(\DP_2.matrix[1] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _468_ (.RESET_B(net73),
    .D(_090_),
    .Q(\DP_2.matrix[16] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _469_ (.RESET_B(net74),
    .D(_091_),
    .Q(\DP_2.matrix[17] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _470_ (.RESET_B(net69),
    .D(_092_),
    .Q(\DP_2.matrix[32] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _471_ (.RESET_B(net69),
    .D(_093_),
    .Q(\DP_2.matrix[33] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _472_ (.RESET_B(net71),
    .D(_094_),
    .Q(\DP_2.matrix[48] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _473_ (.RESET_B(net71),
    .D(_095_),
    .Q(\DP_2.matrix[49] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _474_ (.RESET_B(net77),
    .D(_096_),
    .Q(\DP_2.matrix[64] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _475_ (.RESET_B(net77),
    .D(_097_),
    .Q(\DP_2.matrix[65] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _476_ (.RESET_B(net78),
    .D(_098_),
    .Q(\DP_2.matrix[80] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _477_ (.RESET_B(net78),
    .D(_099_),
    .Q(\DP_2.matrix[81] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _478_ (.RESET_B(net60),
    .D(_100_),
    .Q(\DP_2.matrix[96] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _479_ (.RESET_B(net67),
    .D(_101_),
    .Q(\DP_2.matrix[97] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _480_ (.RESET_B(net60),
    .D(_102_),
    .Q(\DP_2.matrix[112] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _481_ (.RESET_B(net60),
    .D(_103_),
    .Q(\DP_2.matrix[113] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _482_ (.RESET_B(net59),
    .D(_104_),
    .Q(\DP_2.matrix[128] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _483_ (.RESET_B(net59),
    .D(_105_),
    .Q(\DP_2.matrix[129] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _484_ (.RESET_B(net78),
    .D(_106_),
    .Q(\DP_3.matrix[0] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _485_ (.RESET_B(net78),
    .D(_107_),
    .Q(\DP_3.matrix[1] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _486_ (.RESET_B(net79),
    .D(_108_),
    .Q(\DP_3.matrix[16] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _487_ (.RESET_B(net79),
    .D(_109_),
    .Q(\DP_3.matrix[17] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _488_ (.RESET_B(net76),
    .D(_110_),
    .Q(\DP_3.matrix[32] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _489_ (.RESET_B(net76),
    .D(_111_),
    .Q(\DP_3.matrix[33] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _490_ (.RESET_B(net66),
    .D(_112_),
    .Q(\DP_3.matrix[48] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _491_ (.RESET_B(net66),
    .D(_113_),
    .Q(\DP_3.matrix[49] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _492_ (.RESET_B(net68),
    .D(_114_),
    .Q(\DP_3.matrix[64] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _493_ (.RESET_B(net63),
    .D(_115_),
    .Q(\DP_3.matrix[65] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _494_ (.RESET_B(net65),
    .D(_116_),
    .Q(\DP_3.matrix[80] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _495_ (.RESET_B(net65),
    .D(_117_),
    .Q(\DP_3.matrix[81] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _496_ (.RESET_B(net63),
    .D(_118_),
    .Q(\DP_3.matrix[96] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _497_ (.RESET_B(net63),
    .D(_119_),
    .Q(\DP_3.matrix[97] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _498_ (.RESET_B(net64),
    .D(_120_),
    .Q(\DP_3.matrix[112] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _499_ (.RESET_B(net64),
    .D(_121_),
    .Q(\DP_3.matrix[113] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _500_ (.RESET_B(net57),
    .D(_122_),
    .Q(\DP_3.matrix[128] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _501_ (.RESET_B(net57),
    .D(_123_),
    .Q(\DP_3.matrix[129] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _502_ (.RESET_B(net78),
    .D(_124_),
    .Q(\DP_4.matrix[0] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _503_ (.RESET_B(net78),
    .D(_125_),
    .Q(\DP_4.matrix[1] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _504_ (.RESET_B(net79),
    .D(_126_),
    .Q(\DP_4.matrix[16] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _505_ (.RESET_B(net79),
    .D(_127_),
    .Q(\DP_4.matrix[17] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _506_ (.RESET_B(net76),
    .D(_128_),
    .Q(\DP_4.matrix[32] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _507_ (.RESET_B(net76),
    .D(_129_),
    .Q(\DP_4.matrix[33] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _508_ (.RESET_B(net66),
    .D(_130_),
    .Q(\DP_4.matrix[48] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _509_ (.RESET_B(net66),
    .D(_131_),
    .Q(\DP_4.matrix[49] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _510_ (.RESET_B(net68),
    .D(_132_),
    .Q(\DP_4.matrix[64] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _511_ (.RESET_B(net63),
    .D(_133_),
    .Q(\DP_4.matrix[65] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _512_ (.RESET_B(net65),
    .D(_134_),
    .Q(\DP_4.matrix[80] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _513_ (.RESET_B(net65),
    .D(_135_),
    .Q(\DP_4.matrix[81] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _514_ (.RESET_B(net63),
    .D(_136_),
    .Q(\DP_4.matrix[96] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _515_ (.RESET_B(net63),
    .D(_137_),
    .Q(\DP_4.matrix[97] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _516_ (.RESET_B(net64),
    .D(_138_),
    .Q(\DP_4.matrix[112] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _517_ (.RESET_B(net64),
    .D(_139_),
    .Q(\DP_4.matrix[113] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _518_ (.RESET_B(net57),
    .D(_140_),
    .Q(\DP_4.matrix[128] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _519_ (.RESET_B(net57),
    .D(_141_),
    .Q(\DP_4.matrix[129] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _520_ (.RESET_B(net73),
    .D(_048_),
    .Q(\mac1.products_ff[80] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _521_ (.RESET_B(net78),
    .D(_049_),
    .Q(\mac1.products_ff[81] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _522_ (.RESET_B(net77),
    .D(_050_),
    .Q(\mac1.products_ff[64] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _523_ (.RESET_B(net77),
    .D(_051_),
    .Q(\mac1.products_ff[65] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _524_ (.RESET_B(net73),
    .D(net127),
    .Q(\mac1.sum_lvl1_ff[0] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _525_ (.RESET_B(net72),
    .D(net179),
    .Q(\mac1.sum_lvl1_ff[1] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _526_ (.RESET_B(net71),
    .D(net110),
    .Q(\mac1.sum_lvl1_ff[8] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _527_ (.RESET_B(net71),
    .D(net183),
    .Q(\mac1.sum_lvl1_ff[9] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _528_ (.RESET_B(net59),
    .D(_058_),
    .Q(\mac1.products_ff[128] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _529_ (.RESET_B(net61),
    .D(_059_),
    .Q(\mac1.products_ff[129] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _530_ (.RESET_B(net70),
    .D(net98),
    .Q(\mac1.sum_lvl1_ff[16] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _531_ (.RESET_B(net70),
    .D(net190),
    .Q(\mac1.sum_lvl1_ff[17] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _532_ (.RESET_B(net71),
    .D(_052_),
    .Q(\mac1.products_ff[48] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _533_ (.RESET_B(net71),
    .D(_053_),
    .Q(\mac1.products_ff[49] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _534_ (.RESET_B(net70),
    .D(net38),
    .Q(\mac1.sum_lvl1_ff[24] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _535_ (.RESET_B(net70),
    .D(net195),
    .Q(\mac1.sum_lvl1_ff[25] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _536_ (.RESET_B(net61),
    .D(net35),
    .Q(\mac1.sum_lvl1_ff[32] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _537_ (.RESET_B(net61),
    .D(net27),
    .Q(\mac1.sum_lvl1_ff[33] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _538_ (.RESET_B(net62),
    .D(_062_),
    .Q(\mac1.products_ff[112] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _539_ (.RESET_B(net60),
    .D(_063_),
    .Q(\mac1.products_ff[113] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _540_ (.RESET_B(net70),
    .D(_054_),
    .Q(\mac1.products_ff[32] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _541_ (.RESET_B(net69),
    .D(_055_),
    .Q(\mac1.products_ff[33] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _542_ (.RESET_B(net69),
    .D(net130),
    .Q(\mac1.sum_lvl2_ff[0] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _543_ (.RESET_B(net73),
    .D(net192),
    .Q(\mac1.sum_lvl2_ff[1] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _544_ (.RESET_B(net74),
    .D(_056_),
    .Q(\mac1.products_ff[16] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _545_ (.RESET_B(net73),
    .D(_057_),
    .Q(\mac1.products_ff[17] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _546_ (.RESET_B(net70),
    .D(net103),
    .Q(\mac1.sum_lvl2_ff[4] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _547_ (.RESET_B(net70),
    .D(net174),
    .Q(\mac1.sum_lvl2_ff[5] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _548_ (.RESET_B(net61),
    .D(net34),
    .Q(\mac1.sum_lvl2_ff[8] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _549_ (.RESET_B(net61),
    .D(net26),
    .Q(\mac1.sum_lvl2_ff[9] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _550_ (.RESET_B(net72),
    .D(_042_),
    .Q(\mac1.products_ff[0] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _551_ (.RESET_B(net72),
    .D(_043_),
    .Q(\mac1.products_ff[1] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _552_ (.RESET_B(net75),
    .D(_046_),
    .Q(\mac1.products_ff[96] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _553_ (.RESET_B(net75),
    .D(_047_),
    .Q(\mac1.products_ff[97] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _554_ (.RESET_B(net56),
    .D(net166),
    .Q(\mac1.total_sum[0] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _555_ (.RESET_B(net56),
    .D(net206),
    .Q(\mac1.total_sum[1] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _556_ (.RESET_B(net56),
    .D(net169),
    .Q(\mac1.total_sum[2] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _557_ (.RESET_B(net69),
    .D(net116),
    .Q(\mac1.sum_lvl3_ff[0] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _558_ (.RESET_B(net69),
    .D(net204),
    .Q(\mac1.sum_lvl3_ff[1] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _559_ (.RESET_B(net61),
    .D(net31),
    .Q(\mac1.sum_lvl3_ff[2] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _560_ (.RESET_B(net61),
    .D(net29),
    .Q(\mac1.sum_lvl3_ff[3] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _561_ (.RESET_B(net65),
    .D(_038_),
    .Q(\mac2.products_ff[80] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _562_ (.RESET_B(net65),
    .D(_039_),
    .Q(\mac2.products_ff[81] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _563_ (.RESET_B(net63),
    .D(_060_),
    .Q(\mac2.products_ff[64] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _564_ (.RESET_B(net68),
    .D(_061_),
    .Q(\mac2.products_ff[65] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_2 _565_ (.RESET_B(net78),
    .D(net148),
    .Q(\mac2.sum_lvl1_ff[0] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _566_ (.RESET_B(net79),
    .D(net202),
    .Q(\mac2.sum_lvl1_ff[1] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _567_ (.RESET_B(net81),
    .D(net118),
    .Q(\mac2.sum_lvl1_ff[8] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _568_ (.RESET_B(net77),
    .D(net185),
    .Q(\mac2.sum_lvl1_ff[9] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _569_ (.RESET_B(net57),
    .D(_036_),
    .Q(\mac2.products_ff[128] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _570_ (.RESET_B(net57),
    .D(_037_),
    .Q(\mac2.products_ff[129] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _571_ (.RESET_B(net65),
    .D(net112),
    .Q(\mac2.sum_lvl1_ff[16] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _572_ (.RESET_B(net65),
    .D(net177),
    .Q(\mac2.sum_lvl1_ff[17] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _573_ (.RESET_B(net76),
    .D(_064_),
    .Q(\mac2.products_ff[48] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _574_ (.RESET_B(net76),
    .D(_065_),
    .Q(\mac2.products_ff[49] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _575_ (.RESET_B(net67),
    .D(net114),
    .Q(\mac2.sum_lvl1_ff[24] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _576_ (.RESET_B(net67),
    .D(net181),
    .Q(\mac2.sum_lvl1_ff[25] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _577_ (.RESET_B(net57),
    .D(net28),
    .Q(\mac2.sum_lvl1_ff[32] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _578_ (.RESET_B(net58),
    .D(net32),
    .Q(\mac2.sum_lvl1_ff[33] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _579_ (.RESET_B(net64),
    .D(_034_),
    .Q(\mac2.products_ff[112] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _580_ (.RESET_B(net64),
    .D(_035_),
    .Q(\mac2.products_ff[113] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _581_ (.RESET_B(net76),
    .D(_066_),
    .Q(\mac2.products_ff[32] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _582_ (.RESET_B(net76),
    .D(_067_),
    .Q(\mac2.products_ff[33] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _583_ (.RESET_B(net67),
    .D(net122),
    .Q(\mac2.sum_lvl2_ff[0] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _584_ (.RESET_B(net67),
    .D(net200),
    .Q(\mac2.sum_lvl2_ff[1] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _585_ (.RESET_B(net79),
    .D(_068_),
    .Q(\mac2.products_ff[16] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _586_ (.RESET_B(net79),
    .D(_069_),
    .Q(\mac2.products_ff[17] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _587_ (.RESET_B(net67),
    .D(net106),
    .Q(\mac2.sum_lvl2_ff[4] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _588_ (.RESET_B(net67),
    .D(net187),
    .Q(\mac2.sum_lvl2_ff[5] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _589_ (.RESET_B(net57),
    .D(net30),
    .Q(\mac2.sum_lvl2_ff[8] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _590_ (.RESET_B(net58),
    .D(net25),
    .Q(\mac2.sum_lvl2_ff[9] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _591_ (.RESET_B(net79),
    .D(_044_),
    .Q(\mac2.products_ff[0] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _592_ (.RESET_B(net80),
    .D(_045_),
    .Q(\mac2.products_ff[1] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _593_ (.RESET_B(net64),
    .D(_040_),
    .Q(\mac2.products_ff[96] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _594_ (.RESET_B(net63),
    .D(_041_),
    .Q(\mac2.products_ff[97] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _595_ (.RESET_B(net56),
    .D(net108),
    .Q(\mac2.total_sum[0] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _596_ (.RESET_B(net56),
    .D(net208),
    .Q(\mac2.total_sum[1] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _597_ (.RESET_B(net56),
    .D(net172),
    .Q(\mac2.total_sum[2] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _598_ (.RESET_B(net60),
    .D(net153),
    .Q(\mac2.sum_lvl3_ff[0] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_2 _599_ (.RESET_B(net60),
    .D(net197),
    .Q(\mac2.sum_lvl3_ff[1] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _600_ (.RESET_B(net58),
    .D(net36),
    .Q(\mac2.sum_lvl3_ff[2] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _601_ (.RESET_B(net58),
    .D(net33),
    .Q(\mac2.sum_lvl3_ff[3] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_tiehi heichips25_template_18 (.L_HI(net18));
 sg13g2_tiehi heichips25_template_19 (.L_HI(net19));
 sg13g2_tiehi heichips25_template_20 (.L_HI(net20));
 sg13g2_tiehi heichips25_template_21 (.L_HI(net21));
 sg13g2_tiehi heichips25_template_22 (.L_HI(net22));
 sg13g2_tiehi heichips25_template_23 (.L_HI(net23));
 sg13g2_tiehi heichips25_template_24 (.L_HI(net24));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo heichips25_template_6 (.L_LO(net6));
 sg13g2_tielo heichips25_template_7 (.L_LO(net7));
 sg13g2_tielo heichips25_template_8 (.L_LO(net8));
 sg13g2_tielo heichips25_template_9 (.L_LO(net9));
 sg13g2_tielo heichips25_template_10 (.L_LO(net10));
 sg13g2_tielo heichips25_template_11 (.L_LO(net11));
 sg13g2_tielo heichips25_template_12 (.L_LO(net12));
 sg13g2_tielo heichips25_template_13 (.L_LO(net13));
 sg13g2_tielo heichips25_template_14 (.L_LO(net14));
 sg13g2_tielo heichips25_template_15 (.L_LO(net15));
 sg13g2_tielo heichips25_template_16 (.L_LO(net16));
 sg13g2_tiehi heichips25_template_17 (.L_HI(net17));
 sg13g2_buf_8 fanout56 (.A(net59),
    .X(net56));
 sg13g2_buf_8 fanout57 (.A(net59),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(net59),
    .X(net58));
 sg13g2_buf_8 fanout59 (.A(net62),
    .X(net59));
 sg13g2_buf_8 fanout60 (.A(net61),
    .X(net60));
 sg13g2_buf_8 fanout61 (.A(net62),
    .X(net61));
 sg13g2_buf_8 fanout62 (.A(rst_n),
    .X(net62));
 sg13g2_buf_8 fanout63 (.A(net64),
    .X(net63));
 sg13g2_buf_8 fanout64 (.A(net68),
    .X(net64));
 sg13g2_buf_8 fanout65 (.A(net68),
    .X(net65));
 sg13g2_buf_1 fanout66 (.A(net68),
    .X(net66));
 sg13g2_buf_8 fanout67 (.A(net68),
    .X(net67));
 sg13g2_buf_8 fanout68 (.A(rst_n),
    .X(net68));
 sg13g2_buf_8 fanout69 (.A(net70),
    .X(net69));
 sg13g2_buf_8 fanout70 (.A(net75),
    .X(net70));
 sg13g2_buf_8 fanout71 (.A(net74),
    .X(net71));
 sg13g2_buf_8 fanout72 (.A(net74),
    .X(net72));
 sg13g2_buf_8 fanout73 (.A(net74),
    .X(net73));
 sg13g2_buf_8 fanout74 (.A(net75),
    .X(net74));
 sg13g2_buf_8 fanout75 (.A(net81),
    .X(net75));
 sg13g2_buf_8 fanout76 (.A(net77),
    .X(net76));
 sg13g2_buf_8 fanout77 (.A(net81),
    .X(net77));
 sg13g2_buf_8 fanout78 (.A(net80),
    .X(net78));
 sg13g2_buf_8 fanout79 (.A(net80),
    .X(net79));
 sg13g2_buf_8 fanout80 (.A(net81),
    .X(net80));
 sg13g2_buf_8 fanout81 (.A(rst_n),
    .X(net81));
 sg13g2_buf_1 output1 (.A(net1),
    .X(uo_out[0]));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uo_out[1]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[2]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[3]));
 sg13g2_tielo heichips25_template_5 (.L_LO(net5));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_8 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_8 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_8 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_8 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_8 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_8 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_8 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_8 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_8 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_8 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_8 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_8 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_8 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_8 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_8 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_8 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_8 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_8 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_8 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_8 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_8 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_8 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_8 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_8 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_8 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_8 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_8 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_8 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_8 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_8 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_8 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_5_12__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\mac2.sum_lvl1_ff[33] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold2 (.A(\mac1.sum_lvl1_ff[33] ),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold3 (.A(\mac1.products_ff[129] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold4 (.A(\mac2.products_ff[128] ),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold5 (.A(\mac1.sum_lvl2_ff[9] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold6 (.A(\mac2.sum_lvl1_ff[32] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold7 (.A(\mac1.sum_lvl2_ff[8] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold8 (.A(\mac2.products_ff[129] ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold9 (.A(\mac2.sum_lvl2_ff[9] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold10 (.A(\mac1.sum_lvl1_ff[32] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold11 (.A(\mac1.products_ff[128] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold12 (.A(\mac2.sum_lvl2_ff[8] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold13 (.A(\mac1.products_ff[96] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold14 (.A(_006_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold15 (.A(\DP_4.matrix[17] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold16 (.A(\DP_1.matrix[17] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold17 (.A(\DP_4.matrix[113] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold18 (.A(\DP_3.matrix[49] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold19 (.A(\DP_3.matrix[113] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold20 (.A(\DP_4.matrix[65] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold21 (.A(\DP_3.matrix[1] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold22 (.A(\DP_1.matrix[1] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold23 (.A(\DP_1.matrix[113] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold24 (.A(\DP_1.matrix[97] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold25 (.A(\DP_2.matrix[17] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold26 (.A(\DP_4.matrix[81] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold27 (.A(\DP_4.matrix[1] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold28 (.A(\DP_3.matrix[81] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold29 (.A(\DP_2.matrix[33] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold30 (.A(\DP_4.matrix[33] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold31 (.A(\DP_2.matrix[1] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold32 (.A(\DP_3.matrix[17] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold33 (.A(\DP_4.matrix[129] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold34 (.A(\DP_2.matrix[81] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold35 (.A(\DP_3.matrix[97] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold36 (.A(\DP_1.matrix[49] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold37 (.A(\DP_3.matrix[129] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold38 (.A(\DP_2.matrix[113] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold39 (.A(\DP_1.matrix[81] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold40 (.A(\DP_4.matrix[49] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold41 (.A(\DP_2.matrix[65] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold42 (.A(\DP_1.matrix[33] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold43 (.A(\DP_3.matrix[65] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold44 (.A(\DP_4.matrix[97] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold45 (.A(\DP_2.matrix[97] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold46 (.A(\DP_2.matrix[129] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold47 (.A(\mac1.products_ff[64] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold48 (.A(_004_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold49 (.A(\DP_3.matrix[33] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold50 (.A(\DP_2.matrix[49] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold51 (.A(\DP_1.matrix[65] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold52 (.A(\mac1.sum_lvl1_ff[16] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold53 (.A(_010_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold54 (.A(\DP_1.matrix[129] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold55 (.A(\mac2.sum_lvl1_ff[16] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold56 (.A(_027_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold57 (.A(\mac2.sum_lvl3_ff[2] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold58 (.A(_032_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold59 (.A(\mac1.products_ff[48] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold60 (.A(_002_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold61 (.A(\mac2.products_ff[64] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold62 (.A(_021_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold63 (.A(\mac2.products_ff[112] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold64 (.A(_023_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold65 (.A(\mac1.sum_lvl2_ff[0] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold66 (.A(_012_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold67 (.A(\mac2.products_ff[32] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold68 (.A(_019_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold69 (.A(\DP_1.matrix[128] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold70 (.A(\DP_2.matrix[112] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold71 (.A(\mac2.sum_lvl1_ff[8] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold72 (.A(_025_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold73 (.A(\DP_2.matrix[32] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold74 (.A(\DP_4.matrix[128] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold75 (.A(\DP_3.matrix[112] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold76 (.A(\mac1.products_ff[16] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold77 (.A(_000_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold78 (.A(\DP_1.matrix[16] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold79 (.A(\mac1.sum_lvl1_ff[0] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold80 (.A(_008_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold81 (.A(\DP_1.matrix[64] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold82 (.A(\DP_2.matrix[48] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold83 (.A(\DP_4.matrix[16] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold84 (.A(\DP_4.matrix[64] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold85 (.A(\DP_2.matrix[16] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold86 (.A(\DP_4.matrix[96] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold87 (.A(\DP_3.matrix[96] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold88 (.A(\DP_3.matrix[80] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold89 (.A(\DP_4.matrix[32] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold90 (.A(\DP_2.matrix[96] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold91 (.A(\DP_3.matrix[64] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold92 (.A(\DP_3.matrix[128] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold93 (.A(\DP_4.matrix[0] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold94 (.A(\DP_4.matrix[80] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold95 (.A(\DP_4.matrix[48] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold96 (.A(\DP_3.matrix[0] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold97 (.A(\mac2.products_ff[0] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold98 (.A(_017_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold99 (.A(\DP_3.matrix[48] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold100 (.A(\DP_2.matrix[128] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold101 (.A(\DP_1.matrix[96] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold102 (.A(\mac2.sum_lvl2_ff[0] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold103 (.A(_029_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold104 (.A(\DP_1.matrix[0] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold105 (.A(\DP_4.matrix[112] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold106 (.A(\DP_2.matrix[0] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold107 (.A(\DP_2.matrix[64] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold108 (.A(\DP_2.matrix[80] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold109 (.A(\DP_1.matrix[112] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold110 (.A(\DP_1.matrix[32] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold111 (.A(\DP_3.matrix[16] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold112 (.A(\DP_1.matrix[80] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold113 (.A(\DP_3.matrix[32] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold114 (.A(\DP_1.matrix[48] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold115 (.A(\mac1.sum_lvl3_ff[0] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold116 (.A(_015_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold117 (.A(\mac1.sum_lvl3_ff[3] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold118 (.A(_167_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold119 (.A(_014_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold120 (.A(\mac2.sum_lvl3_ff[1] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold121 (.A(_183_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold122 (.A(_031_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold123 (.A(\mac1.sum_lvl1_ff[24] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold124 (.A(_011_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold125 (.A(\mac2.products_ff[81] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold126 (.A(_179_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold127 (.A(_022_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold128 (.A(\mac1.products_ff[0] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold129 (.A(_001_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold130 (.A(\mac2.products_ff[96] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold131 (.A(_024_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold132 (.A(\mac1.products_ff[32] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold133 (.A(_003_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold134 (.A(\mac2.products_ff[48] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold135 (.A(_020_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold136 (.A(\mac2.sum_lvl1_ff[24] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold137 (.A(_028_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold138 (.A(\mac1.products_ff[65] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold139 (.A(_161_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold140 (.A(_005_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold141 (.A(\mac1.sum_lvl1_ff[8] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold142 (.A(_009_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold143 (.A(\mac1.products_ff[97] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold144 (.A(_159_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold145 (.A(_007_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold146 (.A(\mac2.sum_lvl2_ff[4] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold147 (.A(_030_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold148 (.A(\mac2.sum_lvl1_ff[1] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold149 (.A(_175_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold150 (.A(_026_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold151 (.A(\mac2.products_ff[16] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold152 (.A(_018_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold153 (.A(\mac1.sum_lvl2_ff[4] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold154 (.A(_013_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold155 (.A(\mac1.sum_lvl3_ff[2] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold156 (.A(_016_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold157 (.A(\mac2.sum_lvl3_ff[0] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold158 (.A(_033_),
    .X(net208));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_decap_8 FILLER_0_875 ();
 sg13g2_decap_8 FILLER_0_882 ();
 sg13g2_decap_8 FILLER_0_889 ();
 sg13g2_decap_8 FILLER_0_896 ();
 sg13g2_decap_8 FILLER_0_903 ();
 sg13g2_decap_8 FILLER_0_910 ();
 sg13g2_decap_8 FILLER_0_917 ();
 sg13g2_decap_8 FILLER_0_924 ();
 sg13g2_decap_8 FILLER_0_931 ();
 sg13g2_decap_8 FILLER_0_938 ();
 sg13g2_decap_8 FILLER_0_945 ();
 sg13g2_decap_8 FILLER_0_952 ();
 sg13g2_decap_8 FILLER_0_959 ();
 sg13g2_decap_8 FILLER_0_966 ();
 sg13g2_decap_8 FILLER_0_973 ();
 sg13g2_decap_8 FILLER_0_980 ();
 sg13g2_decap_8 FILLER_0_987 ();
 sg13g2_decap_8 FILLER_0_994 ();
 sg13g2_decap_8 FILLER_0_1001 ();
 sg13g2_decap_8 FILLER_0_1008 ();
 sg13g2_decap_8 FILLER_0_1015 ();
 sg13g2_decap_8 FILLER_0_1022 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_4 FILLER_1_126 ();
 sg13g2_fill_2 FILLER_1_130 ();
 sg13g2_decap_8 FILLER_1_136 ();
 sg13g2_decap_8 FILLER_1_143 ();
 sg13g2_decap_8 FILLER_1_150 ();
 sg13g2_decap_8 FILLER_1_157 ();
 sg13g2_decap_8 FILLER_1_164 ();
 sg13g2_decap_8 FILLER_1_171 ();
 sg13g2_decap_8 FILLER_1_178 ();
 sg13g2_decap_8 FILLER_1_185 ();
 sg13g2_decap_8 FILLER_1_192 ();
 sg13g2_decap_8 FILLER_1_199 ();
 sg13g2_decap_8 FILLER_1_206 ();
 sg13g2_decap_8 FILLER_1_213 ();
 sg13g2_decap_8 FILLER_1_220 ();
 sg13g2_decap_8 FILLER_1_227 ();
 sg13g2_decap_8 FILLER_1_234 ();
 sg13g2_decap_8 FILLER_1_241 ();
 sg13g2_decap_8 FILLER_1_248 ();
 sg13g2_decap_8 FILLER_1_255 ();
 sg13g2_decap_8 FILLER_1_262 ();
 sg13g2_decap_8 FILLER_1_269 ();
 sg13g2_decap_8 FILLER_1_276 ();
 sg13g2_decap_8 FILLER_1_283 ();
 sg13g2_decap_8 FILLER_1_290 ();
 sg13g2_decap_8 FILLER_1_297 ();
 sg13g2_decap_8 FILLER_1_304 ();
 sg13g2_decap_8 FILLER_1_311 ();
 sg13g2_decap_8 FILLER_1_318 ();
 sg13g2_decap_8 FILLER_1_325 ();
 sg13g2_decap_8 FILLER_1_332 ();
 sg13g2_decap_8 FILLER_1_339 ();
 sg13g2_decap_8 FILLER_1_346 ();
 sg13g2_decap_8 FILLER_1_353 ();
 sg13g2_decap_8 FILLER_1_360 ();
 sg13g2_decap_8 FILLER_1_367 ();
 sg13g2_decap_8 FILLER_1_374 ();
 sg13g2_decap_8 FILLER_1_381 ();
 sg13g2_decap_8 FILLER_1_388 ();
 sg13g2_decap_8 FILLER_1_395 ();
 sg13g2_decap_8 FILLER_1_402 ();
 sg13g2_decap_8 FILLER_1_409 ();
 sg13g2_decap_8 FILLER_1_416 ();
 sg13g2_decap_8 FILLER_1_423 ();
 sg13g2_decap_8 FILLER_1_430 ();
 sg13g2_decap_8 FILLER_1_437 ();
 sg13g2_decap_8 FILLER_1_444 ();
 sg13g2_decap_8 FILLER_1_451 ();
 sg13g2_decap_8 FILLER_1_458 ();
 sg13g2_decap_8 FILLER_1_465 ();
 sg13g2_decap_8 FILLER_1_472 ();
 sg13g2_decap_8 FILLER_1_479 ();
 sg13g2_decap_8 FILLER_1_486 ();
 sg13g2_decap_8 FILLER_1_493 ();
 sg13g2_decap_8 FILLER_1_500 ();
 sg13g2_decap_8 FILLER_1_507 ();
 sg13g2_decap_8 FILLER_1_514 ();
 sg13g2_decap_8 FILLER_1_521 ();
 sg13g2_decap_8 FILLER_1_528 ();
 sg13g2_decap_8 FILLER_1_535 ();
 sg13g2_decap_8 FILLER_1_542 ();
 sg13g2_decap_8 FILLER_1_549 ();
 sg13g2_decap_8 FILLER_1_556 ();
 sg13g2_decap_8 FILLER_1_563 ();
 sg13g2_decap_8 FILLER_1_570 ();
 sg13g2_decap_8 FILLER_1_577 ();
 sg13g2_decap_8 FILLER_1_584 ();
 sg13g2_decap_8 FILLER_1_591 ();
 sg13g2_decap_8 FILLER_1_598 ();
 sg13g2_decap_8 FILLER_1_605 ();
 sg13g2_decap_8 FILLER_1_612 ();
 sg13g2_decap_8 FILLER_1_619 ();
 sg13g2_decap_8 FILLER_1_626 ();
 sg13g2_decap_8 FILLER_1_633 ();
 sg13g2_decap_8 FILLER_1_640 ();
 sg13g2_decap_8 FILLER_1_647 ();
 sg13g2_decap_8 FILLER_1_654 ();
 sg13g2_decap_8 FILLER_1_661 ();
 sg13g2_decap_8 FILLER_1_668 ();
 sg13g2_decap_8 FILLER_1_675 ();
 sg13g2_decap_8 FILLER_1_682 ();
 sg13g2_decap_8 FILLER_1_689 ();
 sg13g2_decap_8 FILLER_1_696 ();
 sg13g2_decap_8 FILLER_1_703 ();
 sg13g2_decap_8 FILLER_1_710 ();
 sg13g2_decap_8 FILLER_1_717 ();
 sg13g2_decap_8 FILLER_1_724 ();
 sg13g2_decap_8 FILLER_1_731 ();
 sg13g2_decap_8 FILLER_1_738 ();
 sg13g2_decap_8 FILLER_1_745 ();
 sg13g2_decap_8 FILLER_1_752 ();
 sg13g2_decap_8 FILLER_1_759 ();
 sg13g2_decap_8 FILLER_1_766 ();
 sg13g2_decap_8 FILLER_1_773 ();
 sg13g2_decap_8 FILLER_1_780 ();
 sg13g2_decap_8 FILLER_1_787 ();
 sg13g2_decap_8 FILLER_1_794 ();
 sg13g2_decap_8 FILLER_1_801 ();
 sg13g2_decap_8 FILLER_1_808 ();
 sg13g2_decap_8 FILLER_1_815 ();
 sg13g2_decap_8 FILLER_1_822 ();
 sg13g2_decap_8 FILLER_1_829 ();
 sg13g2_decap_8 FILLER_1_836 ();
 sg13g2_decap_8 FILLER_1_843 ();
 sg13g2_decap_8 FILLER_1_850 ();
 sg13g2_decap_8 FILLER_1_857 ();
 sg13g2_decap_8 FILLER_1_864 ();
 sg13g2_decap_8 FILLER_1_871 ();
 sg13g2_decap_8 FILLER_1_878 ();
 sg13g2_decap_8 FILLER_1_885 ();
 sg13g2_decap_8 FILLER_1_892 ();
 sg13g2_decap_8 FILLER_1_899 ();
 sg13g2_decap_8 FILLER_1_906 ();
 sg13g2_decap_8 FILLER_1_913 ();
 sg13g2_decap_8 FILLER_1_920 ();
 sg13g2_decap_8 FILLER_1_927 ();
 sg13g2_decap_8 FILLER_1_934 ();
 sg13g2_decap_8 FILLER_1_941 ();
 sg13g2_decap_8 FILLER_1_948 ();
 sg13g2_decap_8 FILLER_1_955 ();
 sg13g2_decap_8 FILLER_1_962 ();
 sg13g2_decap_8 FILLER_1_969 ();
 sg13g2_decap_8 FILLER_1_976 ();
 sg13g2_decap_8 FILLER_1_983 ();
 sg13g2_decap_8 FILLER_1_990 ();
 sg13g2_decap_8 FILLER_1_997 ();
 sg13g2_decap_8 FILLER_1_1004 ();
 sg13g2_decap_8 FILLER_1_1011 ();
 sg13g2_decap_8 FILLER_1_1018 ();
 sg13g2_decap_4 FILLER_1_1025 ();
 sg13g2_decap_8 FILLER_2_4 ();
 sg13g2_decap_8 FILLER_2_11 ();
 sg13g2_decap_8 FILLER_2_18 ();
 sg13g2_decap_8 FILLER_2_25 ();
 sg13g2_decap_8 FILLER_2_32 ();
 sg13g2_decap_8 FILLER_2_39 ();
 sg13g2_decap_8 FILLER_2_46 ();
 sg13g2_decap_8 FILLER_2_53 ();
 sg13g2_decap_8 FILLER_2_60 ();
 sg13g2_decap_8 FILLER_2_67 ();
 sg13g2_decap_8 FILLER_2_74 ();
 sg13g2_decap_8 FILLER_2_81 ();
 sg13g2_decap_8 FILLER_2_88 ();
 sg13g2_decap_8 FILLER_2_95 ();
 sg13g2_decap_8 FILLER_2_102 ();
 sg13g2_decap_8 FILLER_2_109 ();
 sg13g2_decap_4 FILLER_2_116 ();
 sg13g2_fill_1 FILLER_2_120 ();
 sg13g2_decap_8 FILLER_2_157 ();
 sg13g2_decap_4 FILLER_2_164 ();
 sg13g2_fill_1 FILLER_2_168 ();
 sg13g2_fill_2 FILLER_2_173 ();
 sg13g2_fill_2 FILLER_2_179 ();
 sg13g2_fill_2 FILLER_2_185 ();
 sg13g2_fill_1 FILLER_2_187 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_fill_1 FILLER_2_210 ();
 sg13g2_fill_2 FILLER_2_238 ();
 sg13g2_fill_1 FILLER_2_240 ();
 sg13g2_fill_1 FILLER_2_277 ();
 sg13g2_decap_8 FILLER_2_314 ();
 sg13g2_decap_8 FILLER_2_321 ();
 sg13g2_decap_8 FILLER_2_328 ();
 sg13g2_decap_8 FILLER_2_335 ();
 sg13g2_decap_8 FILLER_2_342 ();
 sg13g2_decap_8 FILLER_2_349 ();
 sg13g2_decap_8 FILLER_2_356 ();
 sg13g2_decap_8 FILLER_2_363 ();
 sg13g2_decap_8 FILLER_2_370 ();
 sg13g2_decap_8 FILLER_2_377 ();
 sg13g2_decap_4 FILLER_2_384 ();
 sg13g2_fill_2 FILLER_2_388 ();
 sg13g2_decap_8 FILLER_2_444 ();
 sg13g2_decap_8 FILLER_2_451 ();
 sg13g2_decap_4 FILLER_2_458 ();
 sg13g2_decap_8 FILLER_2_516 ();
 sg13g2_decap_8 FILLER_2_523 ();
 sg13g2_fill_2 FILLER_2_530 ();
 sg13g2_fill_1 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_564 ();
 sg13g2_decap_8 FILLER_2_571 ();
 sg13g2_decap_8 FILLER_2_578 ();
 sg13g2_decap_8 FILLER_2_585 ();
 sg13g2_decap_8 FILLER_2_592 ();
 sg13g2_decap_8 FILLER_2_599 ();
 sg13g2_decap_8 FILLER_2_606 ();
 sg13g2_decap_8 FILLER_2_613 ();
 sg13g2_decap_8 FILLER_2_620 ();
 sg13g2_decap_8 FILLER_2_627 ();
 sg13g2_decap_8 FILLER_2_634 ();
 sg13g2_decap_8 FILLER_2_641 ();
 sg13g2_decap_8 FILLER_2_648 ();
 sg13g2_decap_8 FILLER_2_655 ();
 sg13g2_decap_8 FILLER_2_662 ();
 sg13g2_decap_8 FILLER_2_669 ();
 sg13g2_decap_8 FILLER_2_676 ();
 sg13g2_decap_8 FILLER_2_683 ();
 sg13g2_decap_8 FILLER_2_690 ();
 sg13g2_decap_8 FILLER_2_697 ();
 sg13g2_decap_8 FILLER_2_704 ();
 sg13g2_decap_8 FILLER_2_711 ();
 sg13g2_decap_8 FILLER_2_718 ();
 sg13g2_decap_8 FILLER_2_725 ();
 sg13g2_decap_8 FILLER_2_732 ();
 sg13g2_decap_8 FILLER_2_739 ();
 sg13g2_decap_8 FILLER_2_746 ();
 sg13g2_decap_8 FILLER_2_753 ();
 sg13g2_decap_8 FILLER_2_760 ();
 sg13g2_decap_8 FILLER_2_767 ();
 sg13g2_decap_8 FILLER_2_774 ();
 sg13g2_decap_8 FILLER_2_781 ();
 sg13g2_decap_8 FILLER_2_788 ();
 sg13g2_decap_8 FILLER_2_795 ();
 sg13g2_decap_8 FILLER_2_802 ();
 sg13g2_decap_8 FILLER_2_809 ();
 sg13g2_decap_8 FILLER_2_816 ();
 sg13g2_decap_8 FILLER_2_823 ();
 sg13g2_decap_8 FILLER_2_830 ();
 sg13g2_decap_8 FILLER_2_837 ();
 sg13g2_decap_8 FILLER_2_844 ();
 sg13g2_decap_8 FILLER_2_851 ();
 sg13g2_decap_8 FILLER_2_858 ();
 sg13g2_decap_8 FILLER_2_865 ();
 sg13g2_decap_8 FILLER_2_872 ();
 sg13g2_decap_8 FILLER_2_879 ();
 sg13g2_decap_8 FILLER_2_886 ();
 sg13g2_decap_8 FILLER_2_893 ();
 sg13g2_decap_8 FILLER_2_900 ();
 sg13g2_decap_8 FILLER_2_907 ();
 sg13g2_decap_8 FILLER_2_914 ();
 sg13g2_decap_8 FILLER_2_921 ();
 sg13g2_decap_8 FILLER_2_928 ();
 sg13g2_decap_8 FILLER_2_935 ();
 sg13g2_decap_8 FILLER_2_942 ();
 sg13g2_decap_8 FILLER_2_949 ();
 sg13g2_decap_8 FILLER_2_956 ();
 sg13g2_decap_8 FILLER_2_963 ();
 sg13g2_decap_8 FILLER_2_970 ();
 sg13g2_decap_8 FILLER_2_977 ();
 sg13g2_decap_8 FILLER_2_984 ();
 sg13g2_decap_8 FILLER_2_991 ();
 sg13g2_decap_8 FILLER_2_998 ();
 sg13g2_decap_8 FILLER_2_1005 ();
 sg13g2_decap_8 FILLER_2_1012 ();
 sg13g2_decap_8 FILLER_2_1019 ();
 sg13g2_fill_2 FILLER_2_1026 ();
 sg13g2_fill_1 FILLER_2_1028 ();
 sg13g2_decap_8 FILLER_3_4 ();
 sg13g2_decap_8 FILLER_3_11 ();
 sg13g2_decap_8 FILLER_3_18 ();
 sg13g2_decap_8 FILLER_3_25 ();
 sg13g2_decap_8 FILLER_3_32 ();
 sg13g2_decap_8 FILLER_3_39 ();
 sg13g2_decap_8 FILLER_3_46 ();
 sg13g2_decap_8 FILLER_3_53 ();
 sg13g2_decap_8 FILLER_3_60 ();
 sg13g2_decap_8 FILLER_3_67 ();
 sg13g2_decap_8 FILLER_3_74 ();
 sg13g2_decap_8 FILLER_3_81 ();
 sg13g2_decap_8 FILLER_3_88 ();
 sg13g2_decap_8 FILLER_3_95 ();
 sg13g2_decap_8 FILLER_3_102 ();
 sg13g2_decap_8 FILLER_3_109 ();
 sg13g2_decap_8 FILLER_3_143 ();
 sg13g2_decap_8 FILLER_3_150 ();
 sg13g2_decap_4 FILLER_3_157 ();
 sg13g2_fill_2 FILLER_3_161 ();
 sg13g2_decap_4 FILLER_3_190 ();
 sg13g2_fill_1 FILLER_3_194 ();
 sg13g2_decap_8 FILLER_3_222 ();
 sg13g2_decap_8 FILLER_3_229 ();
 sg13g2_decap_8 FILLER_3_236 ();
 sg13g2_decap_8 FILLER_3_243 ();
 sg13g2_decap_8 FILLER_3_250 ();
 sg13g2_decap_8 FILLER_3_257 ();
 sg13g2_decap_8 FILLER_3_264 ();
 sg13g2_decap_8 FILLER_3_271 ();
 sg13g2_decap_8 FILLER_3_278 ();
 sg13g2_decap_8 FILLER_3_285 ();
 sg13g2_decap_8 FILLER_3_292 ();
 sg13g2_decap_8 FILLER_3_299 ();
 sg13g2_decap_8 FILLER_3_306 ();
 sg13g2_decap_4 FILLER_3_313 ();
 sg13g2_decap_8 FILLER_3_345 ();
 sg13g2_decap_8 FILLER_3_352 ();
 sg13g2_decap_8 FILLER_3_359 ();
 sg13g2_decap_8 FILLER_3_366 ();
 sg13g2_decap_8 FILLER_3_373 ();
 sg13g2_decap_8 FILLER_3_380 ();
 sg13g2_decap_8 FILLER_3_387 ();
 sg13g2_decap_8 FILLER_3_394 ();
 sg13g2_fill_1 FILLER_3_401 ();
 sg13g2_decap_4 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_410 ();
 sg13g2_decap_8 FILLER_3_433 ();
 sg13g2_decap_8 FILLER_3_440 ();
 sg13g2_decap_8 FILLER_3_447 ();
 sg13g2_decap_8 FILLER_3_454 ();
 sg13g2_decap_8 FILLER_3_461 ();
 sg13g2_fill_2 FILLER_3_468 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_fill_2 FILLER_3_497 ();
 sg13g2_fill_2 FILLER_3_503 ();
 sg13g2_decap_8 FILLER_3_522 ();
 sg13g2_decap_8 FILLER_3_529 ();
 sg13g2_decap_8 FILLER_3_536 ();
 sg13g2_decap_4 FILLER_3_543 ();
 sg13g2_fill_2 FILLER_3_547 ();
 sg13g2_decap_8 FILLER_3_558 ();
 sg13g2_decap_8 FILLER_3_565 ();
 sg13g2_decap_8 FILLER_3_572 ();
 sg13g2_decap_8 FILLER_3_579 ();
 sg13g2_decap_8 FILLER_3_586 ();
 sg13g2_decap_8 FILLER_3_593 ();
 sg13g2_decap_8 FILLER_3_600 ();
 sg13g2_decap_8 FILLER_3_607 ();
 sg13g2_decap_8 FILLER_3_614 ();
 sg13g2_decap_8 FILLER_3_621 ();
 sg13g2_decap_8 FILLER_3_628 ();
 sg13g2_decap_8 FILLER_3_635 ();
 sg13g2_decap_8 FILLER_3_642 ();
 sg13g2_decap_8 FILLER_3_649 ();
 sg13g2_decap_8 FILLER_3_656 ();
 sg13g2_decap_8 FILLER_3_663 ();
 sg13g2_decap_8 FILLER_3_670 ();
 sg13g2_decap_8 FILLER_3_677 ();
 sg13g2_decap_8 FILLER_3_684 ();
 sg13g2_decap_8 FILLER_3_691 ();
 sg13g2_decap_8 FILLER_3_698 ();
 sg13g2_decap_8 FILLER_3_705 ();
 sg13g2_decap_8 FILLER_3_712 ();
 sg13g2_decap_8 FILLER_3_719 ();
 sg13g2_decap_8 FILLER_3_726 ();
 sg13g2_decap_8 FILLER_3_733 ();
 sg13g2_decap_8 FILLER_3_740 ();
 sg13g2_decap_8 FILLER_3_747 ();
 sg13g2_decap_8 FILLER_3_754 ();
 sg13g2_decap_8 FILLER_3_761 ();
 sg13g2_decap_8 FILLER_3_768 ();
 sg13g2_decap_8 FILLER_3_775 ();
 sg13g2_decap_8 FILLER_3_782 ();
 sg13g2_decap_8 FILLER_3_789 ();
 sg13g2_decap_8 FILLER_3_796 ();
 sg13g2_decap_8 FILLER_3_803 ();
 sg13g2_decap_8 FILLER_3_810 ();
 sg13g2_decap_8 FILLER_3_817 ();
 sg13g2_decap_8 FILLER_3_824 ();
 sg13g2_decap_8 FILLER_3_831 ();
 sg13g2_decap_8 FILLER_3_838 ();
 sg13g2_decap_8 FILLER_3_845 ();
 sg13g2_decap_8 FILLER_3_852 ();
 sg13g2_decap_8 FILLER_3_859 ();
 sg13g2_decap_8 FILLER_3_866 ();
 sg13g2_decap_8 FILLER_3_873 ();
 sg13g2_decap_8 FILLER_3_880 ();
 sg13g2_decap_8 FILLER_3_887 ();
 sg13g2_decap_8 FILLER_3_894 ();
 sg13g2_decap_8 FILLER_3_901 ();
 sg13g2_decap_8 FILLER_3_908 ();
 sg13g2_decap_8 FILLER_3_915 ();
 sg13g2_decap_8 FILLER_3_922 ();
 sg13g2_decap_8 FILLER_3_929 ();
 sg13g2_decap_8 FILLER_3_936 ();
 sg13g2_decap_8 FILLER_3_943 ();
 sg13g2_decap_8 FILLER_3_950 ();
 sg13g2_decap_8 FILLER_3_957 ();
 sg13g2_decap_8 FILLER_3_964 ();
 sg13g2_decap_8 FILLER_3_971 ();
 sg13g2_decap_8 FILLER_3_978 ();
 sg13g2_decap_8 FILLER_3_985 ();
 sg13g2_decap_8 FILLER_3_992 ();
 sg13g2_decap_8 FILLER_3_999 ();
 sg13g2_decap_8 FILLER_3_1006 ();
 sg13g2_decap_8 FILLER_3_1013 ();
 sg13g2_decap_8 FILLER_3_1020 ();
 sg13g2_fill_2 FILLER_3_1027 ();
 sg13g2_decap_8 FILLER_4_4 ();
 sg13g2_decap_8 FILLER_4_11 ();
 sg13g2_decap_8 FILLER_4_18 ();
 sg13g2_decap_8 FILLER_4_25 ();
 sg13g2_decap_8 FILLER_4_32 ();
 sg13g2_decap_8 FILLER_4_43 ();
 sg13g2_decap_8 FILLER_4_50 ();
 sg13g2_decap_8 FILLER_4_57 ();
 sg13g2_decap_8 FILLER_4_64 ();
 sg13g2_decap_8 FILLER_4_71 ();
 sg13g2_decap_8 FILLER_4_78 ();
 sg13g2_decap_8 FILLER_4_85 ();
 sg13g2_decap_8 FILLER_4_92 ();
 sg13g2_decap_8 FILLER_4_99 ();
 sg13g2_decap_8 FILLER_4_106 ();
 sg13g2_decap_8 FILLER_4_113 ();
 sg13g2_decap_4 FILLER_4_120 ();
 sg13g2_fill_2 FILLER_4_124 ();
 sg13g2_decap_8 FILLER_4_130 ();
 sg13g2_decap_8 FILLER_4_137 ();
 sg13g2_decap_8 FILLER_4_144 ();
 sg13g2_decap_8 FILLER_4_151 ();
 sg13g2_decap_4 FILLER_4_158 ();
 sg13g2_fill_1 FILLER_4_162 ();
 sg13g2_decap_4 FILLER_4_172 ();
 sg13g2_decap_8 FILLER_4_190 ();
 sg13g2_decap_8 FILLER_4_197 ();
 sg13g2_decap_8 FILLER_4_204 ();
 sg13g2_decap_8 FILLER_4_211 ();
 sg13g2_decap_8 FILLER_4_218 ();
 sg13g2_decap_8 FILLER_4_225 ();
 sg13g2_decap_8 FILLER_4_268 ();
 sg13g2_decap_8 FILLER_4_275 ();
 sg13g2_decap_8 FILLER_4_282 ();
 sg13g2_decap_8 FILLER_4_289 ();
 sg13g2_decap_8 FILLER_4_296 ();
 sg13g2_decap_8 FILLER_4_303 ();
 sg13g2_decap_4 FILLER_4_310 ();
 sg13g2_fill_2 FILLER_4_314 ();
 sg13g2_decap_8 FILLER_4_325 ();
 sg13g2_decap_8 FILLER_4_332 ();
 sg13g2_decap_8 FILLER_4_339 ();
 sg13g2_decap_8 FILLER_4_346 ();
 sg13g2_decap_8 FILLER_4_353 ();
 sg13g2_decap_8 FILLER_4_360 ();
 sg13g2_decap_8 FILLER_4_367 ();
 sg13g2_decap_8 FILLER_4_374 ();
 sg13g2_decap_8 FILLER_4_381 ();
 sg13g2_decap_8 FILLER_4_388 ();
 sg13g2_decap_8 FILLER_4_395 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_4_409 ();
 sg13g2_decap_4 FILLER_4_416 ();
 sg13g2_fill_1 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_425 ();
 sg13g2_decap_8 FILLER_4_432 ();
 sg13g2_decap_8 FILLER_4_439 ();
 sg13g2_decap_8 FILLER_4_446 ();
 sg13g2_decap_8 FILLER_4_453 ();
 sg13g2_decap_8 FILLER_4_460 ();
 sg13g2_decap_8 FILLER_4_467 ();
 sg13g2_decap_8 FILLER_4_474 ();
 sg13g2_decap_8 FILLER_4_481 ();
 sg13g2_decap_8 FILLER_4_488 ();
 sg13g2_decap_8 FILLER_4_495 ();
 sg13g2_fill_2 FILLER_4_502 ();
 sg13g2_decap_8 FILLER_4_512 ();
 sg13g2_decap_8 FILLER_4_519 ();
 sg13g2_decap_8 FILLER_4_526 ();
 sg13g2_fill_1 FILLER_4_533 ();
 sg13g2_decap_8 FILLER_4_538 ();
 sg13g2_decap_8 FILLER_4_545 ();
 sg13g2_decap_8 FILLER_4_552 ();
 sg13g2_decap_8 FILLER_4_559 ();
 sg13g2_decap_8 FILLER_4_566 ();
 sg13g2_decap_8 FILLER_4_573 ();
 sg13g2_decap_8 FILLER_4_580 ();
 sg13g2_decap_8 FILLER_4_587 ();
 sg13g2_decap_8 FILLER_4_594 ();
 sg13g2_decap_8 FILLER_4_601 ();
 sg13g2_decap_8 FILLER_4_608 ();
 sg13g2_decap_8 FILLER_4_615 ();
 sg13g2_decap_8 FILLER_4_622 ();
 sg13g2_decap_8 FILLER_4_629 ();
 sg13g2_decap_8 FILLER_4_636 ();
 sg13g2_decap_8 FILLER_4_643 ();
 sg13g2_decap_8 FILLER_4_650 ();
 sg13g2_decap_8 FILLER_4_657 ();
 sg13g2_decap_8 FILLER_4_664 ();
 sg13g2_decap_8 FILLER_4_671 ();
 sg13g2_decap_8 FILLER_4_678 ();
 sg13g2_decap_8 FILLER_4_685 ();
 sg13g2_decap_8 FILLER_4_692 ();
 sg13g2_decap_8 FILLER_4_699 ();
 sg13g2_decap_8 FILLER_4_706 ();
 sg13g2_decap_8 FILLER_4_713 ();
 sg13g2_decap_8 FILLER_4_720 ();
 sg13g2_decap_8 FILLER_4_727 ();
 sg13g2_decap_8 FILLER_4_734 ();
 sg13g2_decap_8 FILLER_4_741 ();
 sg13g2_decap_8 FILLER_4_748 ();
 sg13g2_decap_8 FILLER_4_755 ();
 sg13g2_decap_8 FILLER_4_762 ();
 sg13g2_decap_8 FILLER_4_769 ();
 sg13g2_decap_8 FILLER_4_776 ();
 sg13g2_decap_8 FILLER_4_783 ();
 sg13g2_decap_8 FILLER_4_790 ();
 sg13g2_decap_8 FILLER_4_797 ();
 sg13g2_decap_8 FILLER_4_804 ();
 sg13g2_decap_8 FILLER_4_811 ();
 sg13g2_decap_8 FILLER_4_818 ();
 sg13g2_decap_8 FILLER_4_825 ();
 sg13g2_decap_8 FILLER_4_832 ();
 sg13g2_decap_8 FILLER_4_839 ();
 sg13g2_decap_8 FILLER_4_846 ();
 sg13g2_decap_8 FILLER_4_853 ();
 sg13g2_decap_8 FILLER_4_860 ();
 sg13g2_decap_8 FILLER_4_867 ();
 sg13g2_decap_8 FILLER_4_874 ();
 sg13g2_decap_8 FILLER_4_881 ();
 sg13g2_decap_8 FILLER_4_888 ();
 sg13g2_decap_8 FILLER_4_895 ();
 sg13g2_decap_8 FILLER_4_902 ();
 sg13g2_decap_8 FILLER_4_909 ();
 sg13g2_decap_8 FILLER_4_916 ();
 sg13g2_decap_8 FILLER_4_923 ();
 sg13g2_decap_8 FILLER_4_930 ();
 sg13g2_decap_8 FILLER_4_937 ();
 sg13g2_decap_8 FILLER_4_944 ();
 sg13g2_decap_8 FILLER_4_951 ();
 sg13g2_decap_8 FILLER_4_958 ();
 sg13g2_decap_8 FILLER_4_965 ();
 sg13g2_decap_8 FILLER_4_972 ();
 sg13g2_decap_8 FILLER_4_979 ();
 sg13g2_decap_8 FILLER_4_986 ();
 sg13g2_decap_8 FILLER_4_993 ();
 sg13g2_decap_8 FILLER_4_1000 ();
 sg13g2_decap_8 FILLER_4_1007 ();
 sg13g2_decap_8 FILLER_4_1014 ();
 sg13g2_decap_8 FILLER_4_1021 ();
 sg13g2_fill_1 FILLER_4_1028 ();
 sg13g2_fill_2 FILLER_5_4 ();
 sg13g2_fill_1 FILLER_5_6 ();
 sg13g2_decap_4 FILLER_5_61 ();
 sg13g2_fill_1 FILLER_5_65 ();
 sg13g2_decap_8 FILLER_5_93 ();
 sg13g2_decap_8 FILLER_5_100 ();
 sg13g2_decap_8 FILLER_5_107 ();
 sg13g2_decap_8 FILLER_5_114 ();
 sg13g2_decap_8 FILLER_5_121 ();
 sg13g2_decap_8 FILLER_5_128 ();
 sg13g2_decap_8 FILLER_5_135 ();
 sg13g2_decap_8 FILLER_5_142 ();
 sg13g2_decap_8 FILLER_5_149 ();
 sg13g2_decap_8 FILLER_5_156 ();
 sg13g2_decap_8 FILLER_5_163 ();
 sg13g2_decap_8 FILLER_5_170 ();
 sg13g2_decap_8 FILLER_5_177 ();
 sg13g2_decap_8 FILLER_5_184 ();
 sg13g2_decap_8 FILLER_5_191 ();
 sg13g2_decap_8 FILLER_5_198 ();
 sg13g2_decap_8 FILLER_5_205 ();
 sg13g2_decap_8 FILLER_5_212 ();
 sg13g2_decap_8 FILLER_5_219 ();
 sg13g2_decap_8 FILLER_5_226 ();
 sg13g2_decap_8 FILLER_5_233 ();
 sg13g2_decap_8 FILLER_5_240 ();
 sg13g2_decap_8 FILLER_5_247 ();
 sg13g2_decap_8 FILLER_5_254 ();
 sg13g2_decap_8 FILLER_5_261 ();
 sg13g2_decap_4 FILLER_5_268 ();
 sg13g2_fill_1 FILLER_5_272 ();
 sg13g2_decap_8 FILLER_5_309 ();
 sg13g2_decap_8 FILLER_5_316 ();
 sg13g2_decap_8 FILLER_5_323 ();
 sg13g2_decap_8 FILLER_5_330 ();
 sg13g2_decap_8 FILLER_5_337 ();
 sg13g2_decap_8 FILLER_5_344 ();
 sg13g2_decap_8 FILLER_5_351 ();
 sg13g2_decap_8 FILLER_5_358 ();
 sg13g2_fill_2 FILLER_5_365 ();
 sg13g2_fill_1 FILLER_5_367 ();
 sg13g2_decap_8 FILLER_5_395 ();
 sg13g2_fill_2 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_5_436 ();
 sg13g2_decap_8 FILLER_5_443 ();
 sg13g2_decap_8 FILLER_5_450 ();
 sg13g2_decap_8 FILLER_5_457 ();
 sg13g2_decap_8 FILLER_5_464 ();
 sg13g2_decap_8 FILLER_5_471 ();
 sg13g2_decap_8 FILLER_5_478 ();
 sg13g2_decap_8 FILLER_5_485 ();
 sg13g2_decap_8 FILLER_5_492 ();
 sg13g2_decap_8 FILLER_5_499 ();
 sg13g2_decap_8 FILLER_5_506 ();
 sg13g2_fill_2 FILLER_5_513 ();
 sg13g2_decap_8 FILLER_5_520 ();
 sg13g2_decap_8 FILLER_5_527 ();
 sg13g2_decap_8 FILLER_5_561 ();
 sg13g2_decap_8 FILLER_5_568 ();
 sg13g2_decap_8 FILLER_5_575 ();
 sg13g2_decap_8 FILLER_5_582 ();
 sg13g2_decap_8 FILLER_5_589 ();
 sg13g2_decap_8 FILLER_5_596 ();
 sg13g2_decap_8 FILLER_5_603 ();
 sg13g2_decap_8 FILLER_5_610 ();
 sg13g2_decap_8 FILLER_5_617 ();
 sg13g2_decap_8 FILLER_5_624 ();
 sg13g2_decap_8 FILLER_5_631 ();
 sg13g2_decap_8 FILLER_5_638 ();
 sg13g2_decap_8 FILLER_5_645 ();
 sg13g2_decap_8 FILLER_5_652 ();
 sg13g2_decap_8 FILLER_5_659 ();
 sg13g2_decap_8 FILLER_5_666 ();
 sg13g2_decap_8 FILLER_5_673 ();
 sg13g2_decap_8 FILLER_5_680 ();
 sg13g2_decap_8 FILLER_5_687 ();
 sg13g2_decap_8 FILLER_5_694 ();
 sg13g2_decap_8 FILLER_5_701 ();
 sg13g2_decap_8 FILLER_5_708 ();
 sg13g2_decap_8 FILLER_5_715 ();
 sg13g2_decap_8 FILLER_5_722 ();
 sg13g2_decap_8 FILLER_5_729 ();
 sg13g2_decap_8 FILLER_5_736 ();
 sg13g2_decap_8 FILLER_5_743 ();
 sg13g2_decap_8 FILLER_5_750 ();
 sg13g2_decap_8 FILLER_5_757 ();
 sg13g2_decap_8 FILLER_5_764 ();
 sg13g2_decap_8 FILLER_5_771 ();
 sg13g2_decap_8 FILLER_5_778 ();
 sg13g2_decap_8 FILLER_5_785 ();
 sg13g2_decap_8 FILLER_5_792 ();
 sg13g2_decap_8 FILLER_5_799 ();
 sg13g2_decap_8 FILLER_5_806 ();
 sg13g2_decap_8 FILLER_5_813 ();
 sg13g2_decap_8 FILLER_5_820 ();
 sg13g2_decap_8 FILLER_5_827 ();
 sg13g2_decap_8 FILLER_5_834 ();
 sg13g2_decap_8 FILLER_5_841 ();
 sg13g2_decap_8 FILLER_5_848 ();
 sg13g2_decap_8 FILLER_5_855 ();
 sg13g2_decap_8 FILLER_5_862 ();
 sg13g2_decap_8 FILLER_5_869 ();
 sg13g2_decap_8 FILLER_5_876 ();
 sg13g2_decap_8 FILLER_5_883 ();
 sg13g2_decap_8 FILLER_5_890 ();
 sg13g2_decap_8 FILLER_5_897 ();
 sg13g2_decap_8 FILLER_5_904 ();
 sg13g2_decap_8 FILLER_5_911 ();
 sg13g2_decap_8 FILLER_5_918 ();
 sg13g2_decap_8 FILLER_5_925 ();
 sg13g2_decap_8 FILLER_5_932 ();
 sg13g2_decap_8 FILLER_5_939 ();
 sg13g2_decap_8 FILLER_5_946 ();
 sg13g2_decap_8 FILLER_5_953 ();
 sg13g2_decap_8 FILLER_5_960 ();
 sg13g2_decap_8 FILLER_5_967 ();
 sg13g2_decap_8 FILLER_5_974 ();
 sg13g2_decap_8 FILLER_5_981 ();
 sg13g2_decap_8 FILLER_5_988 ();
 sg13g2_decap_8 FILLER_5_995 ();
 sg13g2_decap_8 FILLER_5_1002 ();
 sg13g2_decap_8 FILLER_5_1009 ();
 sg13g2_decap_8 FILLER_5_1016 ();
 sg13g2_decap_4 FILLER_5_1023 ();
 sg13g2_fill_2 FILLER_5_1027 ();
 sg13g2_decap_8 FILLER_6_4 ();
 sg13g2_decap_4 FILLER_6_11 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_4 FILLER_6_35 ();
 sg13g2_fill_1 FILLER_6_39 ();
 sg13g2_fill_2 FILLER_6_44 ();
 sg13g2_decap_8 FILLER_6_60 ();
 sg13g2_decap_8 FILLER_6_67 ();
 sg13g2_decap_8 FILLER_6_74 ();
 sg13g2_decap_8 FILLER_6_81 ();
 sg13g2_decap_8 FILLER_6_88 ();
 sg13g2_decap_8 FILLER_6_131 ();
 sg13g2_decap_8 FILLER_6_138 ();
 sg13g2_decap_8 FILLER_6_145 ();
 sg13g2_decap_8 FILLER_6_152 ();
 sg13g2_decap_8 FILLER_6_159 ();
 sg13g2_fill_1 FILLER_6_166 ();
 sg13g2_decap_4 FILLER_6_194 ();
 sg13g2_decap_8 FILLER_6_211 ();
 sg13g2_decap_8 FILLER_6_218 ();
 sg13g2_decap_8 FILLER_6_225 ();
 sg13g2_decap_8 FILLER_6_232 ();
 sg13g2_decap_8 FILLER_6_239 ();
 sg13g2_decap_8 FILLER_6_246 ();
 sg13g2_decap_8 FILLER_6_253 ();
 sg13g2_decap_8 FILLER_6_260 ();
 sg13g2_decap_8 FILLER_6_267 ();
 sg13g2_decap_8 FILLER_6_274 ();
 sg13g2_decap_8 FILLER_6_281 ();
 sg13g2_decap_8 FILLER_6_288 ();
 sg13g2_decap_8 FILLER_6_295 ();
 sg13g2_decap_4 FILLER_6_302 ();
 sg13g2_fill_2 FILLER_6_306 ();
 sg13g2_decap_8 FILLER_6_344 ();
 sg13g2_decap_8 FILLER_6_351 ();
 sg13g2_decap_8 FILLER_6_358 ();
 sg13g2_decap_8 FILLER_6_365 ();
 sg13g2_fill_2 FILLER_6_372 ();
 sg13g2_decap_8 FILLER_6_387 ();
 sg13g2_decap_8 FILLER_6_394 ();
 sg13g2_fill_2 FILLER_6_401 ();
 sg13g2_decap_8 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_6_414 ();
 sg13g2_decap_8 FILLER_6_421 ();
 sg13g2_decap_4 FILLER_6_428 ();
 sg13g2_fill_1 FILLER_6_432 ();
 sg13g2_decap_8 FILLER_6_460 ();
 sg13g2_decap_8 FILLER_6_467 ();
 sg13g2_fill_2 FILLER_6_474 ();
 sg13g2_decap_8 FILLER_6_503 ();
 sg13g2_decap_8 FILLER_6_510 ();
 sg13g2_decap_8 FILLER_6_517 ();
 sg13g2_decap_8 FILLER_6_524 ();
 sg13g2_decap_8 FILLER_6_531 ();
 sg13g2_decap_8 FILLER_6_538 ();
 sg13g2_decap_4 FILLER_6_545 ();
 sg13g2_decap_8 FILLER_6_558 ();
 sg13g2_decap_8 FILLER_6_565 ();
 sg13g2_decap_8 FILLER_6_572 ();
 sg13g2_decap_8 FILLER_6_579 ();
 sg13g2_decap_8 FILLER_6_586 ();
 sg13g2_decap_8 FILLER_6_593 ();
 sg13g2_decap_8 FILLER_6_600 ();
 sg13g2_decap_8 FILLER_6_607 ();
 sg13g2_decap_8 FILLER_6_614 ();
 sg13g2_decap_8 FILLER_6_621 ();
 sg13g2_decap_8 FILLER_6_628 ();
 sg13g2_decap_8 FILLER_6_635 ();
 sg13g2_decap_8 FILLER_6_642 ();
 sg13g2_decap_8 FILLER_6_649 ();
 sg13g2_decap_8 FILLER_6_656 ();
 sg13g2_decap_8 FILLER_6_663 ();
 sg13g2_decap_8 FILLER_6_670 ();
 sg13g2_decap_8 FILLER_6_677 ();
 sg13g2_decap_8 FILLER_6_684 ();
 sg13g2_decap_8 FILLER_6_691 ();
 sg13g2_decap_8 FILLER_6_698 ();
 sg13g2_decap_8 FILLER_6_705 ();
 sg13g2_decap_8 FILLER_6_712 ();
 sg13g2_decap_8 FILLER_6_719 ();
 sg13g2_decap_8 FILLER_6_726 ();
 sg13g2_decap_8 FILLER_6_733 ();
 sg13g2_decap_8 FILLER_6_740 ();
 sg13g2_decap_8 FILLER_6_747 ();
 sg13g2_decap_8 FILLER_6_754 ();
 sg13g2_decap_8 FILLER_6_761 ();
 sg13g2_decap_8 FILLER_6_768 ();
 sg13g2_decap_8 FILLER_6_775 ();
 sg13g2_decap_8 FILLER_6_782 ();
 sg13g2_decap_8 FILLER_6_789 ();
 sg13g2_decap_8 FILLER_6_796 ();
 sg13g2_decap_8 FILLER_6_803 ();
 sg13g2_decap_8 FILLER_6_810 ();
 sg13g2_decap_8 FILLER_6_817 ();
 sg13g2_decap_8 FILLER_6_824 ();
 sg13g2_decap_8 FILLER_6_831 ();
 sg13g2_decap_8 FILLER_6_838 ();
 sg13g2_decap_8 FILLER_6_845 ();
 sg13g2_decap_8 FILLER_6_852 ();
 sg13g2_decap_8 FILLER_6_859 ();
 sg13g2_decap_8 FILLER_6_866 ();
 sg13g2_decap_8 FILLER_6_873 ();
 sg13g2_decap_8 FILLER_6_880 ();
 sg13g2_decap_8 FILLER_6_887 ();
 sg13g2_decap_8 FILLER_6_894 ();
 sg13g2_decap_8 FILLER_6_901 ();
 sg13g2_decap_8 FILLER_6_908 ();
 sg13g2_decap_8 FILLER_6_915 ();
 sg13g2_decap_8 FILLER_6_922 ();
 sg13g2_decap_8 FILLER_6_929 ();
 sg13g2_decap_8 FILLER_6_936 ();
 sg13g2_decap_8 FILLER_6_943 ();
 sg13g2_decap_8 FILLER_6_950 ();
 sg13g2_decap_8 FILLER_6_957 ();
 sg13g2_decap_8 FILLER_6_964 ();
 sg13g2_decap_8 FILLER_6_971 ();
 sg13g2_decap_8 FILLER_6_978 ();
 sg13g2_decap_8 FILLER_6_985 ();
 sg13g2_decap_8 FILLER_6_992 ();
 sg13g2_decap_8 FILLER_6_999 ();
 sg13g2_decap_8 FILLER_6_1006 ();
 sg13g2_decap_8 FILLER_6_1013 ();
 sg13g2_decap_8 FILLER_6_1020 ();
 sg13g2_fill_2 FILLER_6_1027 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_fill_2 FILLER_7_91 ();
 sg13g2_fill_1 FILLER_7_93 ();
 sg13g2_decap_8 FILLER_7_103 ();
 sg13g2_decap_8 FILLER_7_110 ();
 sg13g2_fill_2 FILLER_7_117 ();
 sg13g2_fill_1 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_179 ();
 sg13g2_decap_8 FILLER_7_195 ();
 sg13g2_decap_8 FILLER_7_202 ();
 sg13g2_decap_8 FILLER_7_209 ();
 sg13g2_decap_8 FILLER_7_216 ();
 sg13g2_decap_8 FILLER_7_223 ();
 sg13g2_decap_8 FILLER_7_230 ();
 sg13g2_decap_8 FILLER_7_237 ();
 sg13g2_decap_8 FILLER_7_244 ();
 sg13g2_decap_8 FILLER_7_251 ();
 sg13g2_decap_8 FILLER_7_258 ();
 sg13g2_decap_8 FILLER_7_265 ();
 sg13g2_decap_8 FILLER_7_272 ();
 sg13g2_decap_8 FILLER_7_279 ();
 sg13g2_decap_8 FILLER_7_286 ();
 sg13g2_decap_8 FILLER_7_293 ();
 sg13g2_decap_8 FILLER_7_300 ();
 sg13g2_decap_8 FILLER_7_307 ();
 sg13g2_decap_8 FILLER_7_314 ();
 sg13g2_decap_8 FILLER_7_321 ();
 sg13g2_decap_8 FILLER_7_328 ();
 sg13g2_decap_8 FILLER_7_335 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_fill_2 FILLER_7_385 ();
 sg13g2_fill_1 FILLER_7_387 ();
 sg13g2_fill_2 FILLER_7_415 ();
 sg13g2_decap_8 FILLER_7_422 ();
 sg13g2_decap_8 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_7_436 ();
 sg13g2_decap_8 FILLER_7_443 ();
 sg13g2_decap_8 FILLER_7_450 ();
 sg13g2_decap_8 FILLER_7_457 ();
 sg13g2_decap_8 FILLER_7_464 ();
 sg13g2_decap_4 FILLER_7_471 ();
 sg13g2_fill_2 FILLER_7_475 ();
 sg13g2_decap_8 FILLER_7_485 ();
 sg13g2_decap_8 FILLER_7_492 ();
 sg13g2_decap_8 FILLER_7_499 ();
 sg13g2_decap_8 FILLER_7_506 ();
 sg13g2_decap_8 FILLER_7_513 ();
 sg13g2_decap_8 FILLER_7_520 ();
 sg13g2_decap_8 FILLER_7_527 ();
 sg13g2_decap_8 FILLER_7_534 ();
 sg13g2_decap_8 FILLER_7_541 ();
 sg13g2_decap_8 FILLER_7_548 ();
 sg13g2_decap_8 FILLER_7_555 ();
 sg13g2_decap_8 FILLER_7_562 ();
 sg13g2_decap_8 FILLER_7_569 ();
 sg13g2_decap_8 FILLER_7_576 ();
 sg13g2_decap_8 FILLER_7_583 ();
 sg13g2_decap_8 FILLER_7_590 ();
 sg13g2_decap_8 FILLER_7_597 ();
 sg13g2_decap_8 FILLER_7_604 ();
 sg13g2_decap_8 FILLER_7_611 ();
 sg13g2_decap_8 FILLER_7_618 ();
 sg13g2_decap_8 FILLER_7_625 ();
 sg13g2_decap_8 FILLER_7_632 ();
 sg13g2_decap_8 FILLER_7_639 ();
 sg13g2_decap_8 FILLER_7_646 ();
 sg13g2_decap_8 FILLER_7_653 ();
 sg13g2_decap_8 FILLER_7_660 ();
 sg13g2_decap_8 FILLER_7_667 ();
 sg13g2_decap_8 FILLER_7_674 ();
 sg13g2_decap_8 FILLER_7_681 ();
 sg13g2_decap_8 FILLER_7_688 ();
 sg13g2_decap_8 FILLER_7_695 ();
 sg13g2_decap_8 FILLER_7_702 ();
 sg13g2_decap_8 FILLER_7_709 ();
 sg13g2_decap_8 FILLER_7_716 ();
 sg13g2_decap_8 FILLER_7_723 ();
 sg13g2_decap_8 FILLER_7_730 ();
 sg13g2_decap_8 FILLER_7_737 ();
 sg13g2_decap_8 FILLER_7_744 ();
 sg13g2_decap_8 FILLER_7_751 ();
 sg13g2_decap_8 FILLER_7_758 ();
 sg13g2_decap_8 FILLER_7_765 ();
 sg13g2_decap_8 FILLER_7_772 ();
 sg13g2_decap_8 FILLER_7_779 ();
 sg13g2_decap_8 FILLER_7_786 ();
 sg13g2_decap_8 FILLER_7_793 ();
 sg13g2_decap_8 FILLER_7_800 ();
 sg13g2_decap_8 FILLER_7_807 ();
 sg13g2_decap_8 FILLER_7_814 ();
 sg13g2_decap_8 FILLER_7_821 ();
 sg13g2_decap_8 FILLER_7_828 ();
 sg13g2_decap_8 FILLER_7_835 ();
 sg13g2_decap_8 FILLER_7_842 ();
 sg13g2_decap_8 FILLER_7_849 ();
 sg13g2_decap_8 FILLER_7_856 ();
 sg13g2_decap_8 FILLER_7_863 ();
 sg13g2_decap_8 FILLER_7_870 ();
 sg13g2_decap_8 FILLER_7_877 ();
 sg13g2_decap_8 FILLER_7_884 ();
 sg13g2_decap_8 FILLER_7_891 ();
 sg13g2_decap_8 FILLER_7_898 ();
 sg13g2_decap_8 FILLER_7_905 ();
 sg13g2_decap_8 FILLER_7_912 ();
 sg13g2_decap_8 FILLER_7_919 ();
 sg13g2_decap_8 FILLER_7_926 ();
 sg13g2_decap_8 FILLER_7_933 ();
 sg13g2_decap_8 FILLER_7_940 ();
 sg13g2_decap_8 FILLER_7_947 ();
 sg13g2_decap_8 FILLER_7_954 ();
 sg13g2_decap_8 FILLER_7_961 ();
 sg13g2_decap_8 FILLER_7_968 ();
 sg13g2_decap_8 FILLER_7_975 ();
 sg13g2_decap_8 FILLER_7_982 ();
 sg13g2_decap_8 FILLER_7_989 ();
 sg13g2_decap_8 FILLER_7_996 ();
 sg13g2_decap_8 FILLER_7_1003 ();
 sg13g2_decap_8 FILLER_7_1010 ();
 sg13g2_decap_8 FILLER_7_1017 ();
 sg13g2_decap_4 FILLER_7_1024 ();
 sg13g2_fill_1 FILLER_7_1028 ();
 sg13g2_decap_8 FILLER_8_4 ();
 sg13g2_decap_8 FILLER_8_11 ();
 sg13g2_decap_8 FILLER_8_18 ();
 sg13g2_decap_8 FILLER_8_25 ();
 sg13g2_decap_8 FILLER_8_32 ();
 sg13g2_decap_8 FILLER_8_39 ();
 sg13g2_decap_8 FILLER_8_46 ();
 sg13g2_decap_8 FILLER_8_53 ();
 sg13g2_decap_8 FILLER_8_60 ();
 sg13g2_decap_8 FILLER_8_67 ();
 sg13g2_decap_8 FILLER_8_74 ();
 sg13g2_decap_8 FILLER_8_81 ();
 sg13g2_decap_8 FILLER_8_88 ();
 sg13g2_decap_8 FILLER_8_95 ();
 sg13g2_decap_8 FILLER_8_102 ();
 sg13g2_decap_8 FILLER_8_149 ();
 sg13g2_decap_8 FILLER_8_156 ();
 sg13g2_decap_8 FILLER_8_163 ();
 sg13g2_decap_8 FILLER_8_170 ();
 sg13g2_decap_8 FILLER_8_177 ();
 sg13g2_decap_8 FILLER_8_184 ();
 sg13g2_decap_8 FILLER_8_191 ();
 sg13g2_decap_8 FILLER_8_198 ();
 sg13g2_decap_8 FILLER_8_205 ();
 sg13g2_decap_8 FILLER_8_212 ();
 sg13g2_decap_8 FILLER_8_219 ();
 sg13g2_decap_8 FILLER_8_226 ();
 sg13g2_decap_8 FILLER_8_260 ();
 sg13g2_decap_8 FILLER_8_267 ();
 sg13g2_decap_8 FILLER_8_274 ();
 sg13g2_decap_8 FILLER_8_281 ();
 sg13g2_decap_8 FILLER_8_288 ();
 sg13g2_decap_8 FILLER_8_295 ();
 sg13g2_decap_8 FILLER_8_302 ();
 sg13g2_decap_8 FILLER_8_309 ();
 sg13g2_decap_8 FILLER_8_316 ();
 sg13g2_decap_8 FILLER_8_323 ();
 sg13g2_decap_8 FILLER_8_330 ();
 sg13g2_fill_2 FILLER_8_337 ();
 sg13g2_decap_8 FILLER_8_352 ();
 sg13g2_decap_8 FILLER_8_359 ();
 sg13g2_decap_8 FILLER_8_366 ();
 sg13g2_decap_8 FILLER_8_373 ();
 sg13g2_decap_8 FILLER_8_380 ();
 sg13g2_decap_8 FILLER_8_387 ();
 sg13g2_fill_2 FILLER_8_394 ();
 sg13g2_decap_8 FILLER_8_400 ();
 sg13g2_decap_8 FILLER_8_416 ();
 sg13g2_decap_8 FILLER_8_423 ();
 sg13g2_decap_8 FILLER_8_430 ();
 sg13g2_decap_8 FILLER_8_437 ();
 sg13g2_decap_8 FILLER_8_444 ();
 sg13g2_decap_8 FILLER_8_451 ();
 sg13g2_decap_8 FILLER_8_458 ();
 sg13g2_decap_8 FILLER_8_465 ();
 sg13g2_decap_8 FILLER_8_472 ();
 sg13g2_decap_8 FILLER_8_479 ();
 sg13g2_decap_8 FILLER_8_486 ();
 sg13g2_decap_8 FILLER_8_493 ();
 sg13g2_fill_2 FILLER_8_500 ();
 sg13g2_fill_2 FILLER_8_515 ();
 sg13g2_fill_1 FILLER_8_517 ();
 sg13g2_decap_8 FILLER_8_545 ();
 sg13g2_decap_8 FILLER_8_552 ();
 sg13g2_decap_8 FILLER_8_559 ();
 sg13g2_decap_8 FILLER_8_566 ();
 sg13g2_decap_8 FILLER_8_573 ();
 sg13g2_decap_8 FILLER_8_593 ();
 sg13g2_decap_8 FILLER_8_600 ();
 sg13g2_decap_8 FILLER_8_607 ();
 sg13g2_decap_8 FILLER_8_614 ();
 sg13g2_decap_8 FILLER_8_621 ();
 sg13g2_decap_8 FILLER_8_628 ();
 sg13g2_decap_8 FILLER_8_635 ();
 sg13g2_decap_8 FILLER_8_642 ();
 sg13g2_decap_8 FILLER_8_649 ();
 sg13g2_decap_8 FILLER_8_656 ();
 sg13g2_decap_8 FILLER_8_663 ();
 sg13g2_decap_8 FILLER_8_670 ();
 sg13g2_decap_8 FILLER_8_677 ();
 sg13g2_decap_8 FILLER_8_684 ();
 sg13g2_decap_8 FILLER_8_691 ();
 sg13g2_decap_8 FILLER_8_698 ();
 sg13g2_decap_8 FILLER_8_705 ();
 sg13g2_decap_8 FILLER_8_712 ();
 sg13g2_decap_8 FILLER_8_719 ();
 sg13g2_decap_8 FILLER_8_726 ();
 sg13g2_decap_8 FILLER_8_733 ();
 sg13g2_decap_8 FILLER_8_740 ();
 sg13g2_decap_8 FILLER_8_747 ();
 sg13g2_decap_8 FILLER_8_754 ();
 sg13g2_decap_8 FILLER_8_761 ();
 sg13g2_decap_8 FILLER_8_768 ();
 sg13g2_decap_8 FILLER_8_775 ();
 sg13g2_decap_8 FILLER_8_782 ();
 sg13g2_decap_8 FILLER_8_789 ();
 sg13g2_decap_8 FILLER_8_796 ();
 sg13g2_decap_8 FILLER_8_803 ();
 sg13g2_decap_8 FILLER_8_810 ();
 sg13g2_decap_8 FILLER_8_817 ();
 sg13g2_decap_8 FILLER_8_824 ();
 sg13g2_decap_8 FILLER_8_831 ();
 sg13g2_decap_8 FILLER_8_838 ();
 sg13g2_decap_8 FILLER_8_845 ();
 sg13g2_decap_8 FILLER_8_852 ();
 sg13g2_decap_8 FILLER_8_859 ();
 sg13g2_decap_8 FILLER_8_866 ();
 sg13g2_decap_8 FILLER_8_873 ();
 sg13g2_decap_8 FILLER_8_880 ();
 sg13g2_decap_8 FILLER_8_887 ();
 sg13g2_decap_8 FILLER_8_894 ();
 sg13g2_decap_8 FILLER_8_901 ();
 sg13g2_decap_8 FILLER_8_908 ();
 sg13g2_decap_8 FILLER_8_915 ();
 sg13g2_decap_8 FILLER_8_922 ();
 sg13g2_decap_8 FILLER_8_929 ();
 sg13g2_decap_8 FILLER_8_936 ();
 sg13g2_decap_8 FILLER_8_943 ();
 sg13g2_decap_8 FILLER_8_950 ();
 sg13g2_decap_8 FILLER_8_957 ();
 sg13g2_decap_8 FILLER_8_964 ();
 sg13g2_decap_8 FILLER_8_971 ();
 sg13g2_decap_8 FILLER_8_978 ();
 sg13g2_decap_8 FILLER_8_985 ();
 sg13g2_decap_8 FILLER_8_992 ();
 sg13g2_decap_8 FILLER_8_999 ();
 sg13g2_decap_8 FILLER_8_1006 ();
 sg13g2_decap_8 FILLER_8_1013 ();
 sg13g2_decap_8 FILLER_8_1020 ();
 sg13g2_fill_2 FILLER_8_1027 ();
 sg13g2_decap_8 FILLER_9_4 ();
 sg13g2_decap_8 FILLER_9_11 ();
 sg13g2_decap_8 FILLER_9_18 ();
 sg13g2_decap_8 FILLER_9_25 ();
 sg13g2_fill_2 FILLER_9_36 ();
 sg13g2_fill_1 FILLER_9_38 ();
 sg13g2_fill_2 FILLER_9_60 ();
 sg13g2_decap_8 FILLER_9_75 ();
 sg13g2_decap_8 FILLER_9_82 ();
 sg13g2_decap_8 FILLER_9_89 ();
 sg13g2_decap_8 FILLER_9_96 ();
 sg13g2_decap_8 FILLER_9_103 ();
 sg13g2_decap_8 FILLER_9_110 ();
 sg13g2_decap_8 FILLER_9_117 ();
 sg13g2_decap_8 FILLER_9_124 ();
 sg13g2_decap_8 FILLER_9_131 ();
 sg13g2_decap_8 FILLER_9_138 ();
 sg13g2_decap_8 FILLER_9_145 ();
 sg13g2_decap_4 FILLER_9_152 ();
 sg13g2_fill_2 FILLER_9_156 ();
 sg13g2_decap_8 FILLER_9_167 ();
 sg13g2_decap_4 FILLER_9_174 ();
 sg13g2_fill_2 FILLER_9_178 ();
 sg13g2_decap_8 FILLER_9_193 ();
 sg13g2_decap_8 FILLER_9_200 ();
 sg13g2_decap_8 FILLER_9_207 ();
 sg13g2_decap_8 FILLER_9_214 ();
 sg13g2_fill_1 FILLER_9_221 ();
 sg13g2_decap_8 FILLER_9_249 ();
 sg13g2_decap_8 FILLER_9_264 ();
 sg13g2_decap_8 FILLER_9_271 ();
 sg13g2_fill_2 FILLER_9_278 ();
 sg13g2_fill_1 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_fill_2 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_354 ();
 sg13g2_decap_8 FILLER_9_361 ();
 sg13g2_decap_8 FILLER_9_368 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_8 FILLER_9_403 ();
 sg13g2_decap_8 FILLER_9_410 ();
 sg13g2_decap_8 FILLER_9_417 ();
 sg13g2_decap_8 FILLER_9_424 ();
 sg13g2_decap_8 FILLER_9_431 ();
 sg13g2_decap_8 FILLER_9_438 ();
 sg13g2_decap_8 FILLER_9_445 ();
 sg13g2_decap_8 FILLER_9_452 ();
 sg13g2_decap_8 FILLER_9_459 ();
 sg13g2_decap_8 FILLER_9_466 ();
 sg13g2_decap_4 FILLER_9_473 ();
 sg13g2_fill_1 FILLER_9_477 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_fill_2 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_508 ();
 sg13g2_decap_8 FILLER_9_515 ();
 sg13g2_decap_8 FILLER_9_522 ();
 sg13g2_decap_8 FILLER_9_529 ();
 sg13g2_decap_8 FILLER_9_536 ();
 sg13g2_decap_8 FILLER_9_543 ();
 sg13g2_decap_8 FILLER_9_550 ();
 sg13g2_decap_8 FILLER_9_557 ();
 sg13g2_decap_8 FILLER_9_564 ();
 sg13g2_fill_1 FILLER_9_571 ();
 sg13g2_decap_8 FILLER_9_576 ();
 sg13g2_decap_8 FILLER_9_583 ();
 sg13g2_decap_8 FILLER_9_590 ();
 sg13g2_decap_8 FILLER_9_597 ();
 sg13g2_decap_8 FILLER_9_604 ();
 sg13g2_decap_8 FILLER_9_611 ();
 sg13g2_decap_8 FILLER_9_618 ();
 sg13g2_decap_8 FILLER_9_625 ();
 sg13g2_decap_8 FILLER_9_632 ();
 sg13g2_decap_8 FILLER_9_639 ();
 sg13g2_decap_8 FILLER_9_646 ();
 sg13g2_decap_8 FILLER_9_653 ();
 sg13g2_decap_8 FILLER_9_660 ();
 sg13g2_decap_8 FILLER_9_667 ();
 sg13g2_decap_8 FILLER_9_674 ();
 sg13g2_decap_8 FILLER_9_681 ();
 sg13g2_decap_8 FILLER_9_688 ();
 sg13g2_decap_8 FILLER_9_695 ();
 sg13g2_decap_8 FILLER_9_702 ();
 sg13g2_decap_8 FILLER_9_709 ();
 sg13g2_decap_8 FILLER_9_716 ();
 sg13g2_decap_8 FILLER_9_723 ();
 sg13g2_decap_8 FILLER_9_730 ();
 sg13g2_decap_8 FILLER_9_737 ();
 sg13g2_decap_8 FILLER_9_744 ();
 sg13g2_decap_8 FILLER_9_751 ();
 sg13g2_decap_8 FILLER_9_758 ();
 sg13g2_decap_8 FILLER_9_765 ();
 sg13g2_decap_8 FILLER_9_772 ();
 sg13g2_decap_8 FILLER_9_779 ();
 sg13g2_decap_8 FILLER_9_786 ();
 sg13g2_decap_8 FILLER_9_793 ();
 sg13g2_decap_8 FILLER_9_800 ();
 sg13g2_decap_8 FILLER_9_807 ();
 sg13g2_decap_8 FILLER_9_814 ();
 sg13g2_decap_8 FILLER_9_821 ();
 sg13g2_decap_8 FILLER_9_828 ();
 sg13g2_decap_8 FILLER_9_835 ();
 sg13g2_decap_8 FILLER_9_842 ();
 sg13g2_decap_8 FILLER_9_849 ();
 sg13g2_decap_8 FILLER_9_856 ();
 sg13g2_decap_8 FILLER_9_863 ();
 sg13g2_decap_8 FILLER_9_870 ();
 sg13g2_decap_8 FILLER_9_877 ();
 sg13g2_decap_8 FILLER_9_884 ();
 sg13g2_decap_8 FILLER_9_891 ();
 sg13g2_decap_8 FILLER_9_898 ();
 sg13g2_decap_8 FILLER_9_905 ();
 sg13g2_decap_8 FILLER_9_912 ();
 sg13g2_decap_8 FILLER_9_919 ();
 sg13g2_decap_8 FILLER_9_926 ();
 sg13g2_decap_8 FILLER_9_933 ();
 sg13g2_decap_8 FILLER_9_940 ();
 sg13g2_decap_8 FILLER_9_947 ();
 sg13g2_decap_8 FILLER_9_954 ();
 sg13g2_decap_8 FILLER_9_961 ();
 sg13g2_decap_8 FILLER_9_968 ();
 sg13g2_decap_8 FILLER_9_975 ();
 sg13g2_decap_8 FILLER_9_982 ();
 sg13g2_decap_8 FILLER_9_989 ();
 sg13g2_decap_8 FILLER_9_996 ();
 sg13g2_decap_8 FILLER_9_1003 ();
 sg13g2_decap_8 FILLER_9_1010 ();
 sg13g2_decap_8 FILLER_9_1017 ();
 sg13g2_decap_4 FILLER_9_1024 ();
 sg13g2_fill_1 FILLER_9_1028 ();
 sg13g2_decap_8 FILLER_10_4 ();
 sg13g2_decap_8 FILLER_10_11 ();
 sg13g2_decap_4 FILLER_10_18 ();
 sg13g2_fill_2 FILLER_10_22 ();
 sg13g2_decap_8 FILLER_10_51 ();
 sg13g2_decap_8 FILLER_10_58 ();
 sg13g2_decap_8 FILLER_10_65 ();
 sg13g2_decap_8 FILLER_10_72 ();
 sg13g2_decap_8 FILLER_10_79 ();
 sg13g2_decap_8 FILLER_10_86 ();
 sg13g2_decap_8 FILLER_10_93 ();
 sg13g2_decap_8 FILLER_10_100 ();
 sg13g2_decap_8 FILLER_10_107 ();
 sg13g2_decap_8 FILLER_10_114 ();
 sg13g2_decap_8 FILLER_10_121 ();
 sg13g2_decap_8 FILLER_10_128 ();
 sg13g2_decap_8 FILLER_10_135 ();
 sg13g2_decap_8 FILLER_10_142 ();
 sg13g2_decap_8 FILLER_10_149 ();
 sg13g2_decap_8 FILLER_10_156 ();
 sg13g2_decap_4 FILLER_10_163 ();
 sg13g2_decap_8 FILLER_10_194 ();
 sg13g2_decap_8 FILLER_10_201 ();
 sg13g2_decap_8 FILLER_10_208 ();
 sg13g2_decap_8 FILLER_10_215 ();
 sg13g2_decap_8 FILLER_10_222 ();
 sg13g2_decap_8 FILLER_10_229 ();
 sg13g2_fill_1 FILLER_10_236 ();
 sg13g2_decap_8 FILLER_10_250 ();
 sg13g2_decap_4 FILLER_10_257 ();
 sg13g2_fill_2 FILLER_10_261 ();
 sg13g2_decap_8 FILLER_10_267 ();
 sg13g2_fill_2 FILLER_10_299 ();
 sg13g2_decap_8 FILLER_10_306 ();
 sg13g2_decap_8 FILLER_10_313 ();
 sg13g2_fill_2 FILLER_10_320 ();
 sg13g2_fill_1 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_332 ();
 sg13g2_decap_8 FILLER_10_355 ();
 sg13g2_decap_8 FILLER_10_362 ();
 sg13g2_decap_8 FILLER_10_369 ();
 sg13g2_decap_8 FILLER_10_376 ();
 sg13g2_fill_1 FILLER_10_383 ();
 sg13g2_decap_8 FILLER_10_397 ();
 sg13g2_decap_8 FILLER_10_404 ();
 sg13g2_decap_8 FILLER_10_411 ();
 sg13g2_decap_8 FILLER_10_418 ();
 sg13g2_decap_8 FILLER_10_425 ();
 sg13g2_decap_8 FILLER_10_459 ();
 sg13g2_fill_2 FILLER_10_466 ();
 sg13g2_fill_1 FILLER_10_468 ();
 sg13g2_decap_8 FILLER_10_486 ();
 sg13g2_decap_8 FILLER_10_493 ();
 sg13g2_decap_8 FILLER_10_500 ();
 sg13g2_decap_8 FILLER_10_507 ();
 sg13g2_decap_8 FILLER_10_514 ();
 sg13g2_decap_8 FILLER_10_521 ();
 sg13g2_decap_8 FILLER_10_528 ();
 sg13g2_decap_8 FILLER_10_535 ();
 sg13g2_decap_8 FILLER_10_542 ();
 sg13g2_decap_8 FILLER_10_549 ();
 sg13g2_fill_1 FILLER_10_556 ();
 sg13g2_fill_1 FILLER_10_584 ();
 sg13g2_decap_8 FILLER_10_594 ();
 sg13g2_decap_8 FILLER_10_601 ();
 sg13g2_decap_8 FILLER_10_608 ();
 sg13g2_decap_8 FILLER_10_615 ();
 sg13g2_decap_8 FILLER_10_622 ();
 sg13g2_decap_8 FILLER_10_629 ();
 sg13g2_decap_8 FILLER_10_636 ();
 sg13g2_decap_8 FILLER_10_643 ();
 sg13g2_decap_8 FILLER_10_650 ();
 sg13g2_decap_8 FILLER_10_657 ();
 sg13g2_decap_8 FILLER_10_664 ();
 sg13g2_decap_8 FILLER_10_671 ();
 sg13g2_decap_8 FILLER_10_678 ();
 sg13g2_decap_8 FILLER_10_685 ();
 sg13g2_decap_8 FILLER_10_692 ();
 sg13g2_decap_8 FILLER_10_699 ();
 sg13g2_decap_8 FILLER_10_706 ();
 sg13g2_decap_8 FILLER_10_713 ();
 sg13g2_decap_8 FILLER_10_720 ();
 sg13g2_decap_8 FILLER_10_727 ();
 sg13g2_decap_8 FILLER_10_734 ();
 sg13g2_decap_8 FILLER_10_741 ();
 sg13g2_decap_8 FILLER_10_748 ();
 sg13g2_decap_8 FILLER_10_755 ();
 sg13g2_decap_8 FILLER_10_762 ();
 sg13g2_decap_8 FILLER_10_769 ();
 sg13g2_decap_8 FILLER_10_776 ();
 sg13g2_decap_8 FILLER_10_783 ();
 sg13g2_decap_8 FILLER_10_790 ();
 sg13g2_decap_8 FILLER_10_797 ();
 sg13g2_decap_8 FILLER_10_804 ();
 sg13g2_decap_8 FILLER_10_811 ();
 sg13g2_decap_8 FILLER_10_818 ();
 sg13g2_decap_8 FILLER_10_825 ();
 sg13g2_decap_8 FILLER_10_832 ();
 sg13g2_decap_8 FILLER_10_839 ();
 sg13g2_decap_8 FILLER_10_846 ();
 sg13g2_decap_8 FILLER_10_853 ();
 sg13g2_decap_8 FILLER_10_860 ();
 sg13g2_decap_8 FILLER_10_867 ();
 sg13g2_decap_8 FILLER_10_874 ();
 sg13g2_decap_8 FILLER_10_881 ();
 sg13g2_decap_8 FILLER_10_888 ();
 sg13g2_decap_8 FILLER_10_895 ();
 sg13g2_decap_8 FILLER_10_902 ();
 sg13g2_decap_8 FILLER_10_909 ();
 sg13g2_decap_8 FILLER_10_916 ();
 sg13g2_decap_8 FILLER_10_923 ();
 sg13g2_decap_8 FILLER_10_930 ();
 sg13g2_decap_8 FILLER_10_937 ();
 sg13g2_decap_8 FILLER_10_944 ();
 sg13g2_decap_8 FILLER_10_951 ();
 sg13g2_decap_8 FILLER_10_958 ();
 sg13g2_decap_8 FILLER_10_965 ();
 sg13g2_decap_8 FILLER_10_972 ();
 sg13g2_decap_8 FILLER_10_979 ();
 sg13g2_decap_8 FILLER_10_986 ();
 sg13g2_decap_8 FILLER_10_993 ();
 sg13g2_decap_8 FILLER_10_1000 ();
 sg13g2_decap_8 FILLER_10_1007 ();
 sg13g2_decap_8 FILLER_10_1014 ();
 sg13g2_decap_8 FILLER_10_1021 ();
 sg13g2_fill_1 FILLER_10_1028 ();
 sg13g2_decap_8 FILLER_11_4 ();
 sg13g2_decap_4 FILLER_11_11 ();
 sg13g2_fill_2 FILLER_11_15 ();
 sg13g2_decap_8 FILLER_11_44 ();
 sg13g2_decap_8 FILLER_11_51 ();
 sg13g2_decap_4 FILLER_11_58 ();
 sg13g2_fill_2 FILLER_11_62 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_fill_2 FILLER_11_98 ();
 sg13g2_fill_1 FILLER_11_100 ();
 sg13g2_decap_8 FILLER_11_128 ();
 sg13g2_decap_8 FILLER_11_135 ();
 sg13g2_decap_8 FILLER_11_142 ();
 sg13g2_decap_8 FILLER_11_149 ();
 sg13g2_decap_8 FILLER_11_156 ();
 sg13g2_decap_8 FILLER_11_163 ();
 sg13g2_decap_8 FILLER_11_170 ();
 sg13g2_decap_8 FILLER_11_177 ();
 sg13g2_decap_8 FILLER_11_184 ();
 sg13g2_decap_8 FILLER_11_191 ();
 sg13g2_decap_8 FILLER_11_198 ();
 sg13g2_decap_8 FILLER_11_214 ();
 sg13g2_decap_8 FILLER_11_230 ();
 sg13g2_decap_8 FILLER_11_237 ();
 sg13g2_decap_8 FILLER_11_244 ();
 sg13g2_decap_8 FILLER_11_251 ();
 sg13g2_decap_8 FILLER_11_258 ();
 sg13g2_decap_8 FILLER_11_265 ();
 sg13g2_decap_8 FILLER_11_272 ();
 sg13g2_decap_8 FILLER_11_279 ();
 sg13g2_decap_8 FILLER_11_286 ();
 sg13g2_decap_8 FILLER_11_293 ();
 sg13g2_decap_8 FILLER_11_300 ();
 sg13g2_decap_8 FILLER_11_307 ();
 sg13g2_decap_8 FILLER_11_314 ();
 sg13g2_decap_8 FILLER_11_321 ();
 sg13g2_decap_8 FILLER_11_328 ();
 sg13g2_fill_2 FILLER_11_335 ();
 sg13g2_decap_8 FILLER_11_351 ();
 sg13g2_decap_8 FILLER_11_358 ();
 sg13g2_decap_4 FILLER_11_374 ();
 sg13g2_fill_2 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_11_414 ();
 sg13g2_decap_8 FILLER_11_421 ();
 sg13g2_decap_8 FILLER_11_428 ();
 sg13g2_decap_8 FILLER_11_435 ();
 sg13g2_decap_8 FILLER_11_442 ();
 sg13g2_decap_8 FILLER_11_449 ();
 sg13g2_decap_8 FILLER_11_456 ();
 sg13g2_decap_8 FILLER_11_463 ();
 sg13g2_decap_4 FILLER_11_470 ();
 sg13g2_fill_2 FILLER_11_474 ();
 sg13g2_decap_8 FILLER_11_521 ();
 sg13g2_decap_8 FILLER_11_528 ();
 sg13g2_decap_4 FILLER_11_535 ();
 sg13g2_fill_2 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_554 ();
 sg13g2_fill_2 FILLER_11_561 ();
 sg13g2_fill_2 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_596 ();
 sg13g2_decap_8 FILLER_11_603 ();
 sg13g2_decap_8 FILLER_11_641 ();
 sg13g2_decap_8 FILLER_11_648 ();
 sg13g2_decap_8 FILLER_11_655 ();
 sg13g2_decap_8 FILLER_11_662 ();
 sg13g2_decap_8 FILLER_11_669 ();
 sg13g2_decap_8 FILLER_11_676 ();
 sg13g2_decap_8 FILLER_11_683 ();
 sg13g2_decap_8 FILLER_11_690 ();
 sg13g2_decap_8 FILLER_11_697 ();
 sg13g2_decap_8 FILLER_11_704 ();
 sg13g2_decap_8 FILLER_11_711 ();
 sg13g2_decap_8 FILLER_11_718 ();
 sg13g2_decap_8 FILLER_11_725 ();
 sg13g2_decap_8 FILLER_11_732 ();
 sg13g2_decap_8 FILLER_11_739 ();
 sg13g2_decap_8 FILLER_11_746 ();
 sg13g2_decap_8 FILLER_11_753 ();
 sg13g2_decap_8 FILLER_11_760 ();
 sg13g2_decap_8 FILLER_11_767 ();
 sg13g2_decap_8 FILLER_11_774 ();
 sg13g2_decap_8 FILLER_11_781 ();
 sg13g2_decap_8 FILLER_11_788 ();
 sg13g2_decap_8 FILLER_11_795 ();
 sg13g2_decap_8 FILLER_11_802 ();
 sg13g2_decap_8 FILLER_11_809 ();
 sg13g2_decap_8 FILLER_11_816 ();
 sg13g2_decap_8 FILLER_11_823 ();
 sg13g2_decap_8 FILLER_11_830 ();
 sg13g2_decap_8 FILLER_11_837 ();
 sg13g2_decap_8 FILLER_11_844 ();
 sg13g2_decap_8 FILLER_11_851 ();
 sg13g2_decap_8 FILLER_11_858 ();
 sg13g2_decap_8 FILLER_11_865 ();
 sg13g2_decap_8 FILLER_11_872 ();
 sg13g2_decap_8 FILLER_11_879 ();
 sg13g2_decap_8 FILLER_11_886 ();
 sg13g2_decap_8 FILLER_11_893 ();
 sg13g2_decap_8 FILLER_11_900 ();
 sg13g2_decap_8 FILLER_11_907 ();
 sg13g2_decap_8 FILLER_11_914 ();
 sg13g2_decap_8 FILLER_11_921 ();
 sg13g2_decap_8 FILLER_11_928 ();
 sg13g2_decap_8 FILLER_11_935 ();
 sg13g2_decap_8 FILLER_11_942 ();
 sg13g2_decap_8 FILLER_11_949 ();
 sg13g2_decap_8 FILLER_11_956 ();
 sg13g2_decap_8 FILLER_11_963 ();
 sg13g2_decap_8 FILLER_11_970 ();
 sg13g2_decap_8 FILLER_11_977 ();
 sg13g2_decap_8 FILLER_11_984 ();
 sg13g2_decap_8 FILLER_11_991 ();
 sg13g2_decap_8 FILLER_11_998 ();
 sg13g2_decap_8 FILLER_11_1005 ();
 sg13g2_decap_8 FILLER_11_1012 ();
 sg13g2_decap_8 FILLER_11_1019 ();
 sg13g2_fill_2 FILLER_11_1026 ();
 sg13g2_fill_1 FILLER_11_1028 ();
 sg13g2_decap_8 FILLER_12_4 ();
 sg13g2_decap_8 FILLER_12_11 ();
 sg13g2_decap_8 FILLER_12_18 ();
 sg13g2_fill_1 FILLER_12_25 ();
 sg13g2_decap_4 FILLER_12_30 ();
 sg13g2_fill_2 FILLER_12_34 ();
 sg13g2_decap_8 FILLER_12_45 ();
 sg13g2_decap_8 FILLER_12_52 ();
 sg13g2_decap_8 FILLER_12_59 ();
 sg13g2_decap_8 FILLER_12_66 ();
 sg13g2_decap_8 FILLER_12_73 ();
 sg13g2_decap_8 FILLER_12_80 ();
 sg13g2_decap_8 FILLER_12_87 ();
 sg13g2_fill_2 FILLER_12_94 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_4 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_155 ();
 sg13g2_decap_8 FILLER_12_162 ();
 sg13g2_decap_8 FILLER_12_169 ();
 sg13g2_decap_8 FILLER_12_176 ();
 sg13g2_decap_8 FILLER_12_183 ();
 sg13g2_decap_8 FILLER_12_190 ();
 sg13g2_decap_8 FILLER_12_197 ();
 sg13g2_decap_8 FILLER_12_204 ();
 sg13g2_fill_2 FILLER_12_211 ();
 sg13g2_decap_8 FILLER_12_225 ();
 sg13g2_decap_8 FILLER_12_232 ();
 sg13g2_decap_8 FILLER_12_239 ();
 sg13g2_decap_8 FILLER_12_246 ();
 sg13g2_decap_8 FILLER_12_253 ();
 sg13g2_decap_8 FILLER_12_260 ();
 sg13g2_decap_8 FILLER_12_267 ();
 sg13g2_decap_8 FILLER_12_274 ();
 sg13g2_fill_2 FILLER_12_281 ();
 sg13g2_decap_8 FILLER_12_291 ();
 sg13g2_decap_8 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_305 ();
 sg13g2_decap_8 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_decap_8 FILLER_12_326 ();
 sg13g2_decap_8 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_decap_8 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_fill_2 FILLER_12_375 ();
 sg13g2_fill_1 FILLER_12_377 ();
 sg13g2_decap_8 FILLER_12_404 ();
 sg13g2_decap_8 FILLER_12_411 ();
 sg13g2_decap_4 FILLER_12_418 ();
 sg13g2_decap_8 FILLER_12_430 ();
 sg13g2_decap_8 FILLER_12_437 ();
 sg13g2_decap_8 FILLER_12_444 ();
 sg13g2_decap_8 FILLER_12_451 ();
 sg13g2_decap_8 FILLER_12_458 ();
 sg13g2_decap_8 FILLER_12_465 ();
 sg13g2_decap_8 FILLER_12_472 ();
 sg13g2_fill_2 FILLER_12_479 ();
 sg13g2_decap_8 FILLER_12_508 ();
 sg13g2_decap_8 FILLER_12_515 ();
 sg13g2_decap_8 FILLER_12_522 ();
 sg13g2_decap_8 FILLER_12_529 ();
 sg13g2_decap_8 FILLER_12_536 ();
 sg13g2_decap_8 FILLER_12_543 ();
 sg13g2_decap_8 FILLER_12_550 ();
 sg13g2_decap_8 FILLER_12_557 ();
 sg13g2_decap_4 FILLER_12_564 ();
 sg13g2_fill_2 FILLER_12_573 ();
 sg13g2_decap_8 FILLER_12_584 ();
 sg13g2_decap_8 FILLER_12_591 ();
 sg13g2_decap_4 FILLER_12_598 ();
 sg13g2_decap_4 FILLER_12_610 ();
 sg13g2_fill_2 FILLER_12_614 ();
 sg13g2_decap_4 FILLER_12_620 ();
 sg13g2_fill_2 FILLER_12_624 ();
 sg13g2_decap_8 FILLER_12_635 ();
 sg13g2_decap_8 FILLER_12_642 ();
 sg13g2_decap_8 FILLER_12_649 ();
 sg13g2_decap_8 FILLER_12_656 ();
 sg13g2_decap_8 FILLER_12_663 ();
 sg13g2_decap_8 FILLER_12_670 ();
 sg13g2_decap_8 FILLER_12_677 ();
 sg13g2_decap_8 FILLER_12_684 ();
 sg13g2_decap_8 FILLER_12_691 ();
 sg13g2_decap_8 FILLER_12_698 ();
 sg13g2_decap_8 FILLER_12_705 ();
 sg13g2_decap_8 FILLER_12_712 ();
 sg13g2_decap_8 FILLER_12_719 ();
 sg13g2_decap_8 FILLER_12_726 ();
 sg13g2_decap_8 FILLER_12_733 ();
 sg13g2_decap_8 FILLER_12_740 ();
 sg13g2_decap_8 FILLER_12_747 ();
 sg13g2_decap_8 FILLER_12_754 ();
 sg13g2_decap_8 FILLER_12_761 ();
 sg13g2_decap_8 FILLER_12_768 ();
 sg13g2_decap_8 FILLER_12_775 ();
 sg13g2_decap_8 FILLER_12_782 ();
 sg13g2_decap_8 FILLER_12_789 ();
 sg13g2_decap_8 FILLER_12_796 ();
 sg13g2_decap_8 FILLER_12_803 ();
 sg13g2_decap_8 FILLER_12_810 ();
 sg13g2_decap_8 FILLER_12_817 ();
 sg13g2_decap_8 FILLER_12_824 ();
 sg13g2_decap_8 FILLER_12_831 ();
 sg13g2_decap_8 FILLER_12_838 ();
 sg13g2_decap_8 FILLER_12_845 ();
 sg13g2_decap_8 FILLER_12_852 ();
 sg13g2_decap_8 FILLER_12_859 ();
 sg13g2_decap_8 FILLER_12_866 ();
 sg13g2_decap_8 FILLER_12_873 ();
 sg13g2_decap_8 FILLER_12_880 ();
 sg13g2_decap_8 FILLER_12_887 ();
 sg13g2_decap_8 FILLER_12_894 ();
 sg13g2_decap_8 FILLER_12_901 ();
 sg13g2_decap_8 FILLER_12_908 ();
 sg13g2_decap_8 FILLER_12_915 ();
 sg13g2_decap_8 FILLER_12_922 ();
 sg13g2_decap_8 FILLER_12_929 ();
 sg13g2_decap_8 FILLER_12_936 ();
 sg13g2_decap_8 FILLER_12_943 ();
 sg13g2_decap_8 FILLER_12_950 ();
 sg13g2_decap_8 FILLER_12_957 ();
 sg13g2_decap_8 FILLER_12_964 ();
 sg13g2_decap_8 FILLER_12_971 ();
 sg13g2_decap_8 FILLER_12_978 ();
 sg13g2_decap_8 FILLER_12_985 ();
 sg13g2_decap_8 FILLER_12_992 ();
 sg13g2_decap_8 FILLER_12_999 ();
 sg13g2_decap_8 FILLER_12_1006 ();
 sg13g2_decap_8 FILLER_12_1013 ();
 sg13g2_decap_8 FILLER_12_1020 ();
 sg13g2_fill_2 FILLER_12_1027 ();
 sg13g2_decap_8 FILLER_13_4 ();
 sg13g2_decap_8 FILLER_13_11 ();
 sg13g2_decap_8 FILLER_13_18 ();
 sg13g2_decap_8 FILLER_13_25 ();
 sg13g2_decap_8 FILLER_13_32 ();
 sg13g2_decap_8 FILLER_13_39 ();
 sg13g2_decap_8 FILLER_13_46 ();
 sg13g2_decap_8 FILLER_13_53 ();
 sg13g2_decap_8 FILLER_13_60 ();
 sg13g2_decap_8 FILLER_13_67 ();
 sg13g2_decap_8 FILLER_13_74 ();
 sg13g2_decap_8 FILLER_13_81 ();
 sg13g2_fill_2 FILLER_13_88 ();
 sg13g2_decap_8 FILLER_13_103 ();
 sg13g2_decap_8 FILLER_13_110 ();
 sg13g2_decap_8 FILLER_13_117 ();
 sg13g2_decap_4 FILLER_13_124 ();
 sg13g2_decap_8 FILLER_13_137 ();
 sg13g2_decap_8 FILLER_13_144 ();
 sg13g2_fill_2 FILLER_13_151 ();
 sg13g2_fill_1 FILLER_13_153 ();
 sg13g2_decap_8 FILLER_13_190 ();
 sg13g2_decap_8 FILLER_13_197 ();
 sg13g2_decap_4 FILLER_13_204 ();
 sg13g2_fill_1 FILLER_13_208 ();
 sg13g2_decap_8 FILLER_13_222 ();
 sg13g2_decap_8 FILLER_13_229 ();
 sg13g2_decap_8 FILLER_13_236 ();
 sg13g2_decap_4 FILLER_13_243 ();
 sg13g2_fill_1 FILLER_13_247 ();
 sg13g2_decap_8 FILLER_13_275 ();
 sg13g2_decap_8 FILLER_13_282 ();
 sg13g2_decap_8 FILLER_13_289 ();
 sg13g2_decap_8 FILLER_13_296 ();
 sg13g2_decap_8 FILLER_13_303 ();
 sg13g2_decap_4 FILLER_13_310 ();
 sg13g2_decap_4 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_331 ();
 sg13g2_decap_8 FILLER_13_347 ();
 sg13g2_decap_8 FILLER_13_354 ();
 sg13g2_decap_4 FILLER_13_361 ();
 sg13g2_fill_1 FILLER_13_365 ();
 sg13g2_decap_8 FILLER_13_394 ();
 sg13g2_decap_8 FILLER_13_401 ();
 sg13g2_decap_8 FILLER_13_408 ();
 sg13g2_decap_4 FILLER_13_424 ();
 sg13g2_fill_2 FILLER_13_428 ();
 sg13g2_decap_8 FILLER_13_457 ();
 sg13g2_decap_8 FILLER_13_464 ();
 sg13g2_decap_8 FILLER_13_471 ();
 sg13g2_decap_8 FILLER_13_478 ();
 sg13g2_decap_8 FILLER_13_485 ();
 sg13g2_decap_8 FILLER_13_492 ();
 sg13g2_decap_8 FILLER_13_499 ();
 sg13g2_decap_8 FILLER_13_506 ();
 sg13g2_decap_8 FILLER_13_513 ();
 sg13g2_decap_8 FILLER_13_520 ();
 sg13g2_decap_4 FILLER_13_527 ();
 sg13g2_decap_8 FILLER_13_544 ();
 sg13g2_decap_8 FILLER_13_551 ();
 sg13g2_decap_8 FILLER_13_558 ();
 sg13g2_decap_8 FILLER_13_565 ();
 sg13g2_decap_8 FILLER_13_572 ();
 sg13g2_decap_8 FILLER_13_579 ();
 sg13g2_decap_8 FILLER_13_586 ();
 sg13g2_decap_8 FILLER_13_593 ();
 sg13g2_decap_4 FILLER_13_600 ();
 sg13g2_fill_1 FILLER_13_604 ();
 sg13g2_fill_1 FILLER_13_613 ();
 sg13g2_decap_8 FILLER_13_641 ();
 sg13g2_decap_8 FILLER_13_648 ();
 sg13g2_decap_8 FILLER_13_655 ();
 sg13g2_decap_8 FILLER_13_662 ();
 sg13g2_decap_8 FILLER_13_669 ();
 sg13g2_decap_8 FILLER_13_676 ();
 sg13g2_decap_8 FILLER_13_683 ();
 sg13g2_decap_8 FILLER_13_690 ();
 sg13g2_decap_8 FILLER_13_697 ();
 sg13g2_decap_8 FILLER_13_704 ();
 sg13g2_decap_8 FILLER_13_711 ();
 sg13g2_decap_8 FILLER_13_718 ();
 sg13g2_decap_8 FILLER_13_725 ();
 sg13g2_decap_8 FILLER_13_732 ();
 sg13g2_decap_8 FILLER_13_739 ();
 sg13g2_decap_8 FILLER_13_746 ();
 sg13g2_decap_8 FILLER_13_753 ();
 sg13g2_decap_8 FILLER_13_760 ();
 sg13g2_decap_8 FILLER_13_767 ();
 sg13g2_decap_8 FILLER_13_774 ();
 sg13g2_decap_8 FILLER_13_781 ();
 sg13g2_decap_8 FILLER_13_788 ();
 sg13g2_decap_8 FILLER_13_795 ();
 sg13g2_decap_8 FILLER_13_802 ();
 sg13g2_decap_8 FILLER_13_809 ();
 sg13g2_decap_8 FILLER_13_816 ();
 sg13g2_decap_8 FILLER_13_823 ();
 sg13g2_decap_8 FILLER_13_830 ();
 sg13g2_decap_8 FILLER_13_837 ();
 sg13g2_decap_8 FILLER_13_844 ();
 sg13g2_decap_8 FILLER_13_851 ();
 sg13g2_decap_8 FILLER_13_858 ();
 sg13g2_decap_8 FILLER_13_865 ();
 sg13g2_decap_8 FILLER_13_872 ();
 sg13g2_decap_8 FILLER_13_879 ();
 sg13g2_decap_8 FILLER_13_886 ();
 sg13g2_decap_8 FILLER_13_893 ();
 sg13g2_decap_8 FILLER_13_900 ();
 sg13g2_decap_8 FILLER_13_907 ();
 sg13g2_decap_8 FILLER_13_914 ();
 sg13g2_decap_8 FILLER_13_921 ();
 sg13g2_decap_8 FILLER_13_928 ();
 sg13g2_decap_8 FILLER_13_935 ();
 sg13g2_decap_8 FILLER_13_942 ();
 sg13g2_decap_8 FILLER_13_949 ();
 sg13g2_decap_8 FILLER_13_956 ();
 sg13g2_decap_8 FILLER_13_963 ();
 sg13g2_decap_8 FILLER_13_970 ();
 sg13g2_decap_8 FILLER_13_977 ();
 sg13g2_decap_8 FILLER_13_984 ();
 sg13g2_decap_8 FILLER_13_991 ();
 sg13g2_decap_8 FILLER_13_998 ();
 sg13g2_decap_8 FILLER_13_1005 ();
 sg13g2_decap_8 FILLER_13_1012 ();
 sg13g2_decap_8 FILLER_13_1019 ();
 sg13g2_fill_2 FILLER_13_1026 ();
 sg13g2_fill_1 FILLER_13_1028 ();
 sg13g2_decap_8 FILLER_14_4 ();
 sg13g2_decap_8 FILLER_14_11 ();
 sg13g2_decap_8 FILLER_14_18 ();
 sg13g2_decap_8 FILLER_14_25 ();
 sg13g2_decap_8 FILLER_14_32 ();
 sg13g2_decap_8 FILLER_14_39 ();
 sg13g2_decap_8 FILLER_14_46 ();
 sg13g2_decap_8 FILLER_14_53 ();
 sg13g2_decap_8 FILLER_14_60 ();
 sg13g2_decap_8 FILLER_14_67 ();
 sg13g2_decap_8 FILLER_14_74 ();
 sg13g2_decap_8 FILLER_14_81 ();
 sg13g2_decap_8 FILLER_14_88 ();
 sg13g2_decap_8 FILLER_14_95 ();
 sg13g2_decap_8 FILLER_14_102 ();
 sg13g2_decap_8 FILLER_14_109 ();
 sg13g2_decap_8 FILLER_14_116 ();
 sg13g2_decap_8 FILLER_14_123 ();
 sg13g2_decap_8 FILLER_14_130 ();
 sg13g2_decap_8 FILLER_14_137 ();
 sg13g2_decap_8 FILLER_14_144 ();
 sg13g2_decap_8 FILLER_14_151 ();
 sg13g2_decap_8 FILLER_14_158 ();
 sg13g2_decap_8 FILLER_14_165 ();
 sg13g2_decap_8 FILLER_14_172 ();
 sg13g2_fill_2 FILLER_14_179 ();
 sg13g2_fill_1 FILLER_14_181 ();
 sg13g2_decap_8 FILLER_14_195 ();
 sg13g2_decap_8 FILLER_14_202 ();
 sg13g2_decap_8 FILLER_14_209 ();
 sg13g2_decap_8 FILLER_14_216 ();
 sg13g2_decap_8 FILLER_14_223 ();
 sg13g2_decap_4 FILLER_14_230 ();
 sg13g2_fill_2 FILLER_14_242 ();
 sg13g2_fill_1 FILLER_14_244 ();
 sg13g2_decap_8 FILLER_14_254 ();
 sg13g2_decap_8 FILLER_14_261 ();
 sg13g2_decap_8 FILLER_14_268 ();
 sg13g2_decap_8 FILLER_14_275 ();
 sg13g2_decap_8 FILLER_14_282 ();
 sg13g2_decap_8 FILLER_14_289 ();
 sg13g2_decap_8 FILLER_14_296 ();
 sg13g2_fill_1 FILLER_14_303 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_4 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_447 ();
 sg13g2_decap_8 FILLER_14_454 ();
 sg13g2_decap_8 FILLER_14_461 ();
 sg13g2_decap_8 FILLER_14_468 ();
 sg13g2_decap_4 FILLER_14_475 ();
 sg13g2_decap_8 FILLER_14_488 ();
 sg13g2_decap_4 FILLER_14_495 ();
 sg13g2_fill_2 FILLER_14_499 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_4 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_563 ();
 sg13g2_decap_8 FILLER_14_570 ();
 sg13g2_decap_8 FILLER_14_577 ();
 sg13g2_decap_8 FILLER_14_584 ();
 sg13g2_decap_8 FILLER_14_591 ();
 sg13g2_decap_8 FILLER_14_598 ();
 sg13g2_decap_8 FILLER_14_605 ();
 sg13g2_decap_8 FILLER_14_612 ();
 sg13g2_decap_8 FILLER_14_619 ();
 sg13g2_decap_4 FILLER_14_626 ();
 sg13g2_decap_8 FILLER_14_639 ();
 sg13g2_decap_8 FILLER_14_646 ();
 sg13g2_decap_8 FILLER_14_653 ();
 sg13g2_decap_8 FILLER_14_660 ();
 sg13g2_decap_8 FILLER_14_667 ();
 sg13g2_decap_8 FILLER_14_674 ();
 sg13g2_decap_8 FILLER_14_681 ();
 sg13g2_decap_8 FILLER_14_688 ();
 sg13g2_decap_8 FILLER_14_695 ();
 sg13g2_decap_8 FILLER_14_702 ();
 sg13g2_decap_8 FILLER_14_709 ();
 sg13g2_decap_8 FILLER_14_716 ();
 sg13g2_decap_8 FILLER_14_723 ();
 sg13g2_decap_8 FILLER_14_730 ();
 sg13g2_decap_8 FILLER_14_737 ();
 sg13g2_decap_8 FILLER_14_744 ();
 sg13g2_decap_8 FILLER_14_751 ();
 sg13g2_decap_8 FILLER_14_758 ();
 sg13g2_decap_8 FILLER_14_765 ();
 sg13g2_decap_8 FILLER_14_772 ();
 sg13g2_decap_8 FILLER_14_779 ();
 sg13g2_decap_8 FILLER_14_786 ();
 sg13g2_decap_8 FILLER_14_793 ();
 sg13g2_decap_8 FILLER_14_800 ();
 sg13g2_decap_8 FILLER_14_807 ();
 sg13g2_decap_8 FILLER_14_814 ();
 sg13g2_decap_8 FILLER_14_821 ();
 sg13g2_decap_8 FILLER_14_828 ();
 sg13g2_decap_8 FILLER_14_835 ();
 sg13g2_decap_8 FILLER_14_842 ();
 sg13g2_decap_8 FILLER_14_849 ();
 sg13g2_decap_8 FILLER_14_856 ();
 sg13g2_decap_8 FILLER_14_863 ();
 sg13g2_decap_8 FILLER_14_870 ();
 sg13g2_decap_8 FILLER_14_877 ();
 sg13g2_decap_8 FILLER_14_884 ();
 sg13g2_decap_8 FILLER_14_891 ();
 sg13g2_decap_8 FILLER_14_898 ();
 sg13g2_decap_8 FILLER_14_905 ();
 sg13g2_decap_8 FILLER_14_912 ();
 sg13g2_decap_8 FILLER_14_919 ();
 sg13g2_decap_8 FILLER_14_926 ();
 sg13g2_decap_8 FILLER_14_933 ();
 sg13g2_decap_8 FILLER_14_940 ();
 sg13g2_decap_8 FILLER_14_947 ();
 sg13g2_decap_8 FILLER_14_954 ();
 sg13g2_decap_8 FILLER_14_961 ();
 sg13g2_decap_8 FILLER_14_968 ();
 sg13g2_decap_8 FILLER_14_975 ();
 sg13g2_decap_8 FILLER_14_982 ();
 sg13g2_decap_8 FILLER_14_989 ();
 sg13g2_decap_8 FILLER_14_996 ();
 sg13g2_decap_8 FILLER_14_1003 ();
 sg13g2_decap_8 FILLER_14_1010 ();
 sg13g2_decap_8 FILLER_14_1017 ();
 sg13g2_decap_4 FILLER_14_1024 ();
 sg13g2_fill_1 FILLER_14_1028 ();
 sg13g2_decap_8 FILLER_15_4 ();
 sg13g2_decap_8 FILLER_15_11 ();
 sg13g2_decap_8 FILLER_15_18 ();
 sg13g2_decap_8 FILLER_15_25 ();
 sg13g2_decap_8 FILLER_15_32 ();
 sg13g2_decap_8 FILLER_15_39 ();
 sg13g2_decap_8 FILLER_15_46 ();
 sg13g2_decap_8 FILLER_15_53 ();
 sg13g2_decap_8 FILLER_15_60 ();
 sg13g2_decap_8 FILLER_15_67 ();
 sg13g2_decap_8 FILLER_15_74 ();
 sg13g2_fill_1 FILLER_15_81 ();
 sg13g2_decap_8 FILLER_15_95 ();
 sg13g2_decap_8 FILLER_15_102 ();
 sg13g2_decap_8 FILLER_15_109 ();
 sg13g2_decap_8 FILLER_15_116 ();
 sg13g2_decap_8 FILLER_15_123 ();
 sg13g2_decap_8 FILLER_15_130 ();
 sg13g2_decap_8 FILLER_15_137 ();
 sg13g2_decap_8 FILLER_15_144 ();
 sg13g2_decap_8 FILLER_15_151 ();
 sg13g2_decap_8 FILLER_15_158 ();
 sg13g2_decap_8 FILLER_15_165 ();
 sg13g2_decap_8 FILLER_15_172 ();
 sg13g2_decap_8 FILLER_15_179 ();
 sg13g2_decap_8 FILLER_15_199 ();
 sg13g2_decap_8 FILLER_15_206 ();
 sg13g2_fill_1 FILLER_15_213 ();
 sg13g2_fill_2 FILLER_15_227 ();
 sg13g2_fill_1 FILLER_15_229 ();
 sg13g2_decap_8 FILLER_15_247 ();
 sg13g2_decap_8 FILLER_15_254 ();
 sg13g2_decap_8 FILLER_15_261 ();
 sg13g2_decap_8 FILLER_15_268 ();
 sg13g2_decap_8 FILLER_15_275 ();
 sg13g2_decap_4 FILLER_15_282 ();
 sg13g2_fill_2 FILLER_15_286 ();
 sg13g2_decap_8 FILLER_15_328 ();
 sg13g2_decap_8 FILLER_15_335 ();
 sg13g2_decap_8 FILLER_15_342 ();
 sg13g2_decap_8 FILLER_15_349 ();
 sg13g2_fill_1 FILLER_15_356 ();
 sg13g2_decap_8 FILLER_15_370 ();
 sg13g2_decap_8 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_8 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_15_412 ();
 sg13g2_fill_2 FILLER_15_419 ();
 sg13g2_fill_1 FILLER_15_421 ();
 sg13g2_fill_2 FILLER_15_426 ();
 sg13g2_decap_8 FILLER_15_441 ();
 sg13g2_decap_8 FILLER_15_448 ();
 sg13g2_decap_8 FILLER_15_455 ();
 sg13g2_decap_8 FILLER_15_462 ();
 sg13g2_decap_8 FILLER_15_469 ();
 sg13g2_decap_8 FILLER_15_476 ();
 sg13g2_decap_8 FILLER_15_483 ();
 sg13g2_decap_8 FILLER_15_490 ();
 sg13g2_decap_8 FILLER_15_497 ();
 sg13g2_fill_2 FILLER_15_504 ();
 sg13g2_fill_1 FILLER_15_506 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_526 ();
 sg13g2_decap_8 FILLER_15_533 ();
 sg13g2_decap_4 FILLER_15_540 ();
 sg13g2_fill_2 FILLER_15_544 ();
 sg13g2_fill_1 FILLER_15_559 ();
 sg13g2_decap_8 FILLER_15_587 ();
 sg13g2_decap_8 FILLER_15_594 ();
 sg13g2_decap_8 FILLER_15_601 ();
 sg13g2_decap_8 FILLER_15_608 ();
 sg13g2_decap_8 FILLER_15_615 ();
 sg13g2_decap_8 FILLER_15_622 ();
 sg13g2_decap_8 FILLER_15_629 ();
 sg13g2_decap_8 FILLER_15_636 ();
 sg13g2_decap_8 FILLER_15_643 ();
 sg13g2_decap_8 FILLER_15_650 ();
 sg13g2_decap_8 FILLER_15_657 ();
 sg13g2_decap_8 FILLER_15_664 ();
 sg13g2_decap_8 FILLER_15_671 ();
 sg13g2_decap_8 FILLER_15_678 ();
 sg13g2_decap_8 FILLER_15_685 ();
 sg13g2_decap_8 FILLER_15_692 ();
 sg13g2_decap_8 FILLER_15_699 ();
 sg13g2_decap_8 FILLER_15_706 ();
 sg13g2_decap_8 FILLER_15_713 ();
 sg13g2_decap_8 FILLER_15_720 ();
 sg13g2_decap_8 FILLER_15_727 ();
 sg13g2_decap_8 FILLER_15_734 ();
 sg13g2_decap_8 FILLER_15_741 ();
 sg13g2_decap_8 FILLER_15_748 ();
 sg13g2_decap_8 FILLER_15_755 ();
 sg13g2_decap_8 FILLER_15_762 ();
 sg13g2_decap_8 FILLER_15_769 ();
 sg13g2_decap_8 FILLER_15_776 ();
 sg13g2_decap_8 FILLER_15_783 ();
 sg13g2_decap_8 FILLER_15_790 ();
 sg13g2_decap_8 FILLER_15_797 ();
 sg13g2_decap_8 FILLER_15_804 ();
 sg13g2_decap_8 FILLER_15_811 ();
 sg13g2_decap_8 FILLER_15_818 ();
 sg13g2_decap_8 FILLER_15_825 ();
 sg13g2_decap_8 FILLER_15_832 ();
 sg13g2_decap_8 FILLER_15_839 ();
 sg13g2_decap_8 FILLER_15_846 ();
 sg13g2_decap_8 FILLER_15_853 ();
 sg13g2_decap_8 FILLER_15_860 ();
 sg13g2_decap_8 FILLER_15_867 ();
 sg13g2_decap_8 FILLER_15_874 ();
 sg13g2_decap_8 FILLER_15_881 ();
 sg13g2_decap_8 FILLER_15_888 ();
 sg13g2_decap_8 FILLER_15_895 ();
 sg13g2_decap_8 FILLER_15_902 ();
 sg13g2_decap_8 FILLER_15_909 ();
 sg13g2_decap_8 FILLER_15_916 ();
 sg13g2_decap_8 FILLER_15_923 ();
 sg13g2_decap_8 FILLER_15_930 ();
 sg13g2_decap_8 FILLER_15_937 ();
 sg13g2_decap_8 FILLER_15_944 ();
 sg13g2_decap_8 FILLER_15_951 ();
 sg13g2_decap_8 FILLER_15_958 ();
 sg13g2_decap_8 FILLER_15_965 ();
 sg13g2_decap_8 FILLER_15_972 ();
 sg13g2_decap_8 FILLER_15_979 ();
 sg13g2_decap_8 FILLER_15_986 ();
 sg13g2_decap_8 FILLER_15_993 ();
 sg13g2_decap_8 FILLER_15_1000 ();
 sg13g2_decap_8 FILLER_15_1007 ();
 sg13g2_decap_8 FILLER_15_1014 ();
 sg13g2_decap_8 FILLER_15_1021 ();
 sg13g2_fill_1 FILLER_15_1028 ();
 sg13g2_decap_8 FILLER_16_4 ();
 sg13g2_decap_8 FILLER_16_11 ();
 sg13g2_decap_8 FILLER_16_18 ();
 sg13g2_decap_8 FILLER_16_25 ();
 sg13g2_fill_2 FILLER_16_32 ();
 sg13g2_fill_1 FILLER_16_34 ();
 sg13g2_decap_8 FILLER_16_62 ();
 sg13g2_decap_8 FILLER_16_69 ();
 sg13g2_decap_8 FILLER_16_76 ();
 sg13g2_decap_4 FILLER_16_83 ();
 sg13g2_fill_1 FILLER_16_87 ();
 sg13g2_decap_8 FILLER_16_123 ();
 sg13g2_decap_8 FILLER_16_130 ();
 sg13g2_decap_8 FILLER_16_137 ();
 sg13g2_decap_8 FILLER_16_144 ();
 sg13g2_decap_8 FILLER_16_151 ();
 sg13g2_decap_8 FILLER_16_158 ();
 sg13g2_decap_4 FILLER_16_165 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_fill_2 FILLER_16_231 ();
 sg13g2_fill_1 FILLER_16_237 ();
 sg13g2_decap_8 FILLER_16_247 ();
 sg13g2_decap_8 FILLER_16_254 ();
 sg13g2_decap_4 FILLER_16_261 ();
 sg13g2_decap_8 FILLER_16_274 ();
 sg13g2_decap_8 FILLER_16_281 ();
 sg13g2_decap_8 FILLER_16_288 ();
 sg13g2_decap_8 FILLER_16_295 ();
 sg13g2_decap_8 FILLER_16_302 ();
 sg13g2_decap_8 FILLER_16_309 ();
 sg13g2_decap_8 FILLER_16_316 ();
 sg13g2_decap_8 FILLER_16_323 ();
 sg13g2_decap_8 FILLER_16_330 ();
 sg13g2_decap_8 FILLER_16_337 ();
 sg13g2_decap_8 FILLER_16_344 ();
 sg13g2_decap_8 FILLER_16_351 ();
 sg13g2_decap_8 FILLER_16_358 ();
 sg13g2_decap_8 FILLER_16_365 ();
 sg13g2_decap_8 FILLER_16_372 ();
 sg13g2_decap_8 FILLER_16_379 ();
 sg13g2_decap_8 FILLER_16_386 ();
 sg13g2_fill_1 FILLER_16_393 ();
 sg13g2_decap_4 FILLER_16_421 ();
 sg13g2_fill_2 FILLER_16_425 ();
 sg13g2_decap_8 FILLER_16_436 ();
 sg13g2_decap_8 FILLER_16_443 ();
 sg13g2_decap_8 FILLER_16_450 ();
 sg13g2_decap_8 FILLER_16_457 ();
 sg13g2_decap_8 FILLER_16_464 ();
 sg13g2_decap_8 FILLER_16_471 ();
 sg13g2_decap_8 FILLER_16_478 ();
 sg13g2_decap_8 FILLER_16_485 ();
 sg13g2_decap_8 FILLER_16_492 ();
 sg13g2_fill_1 FILLER_16_499 ();
 sg13g2_decap_8 FILLER_16_517 ();
 sg13g2_decap_8 FILLER_16_524 ();
 sg13g2_decap_8 FILLER_16_531 ();
 sg13g2_decap_8 FILLER_16_538 ();
 sg13g2_decap_8 FILLER_16_545 ();
 sg13g2_decap_4 FILLER_16_579 ();
 sg13g2_decap_8 FILLER_16_586 ();
 sg13g2_decap_8 FILLER_16_593 ();
 sg13g2_decap_8 FILLER_16_600 ();
 sg13g2_decap_8 FILLER_16_607 ();
 sg13g2_decap_8 FILLER_16_614 ();
 sg13g2_decap_8 FILLER_16_621 ();
 sg13g2_decap_8 FILLER_16_628 ();
 sg13g2_decap_8 FILLER_16_635 ();
 sg13g2_decap_8 FILLER_16_642 ();
 sg13g2_decap_8 FILLER_16_649 ();
 sg13g2_decap_8 FILLER_16_656 ();
 sg13g2_decap_8 FILLER_16_663 ();
 sg13g2_decap_8 FILLER_16_670 ();
 sg13g2_decap_8 FILLER_16_677 ();
 sg13g2_decap_8 FILLER_16_684 ();
 sg13g2_decap_8 FILLER_16_691 ();
 sg13g2_decap_8 FILLER_16_698 ();
 sg13g2_decap_8 FILLER_16_705 ();
 sg13g2_decap_8 FILLER_16_712 ();
 sg13g2_decap_8 FILLER_16_719 ();
 sg13g2_decap_8 FILLER_16_726 ();
 sg13g2_decap_8 FILLER_16_733 ();
 sg13g2_decap_8 FILLER_16_740 ();
 sg13g2_decap_8 FILLER_16_747 ();
 sg13g2_decap_8 FILLER_16_754 ();
 sg13g2_decap_8 FILLER_16_761 ();
 sg13g2_decap_8 FILLER_16_768 ();
 sg13g2_decap_8 FILLER_16_775 ();
 sg13g2_decap_8 FILLER_16_782 ();
 sg13g2_decap_8 FILLER_16_789 ();
 sg13g2_decap_8 FILLER_16_796 ();
 sg13g2_decap_8 FILLER_16_803 ();
 sg13g2_decap_8 FILLER_16_810 ();
 sg13g2_decap_8 FILLER_16_817 ();
 sg13g2_decap_8 FILLER_16_824 ();
 sg13g2_decap_8 FILLER_16_831 ();
 sg13g2_decap_8 FILLER_16_838 ();
 sg13g2_decap_8 FILLER_16_845 ();
 sg13g2_decap_8 FILLER_16_852 ();
 sg13g2_decap_8 FILLER_16_859 ();
 sg13g2_decap_8 FILLER_16_866 ();
 sg13g2_decap_8 FILLER_16_873 ();
 sg13g2_decap_8 FILLER_16_880 ();
 sg13g2_decap_8 FILLER_16_887 ();
 sg13g2_decap_8 FILLER_16_894 ();
 sg13g2_decap_8 FILLER_16_901 ();
 sg13g2_decap_8 FILLER_16_908 ();
 sg13g2_decap_8 FILLER_16_915 ();
 sg13g2_decap_8 FILLER_16_922 ();
 sg13g2_decap_8 FILLER_16_929 ();
 sg13g2_decap_8 FILLER_16_936 ();
 sg13g2_decap_8 FILLER_16_943 ();
 sg13g2_decap_8 FILLER_16_950 ();
 sg13g2_decap_8 FILLER_16_957 ();
 sg13g2_decap_8 FILLER_16_964 ();
 sg13g2_decap_8 FILLER_16_971 ();
 sg13g2_decap_8 FILLER_16_978 ();
 sg13g2_decap_8 FILLER_16_985 ();
 sg13g2_decap_8 FILLER_16_992 ();
 sg13g2_decap_8 FILLER_16_999 ();
 sg13g2_decap_8 FILLER_16_1006 ();
 sg13g2_decap_8 FILLER_16_1013 ();
 sg13g2_decap_8 FILLER_16_1020 ();
 sg13g2_fill_2 FILLER_16_1027 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_fill_2 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_23 ();
 sg13g2_fill_2 FILLER_17_55 ();
 sg13g2_fill_1 FILLER_17_57 ();
 sg13g2_decap_8 FILLER_17_71 ();
 sg13g2_decap_8 FILLER_17_78 ();
 sg13g2_fill_2 FILLER_17_85 ();
 sg13g2_fill_1 FILLER_17_87 ();
 sg13g2_decap_8 FILLER_17_128 ();
 sg13g2_decap_8 FILLER_17_135 ();
 sg13g2_decap_8 FILLER_17_142 ();
 sg13g2_decap_8 FILLER_17_149 ();
 sg13g2_decap_8 FILLER_17_156 ();
 sg13g2_decap_8 FILLER_17_163 ();
 sg13g2_decap_4 FILLER_17_170 ();
 sg13g2_decap_8 FILLER_17_178 ();
 sg13g2_fill_1 FILLER_17_185 ();
 sg13g2_decap_8 FILLER_17_195 ();
 sg13g2_decap_8 FILLER_17_202 ();
 sg13g2_decap_8 FILLER_17_209 ();
 sg13g2_decap_8 FILLER_17_216 ();
 sg13g2_decap_8 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_230 ();
 sg13g2_decap_8 FILLER_17_237 ();
 sg13g2_decap_8 FILLER_17_244 ();
 sg13g2_decap_8 FILLER_17_251 ();
 sg13g2_decap_8 FILLER_17_258 ();
 sg13g2_decap_8 FILLER_17_265 ();
 sg13g2_fill_1 FILLER_17_272 ();
 sg13g2_decap_8 FILLER_17_286 ();
 sg13g2_decap_8 FILLER_17_293 ();
 sg13g2_decap_8 FILLER_17_300 ();
 sg13g2_decap_8 FILLER_17_307 ();
 sg13g2_decap_8 FILLER_17_314 ();
 sg13g2_decap_8 FILLER_17_321 ();
 sg13g2_decap_8 FILLER_17_328 ();
 sg13g2_decap_8 FILLER_17_335 ();
 sg13g2_decap_8 FILLER_17_342 ();
 sg13g2_decap_8 FILLER_17_349 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_decap_8 FILLER_17_363 ();
 sg13g2_decap_8 FILLER_17_370 ();
 sg13g2_decap_8 FILLER_17_377 ();
 sg13g2_decap_8 FILLER_17_384 ();
 sg13g2_fill_2 FILLER_17_391 ();
 sg13g2_fill_1 FILLER_17_393 ();
 sg13g2_decap_8 FILLER_17_403 ();
 sg13g2_decap_8 FILLER_17_410 ();
 sg13g2_decap_8 FILLER_17_417 ();
 sg13g2_decap_8 FILLER_17_424 ();
 sg13g2_decap_8 FILLER_17_431 ();
 sg13g2_decap_8 FILLER_17_438 ();
 sg13g2_fill_1 FILLER_17_445 ();
 sg13g2_decap_4 FILLER_17_481 ();
 sg13g2_fill_1 FILLER_17_485 ();
 sg13g2_decap_8 FILLER_17_522 ();
 sg13g2_decap_8 FILLER_17_529 ();
 sg13g2_decap_8 FILLER_17_536 ();
 sg13g2_decap_8 FILLER_17_543 ();
 sg13g2_decap_8 FILLER_17_550 ();
 sg13g2_decap_8 FILLER_17_557 ();
 sg13g2_fill_2 FILLER_17_564 ();
 sg13g2_fill_1 FILLER_17_566 ();
 sg13g2_fill_2 FILLER_17_575 ();
 sg13g2_decap_8 FILLER_17_599 ();
 sg13g2_fill_2 FILLER_17_606 ();
 sg13g2_decap_8 FILLER_17_635 ();
 sg13g2_decap_8 FILLER_17_642 ();
 sg13g2_decap_8 FILLER_17_649 ();
 sg13g2_decap_8 FILLER_17_656 ();
 sg13g2_decap_8 FILLER_17_663 ();
 sg13g2_decap_8 FILLER_17_670 ();
 sg13g2_decap_8 FILLER_17_677 ();
 sg13g2_decap_8 FILLER_17_684 ();
 sg13g2_decap_8 FILLER_17_691 ();
 sg13g2_decap_8 FILLER_17_698 ();
 sg13g2_decap_8 FILLER_17_705 ();
 sg13g2_decap_8 FILLER_17_712 ();
 sg13g2_decap_8 FILLER_17_719 ();
 sg13g2_decap_8 FILLER_17_726 ();
 sg13g2_decap_8 FILLER_17_733 ();
 sg13g2_decap_8 FILLER_17_740 ();
 sg13g2_decap_8 FILLER_17_747 ();
 sg13g2_decap_8 FILLER_17_754 ();
 sg13g2_decap_8 FILLER_17_761 ();
 sg13g2_decap_8 FILLER_17_768 ();
 sg13g2_decap_8 FILLER_17_775 ();
 sg13g2_decap_8 FILLER_17_782 ();
 sg13g2_decap_8 FILLER_17_789 ();
 sg13g2_decap_8 FILLER_17_796 ();
 sg13g2_decap_8 FILLER_17_803 ();
 sg13g2_decap_8 FILLER_17_810 ();
 sg13g2_decap_8 FILLER_17_817 ();
 sg13g2_decap_8 FILLER_17_824 ();
 sg13g2_decap_8 FILLER_17_831 ();
 sg13g2_decap_8 FILLER_17_838 ();
 sg13g2_decap_8 FILLER_17_845 ();
 sg13g2_decap_8 FILLER_17_852 ();
 sg13g2_decap_8 FILLER_17_859 ();
 sg13g2_decap_8 FILLER_17_866 ();
 sg13g2_decap_8 FILLER_17_873 ();
 sg13g2_decap_8 FILLER_17_880 ();
 sg13g2_decap_8 FILLER_17_887 ();
 sg13g2_decap_8 FILLER_17_894 ();
 sg13g2_decap_8 FILLER_17_901 ();
 sg13g2_decap_8 FILLER_17_908 ();
 sg13g2_decap_8 FILLER_17_915 ();
 sg13g2_decap_8 FILLER_17_922 ();
 sg13g2_decap_8 FILLER_17_929 ();
 sg13g2_decap_8 FILLER_17_936 ();
 sg13g2_decap_8 FILLER_17_943 ();
 sg13g2_decap_8 FILLER_17_950 ();
 sg13g2_decap_8 FILLER_17_957 ();
 sg13g2_decap_8 FILLER_17_964 ();
 sg13g2_decap_8 FILLER_17_971 ();
 sg13g2_decap_8 FILLER_17_978 ();
 sg13g2_decap_8 FILLER_17_985 ();
 sg13g2_decap_8 FILLER_17_992 ();
 sg13g2_decap_8 FILLER_17_999 ();
 sg13g2_decap_8 FILLER_17_1006 ();
 sg13g2_decap_8 FILLER_17_1013 ();
 sg13g2_decap_8 FILLER_17_1020 ();
 sg13g2_fill_2 FILLER_17_1027 ();
 sg13g2_decap_8 FILLER_18_4 ();
 sg13g2_decap_8 FILLER_18_11 ();
 sg13g2_decap_8 FILLER_18_18 ();
 sg13g2_decap_8 FILLER_18_25 ();
 sg13g2_fill_1 FILLER_18_32 ();
 sg13g2_fill_2 FILLER_18_37 ();
 sg13g2_fill_1 FILLER_18_39 ();
 sg13g2_decap_8 FILLER_18_62 ();
 sg13g2_decap_8 FILLER_18_69 ();
 sg13g2_fill_1 FILLER_18_76 ();
 sg13g2_decap_8 FILLER_18_90 ();
 sg13g2_decap_8 FILLER_18_97 ();
 sg13g2_decap_8 FILLER_18_113 ();
 sg13g2_decap_8 FILLER_18_120 ();
 sg13g2_decap_8 FILLER_18_127 ();
 sg13g2_decap_8 FILLER_18_134 ();
 sg13g2_decap_8 FILLER_18_141 ();
 sg13g2_decap_8 FILLER_18_148 ();
 sg13g2_decap_8 FILLER_18_155 ();
 sg13g2_decap_8 FILLER_18_162 ();
 sg13g2_decap_8 FILLER_18_169 ();
 sg13g2_decap_8 FILLER_18_176 ();
 sg13g2_decap_8 FILLER_18_183 ();
 sg13g2_decap_8 FILLER_18_190 ();
 sg13g2_decap_8 FILLER_18_197 ();
 sg13g2_decap_8 FILLER_18_204 ();
 sg13g2_decap_4 FILLER_18_211 ();
 sg13g2_decap_8 FILLER_18_242 ();
 sg13g2_decap_8 FILLER_18_249 ();
 sg13g2_decap_8 FILLER_18_256 ();
 sg13g2_decap_8 FILLER_18_263 ();
 sg13g2_decap_8 FILLER_18_270 ();
 sg13g2_decap_8 FILLER_18_277 ();
 sg13g2_decap_8 FILLER_18_284 ();
 sg13g2_decap_8 FILLER_18_291 ();
 sg13g2_decap_8 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_305 ();
 sg13g2_decap_8 FILLER_18_312 ();
 sg13g2_decap_8 FILLER_18_319 ();
 sg13g2_decap_8 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_333 ();
 sg13g2_decap_4 FILLER_18_340 ();
 sg13g2_fill_1 FILLER_18_352 ();
 sg13g2_fill_2 FILLER_18_389 ();
 sg13g2_fill_1 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_400 ();
 sg13g2_decap_8 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_18_414 ();
 sg13g2_decap_8 FILLER_18_421 ();
 sg13g2_decap_8 FILLER_18_428 ();
 sg13g2_decap_8 FILLER_18_435 ();
 sg13g2_decap_8 FILLER_18_442 ();
 sg13g2_decap_8 FILLER_18_449 ();
 sg13g2_decap_8 FILLER_18_456 ();
 sg13g2_decap_8 FILLER_18_463 ();
 sg13g2_decap_8 FILLER_18_470 ();
 sg13g2_decap_8 FILLER_18_477 ();
 sg13g2_decap_8 FILLER_18_484 ();
 sg13g2_decap_8 FILLER_18_491 ();
 sg13g2_decap_8 FILLER_18_498 ();
 sg13g2_decap_8 FILLER_18_505 ();
 sg13g2_decap_8 FILLER_18_512 ();
 sg13g2_decap_8 FILLER_18_519 ();
 sg13g2_fill_1 FILLER_18_526 ();
 sg13g2_decap_4 FILLER_18_540 ();
 sg13g2_fill_1 FILLER_18_544 ();
 sg13g2_decap_8 FILLER_18_554 ();
 sg13g2_decap_8 FILLER_18_561 ();
 sg13g2_fill_2 FILLER_18_568 ();
 sg13g2_decap_8 FILLER_18_591 ();
 sg13g2_decap_8 FILLER_18_598 ();
 sg13g2_decap_4 FILLER_18_605 ();
 sg13g2_fill_1 FILLER_18_609 ();
 sg13g2_decap_8 FILLER_18_618 ();
 sg13g2_decap_8 FILLER_18_625 ();
 sg13g2_decap_8 FILLER_18_632 ();
 sg13g2_decap_8 FILLER_18_639 ();
 sg13g2_decap_8 FILLER_18_646 ();
 sg13g2_decap_8 FILLER_18_653 ();
 sg13g2_decap_8 FILLER_18_660 ();
 sg13g2_decap_8 FILLER_18_667 ();
 sg13g2_decap_8 FILLER_18_674 ();
 sg13g2_decap_8 FILLER_18_681 ();
 sg13g2_decap_8 FILLER_18_688 ();
 sg13g2_decap_8 FILLER_18_695 ();
 sg13g2_decap_8 FILLER_18_702 ();
 sg13g2_decap_8 FILLER_18_709 ();
 sg13g2_decap_8 FILLER_18_716 ();
 sg13g2_decap_8 FILLER_18_723 ();
 sg13g2_decap_8 FILLER_18_730 ();
 sg13g2_decap_8 FILLER_18_737 ();
 sg13g2_decap_8 FILLER_18_744 ();
 sg13g2_decap_8 FILLER_18_751 ();
 sg13g2_decap_8 FILLER_18_758 ();
 sg13g2_decap_8 FILLER_18_765 ();
 sg13g2_decap_8 FILLER_18_772 ();
 sg13g2_decap_8 FILLER_18_779 ();
 sg13g2_decap_8 FILLER_18_786 ();
 sg13g2_decap_8 FILLER_18_793 ();
 sg13g2_decap_8 FILLER_18_800 ();
 sg13g2_decap_8 FILLER_18_807 ();
 sg13g2_decap_8 FILLER_18_814 ();
 sg13g2_decap_8 FILLER_18_821 ();
 sg13g2_decap_8 FILLER_18_828 ();
 sg13g2_decap_8 FILLER_18_835 ();
 sg13g2_decap_8 FILLER_18_842 ();
 sg13g2_decap_8 FILLER_18_849 ();
 sg13g2_decap_8 FILLER_18_856 ();
 sg13g2_decap_8 FILLER_18_863 ();
 sg13g2_decap_8 FILLER_18_870 ();
 sg13g2_decap_8 FILLER_18_877 ();
 sg13g2_decap_8 FILLER_18_884 ();
 sg13g2_decap_8 FILLER_18_891 ();
 sg13g2_decap_8 FILLER_18_898 ();
 sg13g2_decap_8 FILLER_18_905 ();
 sg13g2_decap_8 FILLER_18_912 ();
 sg13g2_decap_8 FILLER_18_919 ();
 sg13g2_decap_8 FILLER_18_926 ();
 sg13g2_decap_8 FILLER_18_933 ();
 sg13g2_decap_8 FILLER_18_940 ();
 sg13g2_decap_8 FILLER_18_947 ();
 sg13g2_decap_8 FILLER_18_954 ();
 sg13g2_decap_8 FILLER_18_961 ();
 sg13g2_decap_8 FILLER_18_968 ();
 sg13g2_decap_8 FILLER_18_975 ();
 sg13g2_decap_8 FILLER_18_982 ();
 sg13g2_decap_8 FILLER_18_989 ();
 sg13g2_decap_8 FILLER_18_996 ();
 sg13g2_decap_8 FILLER_18_1003 ();
 sg13g2_decap_8 FILLER_18_1010 ();
 sg13g2_decap_8 FILLER_18_1017 ();
 sg13g2_decap_4 FILLER_18_1024 ();
 sg13g2_fill_1 FILLER_18_1028 ();
 sg13g2_decap_8 FILLER_19_4 ();
 sg13g2_decap_8 FILLER_19_11 ();
 sg13g2_decap_8 FILLER_19_18 ();
 sg13g2_decap_8 FILLER_19_25 ();
 sg13g2_decap_8 FILLER_19_32 ();
 sg13g2_decap_8 FILLER_19_39 ();
 sg13g2_decap_8 FILLER_19_46 ();
 sg13g2_decap_8 FILLER_19_53 ();
 sg13g2_decap_8 FILLER_19_60 ();
 sg13g2_decap_8 FILLER_19_67 ();
 sg13g2_decap_8 FILLER_19_74 ();
 sg13g2_decap_8 FILLER_19_81 ();
 sg13g2_decap_8 FILLER_19_88 ();
 sg13g2_decap_8 FILLER_19_95 ();
 sg13g2_decap_8 FILLER_19_102 ();
 sg13g2_decap_8 FILLER_19_109 ();
 sg13g2_decap_8 FILLER_19_116 ();
 sg13g2_decap_8 FILLER_19_123 ();
 sg13g2_decap_8 FILLER_19_130 ();
 sg13g2_decap_8 FILLER_19_137 ();
 sg13g2_decap_8 FILLER_19_144 ();
 sg13g2_decap_4 FILLER_19_151 ();
 sg13g2_fill_1 FILLER_19_155 ();
 sg13g2_fill_2 FILLER_19_173 ();
 sg13g2_decap_8 FILLER_19_191 ();
 sg13g2_fill_2 FILLER_19_198 ();
 sg13g2_fill_1 FILLER_19_200 ();
 sg13g2_decap_8 FILLER_19_209 ();
 sg13g2_decap_8 FILLER_19_216 ();
 sg13g2_fill_2 FILLER_19_223 ();
 sg13g2_decap_8 FILLER_19_234 ();
 sg13g2_decap_8 FILLER_19_241 ();
 sg13g2_decap_8 FILLER_19_248 ();
 sg13g2_fill_2 FILLER_19_255 ();
 sg13g2_decap_8 FILLER_19_284 ();
 sg13g2_decap_8 FILLER_19_291 ();
 sg13g2_decap_8 FILLER_19_298 ();
 sg13g2_decap_8 FILLER_19_305 ();
 sg13g2_decap_8 FILLER_19_312 ();
 sg13g2_decap_8 FILLER_19_319 ();
 sg13g2_decap_8 FILLER_19_326 ();
 sg13g2_decap_8 FILLER_19_333 ();
 sg13g2_fill_2 FILLER_19_340 ();
 sg13g2_decap_8 FILLER_19_355 ();
 sg13g2_decap_8 FILLER_19_362 ();
 sg13g2_decap_8 FILLER_19_369 ();
 sg13g2_decap_8 FILLER_19_376 ();
 sg13g2_decap_8 FILLER_19_383 ();
 sg13g2_decap_4 FILLER_19_390 ();
 sg13g2_fill_2 FILLER_19_394 ();
 sg13g2_decap_4 FILLER_19_409 ();
 sg13g2_fill_1 FILLER_19_413 ();
 sg13g2_decap_4 FILLER_19_422 ();
 sg13g2_fill_2 FILLER_19_426 ();
 sg13g2_decap_8 FILLER_19_455 ();
 sg13g2_decap_8 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_490 ();
 sg13g2_decap_8 FILLER_19_497 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_532 ();
 sg13g2_decap_8 FILLER_19_539 ();
 sg13g2_decap_8 FILLER_19_546 ();
 sg13g2_decap_8 FILLER_19_553 ();
 sg13g2_decap_8 FILLER_19_560 ();
 sg13g2_decap_8 FILLER_19_567 ();
 sg13g2_decap_8 FILLER_19_574 ();
 sg13g2_decap_8 FILLER_19_581 ();
 sg13g2_decap_8 FILLER_19_588 ();
 sg13g2_decap_8 FILLER_19_595 ();
 sg13g2_decap_8 FILLER_19_602 ();
 sg13g2_decap_8 FILLER_19_609 ();
 sg13g2_decap_8 FILLER_19_616 ();
 sg13g2_decap_8 FILLER_19_623 ();
 sg13g2_decap_8 FILLER_19_630 ();
 sg13g2_decap_8 FILLER_19_637 ();
 sg13g2_decap_8 FILLER_19_644 ();
 sg13g2_decap_8 FILLER_19_651 ();
 sg13g2_decap_8 FILLER_19_658 ();
 sg13g2_decap_8 FILLER_19_665 ();
 sg13g2_decap_8 FILLER_19_672 ();
 sg13g2_decap_8 FILLER_19_679 ();
 sg13g2_decap_8 FILLER_19_686 ();
 sg13g2_decap_8 FILLER_19_693 ();
 sg13g2_decap_8 FILLER_19_700 ();
 sg13g2_decap_8 FILLER_19_707 ();
 sg13g2_decap_8 FILLER_19_714 ();
 sg13g2_decap_8 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_784 ();
 sg13g2_decap_8 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_798 ();
 sg13g2_decap_8 FILLER_19_805 ();
 sg13g2_decap_8 FILLER_19_812 ();
 sg13g2_decap_8 FILLER_19_819 ();
 sg13g2_decap_8 FILLER_19_826 ();
 sg13g2_decap_8 FILLER_19_833 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_decap_8 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_854 ();
 sg13g2_decap_8 FILLER_19_861 ();
 sg13g2_decap_8 FILLER_19_868 ();
 sg13g2_decap_8 FILLER_19_875 ();
 sg13g2_decap_8 FILLER_19_882 ();
 sg13g2_decap_8 FILLER_19_889 ();
 sg13g2_decap_8 FILLER_19_896 ();
 sg13g2_decap_8 FILLER_19_903 ();
 sg13g2_decap_8 FILLER_19_910 ();
 sg13g2_decap_8 FILLER_19_917 ();
 sg13g2_decap_8 FILLER_19_924 ();
 sg13g2_decap_8 FILLER_19_931 ();
 sg13g2_decap_8 FILLER_19_938 ();
 sg13g2_decap_8 FILLER_19_945 ();
 sg13g2_decap_8 FILLER_19_952 ();
 sg13g2_decap_8 FILLER_19_959 ();
 sg13g2_decap_8 FILLER_19_966 ();
 sg13g2_decap_8 FILLER_19_973 ();
 sg13g2_decap_8 FILLER_19_980 ();
 sg13g2_decap_8 FILLER_19_987 ();
 sg13g2_decap_8 FILLER_19_994 ();
 sg13g2_decap_8 FILLER_19_1001 ();
 sg13g2_decap_8 FILLER_19_1008 ();
 sg13g2_decap_8 FILLER_19_1015 ();
 sg13g2_decap_8 FILLER_19_1022 ();
 sg13g2_decap_8 FILLER_20_4 ();
 sg13g2_decap_8 FILLER_20_11 ();
 sg13g2_decap_8 FILLER_20_18 ();
 sg13g2_decap_8 FILLER_20_25 ();
 sg13g2_decap_8 FILLER_20_32 ();
 sg13g2_decap_8 FILLER_20_39 ();
 sg13g2_decap_8 FILLER_20_46 ();
 sg13g2_decap_8 FILLER_20_53 ();
 sg13g2_decap_8 FILLER_20_60 ();
 sg13g2_decap_8 FILLER_20_67 ();
 sg13g2_decap_8 FILLER_20_74 ();
 sg13g2_decap_8 FILLER_20_81 ();
 sg13g2_decap_8 FILLER_20_88 ();
 sg13g2_decap_4 FILLER_20_95 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_4 FILLER_20_140 ();
 sg13g2_fill_1 FILLER_20_144 ();
 sg13g2_decap_4 FILLER_20_181 ();
 sg13g2_fill_1 FILLER_20_185 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_fill_2 FILLER_20_315 ();
 sg13g2_fill_1 FILLER_20_344 ();
 sg13g2_decap_8 FILLER_20_353 ();
 sg13g2_decap_8 FILLER_20_360 ();
 sg13g2_decap_8 FILLER_20_367 ();
 sg13g2_decap_8 FILLER_20_374 ();
 sg13g2_decap_8 FILLER_20_381 ();
 sg13g2_decap_8 FILLER_20_388 ();
 sg13g2_decap_8 FILLER_20_395 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_20_409 ();
 sg13g2_decap_8 FILLER_20_416 ();
 sg13g2_fill_2 FILLER_20_423 ();
 sg13g2_decap_8 FILLER_20_434 ();
 sg13g2_decap_8 FILLER_20_441 ();
 sg13g2_decap_8 FILLER_20_448 ();
 sg13g2_decap_8 FILLER_20_455 ();
 sg13g2_decap_8 FILLER_20_462 ();
 sg13g2_fill_1 FILLER_20_469 ();
 sg13g2_decap_8 FILLER_20_483 ();
 sg13g2_decap_8 FILLER_20_490 ();
 sg13g2_decap_8 FILLER_20_497 ();
 sg13g2_decap_8 FILLER_20_504 ();
 sg13g2_decap_8 FILLER_20_511 ();
 sg13g2_decap_8 FILLER_20_518 ();
 sg13g2_decap_8 FILLER_20_525 ();
 sg13g2_decap_8 FILLER_20_532 ();
 sg13g2_decap_8 FILLER_20_539 ();
 sg13g2_decap_8 FILLER_20_546 ();
 sg13g2_decap_8 FILLER_20_553 ();
 sg13g2_decap_8 FILLER_20_560 ();
 sg13g2_fill_2 FILLER_20_567 ();
 sg13g2_fill_1 FILLER_20_569 ();
 sg13g2_decap_8 FILLER_20_579 ();
 sg13g2_decap_8 FILLER_20_586 ();
 sg13g2_decap_8 FILLER_20_593 ();
 sg13g2_decap_8 FILLER_20_600 ();
 sg13g2_decap_8 FILLER_20_607 ();
 sg13g2_decap_8 FILLER_20_614 ();
 sg13g2_decap_8 FILLER_20_621 ();
 sg13g2_decap_8 FILLER_20_628 ();
 sg13g2_decap_8 FILLER_20_635 ();
 sg13g2_decap_8 FILLER_20_642 ();
 sg13g2_decap_8 FILLER_20_649 ();
 sg13g2_decap_8 FILLER_20_656 ();
 sg13g2_decap_8 FILLER_20_663 ();
 sg13g2_decap_8 FILLER_20_670 ();
 sg13g2_decap_8 FILLER_20_677 ();
 sg13g2_decap_8 FILLER_20_684 ();
 sg13g2_decap_8 FILLER_20_691 ();
 sg13g2_decap_8 FILLER_20_698 ();
 sg13g2_decap_8 FILLER_20_705 ();
 sg13g2_decap_8 FILLER_20_712 ();
 sg13g2_decap_8 FILLER_20_719 ();
 sg13g2_decap_8 FILLER_20_726 ();
 sg13g2_decap_8 FILLER_20_733 ();
 sg13g2_decap_8 FILLER_20_740 ();
 sg13g2_decap_8 FILLER_20_747 ();
 sg13g2_decap_8 FILLER_20_754 ();
 sg13g2_decap_8 FILLER_20_761 ();
 sg13g2_decap_8 FILLER_20_768 ();
 sg13g2_decap_8 FILLER_20_775 ();
 sg13g2_decap_8 FILLER_20_782 ();
 sg13g2_decap_8 FILLER_20_789 ();
 sg13g2_decap_8 FILLER_20_796 ();
 sg13g2_decap_8 FILLER_20_803 ();
 sg13g2_decap_8 FILLER_20_810 ();
 sg13g2_decap_8 FILLER_20_817 ();
 sg13g2_decap_8 FILLER_20_824 ();
 sg13g2_decap_8 FILLER_20_831 ();
 sg13g2_decap_8 FILLER_20_838 ();
 sg13g2_decap_8 FILLER_20_845 ();
 sg13g2_decap_8 FILLER_20_852 ();
 sg13g2_decap_8 FILLER_20_859 ();
 sg13g2_decap_8 FILLER_20_866 ();
 sg13g2_decap_8 FILLER_20_873 ();
 sg13g2_decap_8 FILLER_20_880 ();
 sg13g2_decap_8 FILLER_20_887 ();
 sg13g2_decap_8 FILLER_20_894 ();
 sg13g2_decap_8 FILLER_20_901 ();
 sg13g2_decap_8 FILLER_20_908 ();
 sg13g2_decap_8 FILLER_20_915 ();
 sg13g2_decap_8 FILLER_20_922 ();
 sg13g2_decap_8 FILLER_20_929 ();
 sg13g2_decap_8 FILLER_20_936 ();
 sg13g2_decap_8 FILLER_20_943 ();
 sg13g2_decap_8 FILLER_20_950 ();
 sg13g2_decap_8 FILLER_20_957 ();
 sg13g2_decap_8 FILLER_20_964 ();
 sg13g2_decap_8 FILLER_20_971 ();
 sg13g2_decap_8 FILLER_20_978 ();
 sg13g2_decap_8 FILLER_20_985 ();
 sg13g2_decap_8 FILLER_20_992 ();
 sg13g2_decap_8 FILLER_20_999 ();
 sg13g2_decap_8 FILLER_20_1006 ();
 sg13g2_decap_8 FILLER_20_1013 ();
 sg13g2_decap_8 FILLER_20_1020 ();
 sg13g2_fill_2 FILLER_20_1027 ();
 sg13g2_decap_8 FILLER_21_4 ();
 sg13g2_decap_8 FILLER_21_11 ();
 sg13g2_decap_8 FILLER_21_18 ();
 sg13g2_decap_4 FILLER_21_29 ();
 sg13g2_fill_2 FILLER_21_33 ();
 sg13g2_decap_8 FILLER_21_44 ();
 sg13g2_decap_8 FILLER_21_51 ();
 sg13g2_decap_8 FILLER_21_58 ();
 sg13g2_decap_8 FILLER_21_65 ();
 sg13g2_decap_8 FILLER_21_72 ();
 sg13g2_decap_8 FILLER_21_79 ();
 sg13g2_decap_8 FILLER_21_86 ();
 sg13g2_decap_8 FILLER_21_120 ();
 sg13g2_decap_8 FILLER_21_127 ();
 sg13g2_decap_8 FILLER_21_134 ();
 sg13g2_decap_8 FILLER_21_141 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_218 ();
 sg13g2_decap_8 FILLER_21_225 ();
 sg13g2_decap_4 FILLER_21_232 ();
 sg13g2_fill_1 FILLER_21_236 ();
 sg13g2_decap_8 FILLER_21_246 ();
 sg13g2_decap_8 FILLER_21_253 ();
 sg13g2_decap_4 FILLER_21_260 ();
 sg13g2_fill_2 FILLER_21_264 ();
 sg13g2_decap_8 FILLER_21_293 ();
 sg13g2_decap_8 FILLER_21_300 ();
 sg13g2_decap_8 FILLER_21_307 ();
 sg13g2_decap_8 FILLER_21_314 ();
 sg13g2_decap_8 FILLER_21_321 ();
 sg13g2_decap_4 FILLER_21_328 ();
 sg13g2_fill_2 FILLER_21_332 ();
 sg13g2_fill_2 FILLER_21_342 ();
 sg13g2_fill_1 FILLER_21_344 ();
 sg13g2_decap_8 FILLER_21_354 ();
 sg13g2_fill_1 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_decap_8 FILLER_21_405 ();
 sg13g2_fill_2 FILLER_21_412 ();
 sg13g2_decap_8 FILLER_21_422 ();
 sg13g2_decap_8 FILLER_21_429 ();
 sg13g2_decap_8 FILLER_21_436 ();
 sg13g2_decap_8 FILLER_21_443 ();
 sg13g2_decap_8 FILLER_21_450 ();
 sg13g2_decap_4 FILLER_21_457 ();
 sg13g2_fill_1 FILLER_21_461 ();
 sg13g2_decap_8 FILLER_21_475 ();
 sg13g2_decap_8 FILLER_21_482 ();
 sg13g2_fill_2 FILLER_21_489 ();
 sg13g2_decap_8 FILLER_21_518 ();
 sg13g2_decap_8 FILLER_21_525 ();
 sg13g2_decap_8 FILLER_21_532 ();
 sg13g2_decap_4 FILLER_21_539 ();
 sg13g2_decap_8 FILLER_21_570 ();
 sg13g2_decap_4 FILLER_21_577 ();
 sg13g2_fill_2 FILLER_21_581 ();
 sg13g2_decap_8 FILLER_21_610 ();
 sg13g2_decap_8 FILLER_21_617 ();
 sg13g2_decap_8 FILLER_21_624 ();
 sg13g2_decap_8 FILLER_21_631 ();
 sg13g2_decap_8 FILLER_21_638 ();
 sg13g2_decap_8 FILLER_21_645 ();
 sg13g2_decap_8 FILLER_21_652 ();
 sg13g2_decap_8 FILLER_21_659 ();
 sg13g2_decap_8 FILLER_21_666 ();
 sg13g2_decap_8 FILLER_21_673 ();
 sg13g2_decap_8 FILLER_21_680 ();
 sg13g2_decap_8 FILLER_21_687 ();
 sg13g2_decap_8 FILLER_21_694 ();
 sg13g2_decap_8 FILLER_21_701 ();
 sg13g2_decap_8 FILLER_21_708 ();
 sg13g2_decap_8 FILLER_21_715 ();
 sg13g2_decap_8 FILLER_21_722 ();
 sg13g2_decap_8 FILLER_21_729 ();
 sg13g2_decap_8 FILLER_21_736 ();
 sg13g2_decap_8 FILLER_21_743 ();
 sg13g2_decap_8 FILLER_21_750 ();
 sg13g2_decap_8 FILLER_21_757 ();
 sg13g2_decap_8 FILLER_21_764 ();
 sg13g2_decap_8 FILLER_21_771 ();
 sg13g2_decap_8 FILLER_21_778 ();
 sg13g2_decap_8 FILLER_21_785 ();
 sg13g2_decap_8 FILLER_21_792 ();
 sg13g2_decap_8 FILLER_21_799 ();
 sg13g2_decap_8 FILLER_21_806 ();
 sg13g2_decap_8 FILLER_21_813 ();
 sg13g2_decap_8 FILLER_21_820 ();
 sg13g2_decap_8 FILLER_21_827 ();
 sg13g2_decap_8 FILLER_21_834 ();
 sg13g2_decap_8 FILLER_21_841 ();
 sg13g2_decap_8 FILLER_21_848 ();
 sg13g2_decap_8 FILLER_21_855 ();
 sg13g2_decap_8 FILLER_21_862 ();
 sg13g2_decap_8 FILLER_21_869 ();
 sg13g2_decap_8 FILLER_21_876 ();
 sg13g2_decap_8 FILLER_21_883 ();
 sg13g2_decap_8 FILLER_21_890 ();
 sg13g2_decap_8 FILLER_21_897 ();
 sg13g2_decap_8 FILLER_21_904 ();
 sg13g2_decap_8 FILLER_21_911 ();
 sg13g2_decap_8 FILLER_21_918 ();
 sg13g2_decap_8 FILLER_21_925 ();
 sg13g2_decap_8 FILLER_21_932 ();
 sg13g2_decap_8 FILLER_21_939 ();
 sg13g2_decap_8 FILLER_21_946 ();
 sg13g2_decap_8 FILLER_21_953 ();
 sg13g2_decap_8 FILLER_21_960 ();
 sg13g2_decap_8 FILLER_21_967 ();
 sg13g2_decap_8 FILLER_21_974 ();
 sg13g2_decap_8 FILLER_21_981 ();
 sg13g2_decap_8 FILLER_21_988 ();
 sg13g2_decap_8 FILLER_21_995 ();
 sg13g2_decap_8 FILLER_21_1002 ();
 sg13g2_decap_8 FILLER_21_1009 ();
 sg13g2_decap_8 FILLER_21_1016 ();
 sg13g2_decap_4 FILLER_21_1023 ();
 sg13g2_fill_2 FILLER_21_1027 ();
 sg13g2_decap_8 FILLER_22_4 ();
 sg13g2_decap_4 FILLER_22_11 ();
 sg13g2_fill_1 FILLER_22_15 ();
 sg13g2_decap_8 FILLER_22_43 ();
 sg13g2_decap_8 FILLER_22_50 ();
 sg13g2_decap_8 FILLER_22_57 ();
 sg13g2_decap_8 FILLER_22_64 ();
 sg13g2_decap_8 FILLER_22_71 ();
 sg13g2_decap_4 FILLER_22_78 ();
 sg13g2_fill_1 FILLER_22_82 ();
 sg13g2_decap_8 FILLER_22_110 ();
 sg13g2_decap_8 FILLER_22_117 ();
 sg13g2_decap_8 FILLER_22_124 ();
 sg13g2_decap_8 FILLER_22_131 ();
 sg13g2_decap_8 FILLER_22_138 ();
 sg13g2_decap_8 FILLER_22_145 ();
 sg13g2_decap_4 FILLER_22_152 ();
 sg13g2_fill_2 FILLER_22_156 ();
 sg13g2_decap_4 FILLER_22_162 ();
 sg13g2_fill_2 FILLER_22_166 ();
 sg13g2_decap_8 FILLER_22_177 ();
 sg13g2_decap_8 FILLER_22_184 ();
 sg13g2_decap_8 FILLER_22_191 ();
 sg13g2_decap_8 FILLER_22_198 ();
 sg13g2_decap_8 FILLER_22_205 ();
 sg13g2_decap_8 FILLER_22_212 ();
 sg13g2_decap_8 FILLER_22_219 ();
 sg13g2_decap_8 FILLER_22_226 ();
 sg13g2_decap_8 FILLER_22_233 ();
 sg13g2_decap_8 FILLER_22_240 ();
 sg13g2_decap_8 FILLER_22_247 ();
 sg13g2_decap_8 FILLER_22_254 ();
 sg13g2_decap_8 FILLER_22_302 ();
 sg13g2_decap_8 FILLER_22_309 ();
 sg13g2_decap_8 FILLER_22_316 ();
 sg13g2_decap_8 FILLER_22_323 ();
 sg13g2_decap_8 FILLER_22_330 ();
 sg13g2_decap_8 FILLER_22_337 ();
 sg13g2_decap_8 FILLER_22_344 ();
 sg13g2_decap_8 FILLER_22_351 ();
 sg13g2_decap_8 FILLER_22_358 ();
 sg13g2_decap_8 FILLER_22_365 ();
 sg13g2_decap_8 FILLER_22_372 ();
 sg13g2_decap_8 FILLER_22_379 ();
 sg13g2_fill_2 FILLER_22_386 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_decap_8 FILLER_22_404 ();
 sg13g2_decap_8 FILLER_22_411 ();
 sg13g2_decap_8 FILLER_22_418 ();
 sg13g2_decap_8 FILLER_22_425 ();
 sg13g2_decap_4 FILLER_22_432 ();
 sg13g2_fill_2 FILLER_22_436 ();
 sg13g2_decap_8 FILLER_22_451 ();
 sg13g2_decap_8 FILLER_22_458 ();
 sg13g2_decap_8 FILLER_22_465 ();
 sg13g2_decap_8 FILLER_22_472 ();
 sg13g2_decap_8 FILLER_22_479 ();
 sg13g2_decap_8 FILLER_22_486 ();
 sg13g2_decap_8 FILLER_22_493 ();
 sg13g2_fill_2 FILLER_22_500 ();
 sg13g2_fill_1 FILLER_22_506 ();
 sg13g2_decap_4 FILLER_22_520 ();
 sg13g2_fill_2 FILLER_22_524 ();
 sg13g2_decap_8 FILLER_22_530 ();
 sg13g2_fill_1 FILLER_22_537 ();
 sg13g2_decap_8 FILLER_22_543 ();
 sg13g2_decap_8 FILLER_22_550 ();
 sg13g2_decap_8 FILLER_22_557 ();
 sg13g2_decap_4 FILLER_22_564 ();
 sg13g2_decap_8 FILLER_22_576 ();
 sg13g2_decap_8 FILLER_22_583 ();
 sg13g2_decap_8 FILLER_22_590 ();
 sg13g2_decap_8 FILLER_22_597 ();
 sg13g2_decap_8 FILLER_22_604 ();
 sg13g2_decap_8 FILLER_22_611 ();
 sg13g2_decap_8 FILLER_22_618 ();
 sg13g2_decap_8 FILLER_22_625 ();
 sg13g2_decap_8 FILLER_22_632 ();
 sg13g2_decap_8 FILLER_22_639 ();
 sg13g2_decap_8 FILLER_22_646 ();
 sg13g2_decap_8 FILLER_22_653 ();
 sg13g2_decap_8 FILLER_22_660 ();
 sg13g2_decap_8 FILLER_22_667 ();
 sg13g2_decap_8 FILLER_22_674 ();
 sg13g2_decap_8 FILLER_22_681 ();
 sg13g2_decap_8 FILLER_22_688 ();
 sg13g2_decap_8 FILLER_22_695 ();
 sg13g2_decap_8 FILLER_22_702 ();
 sg13g2_decap_8 FILLER_22_709 ();
 sg13g2_decap_8 FILLER_22_716 ();
 sg13g2_decap_8 FILLER_22_723 ();
 sg13g2_decap_8 FILLER_22_730 ();
 sg13g2_decap_8 FILLER_22_737 ();
 sg13g2_decap_8 FILLER_22_744 ();
 sg13g2_decap_8 FILLER_22_751 ();
 sg13g2_decap_8 FILLER_22_758 ();
 sg13g2_decap_8 FILLER_22_765 ();
 sg13g2_decap_8 FILLER_22_772 ();
 sg13g2_decap_8 FILLER_22_779 ();
 sg13g2_decap_8 FILLER_22_786 ();
 sg13g2_decap_8 FILLER_22_793 ();
 sg13g2_decap_8 FILLER_22_800 ();
 sg13g2_decap_8 FILLER_22_807 ();
 sg13g2_decap_8 FILLER_22_814 ();
 sg13g2_decap_8 FILLER_22_821 ();
 sg13g2_decap_8 FILLER_22_828 ();
 sg13g2_decap_8 FILLER_22_835 ();
 sg13g2_decap_8 FILLER_22_842 ();
 sg13g2_decap_8 FILLER_22_849 ();
 sg13g2_decap_8 FILLER_22_856 ();
 sg13g2_decap_8 FILLER_22_863 ();
 sg13g2_decap_8 FILLER_22_870 ();
 sg13g2_decap_8 FILLER_22_877 ();
 sg13g2_decap_8 FILLER_22_884 ();
 sg13g2_decap_8 FILLER_22_891 ();
 sg13g2_decap_8 FILLER_22_898 ();
 sg13g2_decap_8 FILLER_22_905 ();
 sg13g2_decap_8 FILLER_22_912 ();
 sg13g2_decap_8 FILLER_22_919 ();
 sg13g2_decap_8 FILLER_22_926 ();
 sg13g2_decap_8 FILLER_22_933 ();
 sg13g2_decap_8 FILLER_22_940 ();
 sg13g2_decap_8 FILLER_22_947 ();
 sg13g2_decap_8 FILLER_22_954 ();
 sg13g2_decap_8 FILLER_22_961 ();
 sg13g2_decap_8 FILLER_22_968 ();
 sg13g2_decap_8 FILLER_22_975 ();
 sg13g2_decap_8 FILLER_22_982 ();
 sg13g2_decap_8 FILLER_22_989 ();
 sg13g2_decap_8 FILLER_22_996 ();
 sg13g2_decap_8 FILLER_22_1003 ();
 sg13g2_decap_8 FILLER_22_1010 ();
 sg13g2_decap_8 FILLER_22_1017 ();
 sg13g2_decap_4 FILLER_22_1024 ();
 sg13g2_fill_1 FILLER_22_1028 ();
 sg13g2_decap_8 FILLER_23_4 ();
 sg13g2_decap_4 FILLER_23_11 ();
 sg13g2_fill_2 FILLER_23_15 ();
 sg13g2_decap_8 FILLER_23_44 ();
 sg13g2_decap_8 FILLER_23_51 ();
 sg13g2_decap_8 FILLER_23_58 ();
 sg13g2_decap_8 FILLER_23_65 ();
 sg13g2_decap_8 FILLER_23_72 ();
 sg13g2_decap_8 FILLER_23_79 ();
 sg13g2_decap_8 FILLER_23_86 ();
 sg13g2_decap_8 FILLER_23_93 ();
 sg13g2_decap_4 FILLER_23_100 ();
 sg13g2_fill_1 FILLER_23_104 ();
 sg13g2_decap_8 FILLER_23_113 ();
 sg13g2_decap_8 FILLER_23_120 ();
 sg13g2_decap_8 FILLER_23_127 ();
 sg13g2_decap_8 FILLER_23_134 ();
 sg13g2_decap_8 FILLER_23_141 ();
 sg13g2_decap_8 FILLER_23_148 ();
 sg13g2_decap_8 FILLER_23_155 ();
 sg13g2_decap_8 FILLER_23_162 ();
 sg13g2_decap_8 FILLER_23_169 ();
 sg13g2_decap_8 FILLER_23_176 ();
 sg13g2_decap_8 FILLER_23_183 ();
 sg13g2_decap_8 FILLER_23_190 ();
 sg13g2_decap_8 FILLER_23_197 ();
 sg13g2_decap_8 FILLER_23_204 ();
 sg13g2_decap_8 FILLER_23_211 ();
 sg13g2_decap_8 FILLER_23_218 ();
 sg13g2_decap_8 FILLER_23_225 ();
 sg13g2_decap_8 FILLER_23_232 ();
 sg13g2_decap_8 FILLER_23_239 ();
 sg13g2_decap_8 FILLER_23_246 ();
 sg13g2_decap_8 FILLER_23_253 ();
 sg13g2_decap_8 FILLER_23_260 ();
 sg13g2_decap_4 FILLER_23_267 ();
 sg13g2_fill_2 FILLER_23_279 ();
 sg13g2_decap_8 FILLER_23_290 ();
 sg13g2_decap_8 FILLER_23_297 ();
 sg13g2_decap_8 FILLER_23_304 ();
 sg13g2_decap_8 FILLER_23_311 ();
 sg13g2_decap_8 FILLER_23_318 ();
 sg13g2_decap_8 FILLER_23_325 ();
 sg13g2_decap_8 FILLER_23_332 ();
 sg13g2_fill_2 FILLER_23_339 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_fill_1 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_406 ();
 sg13g2_decap_4 FILLER_23_413 ();
 sg13g2_decap_8 FILLER_23_444 ();
 sg13g2_decap_8 FILLER_23_451 ();
 sg13g2_decap_8 FILLER_23_458 ();
 sg13g2_decap_8 FILLER_23_465 ();
 sg13g2_decap_8 FILLER_23_472 ();
 sg13g2_decap_8 FILLER_23_479 ();
 sg13g2_decap_8 FILLER_23_486 ();
 sg13g2_decap_8 FILLER_23_493 ();
 sg13g2_fill_1 FILLER_23_500 ();
 sg13g2_decap_8 FILLER_23_537 ();
 sg13g2_decap_8 FILLER_23_544 ();
 sg13g2_decap_8 FILLER_23_551 ();
 sg13g2_decap_8 FILLER_23_558 ();
 sg13g2_fill_2 FILLER_23_565 ();
 sg13g2_fill_1 FILLER_23_567 ();
 sg13g2_decap_8 FILLER_23_572 ();
 sg13g2_decap_8 FILLER_23_579 ();
 sg13g2_decap_8 FILLER_23_586 ();
 sg13g2_decap_8 FILLER_23_593 ();
 sg13g2_decap_8 FILLER_23_600 ();
 sg13g2_decap_8 FILLER_23_607 ();
 sg13g2_decap_8 FILLER_23_614 ();
 sg13g2_decap_8 FILLER_23_621 ();
 sg13g2_decap_8 FILLER_23_628 ();
 sg13g2_decap_8 FILLER_23_635 ();
 sg13g2_decap_8 FILLER_23_642 ();
 sg13g2_decap_8 FILLER_23_649 ();
 sg13g2_decap_8 FILLER_23_656 ();
 sg13g2_decap_8 FILLER_23_663 ();
 sg13g2_decap_8 FILLER_23_670 ();
 sg13g2_decap_8 FILLER_23_677 ();
 sg13g2_decap_8 FILLER_23_684 ();
 sg13g2_decap_8 FILLER_23_691 ();
 sg13g2_decap_8 FILLER_23_698 ();
 sg13g2_decap_8 FILLER_23_705 ();
 sg13g2_decap_8 FILLER_23_712 ();
 sg13g2_decap_8 FILLER_23_719 ();
 sg13g2_decap_8 FILLER_23_726 ();
 sg13g2_decap_8 FILLER_23_733 ();
 sg13g2_decap_8 FILLER_23_740 ();
 sg13g2_decap_8 FILLER_23_747 ();
 sg13g2_decap_8 FILLER_23_754 ();
 sg13g2_decap_8 FILLER_23_761 ();
 sg13g2_decap_8 FILLER_23_768 ();
 sg13g2_decap_8 FILLER_23_775 ();
 sg13g2_decap_8 FILLER_23_782 ();
 sg13g2_decap_8 FILLER_23_789 ();
 sg13g2_decap_8 FILLER_23_796 ();
 sg13g2_decap_8 FILLER_23_803 ();
 sg13g2_decap_8 FILLER_23_810 ();
 sg13g2_decap_8 FILLER_23_817 ();
 sg13g2_decap_8 FILLER_23_824 ();
 sg13g2_decap_8 FILLER_23_831 ();
 sg13g2_decap_8 FILLER_23_838 ();
 sg13g2_decap_8 FILLER_23_845 ();
 sg13g2_decap_8 FILLER_23_852 ();
 sg13g2_decap_8 FILLER_23_859 ();
 sg13g2_decap_8 FILLER_23_866 ();
 sg13g2_decap_8 FILLER_23_873 ();
 sg13g2_decap_8 FILLER_23_880 ();
 sg13g2_decap_8 FILLER_23_887 ();
 sg13g2_decap_8 FILLER_23_894 ();
 sg13g2_decap_8 FILLER_23_901 ();
 sg13g2_decap_8 FILLER_23_908 ();
 sg13g2_decap_8 FILLER_23_915 ();
 sg13g2_decap_8 FILLER_23_922 ();
 sg13g2_decap_8 FILLER_23_929 ();
 sg13g2_decap_8 FILLER_23_936 ();
 sg13g2_decap_8 FILLER_23_943 ();
 sg13g2_decap_8 FILLER_23_950 ();
 sg13g2_decap_8 FILLER_23_957 ();
 sg13g2_decap_8 FILLER_23_964 ();
 sg13g2_decap_8 FILLER_23_971 ();
 sg13g2_decap_8 FILLER_23_978 ();
 sg13g2_decap_8 FILLER_23_985 ();
 sg13g2_decap_8 FILLER_23_992 ();
 sg13g2_decap_8 FILLER_23_999 ();
 sg13g2_decap_8 FILLER_23_1006 ();
 sg13g2_decap_8 FILLER_23_1013 ();
 sg13g2_decap_8 FILLER_23_1020 ();
 sg13g2_fill_2 FILLER_23_1027 ();
 sg13g2_decap_8 FILLER_24_4 ();
 sg13g2_decap_8 FILLER_24_11 ();
 sg13g2_decap_4 FILLER_24_18 ();
 sg13g2_fill_2 FILLER_24_22 ();
 sg13g2_decap_8 FILLER_24_50 ();
 sg13g2_decap_8 FILLER_24_57 ();
 sg13g2_decap_4 FILLER_24_64 ();
 sg13g2_fill_2 FILLER_24_68 ();
 sg13g2_decap_8 FILLER_24_97 ();
 sg13g2_decap_8 FILLER_24_104 ();
 sg13g2_decap_8 FILLER_24_111 ();
 sg13g2_fill_2 FILLER_24_118 ();
 sg13g2_decap_8 FILLER_24_129 ();
 sg13g2_decap_8 FILLER_24_136 ();
 sg13g2_decap_8 FILLER_24_143 ();
 sg13g2_decap_8 FILLER_24_150 ();
 sg13g2_decap_8 FILLER_24_157 ();
 sg13g2_decap_8 FILLER_24_164 ();
 sg13g2_decap_8 FILLER_24_171 ();
 sg13g2_decap_8 FILLER_24_178 ();
 sg13g2_decap_8 FILLER_24_185 ();
 sg13g2_decap_8 FILLER_24_192 ();
 sg13g2_fill_2 FILLER_24_199 ();
 sg13g2_decap_8 FILLER_24_229 ();
 sg13g2_decap_8 FILLER_24_236 ();
 sg13g2_decap_8 FILLER_24_243 ();
 sg13g2_decap_8 FILLER_24_250 ();
 sg13g2_decap_8 FILLER_24_257 ();
 sg13g2_decap_8 FILLER_24_264 ();
 sg13g2_decap_8 FILLER_24_271 ();
 sg13g2_decap_8 FILLER_24_278 ();
 sg13g2_decap_8 FILLER_24_285 ();
 sg13g2_fill_2 FILLER_24_292 ();
 sg13g2_decap_8 FILLER_24_302 ();
 sg13g2_decap_8 FILLER_24_309 ();
 sg13g2_fill_1 FILLER_24_316 ();
 sg13g2_decap_8 FILLER_24_344 ();
 sg13g2_decap_4 FILLER_24_351 ();
 sg13g2_fill_1 FILLER_24_355 ();
 sg13g2_decap_8 FILLER_24_369 ();
 sg13g2_decap_8 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_24_383 ();
 sg13g2_decap_8 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_8 FILLER_24_404 ();
 sg13g2_decap_8 FILLER_24_411 ();
 sg13g2_decap_8 FILLER_24_418 ();
 sg13g2_decap_8 FILLER_24_425 ();
 sg13g2_decap_8 FILLER_24_432 ();
 sg13g2_decap_8 FILLER_24_439 ();
 sg13g2_decap_8 FILLER_24_446 ();
 sg13g2_decap_8 FILLER_24_453 ();
 sg13g2_decap_8 FILLER_24_460 ();
 sg13g2_decap_8 FILLER_24_467 ();
 sg13g2_decap_8 FILLER_24_474 ();
 sg13g2_decap_8 FILLER_24_481 ();
 sg13g2_decap_8 FILLER_24_488 ();
 sg13g2_decap_8 FILLER_24_495 ();
 sg13g2_decap_8 FILLER_24_502 ();
 sg13g2_decap_8 FILLER_24_509 ();
 sg13g2_decap_8 FILLER_24_516 ();
 sg13g2_decap_8 FILLER_24_523 ();
 sg13g2_decap_8 FILLER_24_530 ();
 sg13g2_decap_8 FILLER_24_537 ();
 sg13g2_decap_8 FILLER_24_544 ();
 sg13g2_decap_8 FILLER_24_560 ();
 sg13g2_fill_2 FILLER_24_567 ();
 sg13g2_decap_8 FILLER_24_600 ();
 sg13g2_decap_8 FILLER_24_607 ();
 sg13g2_decap_8 FILLER_24_614 ();
 sg13g2_decap_8 FILLER_24_621 ();
 sg13g2_decap_8 FILLER_24_628 ();
 sg13g2_decap_8 FILLER_24_635 ();
 sg13g2_decap_8 FILLER_24_642 ();
 sg13g2_decap_8 FILLER_24_649 ();
 sg13g2_decap_8 FILLER_24_656 ();
 sg13g2_decap_8 FILLER_24_663 ();
 sg13g2_decap_8 FILLER_24_670 ();
 sg13g2_decap_8 FILLER_24_677 ();
 sg13g2_decap_8 FILLER_24_684 ();
 sg13g2_decap_8 FILLER_24_691 ();
 sg13g2_decap_8 FILLER_24_698 ();
 sg13g2_decap_8 FILLER_24_705 ();
 sg13g2_decap_8 FILLER_24_712 ();
 sg13g2_decap_8 FILLER_24_719 ();
 sg13g2_decap_8 FILLER_24_726 ();
 sg13g2_decap_8 FILLER_24_733 ();
 sg13g2_decap_8 FILLER_24_740 ();
 sg13g2_decap_8 FILLER_24_747 ();
 sg13g2_decap_8 FILLER_24_754 ();
 sg13g2_decap_8 FILLER_24_761 ();
 sg13g2_decap_8 FILLER_24_768 ();
 sg13g2_decap_8 FILLER_24_775 ();
 sg13g2_decap_8 FILLER_24_782 ();
 sg13g2_decap_8 FILLER_24_789 ();
 sg13g2_decap_8 FILLER_24_796 ();
 sg13g2_decap_8 FILLER_24_803 ();
 sg13g2_decap_8 FILLER_24_810 ();
 sg13g2_decap_8 FILLER_24_817 ();
 sg13g2_decap_8 FILLER_24_824 ();
 sg13g2_decap_8 FILLER_24_831 ();
 sg13g2_decap_8 FILLER_24_838 ();
 sg13g2_decap_8 FILLER_24_845 ();
 sg13g2_decap_8 FILLER_24_852 ();
 sg13g2_decap_8 FILLER_24_859 ();
 sg13g2_decap_8 FILLER_24_866 ();
 sg13g2_decap_8 FILLER_24_873 ();
 sg13g2_decap_8 FILLER_24_880 ();
 sg13g2_decap_8 FILLER_24_887 ();
 sg13g2_decap_8 FILLER_24_894 ();
 sg13g2_decap_8 FILLER_24_901 ();
 sg13g2_decap_8 FILLER_24_908 ();
 sg13g2_decap_8 FILLER_24_915 ();
 sg13g2_decap_8 FILLER_24_922 ();
 sg13g2_decap_8 FILLER_24_929 ();
 sg13g2_decap_8 FILLER_24_936 ();
 sg13g2_decap_8 FILLER_24_943 ();
 sg13g2_decap_8 FILLER_24_950 ();
 sg13g2_decap_8 FILLER_24_957 ();
 sg13g2_decap_8 FILLER_24_964 ();
 sg13g2_decap_8 FILLER_24_971 ();
 sg13g2_decap_8 FILLER_24_978 ();
 sg13g2_decap_8 FILLER_24_985 ();
 sg13g2_decap_8 FILLER_24_992 ();
 sg13g2_decap_8 FILLER_24_999 ();
 sg13g2_decap_8 FILLER_24_1006 ();
 sg13g2_decap_8 FILLER_24_1013 ();
 sg13g2_decap_8 FILLER_24_1020 ();
 sg13g2_fill_2 FILLER_24_1027 ();
 sg13g2_decap_8 FILLER_25_4 ();
 sg13g2_decap_8 FILLER_25_11 ();
 sg13g2_decap_8 FILLER_25_18 ();
 sg13g2_decap_8 FILLER_25_25 ();
 sg13g2_decap_8 FILLER_25_32 ();
 sg13g2_fill_1 FILLER_25_39 ();
 sg13g2_decap_8 FILLER_25_52 ();
 sg13g2_decap_8 FILLER_25_59 ();
 sg13g2_decap_8 FILLER_25_66 ();
 sg13g2_decap_8 FILLER_25_73 ();
 sg13g2_decap_8 FILLER_25_80 ();
 sg13g2_decap_8 FILLER_25_87 ();
 sg13g2_decap_8 FILLER_25_94 ();
 sg13g2_decap_8 FILLER_25_101 ();
 sg13g2_decap_8 FILLER_25_108 ();
 sg13g2_fill_2 FILLER_25_115 ();
 sg13g2_decap_8 FILLER_25_125 ();
 sg13g2_decap_8 FILLER_25_132 ();
 sg13g2_decap_8 FILLER_25_139 ();
 sg13g2_decap_8 FILLER_25_146 ();
 sg13g2_decap_8 FILLER_25_153 ();
 sg13g2_decap_8 FILLER_25_160 ();
 sg13g2_decap_8 FILLER_25_167 ();
 sg13g2_decap_8 FILLER_25_174 ();
 sg13g2_decap_8 FILLER_25_181 ();
 sg13g2_decap_8 FILLER_25_188 ();
 sg13g2_decap_4 FILLER_25_195 ();
 sg13g2_decap_8 FILLER_25_240 ();
 sg13g2_decap_8 FILLER_25_247 ();
 sg13g2_decap_8 FILLER_25_254 ();
 sg13g2_decap_8 FILLER_25_261 ();
 sg13g2_decap_8 FILLER_25_268 ();
 sg13g2_decap_8 FILLER_25_275 ();
 sg13g2_fill_2 FILLER_25_282 ();
 sg13g2_decap_8 FILLER_25_292 ();
 sg13g2_decap_8 FILLER_25_299 ();
 sg13g2_decap_8 FILLER_25_306 ();
 sg13g2_decap_4 FILLER_25_313 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_4 FILLER_25_392 ();
 sg13g2_decap_4 FILLER_25_413 ();
 sg13g2_fill_1 FILLER_25_417 ();
 sg13g2_decap_8 FILLER_25_427 ();
 sg13g2_decap_8 FILLER_25_434 ();
 sg13g2_decap_8 FILLER_25_441 ();
 sg13g2_decap_8 FILLER_25_448 ();
 sg13g2_decap_4 FILLER_25_455 ();
 sg13g2_fill_1 FILLER_25_459 ();
 sg13g2_decap_8 FILLER_25_464 ();
 sg13g2_fill_2 FILLER_25_471 ();
 sg13g2_decap_8 FILLER_25_482 ();
 sg13g2_decap_8 FILLER_25_489 ();
 sg13g2_decap_8 FILLER_25_496 ();
 sg13g2_decap_8 FILLER_25_503 ();
 sg13g2_decap_8 FILLER_25_510 ();
 sg13g2_decap_8 FILLER_25_517 ();
 sg13g2_decap_8 FILLER_25_524 ();
 sg13g2_decap_4 FILLER_25_531 ();
 sg13g2_fill_1 FILLER_25_535 ();
 sg13g2_decap_8 FILLER_25_563 ();
 sg13g2_decap_8 FILLER_25_570 ();
 sg13g2_decap_8 FILLER_25_577 ();
 sg13g2_fill_1 FILLER_25_584 ();
 sg13g2_decap_8 FILLER_25_594 ();
 sg13g2_decap_8 FILLER_25_601 ();
 sg13g2_decap_8 FILLER_25_608 ();
 sg13g2_decap_8 FILLER_25_615 ();
 sg13g2_decap_8 FILLER_25_622 ();
 sg13g2_decap_8 FILLER_25_629 ();
 sg13g2_decap_8 FILLER_25_636 ();
 sg13g2_decap_8 FILLER_25_643 ();
 sg13g2_decap_8 FILLER_25_650 ();
 sg13g2_decap_8 FILLER_25_657 ();
 sg13g2_decap_8 FILLER_25_664 ();
 sg13g2_decap_8 FILLER_25_671 ();
 sg13g2_decap_8 FILLER_25_678 ();
 sg13g2_decap_8 FILLER_25_685 ();
 sg13g2_decap_8 FILLER_25_692 ();
 sg13g2_decap_8 FILLER_25_699 ();
 sg13g2_decap_8 FILLER_25_706 ();
 sg13g2_decap_8 FILLER_25_713 ();
 sg13g2_decap_8 FILLER_25_720 ();
 sg13g2_decap_8 FILLER_25_727 ();
 sg13g2_decap_8 FILLER_25_734 ();
 sg13g2_decap_8 FILLER_25_741 ();
 sg13g2_decap_8 FILLER_25_748 ();
 sg13g2_decap_8 FILLER_25_755 ();
 sg13g2_decap_8 FILLER_25_762 ();
 sg13g2_decap_8 FILLER_25_769 ();
 sg13g2_decap_8 FILLER_25_776 ();
 sg13g2_decap_8 FILLER_25_783 ();
 sg13g2_decap_8 FILLER_25_790 ();
 sg13g2_decap_8 FILLER_25_797 ();
 sg13g2_decap_8 FILLER_25_804 ();
 sg13g2_decap_8 FILLER_25_811 ();
 sg13g2_decap_8 FILLER_25_818 ();
 sg13g2_decap_8 FILLER_25_825 ();
 sg13g2_decap_8 FILLER_25_832 ();
 sg13g2_decap_8 FILLER_25_839 ();
 sg13g2_decap_8 FILLER_25_846 ();
 sg13g2_decap_8 FILLER_25_853 ();
 sg13g2_decap_8 FILLER_25_860 ();
 sg13g2_decap_8 FILLER_25_867 ();
 sg13g2_decap_8 FILLER_25_874 ();
 sg13g2_decap_8 FILLER_25_881 ();
 sg13g2_decap_8 FILLER_25_888 ();
 sg13g2_decap_8 FILLER_25_895 ();
 sg13g2_decap_8 FILLER_25_902 ();
 sg13g2_decap_8 FILLER_25_909 ();
 sg13g2_decap_8 FILLER_25_916 ();
 sg13g2_decap_8 FILLER_25_923 ();
 sg13g2_decap_8 FILLER_25_930 ();
 sg13g2_decap_8 FILLER_25_937 ();
 sg13g2_decap_8 FILLER_25_944 ();
 sg13g2_decap_8 FILLER_25_951 ();
 sg13g2_decap_8 FILLER_25_958 ();
 sg13g2_decap_8 FILLER_25_965 ();
 sg13g2_decap_8 FILLER_25_972 ();
 sg13g2_decap_8 FILLER_25_979 ();
 sg13g2_decap_8 FILLER_25_986 ();
 sg13g2_decap_8 FILLER_25_993 ();
 sg13g2_decap_8 FILLER_25_1000 ();
 sg13g2_decap_8 FILLER_25_1007 ();
 sg13g2_decap_8 FILLER_25_1014 ();
 sg13g2_decap_8 FILLER_25_1021 ();
 sg13g2_fill_1 FILLER_25_1028 ();
 sg13g2_decap_8 FILLER_26_4 ();
 sg13g2_decap_8 FILLER_26_11 ();
 sg13g2_decap_8 FILLER_26_18 ();
 sg13g2_decap_8 FILLER_26_25 ();
 sg13g2_decap_8 FILLER_26_32 ();
 sg13g2_decap_8 FILLER_26_39 ();
 sg13g2_decap_4 FILLER_26_46 ();
 sg13g2_fill_1 FILLER_26_50 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_fill_2 FILLER_26_124 ();
 sg13g2_decap_8 FILLER_26_162 ();
 sg13g2_decap_8 FILLER_26_169 ();
 sg13g2_decap_8 FILLER_26_176 ();
 sg13g2_decap_8 FILLER_26_183 ();
 sg13g2_decap_8 FILLER_26_190 ();
 sg13g2_fill_1 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_fill_2 FILLER_26_266 ();
 sg13g2_fill_1 FILLER_26_268 ();
 sg13g2_decap_8 FILLER_26_277 ();
 sg13g2_decap_8 FILLER_26_284 ();
 sg13g2_decap_8 FILLER_26_291 ();
 sg13g2_decap_8 FILLER_26_298 ();
 sg13g2_decap_8 FILLER_26_305 ();
 sg13g2_decap_8 FILLER_26_312 ();
 sg13g2_decap_8 FILLER_26_319 ();
 sg13g2_decap_8 FILLER_26_326 ();
 sg13g2_decap_8 FILLER_26_333 ();
 sg13g2_decap_8 FILLER_26_340 ();
 sg13g2_decap_8 FILLER_26_347 ();
 sg13g2_decap_8 FILLER_26_354 ();
 sg13g2_decap_8 FILLER_26_361 ();
 sg13g2_decap_8 FILLER_26_368 ();
 sg13g2_decap_8 FILLER_26_375 ();
 sg13g2_decap_8 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_decap_8 FILLER_26_419 ();
 sg13g2_decap_8 FILLER_26_426 ();
 sg13g2_decap_8 FILLER_26_433 ();
 sg13g2_decap_8 FILLER_26_440 ();
 sg13g2_decap_8 FILLER_26_447 ();
 sg13g2_fill_2 FILLER_26_454 ();
 sg13g2_decap_8 FILLER_26_483 ();
 sg13g2_decap_8 FILLER_26_490 ();
 sg13g2_decap_8 FILLER_26_497 ();
 sg13g2_decap_8 FILLER_26_504 ();
 sg13g2_decap_8 FILLER_26_511 ();
 sg13g2_decap_8 FILLER_26_518 ();
 sg13g2_decap_8 FILLER_26_525 ();
 sg13g2_decap_8 FILLER_26_532 ();
 sg13g2_fill_1 FILLER_26_539 ();
 sg13g2_decap_8 FILLER_26_544 ();
 sg13g2_decap_8 FILLER_26_551 ();
 sg13g2_decap_8 FILLER_26_558 ();
 sg13g2_decap_8 FILLER_26_565 ();
 sg13g2_decap_8 FILLER_26_572 ();
 sg13g2_decap_8 FILLER_26_579 ();
 sg13g2_decap_8 FILLER_26_586 ();
 sg13g2_decap_8 FILLER_26_593 ();
 sg13g2_decap_8 FILLER_26_600 ();
 sg13g2_decap_8 FILLER_26_607 ();
 sg13g2_decap_8 FILLER_26_614 ();
 sg13g2_decap_8 FILLER_26_621 ();
 sg13g2_decap_8 FILLER_26_628 ();
 sg13g2_decap_8 FILLER_26_635 ();
 sg13g2_decap_8 FILLER_26_642 ();
 sg13g2_decap_8 FILLER_26_649 ();
 sg13g2_decap_8 FILLER_26_656 ();
 sg13g2_decap_8 FILLER_26_663 ();
 sg13g2_decap_8 FILLER_26_670 ();
 sg13g2_decap_8 FILLER_26_677 ();
 sg13g2_decap_8 FILLER_26_684 ();
 sg13g2_decap_8 FILLER_26_691 ();
 sg13g2_decap_8 FILLER_26_698 ();
 sg13g2_decap_8 FILLER_26_705 ();
 sg13g2_decap_8 FILLER_26_712 ();
 sg13g2_decap_8 FILLER_26_719 ();
 sg13g2_decap_8 FILLER_26_726 ();
 sg13g2_decap_8 FILLER_26_733 ();
 sg13g2_decap_8 FILLER_26_740 ();
 sg13g2_decap_8 FILLER_26_747 ();
 sg13g2_decap_8 FILLER_26_754 ();
 sg13g2_decap_8 FILLER_26_761 ();
 sg13g2_decap_8 FILLER_26_768 ();
 sg13g2_decap_8 FILLER_26_775 ();
 sg13g2_decap_8 FILLER_26_782 ();
 sg13g2_decap_8 FILLER_26_789 ();
 sg13g2_decap_8 FILLER_26_796 ();
 sg13g2_decap_8 FILLER_26_803 ();
 sg13g2_decap_8 FILLER_26_810 ();
 sg13g2_decap_8 FILLER_26_817 ();
 sg13g2_decap_8 FILLER_26_824 ();
 sg13g2_decap_8 FILLER_26_831 ();
 sg13g2_decap_8 FILLER_26_838 ();
 sg13g2_decap_8 FILLER_26_845 ();
 sg13g2_decap_8 FILLER_26_852 ();
 sg13g2_decap_8 FILLER_26_859 ();
 sg13g2_decap_8 FILLER_26_866 ();
 sg13g2_decap_8 FILLER_26_873 ();
 sg13g2_decap_8 FILLER_26_880 ();
 sg13g2_decap_8 FILLER_26_887 ();
 sg13g2_decap_8 FILLER_26_894 ();
 sg13g2_decap_8 FILLER_26_901 ();
 sg13g2_decap_8 FILLER_26_908 ();
 sg13g2_decap_8 FILLER_26_915 ();
 sg13g2_decap_8 FILLER_26_922 ();
 sg13g2_decap_8 FILLER_26_929 ();
 sg13g2_decap_8 FILLER_26_936 ();
 sg13g2_decap_8 FILLER_26_943 ();
 sg13g2_decap_8 FILLER_26_950 ();
 sg13g2_decap_8 FILLER_26_957 ();
 sg13g2_decap_8 FILLER_26_964 ();
 sg13g2_decap_8 FILLER_26_971 ();
 sg13g2_decap_8 FILLER_26_978 ();
 sg13g2_decap_8 FILLER_26_985 ();
 sg13g2_decap_8 FILLER_26_992 ();
 sg13g2_decap_8 FILLER_26_999 ();
 sg13g2_decap_8 FILLER_26_1006 ();
 sg13g2_decap_8 FILLER_26_1013 ();
 sg13g2_decap_8 FILLER_26_1020 ();
 sg13g2_fill_2 FILLER_26_1027 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_4 FILLER_27_35 ();
 sg13g2_fill_1 FILLER_27_39 ();
 sg13g2_decap_8 FILLER_27_44 ();
 sg13g2_decap_8 FILLER_27_51 ();
 sg13g2_decap_8 FILLER_27_58 ();
 sg13g2_decap_8 FILLER_27_65 ();
 sg13g2_decap_4 FILLER_27_72 ();
 sg13g2_fill_1 FILLER_27_76 ();
 sg13g2_decap_4 FILLER_27_104 ();
 sg13g2_decap_8 FILLER_27_117 ();
 sg13g2_decap_4 FILLER_27_124 ();
 sg13g2_fill_1 FILLER_27_128 ();
 sg13g2_decap_8 FILLER_27_138 ();
 sg13g2_fill_1 FILLER_27_145 ();
 sg13g2_decap_8 FILLER_27_159 ();
 sg13g2_decap_8 FILLER_27_166 ();
 sg13g2_decap_8 FILLER_27_173 ();
 sg13g2_decap_8 FILLER_27_180 ();
 sg13g2_decap_8 FILLER_27_187 ();
 sg13g2_decap_8 FILLER_27_194 ();
 sg13g2_decap_4 FILLER_27_201 ();
 sg13g2_decap_8 FILLER_27_214 ();
 sg13g2_decap_8 FILLER_27_221 ();
 sg13g2_decap_8 FILLER_27_228 ();
 sg13g2_decap_8 FILLER_27_235 ();
 sg13g2_decap_8 FILLER_27_242 ();
 sg13g2_decap_8 FILLER_27_249 ();
 sg13g2_decap_4 FILLER_27_256 ();
 sg13g2_fill_2 FILLER_27_260 ();
 sg13g2_decap_8 FILLER_27_298 ();
 sg13g2_decap_8 FILLER_27_305 ();
 sg13g2_decap_4 FILLER_27_312 ();
 sg13g2_fill_2 FILLER_27_316 ();
 sg13g2_decap_8 FILLER_27_358 ();
 sg13g2_decap_4 FILLER_27_365 ();
 sg13g2_fill_2 FILLER_27_369 ();
 sg13g2_fill_1 FILLER_27_398 ();
 sg13g2_decap_8 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_27_415 ();
 sg13g2_decap_8 FILLER_27_422 ();
 sg13g2_decap_8 FILLER_27_429 ();
 sg13g2_decap_4 FILLER_27_436 ();
 sg13g2_fill_2 FILLER_27_440 ();
 sg13g2_fill_1 FILLER_27_455 ();
 sg13g2_decap_8 FILLER_27_483 ();
 sg13g2_decap_8 FILLER_27_490 ();
 sg13g2_decap_8 FILLER_27_497 ();
 sg13g2_decap_8 FILLER_27_504 ();
 sg13g2_decap_8 FILLER_27_511 ();
 sg13g2_decap_8 FILLER_27_518 ();
 sg13g2_decap_8 FILLER_27_525 ();
 sg13g2_decap_8 FILLER_27_532 ();
 sg13g2_decap_8 FILLER_27_539 ();
 sg13g2_decap_8 FILLER_27_546 ();
 sg13g2_decap_8 FILLER_27_553 ();
 sg13g2_decap_8 FILLER_27_560 ();
 sg13g2_decap_8 FILLER_27_567 ();
 sg13g2_decap_8 FILLER_27_574 ();
 sg13g2_decap_8 FILLER_27_581 ();
 sg13g2_decap_8 FILLER_27_588 ();
 sg13g2_decap_8 FILLER_27_595 ();
 sg13g2_decap_8 FILLER_27_602 ();
 sg13g2_decap_8 FILLER_27_609 ();
 sg13g2_decap_8 FILLER_27_616 ();
 sg13g2_decap_8 FILLER_27_623 ();
 sg13g2_decap_8 FILLER_27_630 ();
 sg13g2_decap_8 FILLER_27_637 ();
 sg13g2_decap_8 FILLER_27_644 ();
 sg13g2_decap_8 FILLER_27_651 ();
 sg13g2_decap_8 FILLER_27_658 ();
 sg13g2_decap_8 FILLER_27_665 ();
 sg13g2_decap_8 FILLER_27_672 ();
 sg13g2_decap_8 FILLER_27_679 ();
 sg13g2_decap_8 FILLER_27_686 ();
 sg13g2_decap_8 FILLER_27_693 ();
 sg13g2_decap_8 FILLER_27_700 ();
 sg13g2_decap_8 FILLER_27_707 ();
 sg13g2_decap_8 FILLER_27_714 ();
 sg13g2_decap_8 FILLER_27_721 ();
 sg13g2_decap_8 FILLER_27_728 ();
 sg13g2_decap_8 FILLER_27_735 ();
 sg13g2_decap_8 FILLER_27_742 ();
 sg13g2_decap_8 FILLER_27_749 ();
 sg13g2_decap_8 FILLER_27_756 ();
 sg13g2_decap_8 FILLER_27_763 ();
 sg13g2_decap_8 FILLER_27_770 ();
 sg13g2_decap_8 FILLER_27_777 ();
 sg13g2_decap_8 FILLER_27_784 ();
 sg13g2_decap_8 FILLER_27_791 ();
 sg13g2_decap_8 FILLER_27_798 ();
 sg13g2_decap_8 FILLER_27_805 ();
 sg13g2_decap_8 FILLER_27_812 ();
 sg13g2_decap_8 FILLER_27_819 ();
 sg13g2_decap_8 FILLER_27_826 ();
 sg13g2_decap_8 FILLER_27_833 ();
 sg13g2_decap_8 FILLER_27_840 ();
 sg13g2_decap_8 FILLER_27_847 ();
 sg13g2_decap_8 FILLER_27_854 ();
 sg13g2_decap_8 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_27_868 ();
 sg13g2_decap_8 FILLER_27_875 ();
 sg13g2_decap_8 FILLER_27_882 ();
 sg13g2_decap_8 FILLER_27_889 ();
 sg13g2_decap_8 FILLER_27_896 ();
 sg13g2_decap_8 FILLER_27_903 ();
 sg13g2_decap_8 FILLER_27_910 ();
 sg13g2_decap_8 FILLER_27_917 ();
 sg13g2_decap_8 FILLER_27_924 ();
 sg13g2_decap_8 FILLER_27_931 ();
 sg13g2_decap_8 FILLER_27_938 ();
 sg13g2_decap_8 FILLER_27_945 ();
 sg13g2_decap_8 FILLER_27_952 ();
 sg13g2_decap_8 FILLER_27_959 ();
 sg13g2_decap_8 FILLER_27_966 ();
 sg13g2_decap_8 FILLER_27_973 ();
 sg13g2_decap_8 FILLER_27_980 ();
 sg13g2_decap_8 FILLER_27_987 ();
 sg13g2_decap_8 FILLER_27_994 ();
 sg13g2_decap_8 FILLER_27_1001 ();
 sg13g2_decap_8 FILLER_27_1008 ();
 sg13g2_decap_8 FILLER_27_1015 ();
 sg13g2_decap_8 FILLER_27_1022 ();
 sg13g2_fill_2 FILLER_28_4 ();
 sg13g2_decap_8 FILLER_28_60 ();
 sg13g2_decap_8 FILLER_28_67 ();
 sg13g2_decap_8 FILLER_28_74 ();
 sg13g2_decap_4 FILLER_28_81 ();
 sg13g2_fill_2 FILLER_28_85 ();
 sg13g2_decap_8 FILLER_28_100 ();
 sg13g2_decap_8 FILLER_28_107 ();
 sg13g2_decap_8 FILLER_28_114 ();
 sg13g2_decap_8 FILLER_28_121 ();
 sg13g2_decap_8 FILLER_28_128 ();
 sg13g2_decap_8 FILLER_28_162 ();
 sg13g2_decap_8 FILLER_28_169 ();
 sg13g2_decap_8 FILLER_28_176 ();
 sg13g2_decap_8 FILLER_28_183 ();
 sg13g2_decap_8 FILLER_28_190 ();
 sg13g2_decap_8 FILLER_28_197 ();
 sg13g2_decap_8 FILLER_28_204 ();
 sg13g2_decap_4 FILLER_28_211 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_8 FILLER_28_245 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_fill_2 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_288 ();
 sg13g2_decap_8 FILLER_28_295 ();
 sg13g2_decap_8 FILLER_28_302 ();
 sg13g2_decap_8 FILLER_28_309 ();
 sg13g2_decap_8 FILLER_28_316 ();
 sg13g2_decap_8 FILLER_28_323 ();
 sg13g2_decap_8 FILLER_28_330 ();
 sg13g2_fill_2 FILLER_28_337 ();
 sg13g2_fill_1 FILLER_28_339 ();
 sg13g2_decap_4 FILLER_28_344 ();
 sg13g2_fill_2 FILLER_28_348 ();
 sg13g2_decap_8 FILLER_28_364 ();
 sg13g2_decap_8 FILLER_28_371 ();
 sg13g2_decap_8 FILLER_28_378 ();
 sg13g2_decap_8 FILLER_28_385 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_decap_8 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_413 ();
 sg13g2_decap_8 FILLER_28_423 ();
 sg13g2_decap_8 FILLER_28_430 ();
 sg13g2_decap_8 FILLER_28_437 ();
 sg13g2_decap_8 FILLER_28_444 ();
 sg13g2_decap_8 FILLER_28_451 ();
 sg13g2_fill_2 FILLER_28_458 ();
 sg13g2_fill_1 FILLER_28_460 ();
 sg13g2_decap_8 FILLER_28_466 ();
 sg13g2_decap_8 FILLER_28_473 ();
 sg13g2_decap_8 FILLER_28_480 ();
 sg13g2_decap_8 FILLER_28_487 ();
 sg13g2_decap_8 FILLER_28_494 ();
 sg13g2_decap_4 FILLER_28_501 ();
 sg13g2_fill_1 FILLER_28_505 ();
 sg13g2_decap_8 FILLER_28_519 ();
 sg13g2_decap_8 FILLER_28_526 ();
 sg13g2_decap_8 FILLER_28_533 ();
 sg13g2_decap_8 FILLER_28_540 ();
 sg13g2_decap_8 FILLER_28_547 ();
 sg13g2_decap_8 FILLER_28_554 ();
 sg13g2_decap_8 FILLER_28_561 ();
 sg13g2_decap_8 FILLER_28_568 ();
 sg13g2_decap_8 FILLER_28_575 ();
 sg13g2_decap_8 FILLER_28_582 ();
 sg13g2_decap_8 FILLER_28_589 ();
 sg13g2_decap_8 FILLER_28_596 ();
 sg13g2_decap_8 FILLER_28_603 ();
 sg13g2_decap_8 FILLER_28_610 ();
 sg13g2_decap_8 FILLER_28_617 ();
 sg13g2_decap_8 FILLER_28_624 ();
 sg13g2_decap_8 FILLER_28_631 ();
 sg13g2_decap_8 FILLER_28_638 ();
 sg13g2_decap_8 FILLER_28_645 ();
 sg13g2_decap_8 FILLER_28_652 ();
 sg13g2_decap_8 FILLER_28_659 ();
 sg13g2_decap_8 FILLER_28_666 ();
 sg13g2_decap_8 FILLER_28_673 ();
 sg13g2_decap_8 FILLER_28_680 ();
 sg13g2_decap_8 FILLER_28_687 ();
 sg13g2_decap_8 FILLER_28_694 ();
 sg13g2_decap_8 FILLER_28_701 ();
 sg13g2_decap_8 FILLER_28_708 ();
 sg13g2_decap_8 FILLER_28_715 ();
 sg13g2_decap_8 FILLER_28_722 ();
 sg13g2_decap_8 FILLER_28_729 ();
 sg13g2_decap_8 FILLER_28_736 ();
 sg13g2_decap_8 FILLER_28_743 ();
 sg13g2_decap_8 FILLER_28_750 ();
 sg13g2_decap_8 FILLER_28_757 ();
 sg13g2_decap_8 FILLER_28_764 ();
 sg13g2_decap_8 FILLER_28_771 ();
 sg13g2_decap_8 FILLER_28_778 ();
 sg13g2_decap_8 FILLER_28_785 ();
 sg13g2_decap_8 FILLER_28_792 ();
 sg13g2_decap_8 FILLER_28_799 ();
 sg13g2_decap_8 FILLER_28_806 ();
 sg13g2_decap_8 FILLER_28_813 ();
 sg13g2_decap_8 FILLER_28_820 ();
 sg13g2_decap_8 FILLER_28_827 ();
 sg13g2_decap_8 FILLER_28_834 ();
 sg13g2_decap_8 FILLER_28_841 ();
 sg13g2_decap_8 FILLER_28_848 ();
 sg13g2_decap_8 FILLER_28_855 ();
 sg13g2_decap_8 FILLER_28_862 ();
 sg13g2_decap_8 FILLER_28_869 ();
 sg13g2_decap_8 FILLER_28_876 ();
 sg13g2_decap_8 FILLER_28_883 ();
 sg13g2_decap_8 FILLER_28_890 ();
 sg13g2_decap_8 FILLER_28_897 ();
 sg13g2_decap_8 FILLER_28_904 ();
 sg13g2_decap_8 FILLER_28_911 ();
 sg13g2_decap_8 FILLER_28_918 ();
 sg13g2_decap_8 FILLER_28_925 ();
 sg13g2_decap_8 FILLER_28_932 ();
 sg13g2_decap_8 FILLER_28_939 ();
 sg13g2_decap_8 FILLER_28_946 ();
 sg13g2_decap_8 FILLER_28_953 ();
 sg13g2_decap_8 FILLER_28_960 ();
 sg13g2_decap_8 FILLER_28_967 ();
 sg13g2_decap_8 FILLER_28_974 ();
 sg13g2_decap_8 FILLER_28_981 ();
 sg13g2_decap_8 FILLER_28_988 ();
 sg13g2_decap_8 FILLER_28_995 ();
 sg13g2_decap_8 FILLER_28_1002 ();
 sg13g2_decap_8 FILLER_28_1009 ();
 sg13g2_decap_8 FILLER_28_1016 ();
 sg13g2_decap_4 FILLER_28_1023 ();
 sg13g2_fill_2 FILLER_28_1027 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_fill_2 FILLER_29_35 ();
 sg13g2_fill_1 FILLER_29_37 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_fill_1 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_59 ();
 sg13g2_decap_8 FILLER_29_66 ();
 sg13g2_decap_8 FILLER_29_73 ();
 sg13g2_decap_8 FILLER_29_80 ();
 sg13g2_decap_8 FILLER_29_87 ();
 sg13g2_decap_8 FILLER_29_94 ();
 sg13g2_decap_8 FILLER_29_101 ();
 sg13g2_decap_8 FILLER_29_108 ();
 sg13g2_decap_8 FILLER_29_115 ();
 sg13g2_decap_8 FILLER_29_122 ();
 sg13g2_decap_8 FILLER_29_129 ();
 sg13g2_decap_8 FILLER_29_136 ();
 sg13g2_decap_8 FILLER_29_143 ();
 sg13g2_decap_8 FILLER_29_150 ();
 sg13g2_decap_8 FILLER_29_157 ();
 sg13g2_decap_8 FILLER_29_164 ();
 sg13g2_decap_8 FILLER_29_171 ();
 sg13g2_decap_8 FILLER_29_178 ();
 sg13g2_decap_8 FILLER_29_185 ();
 sg13g2_decap_8 FILLER_29_192 ();
 sg13g2_decap_8 FILLER_29_199 ();
 sg13g2_fill_2 FILLER_29_206 ();
 sg13g2_decap_8 FILLER_29_216 ();
 sg13g2_decap_8 FILLER_29_223 ();
 sg13g2_decap_8 FILLER_29_230 ();
 sg13g2_decap_8 FILLER_29_237 ();
 sg13g2_decap_8 FILLER_29_244 ();
 sg13g2_decap_8 FILLER_29_251 ();
 sg13g2_decap_8 FILLER_29_258 ();
 sg13g2_decap_8 FILLER_29_265 ();
 sg13g2_decap_8 FILLER_29_272 ();
 sg13g2_fill_1 FILLER_29_279 ();
 sg13g2_decap_8 FILLER_29_289 ();
 sg13g2_decap_8 FILLER_29_296 ();
 sg13g2_decap_8 FILLER_29_303 ();
 sg13g2_decap_8 FILLER_29_310 ();
 sg13g2_decap_8 FILLER_29_317 ();
 sg13g2_decap_8 FILLER_29_324 ();
 sg13g2_decap_8 FILLER_29_331 ();
 sg13g2_decap_8 FILLER_29_338 ();
 sg13g2_decap_8 FILLER_29_354 ();
 sg13g2_decap_8 FILLER_29_361 ();
 sg13g2_decap_8 FILLER_29_368 ();
 sg13g2_fill_2 FILLER_29_375 ();
 sg13g2_decap_8 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_411 ();
 sg13g2_decap_8 FILLER_29_420 ();
 sg13g2_decap_8 FILLER_29_427 ();
 sg13g2_decap_8 FILLER_29_434 ();
 sg13g2_decap_8 FILLER_29_441 ();
 sg13g2_decap_8 FILLER_29_448 ();
 sg13g2_decap_8 FILLER_29_455 ();
 sg13g2_decap_8 FILLER_29_462 ();
 sg13g2_decap_8 FILLER_29_469 ();
 sg13g2_decap_8 FILLER_29_476 ();
 sg13g2_decap_8 FILLER_29_483 ();
 sg13g2_decap_8 FILLER_29_490 ();
 sg13g2_decap_8 FILLER_29_497 ();
 sg13g2_decap_8 FILLER_29_504 ();
 sg13g2_decap_8 FILLER_29_511 ();
 sg13g2_decap_8 FILLER_29_518 ();
 sg13g2_decap_8 FILLER_29_525 ();
 sg13g2_decap_8 FILLER_29_532 ();
 sg13g2_decap_8 FILLER_29_539 ();
 sg13g2_decap_8 FILLER_29_546 ();
 sg13g2_decap_8 FILLER_29_553 ();
 sg13g2_decap_8 FILLER_29_560 ();
 sg13g2_decap_8 FILLER_29_567 ();
 sg13g2_decap_8 FILLER_29_574 ();
 sg13g2_decap_8 FILLER_29_581 ();
 sg13g2_decap_8 FILLER_29_588 ();
 sg13g2_decap_8 FILLER_29_595 ();
 sg13g2_decap_8 FILLER_29_602 ();
 sg13g2_decap_8 FILLER_29_609 ();
 sg13g2_decap_8 FILLER_29_616 ();
 sg13g2_decap_8 FILLER_29_623 ();
 sg13g2_decap_8 FILLER_29_630 ();
 sg13g2_decap_8 FILLER_29_637 ();
 sg13g2_decap_8 FILLER_29_644 ();
 sg13g2_decap_8 FILLER_29_651 ();
 sg13g2_decap_8 FILLER_29_658 ();
 sg13g2_decap_8 FILLER_29_665 ();
 sg13g2_decap_8 FILLER_29_672 ();
 sg13g2_decap_8 FILLER_29_679 ();
 sg13g2_decap_8 FILLER_29_686 ();
 sg13g2_decap_8 FILLER_29_693 ();
 sg13g2_decap_8 FILLER_29_700 ();
 sg13g2_decap_8 FILLER_29_707 ();
 sg13g2_decap_8 FILLER_29_714 ();
 sg13g2_decap_8 FILLER_29_721 ();
 sg13g2_decap_8 FILLER_29_728 ();
 sg13g2_decap_8 FILLER_29_735 ();
 sg13g2_decap_8 FILLER_29_742 ();
 sg13g2_decap_8 FILLER_29_749 ();
 sg13g2_decap_8 FILLER_29_756 ();
 sg13g2_decap_8 FILLER_29_763 ();
 sg13g2_decap_8 FILLER_29_770 ();
 sg13g2_decap_8 FILLER_29_777 ();
 sg13g2_decap_8 FILLER_29_784 ();
 sg13g2_decap_8 FILLER_29_791 ();
 sg13g2_decap_8 FILLER_29_798 ();
 sg13g2_decap_8 FILLER_29_805 ();
 sg13g2_decap_8 FILLER_29_812 ();
 sg13g2_decap_8 FILLER_29_819 ();
 sg13g2_decap_8 FILLER_29_826 ();
 sg13g2_decap_8 FILLER_29_833 ();
 sg13g2_decap_8 FILLER_29_840 ();
 sg13g2_decap_8 FILLER_29_847 ();
 sg13g2_decap_8 FILLER_29_854 ();
 sg13g2_decap_8 FILLER_29_861 ();
 sg13g2_decap_8 FILLER_29_868 ();
 sg13g2_decap_8 FILLER_29_875 ();
 sg13g2_decap_8 FILLER_29_882 ();
 sg13g2_decap_8 FILLER_29_889 ();
 sg13g2_decap_8 FILLER_29_896 ();
 sg13g2_decap_8 FILLER_29_903 ();
 sg13g2_decap_8 FILLER_29_910 ();
 sg13g2_decap_8 FILLER_29_917 ();
 sg13g2_decap_8 FILLER_29_924 ();
 sg13g2_decap_8 FILLER_29_931 ();
 sg13g2_decap_8 FILLER_29_938 ();
 sg13g2_decap_8 FILLER_29_945 ();
 sg13g2_decap_8 FILLER_29_952 ();
 sg13g2_decap_8 FILLER_29_959 ();
 sg13g2_decap_8 FILLER_29_966 ();
 sg13g2_decap_8 FILLER_29_973 ();
 sg13g2_decap_8 FILLER_29_980 ();
 sg13g2_decap_8 FILLER_29_987 ();
 sg13g2_decap_8 FILLER_29_994 ();
 sg13g2_decap_8 FILLER_29_1001 ();
 sg13g2_decap_8 FILLER_29_1008 ();
 sg13g2_decap_8 FILLER_29_1015 ();
 sg13g2_decap_8 FILLER_29_1022 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_fill_2 FILLER_30_207 ();
 sg13g2_fill_1 FILLER_30_209 ();
 sg13g2_decap_8 FILLER_30_227 ();
 sg13g2_decap_8 FILLER_30_234 ();
 sg13g2_decap_8 FILLER_30_241 ();
 sg13g2_decap_8 FILLER_30_248 ();
 sg13g2_decap_8 FILLER_30_255 ();
 sg13g2_decap_8 FILLER_30_262 ();
 sg13g2_decap_8 FILLER_30_269 ();
 sg13g2_decap_8 FILLER_30_276 ();
 sg13g2_decap_8 FILLER_30_283 ();
 sg13g2_decap_8 FILLER_30_290 ();
 sg13g2_decap_8 FILLER_30_297 ();
 sg13g2_decap_4 FILLER_30_304 ();
 sg13g2_decap_8 FILLER_30_335 ();
 sg13g2_decap_8 FILLER_30_342 ();
 sg13g2_decap_8 FILLER_30_349 ();
 sg13g2_decap_8 FILLER_30_368 ();
 sg13g2_decap_8 FILLER_30_375 ();
 sg13g2_decap_8 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_30_389 ();
 sg13g2_decap_8 FILLER_30_396 ();
 sg13g2_decap_4 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_fill_1 FILLER_30_418 ();
 sg13g2_decap_8 FILLER_30_454 ();
 sg13g2_decap_4 FILLER_30_461 ();
 sg13g2_fill_2 FILLER_30_465 ();
 sg13g2_fill_2 FILLER_30_471 ();
 sg13g2_fill_1 FILLER_30_473 ();
 sg13g2_decap_8 FILLER_30_478 ();
 sg13g2_decap_4 FILLER_30_485 ();
 sg13g2_fill_1 FILLER_30_489 ();
 sg13g2_decap_8 FILLER_30_499 ();
 sg13g2_decap_8 FILLER_30_506 ();
 sg13g2_decap_8 FILLER_30_513 ();
 sg13g2_decap_8 FILLER_30_520 ();
 sg13g2_decap_8 FILLER_30_527 ();
 sg13g2_decap_8 FILLER_30_534 ();
 sg13g2_decap_8 FILLER_30_541 ();
 sg13g2_decap_8 FILLER_30_548 ();
 sg13g2_decap_8 FILLER_30_555 ();
 sg13g2_decap_8 FILLER_30_562 ();
 sg13g2_decap_8 FILLER_30_569 ();
 sg13g2_decap_8 FILLER_30_576 ();
 sg13g2_decap_8 FILLER_30_583 ();
 sg13g2_decap_8 FILLER_30_590 ();
 sg13g2_decap_8 FILLER_30_597 ();
 sg13g2_decap_8 FILLER_30_604 ();
 sg13g2_decap_8 FILLER_30_611 ();
 sg13g2_decap_8 FILLER_30_618 ();
 sg13g2_decap_8 FILLER_30_625 ();
 sg13g2_decap_8 FILLER_30_632 ();
 sg13g2_decap_8 FILLER_30_639 ();
 sg13g2_decap_8 FILLER_30_646 ();
 sg13g2_decap_8 FILLER_30_653 ();
 sg13g2_decap_8 FILLER_30_660 ();
 sg13g2_decap_8 FILLER_30_667 ();
 sg13g2_decap_8 FILLER_30_674 ();
 sg13g2_decap_8 FILLER_30_681 ();
 sg13g2_decap_8 FILLER_30_688 ();
 sg13g2_decap_8 FILLER_30_695 ();
 sg13g2_decap_8 FILLER_30_702 ();
 sg13g2_decap_8 FILLER_30_709 ();
 sg13g2_decap_8 FILLER_30_716 ();
 sg13g2_decap_8 FILLER_30_723 ();
 sg13g2_decap_8 FILLER_30_730 ();
 sg13g2_decap_8 FILLER_30_737 ();
 sg13g2_decap_8 FILLER_30_744 ();
 sg13g2_decap_8 FILLER_30_751 ();
 sg13g2_decap_8 FILLER_30_758 ();
 sg13g2_decap_8 FILLER_30_765 ();
 sg13g2_decap_8 FILLER_30_772 ();
 sg13g2_decap_8 FILLER_30_779 ();
 sg13g2_decap_8 FILLER_30_786 ();
 sg13g2_decap_8 FILLER_30_793 ();
 sg13g2_decap_8 FILLER_30_800 ();
 sg13g2_decap_8 FILLER_30_807 ();
 sg13g2_decap_8 FILLER_30_814 ();
 sg13g2_decap_8 FILLER_30_821 ();
 sg13g2_decap_8 FILLER_30_828 ();
 sg13g2_decap_8 FILLER_30_835 ();
 sg13g2_decap_8 FILLER_30_842 ();
 sg13g2_decap_8 FILLER_30_849 ();
 sg13g2_decap_8 FILLER_30_856 ();
 sg13g2_decap_8 FILLER_30_863 ();
 sg13g2_decap_8 FILLER_30_870 ();
 sg13g2_decap_8 FILLER_30_877 ();
 sg13g2_decap_8 FILLER_30_884 ();
 sg13g2_decap_8 FILLER_30_891 ();
 sg13g2_decap_8 FILLER_30_898 ();
 sg13g2_decap_8 FILLER_30_905 ();
 sg13g2_decap_8 FILLER_30_912 ();
 sg13g2_decap_8 FILLER_30_919 ();
 sg13g2_decap_8 FILLER_30_926 ();
 sg13g2_decap_8 FILLER_30_933 ();
 sg13g2_decap_8 FILLER_30_940 ();
 sg13g2_decap_8 FILLER_30_947 ();
 sg13g2_decap_8 FILLER_30_954 ();
 sg13g2_decap_8 FILLER_30_961 ();
 sg13g2_decap_8 FILLER_30_968 ();
 sg13g2_decap_8 FILLER_30_975 ();
 sg13g2_decap_8 FILLER_30_982 ();
 sg13g2_decap_8 FILLER_30_989 ();
 sg13g2_decap_8 FILLER_30_996 ();
 sg13g2_decap_8 FILLER_30_1003 ();
 sg13g2_decap_8 FILLER_30_1010 ();
 sg13g2_decap_8 FILLER_30_1017 ();
 sg13g2_decap_4 FILLER_30_1024 ();
 sg13g2_fill_1 FILLER_30_1028 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_4 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_129 ();
 sg13g2_decap_8 FILLER_31_136 ();
 sg13g2_decap_8 FILLER_31_143 ();
 sg13g2_fill_2 FILLER_31_150 ();
 sg13g2_decap_8 FILLER_31_173 ();
 sg13g2_decap_8 FILLER_31_180 ();
 sg13g2_decap_8 FILLER_31_187 ();
 sg13g2_decap_8 FILLER_31_194 ();
 sg13g2_decap_8 FILLER_31_201 ();
 sg13g2_fill_2 FILLER_31_208 ();
 sg13g2_fill_1 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_215 ();
 sg13g2_decap_8 FILLER_31_222 ();
 sg13g2_fill_2 FILLER_31_229 ();
 sg13g2_fill_1 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_241 ();
 sg13g2_fill_2 FILLER_31_248 ();
 sg13g2_fill_1 FILLER_31_250 ();
 sg13g2_decap_8 FILLER_31_278 ();
 sg13g2_decap_8 FILLER_31_285 ();
 sg13g2_decap_8 FILLER_31_292 ();
 sg13g2_decap_8 FILLER_31_299 ();
 sg13g2_decap_8 FILLER_31_306 ();
 sg13g2_decap_4 FILLER_31_313 ();
 sg13g2_fill_2 FILLER_31_317 ();
 sg13g2_decap_8 FILLER_31_323 ();
 sg13g2_decap_8 FILLER_31_330 ();
 sg13g2_decap_8 FILLER_31_337 ();
 sg13g2_fill_2 FILLER_31_344 ();
 sg13g2_decap_8 FILLER_31_363 ();
 sg13g2_decap_8 FILLER_31_370 ();
 sg13g2_decap_8 FILLER_31_377 ();
 sg13g2_decap_8 FILLER_31_384 ();
 sg13g2_decap_8 FILLER_31_391 ();
 sg13g2_decap_8 FILLER_31_398 ();
 sg13g2_decap_8 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_31_412 ();
 sg13g2_decap_8 FILLER_31_419 ();
 sg13g2_decap_8 FILLER_31_426 ();
 sg13g2_decap_8 FILLER_31_433 ();
 sg13g2_decap_4 FILLER_31_440 ();
 sg13g2_fill_1 FILLER_31_444 ();
 sg13g2_decap_8 FILLER_31_449 ();
 sg13g2_decap_4 FILLER_31_456 ();
 sg13g2_fill_1 FILLER_31_460 ();
 sg13g2_decap_8 FILLER_31_505 ();
 sg13g2_decap_8 FILLER_31_512 ();
 sg13g2_decap_8 FILLER_31_519 ();
 sg13g2_decap_8 FILLER_31_526 ();
 sg13g2_decap_8 FILLER_31_533 ();
 sg13g2_decap_8 FILLER_31_540 ();
 sg13g2_decap_8 FILLER_31_547 ();
 sg13g2_decap_8 FILLER_31_554 ();
 sg13g2_decap_8 FILLER_31_561 ();
 sg13g2_decap_8 FILLER_31_568 ();
 sg13g2_decap_8 FILLER_31_575 ();
 sg13g2_decap_8 FILLER_31_582 ();
 sg13g2_decap_8 FILLER_31_589 ();
 sg13g2_decap_8 FILLER_31_596 ();
 sg13g2_decap_8 FILLER_31_603 ();
 sg13g2_decap_8 FILLER_31_610 ();
 sg13g2_decap_8 FILLER_31_617 ();
 sg13g2_decap_8 FILLER_31_624 ();
 sg13g2_decap_8 FILLER_31_631 ();
 sg13g2_decap_8 FILLER_31_638 ();
 sg13g2_decap_8 FILLER_31_645 ();
 sg13g2_decap_8 FILLER_31_652 ();
 sg13g2_decap_8 FILLER_31_659 ();
 sg13g2_decap_8 FILLER_31_666 ();
 sg13g2_decap_8 FILLER_31_673 ();
 sg13g2_decap_8 FILLER_31_680 ();
 sg13g2_decap_8 FILLER_31_687 ();
 sg13g2_decap_8 FILLER_31_694 ();
 sg13g2_decap_8 FILLER_31_701 ();
 sg13g2_decap_8 FILLER_31_708 ();
 sg13g2_decap_8 FILLER_31_715 ();
 sg13g2_decap_8 FILLER_31_722 ();
 sg13g2_decap_8 FILLER_31_729 ();
 sg13g2_decap_8 FILLER_31_736 ();
 sg13g2_decap_8 FILLER_31_743 ();
 sg13g2_decap_8 FILLER_31_750 ();
 sg13g2_decap_8 FILLER_31_757 ();
 sg13g2_decap_8 FILLER_31_764 ();
 sg13g2_decap_8 FILLER_31_771 ();
 sg13g2_decap_8 FILLER_31_778 ();
 sg13g2_decap_8 FILLER_31_785 ();
 sg13g2_decap_8 FILLER_31_792 ();
 sg13g2_decap_8 FILLER_31_799 ();
 sg13g2_decap_8 FILLER_31_806 ();
 sg13g2_decap_8 FILLER_31_813 ();
 sg13g2_decap_8 FILLER_31_820 ();
 sg13g2_decap_8 FILLER_31_827 ();
 sg13g2_decap_8 FILLER_31_834 ();
 sg13g2_decap_8 FILLER_31_841 ();
 sg13g2_decap_8 FILLER_31_848 ();
 sg13g2_decap_8 FILLER_31_855 ();
 sg13g2_decap_8 FILLER_31_862 ();
 sg13g2_decap_8 FILLER_31_869 ();
 sg13g2_decap_8 FILLER_31_876 ();
 sg13g2_decap_8 FILLER_31_883 ();
 sg13g2_decap_8 FILLER_31_890 ();
 sg13g2_decap_8 FILLER_31_897 ();
 sg13g2_decap_8 FILLER_31_904 ();
 sg13g2_decap_8 FILLER_31_911 ();
 sg13g2_decap_8 FILLER_31_918 ();
 sg13g2_decap_8 FILLER_31_925 ();
 sg13g2_decap_8 FILLER_31_932 ();
 sg13g2_decap_8 FILLER_31_939 ();
 sg13g2_decap_8 FILLER_31_946 ();
 sg13g2_decap_8 FILLER_31_953 ();
 sg13g2_decap_8 FILLER_31_960 ();
 sg13g2_decap_8 FILLER_31_967 ();
 sg13g2_decap_8 FILLER_31_974 ();
 sg13g2_decap_8 FILLER_31_981 ();
 sg13g2_decap_8 FILLER_31_988 ();
 sg13g2_decap_8 FILLER_31_995 ();
 sg13g2_decap_8 FILLER_31_1002 ();
 sg13g2_decap_8 FILLER_31_1009 ();
 sg13g2_decap_8 FILLER_31_1016 ();
 sg13g2_decap_4 FILLER_31_1023 ();
 sg13g2_fill_2 FILLER_31_1027 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_4 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_45 ();
 sg13g2_fill_2 FILLER_32_52 ();
 sg13g2_decap_8 FILLER_32_67 ();
 sg13g2_decap_8 FILLER_32_74 ();
 sg13g2_decap_8 FILLER_32_81 ();
 sg13g2_decap_8 FILLER_32_88 ();
 sg13g2_decap_8 FILLER_32_95 ();
 sg13g2_decap_8 FILLER_32_102 ();
 sg13g2_fill_2 FILLER_32_109 ();
 sg13g2_fill_1 FILLER_32_111 ();
 sg13g2_decap_8 FILLER_32_139 ();
 sg13g2_decap_8 FILLER_32_146 ();
 sg13g2_decap_8 FILLER_32_153 ();
 sg13g2_decap_4 FILLER_32_160 ();
 sg13g2_decap_8 FILLER_32_172 ();
 sg13g2_decap_8 FILLER_32_179 ();
 sg13g2_decap_8 FILLER_32_186 ();
 sg13g2_decap_8 FILLER_32_193 ();
 sg13g2_decap_8 FILLER_32_200 ();
 sg13g2_decap_8 FILLER_32_207 ();
 sg13g2_decap_4 FILLER_32_214 ();
 sg13g2_fill_2 FILLER_32_218 ();
 sg13g2_decap_8 FILLER_32_228 ();
 sg13g2_decap_8 FILLER_32_235 ();
 sg13g2_fill_2 FILLER_32_242 ();
 sg13g2_fill_1 FILLER_32_244 ();
 sg13g2_decap_8 FILLER_32_258 ();
 sg13g2_decap_8 FILLER_32_265 ();
 sg13g2_decap_8 FILLER_32_272 ();
 sg13g2_decap_8 FILLER_32_279 ();
 sg13g2_decap_4 FILLER_32_286 ();
 sg13g2_fill_1 FILLER_32_290 ();
 sg13g2_decap_8 FILLER_32_304 ();
 sg13g2_decap_8 FILLER_32_311 ();
 sg13g2_decap_8 FILLER_32_318 ();
 sg13g2_decap_8 FILLER_32_325 ();
 sg13g2_decap_8 FILLER_32_332 ();
 sg13g2_decap_8 FILLER_32_339 ();
 sg13g2_decap_8 FILLER_32_346 ();
 sg13g2_decap_8 FILLER_32_353 ();
 sg13g2_decap_8 FILLER_32_360 ();
 sg13g2_decap_8 FILLER_32_367 ();
 sg13g2_decap_8 FILLER_32_374 ();
 sg13g2_decap_8 FILLER_32_381 ();
 sg13g2_decap_8 FILLER_32_388 ();
 sg13g2_decap_8 FILLER_32_395 ();
 sg13g2_decap_8 FILLER_32_402 ();
 sg13g2_decap_8 FILLER_32_409 ();
 sg13g2_decap_8 FILLER_32_416 ();
 sg13g2_decap_8 FILLER_32_423 ();
 sg13g2_decap_8 FILLER_32_430 ();
 sg13g2_decap_8 FILLER_32_437 ();
 sg13g2_decap_8 FILLER_32_444 ();
 sg13g2_decap_8 FILLER_32_451 ();
 sg13g2_decap_4 FILLER_32_458 ();
 sg13g2_fill_2 FILLER_32_462 ();
 sg13g2_decap_8 FILLER_32_491 ();
 sg13g2_decap_8 FILLER_32_498 ();
 sg13g2_decap_8 FILLER_32_505 ();
 sg13g2_decap_8 FILLER_32_512 ();
 sg13g2_decap_8 FILLER_32_519 ();
 sg13g2_decap_8 FILLER_32_526 ();
 sg13g2_decap_8 FILLER_32_533 ();
 sg13g2_decap_8 FILLER_32_540 ();
 sg13g2_decap_8 FILLER_32_547 ();
 sg13g2_decap_8 FILLER_32_554 ();
 sg13g2_decap_8 FILLER_32_561 ();
 sg13g2_decap_8 FILLER_32_568 ();
 sg13g2_decap_8 FILLER_32_575 ();
 sg13g2_decap_8 FILLER_32_582 ();
 sg13g2_decap_8 FILLER_32_589 ();
 sg13g2_decap_8 FILLER_32_596 ();
 sg13g2_decap_8 FILLER_32_603 ();
 sg13g2_decap_8 FILLER_32_610 ();
 sg13g2_decap_8 FILLER_32_617 ();
 sg13g2_decap_8 FILLER_32_624 ();
 sg13g2_decap_8 FILLER_32_631 ();
 sg13g2_decap_8 FILLER_32_638 ();
 sg13g2_decap_8 FILLER_32_645 ();
 sg13g2_decap_8 FILLER_32_652 ();
 sg13g2_decap_8 FILLER_32_659 ();
 sg13g2_decap_8 FILLER_32_666 ();
 sg13g2_decap_8 FILLER_32_673 ();
 sg13g2_decap_8 FILLER_32_680 ();
 sg13g2_decap_8 FILLER_32_687 ();
 sg13g2_decap_8 FILLER_32_694 ();
 sg13g2_decap_8 FILLER_32_701 ();
 sg13g2_decap_8 FILLER_32_708 ();
 sg13g2_decap_8 FILLER_32_715 ();
 sg13g2_decap_8 FILLER_32_722 ();
 sg13g2_decap_8 FILLER_32_729 ();
 sg13g2_decap_8 FILLER_32_736 ();
 sg13g2_decap_8 FILLER_32_743 ();
 sg13g2_decap_8 FILLER_32_750 ();
 sg13g2_decap_8 FILLER_32_757 ();
 sg13g2_decap_8 FILLER_32_764 ();
 sg13g2_decap_8 FILLER_32_771 ();
 sg13g2_decap_8 FILLER_32_778 ();
 sg13g2_decap_8 FILLER_32_785 ();
 sg13g2_decap_8 FILLER_32_792 ();
 sg13g2_decap_8 FILLER_32_799 ();
 sg13g2_decap_8 FILLER_32_806 ();
 sg13g2_decap_8 FILLER_32_813 ();
 sg13g2_decap_8 FILLER_32_820 ();
 sg13g2_decap_8 FILLER_32_827 ();
 sg13g2_decap_8 FILLER_32_834 ();
 sg13g2_decap_8 FILLER_32_841 ();
 sg13g2_decap_8 FILLER_32_848 ();
 sg13g2_decap_8 FILLER_32_855 ();
 sg13g2_decap_8 FILLER_32_862 ();
 sg13g2_decap_8 FILLER_32_869 ();
 sg13g2_decap_8 FILLER_32_876 ();
 sg13g2_decap_8 FILLER_32_883 ();
 sg13g2_decap_8 FILLER_32_890 ();
 sg13g2_decap_8 FILLER_32_897 ();
 sg13g2_decap_8 FILLER_32_904 ();
 sg13g2_decap_8 FILLER_32_911 ();
 sg13g2_decap_8 FILLER_32_918 ();
 sg13g2_decap_8 FILLER_32_925 ();
 sg13g2_decap_8 FILLER_32_932 ();
 sg13g2_decap_8 FILLER_32_939 ();
 sg13g2_decap_8 FILLER_32_946 ();
 sg13g2_decap_8 FILLER_32_953 ();
 sg13g2_decap_8 FILLER_32_960 ();
 sg13g2_decap_8 FILLER_32_967 ();
 sg13g2_decap_8 FILLER_32_974 ();
 sg13g2_decap_8 FILLER_32_981 ();
 sg13g2_decap_8 FILLER_32_988 ();
 sg13g2_decap_8 FILLER_32_995 ();
 sg13g2_decap_8 FILLER_32_1002 ();
 sg13g2_decap_8 FILLER_32_1009 ();
 sg13g2_decap_8 FILLER_32_1016 ();
 sg13g2_decap_4 FILLER_32_1023 ();
 sg13g2_fill_2 FILLER_32_1027 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_4 FILLER_33_14 ();
 sg13g2_fill_1 FILLER_33_18 ();
 sg13g2_decap_8 FILLER_33_46 ();
 sg13g2_decap_8 FILLER_33_53 ();
 sg13g2_decap_8 FILLER_33_60 ();
 sg13g2_decap_4 FILLER_33_94 ();
 sg13g2_decap_8 FILLER_33_142 ();
 sg13g2_decap_8 FILLER_33_149 ();
 sg13g2_decap_8 FILLER_33_156 ();
 sg13g2_decap_8 FILLER_33_163 ();
 sg13g2_decap_8 FILLER_33_170 ();
 sg13g2_fill_2 FILLER_33_177 ();
 sg13g2_fill_2 FILLER_33_215 ();
 sg13g2_fill_1 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_273 ();
 sg13g2_fill_2 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_299 ();
 sg13g2_decap_8 FILLER_33_306 ();
 sg13g2_decap_8 FILLER_33_313 ();
 sg13g2_decap_8 FILLER_33_320 ();
 sg13g2_decap_8 FILLER_33_327 ();
 sg13g2_decap_8 FILLER_33_334 ();
 sg13g2_fill_2 FILLER_33_345 ();
 sg13g2_fill_1 FILLER_33_347 ();
 sg13g2_fill_2 FILLER_33_361 ();
 sg13g2_fill_1 FILLER_33_363 ();
 sg13g2_decap_8 FILLER_33_377 ();
 sg13g2_decap_8 FILLER_33_384 ();
 sg13g2_decap_8 FILLER_33_391 ();
 sg13g2_decap_8 FILLER_33_398 ();
 sg13g2_decap_8 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_33_412 ();
 sg13g2_decap_4 FILLER_33_419 ();
 sg13g2_fill_2 FILLER_33_423 ();
 sg13g2_decap_8 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_33_436 ();
 sg13g2_fill_2 FILLER_33_443 ();
 sg13g2_fill_1 FILLER_33_445 ();
 sg13g2_decap_8 FILLER_33_459 ();
 sg13g2_decap_8 FILLER_33_466 ();
 sg13g2_fill_2 FILLER_33_473 ();
 sg13g2_fill_1 FILLER_33_475 ();
 sg13g2_decap_8 FILLER_33_485 ();
 sg13g2_decap_8 FILLER_33_492 ();
 sg13g2_decap_8 FILLER_33_499 ();
 sg13g2_decap_8 FILLER_33_506 ();
 sg13g2_decap_8 FILLER_33_513 ();
 sg13g2_decap_8 FILLER_33_520 ();
 sg13g2_decap_8 FILLER_33_527 ();
 sg13g2_decap_8 FILLER_33_534 ();
 sg13g2_decap_8 FILLER_33_541 ();
 sg13g2_decap_8 FILLER_33_548 ();
 sg13g2_decap_8 FILLER_33_555 ();
 sg13g2_decap_8 FILLER_33_562 ();
 sg13g2_decap_8 FILLER_33_569 ();
 sg13g2_decap_8 FILLER_33_576 ();
 sg13g2_decap_8 FILLER_33_583 ();
 sg13g2_decap_8 FILLER_33_590 ();
 sg13g2_decap_8 FILLER_33_597 ();
 sg13g2_decap_8 FILLER_33_604 ();
 sg13g2_decap_8 FILLER_33_611 ();
 sg13g2_decap_8 FILLER_33_618 ();
 sg13g2_decap_8 FILLER_33_625 ();
 sg13g2_decap_8 FILLER_33_632 ();
 sg13g2_decap_8 FILLER_33_639 ();
 sg13g2_decap_8 FILLER_33_646 ();
 sg13g2_decap_8 FILLER_33_653 ();
 sg13g2_decap_8 FILLER_33_660 ();
 sg13g2_decap_8 FILLER_33_667 ();
 sg13g2_decap_8 FILLER_33_674 ();
 sg13g2_decap_8 FILLER_33_681 ();
 sg13g2_decap_8 FILLER_33_688 ();
 sg13g2_decap_8 FILLER_33_695 ();
 sg13g2_decap_8 FILLER_33_702 ();
 sg13g2_decap_8 FILLER_33_709 ();
 sg13g2_decap_8 FILLER_33_716 ();
 sg13g2_decap_8 FILLER_33_723 ();
 sg13g2_decap_8 FILLER_33_730 ();
 sg13g2_decap_8 FILLER_33_737 ();
 sg13g2_decap_8 FILLER_33_744 ();
 sg13g2_decap_8 FILLER_33_751 ();
 sg13g2_decap_8 FILLER_33_758 ();
 sg13g2_decap_8 FILLER_33_765 ();
 sg13g2_decap_8 FILLER_33_772 ();
 sg13g2_decap_8 FILLER_33_779 ();
 sg13g2_decap_8 FILLER_33_786 ();
 sg13g2_decap_8 FILLER_33_793 ();
 sg13g2_decap_8 FILLER_33_800 ();
 sg13g2_decap_8 FILLER_33_807 ();
 sg13g2_decap_8 FILLER_33_814 ();
 sg13g2_decap_8 FILLER_33_821 ();
 sg13g2_decap_8 FILLER_33_828 ();
 sg13g2_decap_8 FILLER_33_835 ();
 sg13g2_decap_8 FILLER_33_842 ();
 sg13g2_decap_8 FILLER_33_849 ();
 sg13g2_decap_8 FILLER_33_856 ();
 sg13g2_decap_8 FILLER_33_863 ();
 sg13g2_decap_8 FILLER_33_870 ();
 sg13g2_decap_8 FILLER_33_877 ();
 sg13g2_decap_8 FILLER_33_884 ();
 sg13g2_decap_8 FILLER_33_891 ();
 sg13g2_decap_8 FILLER_33_898 ();
 sg13g2_decap_8 FILLER_33_905 ();
 sg13g2_decap_8 FILLER_33_912 ();
 sg13g2_decap_8 FILLER_33_919 ();
 sg13g2_decap_8 FILLER_33_926 ();
 sg13g2_decap_8 FILLER_33_933 ();
 sg13g2_decap_8 FILLER_33_940 ();
 sg13g2_decap_8 FILLER_33_947 ();
 sg13g2_decap_8 FILLER_33_954 ();
 sg13g2_decap_8 FILLER_33_961 ();
 sg13g2_decap_8 FILLER_33_968 ();
 sg13g2_decap_8 FILLER_33_975 ();
 sg13g2_decap_8 FILLER_33_982 ();
 sg13g2_decap_8 FILLER_33_989 ();
 sg13g2_decap_8 FILLER_33_996 ();
 sg13g2_decap_8 FILLER_33_1003 ();
 sg13g2_decap_8 FILLER_33_1010 ();
 sg13g2_decap_8 FILLER_33_1017 ();
 sg13g2_decap_4 FILLER_33_1024 ();
 sg13g2_fill_1 FILLER_33_1028 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_4 FILLER_34_21 ();
 sg13g2_fill_2 FILLER_34_25 ();
 sg13g2_fill_2 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_55 ();
 sg13g2_decap_8 FILLER_34_62 ();
 sg13g2_decap_8 FILLER_34_69 ();
 sg13g2_decap_8 FILLER_34_76 ();
 sg13g2_decap_8 FILLER_34_83 ();
 sg13g2_decap_8 FILLER_34_90 ();
 sg13g2_fill_2 FILLER_34_97 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_280 ();
 sg13g2_decap_4 FILLER_34_287 ();
 sg13g2_fill_1 FILLER_34_291 ();
 sg13g2_decap_8 FILLER_34_296 ();
 sg13g2_decap_8 FILLER_34_303 ();
 sg13g2_decap_8 FILLER_34_310 ();
 sg13g2_decap_8 FILLER_34_317 ();
 sg13g2_decap_8 FILLER_34_324 ();
 sg13g2_decap_8 FILLER_34_331 ();
 sg13g2_fill_1 FILLER_34_338 ();
 sg13g2_decap_8 FILLER_34_375 ();
 sg13g2_decap_8 FILLER_34_382 ();
 sg13g2_decap_8 FILLER_34_389 ();
 sg13g2_decap_8 FILLER_34_396 ();
 sg13g2_decap_8 FILLER_34_403 ();
 sg13g2_fill_2 FILLER_34_410 ();
 sg13g2_fill_1 FILLER_34_412 ();
 sg13g2_decap_8 FILLER_34_449 ();
 sg13g2_decap_8 FILLER_34_456 ();
 sg13g2_decap_8 FILLER_34_463 ();
 sg13g2_decap_8 FILLER_34_470 ();
 sg13g2_decap_8 FILLER_34_477 ();
 sg13g2_decap_8 FILLER_34_484 ();
 sg13g2_decap_8 FILLER_34_491 ();
 sg13g2_decap_8 FILLER_34_498 ();
 sg13g2_decap_8 FILLER_34_505 ();
 sg13g2_decap_8 FILLER_34_512 ();
 sg13g2_decap_8 FILLER_34_519 ();
 sg13g2_decap_8 FILLER_34_526 ();
 sg13g2_decap_8 FILLER_34_533 ();
 sg13g2_decap_8 FILLER_34_540 ();
 sg13g2_decap_8 FILLER_34_547 ();
 sg13g2_decap_8 FILLER_34_554 ();
 sg13g2_decap_8 FILLER_34_561 ();
 sg13g2_decap_8 FILLER_34_568 ();
 sg13g2_decap_8 FILLER_34_575 ();
 sg13g2_decap_8 FILLER_34_582 ();
 sg13g2_decap_8 FILLER_34_589 ();
 sg13g2_decap_8 FILLER_34_596 ();
 sg13g2_decap_8 FILLER_34_603 ();
 sg13g2_decap_8 FILLER_34_610 ();
 sg13g2_decap_8 FILLER_34_617 ();
 sg13g2_decap_8 FILLER_34_624 ();
 sg13g2_decap_8 FILLER_34_631 ();
 sg13g2_decap_8 FILLER_34_638 ();
 sg13g2_decap_8 FILLER_34_645 ();
 sg13g2_decap_8 FILLER_34_652 ();
 sg13g2_decap_8 FILLER_34_659 ();
 sg13g2_decap_8 FILLER_34_666 ();
 sg13g2_decap_8 FILLER_34_673 ();
 sg13g2_decap_8 FILLER_34_680 ();
 sg13g2_decap_8 FILLER_34_687 ();
 sg13g2_decap_8 FILLER_34_694 ();
 sg13g2_decap_8 FILLER_34_701 ();
 sg13g2_decap_8 FILLER_34_708 ();
 sg13g2_decap_8 FILLER_34_715 ();
 sg13g2_decap_8 FILLER_34_722 ();
 sg13g2_decap_8 FILLER_34_729 ();
 sg13g2_decap_8 FILLER_34_736 ();
 sg13g2_decap_8 FILLER_34_743 ();
 sg13g2_decap_8 FILLER_34_750 ();
 sg13g2_decap_8 FILLER_34_757 ();
 sg13g2_decap_8 FILLER_34_764 ();
 sg13g2_decap_8 FILLER_34_771 ();
 sg13g2_decap_8 FILLER_34_778 ();
 sg13g2_decap_8 FILLER_34_785 ();
 sg13g2_decap_8 FILLER_34_792 ();
 sg13g2_decap_8 FILLER_34_799 ();
 sg13g2_decap_8 FILLER_34_806 ();
 sg13g2_decap_8 FILLER_34_813 ();
 sg13g2_decap_8 FILLER_34_820 ();
 sg13g2_decap_8 FILLER_34_827 ();
 sg13g2_decap_8 FILLER_34_834 ();
 sg13g2_decap_8 FILLER_34_841 ();
 sg13g2_decap_8 FILLER_34_848 ();
 sg13g2_decap_8 FILLER_34_855 ();
 sg13g2_decap_8 FILLER_34_862 ();
 sg13g2_decap_8 FILLER_34_869 ();
 sg13g2_decap_8 FILLER_34_876 ();
 sg13g2_decap_8 FILLER_34_883 ();
 sg13g2_decap_8 FILLER_34_890 ();
 sg13g2_decap_8 FILLER_34_897 ();
 sg13g2_decap_8 FILLER_34_904 ();
 sg13g2_decap_8 FILLER_34_911 ();
 sg13g2_decap_8 FILLER_34_918 ();
 sg13g2_decap_8 FILLER_34_925 ();
 sg13g2_decap_8 FILLER_34_932 ();
 sg13g2_decap_8 FILLER_34_939 ();
 sg13g2_decap_8 FILLER_34_946 ();
 sg13g2_decap_8 FILLER_34_953 ();
 sg13g2_decap_8 FILLER_34_960 ();
 sg13g2_decap_8 FILLER_34_967 ();
 sg13g2_decap_8 FILLER_34_974 ();
 sg13g2_decap_8 FILLER_34_981 ();
 sg13g2_decap_8 FILLER_34_988 ();
 sg13g2_decap_8 FILLER_34_995 ();
 sg13g2_decap_8 FILLER_34_1002 ();
 sg13g2_decap_8 FILLER_34_1009 ();
 sg13g2_decap_8 FILLER_34_1016 ();
 sg13g2_decap_4 FILLER_34_1023 ();
 sg13g2_fill_2 FILLER_34_1027 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_58 ();
 sg13g2_decap_8 FILLER_35_65 ();
 sg13g2_decap_8 FILLER_35_72 ();
 sg13g2_decap_4 FILLER_35_79 ();
 sg13g2_fill_2 FILLER_35_83 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_fill_1 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_123 ();
 sg13g2_decap_8 FILLER_35_130 ();
 sg13g2_decap_8 FILLER_35_137 ();
 sg13g2_decap_8 FILLER_35_144 ();
 sg13g2_decap_8 FILLER_35_151 ();
 sg13g2_decap_8 FILLER_35_158 ();
 sg13g2_decap_8 FILLER_35_165 ();
 sg13g2_decap_8 FILLER_35_172 ();
 sg13g2_decap_8 FILLER_35_179 ();
 sg13g2_decap_8 FILLER_35_186 ();
 sg13g2_decap_8 FILLER_35_193 ();
 sg13g2_decap_8 FILLER_35_200 ();
 sg13g2_decap_8 FILLER_35_207 ();
 sg13g2_decap_8 FILLER_35_214 ();
 sg13g2_decap_8 FILLER_35_221 ();
 sg13g2_decap_8 FILLER_35_228 ();
 sg13g2_decap_8 FILLER_35_235 ();
 sg13g2_decap_8 FILLER_35_242 ();
 sg13g2_decap_8 FILLER_35_249 ();
 sg13g2_decap_8 FILLER_35_256 ();
 sg13g2_fill_2 FILLER_35_263 ();
 sg13g2_fill_1 FILLER_35_265 ();
 sg13g2_decap_8 FILLER_35_302 ();
 sg13g2_decap_8 FILLER_35_309 ();
 sg13g2_decap_8 FILLER_35_316 ();
 sg13g2_decap_8 FILLER_35_323 ();
 sg13g2_fill_2 FILLER_35_330 ();
 sg13g2_decap_8 FILLER_35_359 ();
 sg13g2_decap_8 FILLER_35_366 ();
 sg13g2_decap_8 FILLER_35_373 ();
 sg13g2_decap_8 FILLER_35_380 ();
 sg13g2_decap_4 FILLER_35_387 ();
 sg13g2_fill_2 FILLER_35_391 ();
 sg13g2_decap_8 FILLER_35_421 ();
 sg13g2_decap_8 FILLER_35_428 ();
 sg13g2_decap_8 FILLER_35_435 ();
 sg13g2_decap_8 FILLER_35_442 ();
 sg13g2_decap_8 FILLER_35_449 ();
 sg13g2_decap_8 FILLER_35_456 ();
 sg13g2_decap_8 FILLER_35_463 ();
 sg13g2_decap_8 FILLER_35_470 ();
 sg13g2_decap_8 FILLER_35_477 ();
 sg13g2_decap_8 FILLER_35_484 ();
 sg13g2_decap_8 FILLER_35_491 ();
 sg13g2_decap_8 FILLER_35_498 ();
 sg13g2_decap_8 FILLER_35_505 ();
 sg13g2_decap_8 FILLER_35_512 ();
 sg13g2_decap_8 FILLER_35_519 ();
 sg13g2_decap_8 FILLER_35_526 ();
 sg13g2_decap_8 FILLER_35_533 ();
 sg13g2_decap_8 FILLER_35_540 ();
 sg13g2_decap_8 FILLER_35_547 ();
 sg13g2_decap_8 FILLER_35_554 ();
 sg13g2_decap_8 FILLER_35_561 ();
 sg13g2_decap_8 FILLER_35_568 ();
 sg13g2_decap_8 FILLER_35_575 ();
 sg13g2_decap_8 FILLER_35_582 ();
 sg13g2_decap_8 FILLER_35_589 ();
 sg13g2_decap_8 FILLER_35_596 ();
 sg13g2_decap_8 FILLER_35_603 ();
 sg13g2_decap_8 FILLER_35_610 ();
 sg13g2_decap_8 FILLER_35_617 ();
 sg13g2_decap_8 FILLER_35_624 ();
 sg13g2_decap_8 FILLER_35_631 ();
 sg13g2_decap_8 FILLER_35_638 ();
 sg13g2_decap_8 FILLER_35_645 ();
 sg13g2_decap_8 FILLER_35_652 ();
 sg13g2_decap_8 FILLER_35_659 ();
 sg13g2_decap_8 FILLER_35_666 ();
 sg13g2_decap_8 FILLER_35_673 ();
 sg13g2_decap_8 FILLER_35_680 ();
 sg13g2_decap_8 FILLER_35_687 ();
 sg13g2_decap_8 FILLER_35_694 ();
 sg13g2_decap_8 FILLER_35_701 ();
 sg13g2_decap_8 FILLER_35_708 ();
 sg13g2_decap_8 FILLER_35_715 ();
 sg13g2_decap_8 FILLER_35_722 ();
 sg13g2_decap_8 FILLER_35_729 ();
 sg13g2_decap_8 FILLER_35_736 ();
 sg13g2_decap_8 FILLER_35_743 ();
 sg13g2_decap_8 FILLER_35_750 ();
 sg13g2_decap_8 FILLER_35_757 ();
 sg13g2_decap_8 FILLER_35_764 ();
 sg13g2_decap_8 FILLER_35_771 ();
 sg13g2_decap_8 FILLER_35_778 ();
 sg13g2_decap_8 FILLER_35_785 ();
 sg13g2_decap_8 FILLER_35_792 ();
 sg13g2_decap_8 FILLER_35_799 ();
 sg13g2_decap_8 FILLER_35_806 ();
 sg13g2_decap_8 FILLER_35_813 ();
 sg13g2_decap_8 FILLER_35_820 ();
 sg13g2_decap_8 FILLER_35_827 ();
 sg13g2_decap_8 FILLER_35_834 ();
 sg13g2_decap_8 FILLER_35_841 ();
 sg13g2_decap_8 FILLER_35_848 ();
 sg13g2_decap_8 FILLER_35_855 ();
 sg13g2_decap_8 FILLER_35_862 ();
 sg13g2_decap_8 FILLER_35_869 ();
 sg13g2_decap_8 FILLER_35_876 ();
 sg13g2_decap_8 FILLER_35_883 ();
 sg13g2_decap_8 FILLER_35_890 ();
 sg13g2_decap_8 FILLER_35_897 ();
 sg13g2_decap_8 FILLER_35_904 ();
 sg13g2_decap_8 FILLER_35_911 ();
 sg13g2_decap_8 FILLER_35_918 ();
 sg13g2_decap_8 FILLER_35_925 ();
 sg13g2_decap_8 FILLER_35_932 ();
 sg13g2_decap_8 FILLER_35_939 ();
 sg13g2_decap_8 FILLER_35_946 ();
 sg13g2_decap_8 FILLER_35_953 ();
 sg13g2_decap_8 FILLER_35_960 ();
 sg13g2_decap_8 FILLER_35_967 ();
 sg13g2_decap_8 FILLER_35_974 ();
 sg13g2_decap_8 FILLER_35_981 ();
 sg13g2_decap_8 FILLER_35_988 ();
 sg13g2_decap_8 FILLER_35_995 ();
 sg13g2_decap_8 FILLER_35_1002 ();
 sg13g2_decap_8 FILLER_35_1009 ();
 sg13g2_decap_8 FILLER_35_1016 ();
 sg13g2_decap_4 FILLER_35_1023 ();
 sg13g2_fill_2 FILLER_35_1027 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_fill_1 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_166 ();
 sg13g2_decap_8 FILLER_36_173 ();
 sg13g2_decap_8 FILLER_36_180 ();
 sg13g2_decap_8 FILLER_36_187 ();
 sg13g2_decap_8 FILLER_36_211 ();
 sg13g2_decap_8 FILLER_36_218 ();
 sg13g2_decap_8 FILLER_36_225 ();
 sg13g2_decap_8 FILLER_36_232 ();
 sg13g2_decap_8 FILLER_36_239 ();
 sg13g2_decap_8 FILLER_36_246 ();
 sg13g2_decap_8 FILLER_36_253 ();
 sg13g2_decap_8 FILLER_36_260 ();
 sg13g2_fill_2 FILLER_36_267 ();
 sg13g2_decap_8 FILLER_36_278 ();
 sg13g2_decap_8 FILLER_36_285 ();
 sg13g2_fill_1 FILLER_36_292 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_decap_8 FILLER_36_315 ();
 sg13g2_decap_8 FILLER_36_322 ();
 sg13g2_decap_4 FILLER_36_329 ();
 sg13g2_fill_2 FILLER_36_333 ();
 sg13g2_decap_8 FILLER_36_348 ();
 sg13g2_decap_8 FILLER_36_355 ();
 sg13g2_decap_8 FILLER_36_362 ();
 sg13g2_decap_8 FILLER_36_369 ();
 sg13g2_decap_8 FILLER_36_376 ();
 sg13g2_decap_8 FILLER_36_383 ();
 sg13g2_decap_8 FILLER_36_390 ();
 sg13g2_decap_8 FILLER_36_397 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_2 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_36_423 ();
 sg13g2_decap_8 FILLER_36_430 ();
 sg13g2_decap_8 FILLER_36_437 ();
 sg13g2_decap_8 FILLER_36_444 ();
 sg13g2_decap_4 FILLER_36_451 ();
 sg13g2_fill_2 FILLER_36_455 ();
 sg13g2_decap_8 FILLER_36_484 ();
 sg13g2_decap_8 FILLER_36_491 ();
 sg13g2_decap_8 FILLER_36_498 ();
 sg13g2_decap_8 FILLER_36_505 ();
 sg13g2_decap_8 FILLER_36_512 ();
 sg13g2_decap_8 FILLER_36_519 ();
 sg13g2_decap_8 FILLER_36_526 ();
 sg13g2_decap_8 FILLER_36_533 ();
 sg13g2_decap_8 FILLER_36_540 ();
 sg13g2_decap_8 FILLER_36_547 ();
 sg13g2_decap_8 FILLER_36_554 ();
 sg13g2_decap_8 FILLER_36_561 ();
 sg13g2_decap_8 FILLER_36_568 ();
 sg13g2_decap_8 FILLER_36_575 ();
 sg13g2_decap_8 FILLER_36_582 ();
 sg13g2_decap_8 FILLER_36_589 ();
 sg13g2_decap_8 FILLER_36_596 ();
 sg13g2_decap_8 FILLER_36_603 ();
 sg13g2_decap_8 FILLER_36_610 ();
 sg13g2_decap_8 FILLER_36_617 ();
 sg13g2_decap_8 FILLER_36_624 ();
 sg13g2_decap_8 FILLER_36_631 ();
 sg13g2_decap_8 FILLER_36_638 ();
 sg13g2_decap_8 FILLER_36_645 ();
 sg13g2_decap_8 FILLER_36_652 ();
 sg13g2_decap_8 FILLER_36_659 ();
 sg13g2_decap_8 FILLER_36_666 ();
 sg13g2_decap_8 FILLER_36_673 ();
 sg13g2_decap_8 FILLER_36_680 ();
 sg13g2_decap_8 FILLER_36_687 ();
 sg13g2_decap_8 FILLER_36_694 ();
 sg13g2_decap_8 FILLER_36_701 ();
 sg13g2_decap_8 FILLER_36_708 ();
 sg13g2_decap_8 FILLER_36_715 ();
 sg13g2_decap_8 FILLER_36_722 ();
 sg13g2_decap_8 FILLER_36_729 ();
 sg13g2_decap_8 FILLER_36_736 ();
 sg13g2_decap_8 FILLER_36_743 ();
 sg13g2_decap_8 FILLER_36_750 ();
 sg13g2_decap_8 FILLER_36_757 ();
 sg13g2_decap_8 FILLER_36_764 ();
 sg13g2_decap_8 FILLER_36_771 ();
 sg13g2_decap_8 FILLER_36_778 ();
 sg13g2_decap_8 FILLER_36_785 ();
 sg13g2_decap_8 FILLER_36_792 ();
 sg13g2_decap_8 FILLER_36_799 ();
 sg13g2_decap_8 FILLER_36_806 ();
 sg13g2_decap_8 FILLER_36_813 ();
 sg13g2_decap_8 FILLER_36_820 ();
 sg13g2_decap_8 FILLER_36_827 ();
 sg13g2_decap_8 FILLER_36_834 ();
 sg13g2_decap_8 FILLER_36_841 ();
 sg13g2_decap_8 FILLER_36_848 ();
 sg13g2_decap_8 FILLER_36_855 ();
 sg13g2_decap_8 FILLER_36_862 ();
 sg13g2_decap_8 FILLER_36_869 ();
 sg13g2_decap_8 FILLER_36_876 ();
 sg13g2_decap_8 FILLER_36_883 ();
 sg13g2_decap_8 FILLER_36_890 ();
 sg13g2_decap_8 FILLER_36_897 ();
 sg13g2_decap_8 FILLER_36_904 ();
 sg13g2_decap_8 FILLER_36_911 ();
 sg13g2_decap_8 FILLER_36_918 ();
 sg13g2_decap_8 FILLER_36_925 ();
 sg13g2_decap_8 FILLER_36_932 ();
 sg13g2_decap_8 FILLER_36_939 ();
 sg13g2_decap_8 FILLER_36_946 ();
 sg13g2_decap_8 FILLER_36_953 ();
 sg13g2_decap_8 FILLER_36_960 ();
 sg13g2_decap_8 FILLER_36_967 ();
 sg13g2_decap_8 FILLER_36_974 ();
 sg13g2_decap_8 FILLER_36_981 ();
 sg13g2_decap_8 FILLER_36_988 ();
 sg13g2_decap_8 FILLER_36_995 ();
 sg13g2_decap_8 FILLER_36_1002 ();
 sg13g2_decap_8 FILLER_36_1009 ();
 sg13g2_decap_8 FILLER_36_1016 ();
 sg13g2_decap_4 FILLER_36_1023 ();
 sg13g2_fill_2 FILLER_36_1027 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_fill_1 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_4 FILLER_37_70 ();
 sg13g2_fill_1 FILLER_37_74 ();
 sg13g2_decap_8 FILLER_37_102 ();
 sg13g2_fill_1 FILLER_37_109 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_fill_2 FILLER_37_147 ();
 sg13g2_fill_1 FILLER_37_149 ();
 sg13g2_decap_8 FILLER_37_181 ();
 sg13g2_decap_8 FILLER_37_188 ();
 sg13g2_decap_8 FILLER_37_195 ();
 sg13g2_decap_8 FILLER_37_202 ();
 sg13g2_decap_8 FILLER_37_209 ();
 sg13g2_decap_8 FILLER_37_216 ();
 sg13g2_fill_1 FILLER_37_223 ();
 sg13g2_decap_8 FILLER_37_237 ();
 sg13g2_decap_8 FILLER_37_244 ();
 sg13g2_decap_8 FILLER_37_251 ();
 sg13g2_decap_8 FILLER_37_258 ();
 sg13g2_decap_8 FILLER_37_274 ();
 sg13g2_decap_8 FILLER_37_281 ();
 sg13g2_decap_8 FILLER_37_288 ();
 sg13g2_decap_8 FILLER_37_295 ();
 sg13g2_fill_2 FILLER_37_302 ();
 sg13g2_fill_1 FILLER_37_304 ();
 sg13g2_decap_8 FILLER_37_314 ();
 sg13g2_decap_8 FILLER_37_321 ();
 sg13g2_decap_8 FILLER_37_328 ();
 sg13g2_decap_8 FILLER_37_335 ();
 sg13g2_decap_8 FILLER_37_342 ();
 sg13g2_decap_8 FILLER_37_349 ();
 sg13g2_decap_8 FILLER_37_356 ();
 sg13g2_decap_8 FILLER_37_363 ();
 sg13g2_decap_8 FILLER_37_370 ();
 sg13g2_decap_8 FILLER_37_377 ();
 sg13g2_decap_8 FILLER_37_384 ();
 sg13g2_decap_8 FILLER_37_391 ();
 sg13g2_decap_8 FILLER_37_398 ();
 sg13g2_fill_2 FILLER_37_405 ();
 sg13g2_fill_1 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_37_421 ();
 sg13g2_decap_8 FILLER_37_428 ();
 sg13g2_decap_8 FILLER_37_435 ();
 sg13g2_decap_8 FILLER_37_442 ();
 sg13g2_decap_8 FILLER_37_449 ();
 sg13g2_decap_8 FILLER_37_469 ();
 sg13g2_decap_8 FILLER_37_476 ();
 sg13g2_decap_8 FILLER_37_483 ();
 sg13g2_decap_8 FILLER_37_490 ();
 sg13g2_decap_8 FILLER_37_497 ();
 sg13g2_decap_8 FILLER_37_504 ();
 sg13g2_decap_8 FILLER_37_511 ();
 sg13g2_decap_8 FILLER_37_518 ();
 sg13g2_decap_8 FILLER_37_525 ();
 sg13g2_decap_8 FILLER_37_532 ();
 sg13g2_decap_8 FILLER_37_539 ();
 sg13g2_decap_8 FILLER_37_546 ();
 sg13g2_decap_8 FILLER_37_553 ();
 sg13g2_decap_8 FILLER_37_560 ();
 sg13g2_decap_8 FILLER_37_567 ();
 sg13g2_decap_8 FILLER_37_574 ();
 sg13g2_decap_8 FILLER_37_581 ();
 sg13g2_decap_8 FILLER_37_588 ();
 sg13g2_decap_8 FILLER_37_595 ();
 sg13g2_decap_8 FILLER_37_602 ();
 sg13g2_decap_8 FILLER_37_609 ();
 sg13g2_decap_8 FILLER_37_616 ();
 sg13g2_decap_8 FILLER_37_623 ();
 sg13g2_decap_8 FILLER_37_630 ();
 sg13g2_decap_8 FILLER_37_637 ();
 sg13g2_decap_8 FILLER_37_644 ();
 sg13g2_decap_8 FILLER_37_651 ();
 sg13g2_decap_8 FILLER_37_658 ();
 sg13g2_decap_8 FILLER_37_665 ();
 sg13g2_decap_8 FILLER_37_672 ();
 sg13g2_decap_8 FILLER_37_679 ();
 sg13g2_decap_8 FILLER_37_686 ();
 sg13g2_decap_8 FILLER_37_693 ();
 sg13g2_decap_8 FILLER_37_700 ();
 sg13g2_decap_8 FILLER_37_707 ();
 sg13g2_decap_8 FILLER_37_714 ();
 sg13g2_decap_8 FILLER_37_721 ();
 sg13g2_decap_8 FILLER_37_728 ();
 sg13g2_decap_8 FILLER_37_735 ();
 sg13g2_decap_8 FILLER_37_742 ();
 sg13g2_decap_8 FILLER_37_749 ();
 sg13g2_decap_8 FILLER_37_756 ();
 sg13g2_decap_8 FILLER_37_763 ();
 sg13g2_decap_8 FILLER_37_770 ();
 sg13g2_decap_8 FILLER_37_777 ();
 sg13g2_decap_8 FILLER_37_784 ();
 sg13g2_decap_8 FILLER_37_791 ();
 sg13g2_decap_8 FILLER_37_798 ();
 sg13g2_decap_8 FILLER_37_805 ();
 sg13g2_decap_8 FILLER_37_812 ();
 sg13g2_decap_8 FILLER_37_819 ();
 sg13g2_decap_8 FILLER_37_826 ();
 sg13g2_decap_8 FILLER_37_833 ();
 sg13g2_decap_8 FILLER_37_840 ();
 sg13g2_decap_8 FILLER_37_847 ();
 sg13g2_decap_8 FILLER_37_854 ();
 sg13g2_decap_8 FILLER_37_861 ();
 sg13g2_decap_8 FILLER_37_868 ();
 sg13g2_decap_8 FILLER_37_875 ();
 sg13g2_decap_8 FILLER_37_882 ();
 sg13g2_decap_8 FILLER_37_889 ();
 sg13g2_decap_8 FILLER_37_896 ();
 sg13g2_decap_8 FILLER_37_903 ();
 sg13g2_decap_8 FILLER_37_910 ();
 sg13g2_decap_8 FILLER_37_917 ();
 sg13g2_decap_8 FILLER_37_924 ();
 sg13g2_decap_8 FILLER_37_931 ();
 sg13g2_decap_8 FILLER_37_938 ();
 sg13g2_decap_8 FILLER_37_945 ();
 sg13g2_decap_8 FILLER_37_952 ();
 sg13g2_decap_8 FILLER_37_959 ();
 sg13g2_decap_8 FILLER_37_966 ();
 sg13g2_decap_8 FILLER_37_973 ();
 sg13g2_decap_8 FILLER_37_980 ();
 sg13g2_decap_8 FILLER_37_987 ();
 sg13g2_decap_8 FILLER_37_994 ();
 sg13g2_decap_8 FILLER_37_1001 ();
 sg13g2_decap_8 FILLER_37_1008 ();
 sg13g2_decap_8 FILLER_37_1015 ();
 sg13g2_decap_8 FILLER_37_1022 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_fill_2 FILLER_38_28 ();
 sg13g2_fill_2 FILLER_38_38 ();
 sg13g2_fill_1 FILLER_38_40 ();
 sg13g2_decap_8 FILLER_38_50 ();
 sg13g2_decap_8 FILLER_38_57 ();
 sg13g2_decap_8 FILLER_38_64 ();
 sg13g2_decap_8 FILLER_38_71 ();
 sg13g2_decap_8 FILLER_38_78 ();
 sg13g2_decap_4 FILLER_38_85 ();
 sg13g2_fill_1 FILLER_38_102 ();
 sg13g2_decap_8 FILLER_38_111 ();
 sg13g2_decap_8 FILLER_38_118 ();
 sg13g2_decap_8 FILLER_38_125 ();
 sg13g2_decap_8 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_139 ();
 sg13g2_fill_2 FILLER_38_170 ();
 sg13g2_fill_1 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_237 ();
 sg13g2_decap_8 FILLER_38_244 ();
 sg13g2_decap_4 FILLER_38_251 ();
 sg13g2_fill_2 FILLER_38_255 ();
 sg13g2_fill_1 FILLER_38_305 ();
 sg13g2_decap_8 FILLER_38_314 ();
 sg13g2_decap_8 FILLER_38_321 ();
 sg13g2_decap_8 FILLER_38_328 ();
 sg13g2_decap_8 FILLER_38_335 ();
 sg13g2_decap_8 FILLER_38_342 ();
 sg13g2_decap_8 FILLER_38_349 ();
 sg13g2_decap_8 FILLER_38_356 ();
 sg13g2_decap_8 FILLER_38_363 ();
 sg13g2_decap_8 FILLER_38_370 ();
 sg13g2_decap_8 FILLER_38_377 ();
 sg13g2_decap_8 FILLER_38_384 ();
 sg13g2_decap_8 FILLER_38_391 ();
 sg13g2_decap_8 FILLER_38_398 ();
 sg13g2_fill_1 FILLER_38_405 ();
 sg13g2_decap_8 FILLER_38_415 ();
 sg13g2_decap_8 FILLER_38_422 ();
 sg13g2_decap_8 FILLER_38_429 ();
 sg13g2_decap_8 FILLER_38_436 ();
 sg13g2_decap_8 FILLER_38_443 ();
 sg13g2_decap_8 FILLER_38_450 ();
 sg13g2_decap_4 FILLER_38_477 ();
 sg13g2_fill_1 FILLER_38_481 ();
 sg13g2_decap_8 FILLER_38_509 ();
 sg13g2_decap_8 FILLER_38_516 ();
 sg13g2_decap_8 FILLER_38_523 ();
 sg13g2_decap_8 FILLER_38_530 ();
 sg13g2_decap_8 FILLER_38_537 ();
 sg13g2_decap_8 FILLER_38_544 ();
 sg13g2_decap_8 FILLER_38_551 ();
 sg13g2_decap_8 FILLER_38_558 ();
 sg13g2_decap_8 FILLER_38_565 ();
 sg13g2_decap_8 FILLER_38_572 ();
 sg13g2_decap_8 FILLER_38_579 ();
 sg13g2_decap_8 FILLER_38_586 ();
 sg13g2_decap_8 FILLER_38_593 ();
 sg13g2_decap_8 FILLER_38_600 ();
 sg13g2_decap_8 FILLER_38_607 ();
 sg13g2_decap_8 FILLER_38_614 ();
 sg13g2_decap_8 FILLER_38_621 ();
 sg13g2_decap_8 FILLER_38_628 ();
 sg13g2_decap_8 FILLER_38_635 ();
 sg13g2_decap_8 FILLER_38_642 ();
 sg13g2_decap_8 FILLER_38_649 ();
 sg13g2_decap_8 FILLER_38_656 ();
 sg13g2_decap_8 FILLER_38_663 ();
 sg13g2_decap_8 FILLER_38_670 ();
 sg13g2_decap_8 FILLER_38_677 ();
 sg13g2_decap_8 FILLER_38_684 ();
 sg13g2_decap_8 FILLER_38_691 ();
 sg13g2_decap_8 FILLER_38_698 ();
 sg13g2_decap_8 FILLER_38_705 ();
 sg13g2_decap_8 FILLER_38_712 ();
 sg13g2_decap_8 FILLER_38_719 ();
 sg13g2_decap_8 FILLER_38_726 ();
 sg13g2_decap_8 FILLER_38_733 ();
 sg13g2_decap_8 FILLER_38_740 ();
 sg13g2_decap_8 FILLER_38_747 ();
 sg13g2_decap_8 FILLER_38_754 ();
 sg13g2_decap_8 FILLER_38_761 ();
 sg13g2_decap_8 FILLER_38_768 ();
 sg13g2_decap_8 FILLER_38_775 ();
 sg13g2_decap_8 FILLER_38_782 ();
 sg13g2_decap_8 FILLER_38_789 ();
 sg13g2_decap_8 FILLER_38_796 ();
 sg13g2_decap_8 FILLER_38_803 ();
 sg13g2_decap_8 FILLER_38_810 ();
 sg13g2_decap_8 FILLER_38_817 ();
 sg13g2_decap_8 FILLER_38_824 ();
 sg13g2_decap_8 FILLER_38_831 ();
 sg13g2_decap_8 FILLER_38_838 ();
 sg13g2_decap_8 FILLER_38_845 ();
 sg13g2_decap_8 FILLER_38_852 ();
 sg13g2_decap_8 FILLER_38_859 ();
 sg13g2_decap_8 FILLER_38_866 ();
 sg13g2_decap_8 FILLER_38_873 ();
 sg13g2_decap_8 FILLER_38_880 ();
 sg13g2_decap_8 FILLER_38_887 ();
 sg13g2_decap_8 FILLER_38_894 ();
 sg13g2_decap_8 FILLER_38_901 ();
 sg13g2_decap_8 FILLER_38_908 ();
 sg13g2_decap_8 FILLER_38_915 ();
 sg13g2_decap_8 FILLER_38_922 ();
 sg13g2_decap_8 FILLER_38_929 ();
 sg13g2_decap_8 FILLER_38_936 ();
 sg13g2_decap_8 FILLER_38_943 ();
 sg13g2_decap_8 FILLER_38_950 ();
 sg13g2_decap_8 FILLER_38_957 ();
 sg13g2_decap_8 FILLER_38_964 ();
 sg13g2_decap_8 FILLER_38_971 ();
 sg13g2_decap_8 FILLER_38_978 ();
 sg13g2_decap_8 FILLER_38_985 ();
 sg13g2_decap_8 FILLER_38_992 ();
 sg13g2_decap_8 FILLER_38_999 ();
 sg13g2_decap_8 FILLER_38_1006 ();
 sg13g2_decap_8 FILLER_38_1013 ();
 sg13g2_decap_8 FILLER_38_1020 ();
 sg13g2_fill_2 FILLER_38_1027 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_fill_2 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_59 ();
 sg13g2_decap_8 FILLER_39_66 ();
 sg13g2_decap_8 FILLER_39_73 ();
 sg13g2_decap_8 FILLER_39_80 ();
 sg13g2_decap_8 FILLER_39_87 ();
 sg13g2_decap_8 FILLER_39_94 ();
 sg13g2_decap_8 FILLER_39_101 ();
 sg13g2_decap_8 FILLER_39_108 ();
 sg13g2_decap_8 FILLER_39_115 ();
 sg13g2_decap_8 FILLER_39_122 ();
 sg13g2_decap_8 FILLER_39_129 ();
 sg13g2_decap_8 FILLER_39_136 ();
 sg13g2_decap_8 FILLER_39_143 ();
 sg13g2_fill_2 FILLER_39_150 ();
 sg13g2_decap_4 FILLER_39_156 ();
 sg13g2_fill_2 FILLER_39_160 ();
 sg13g2_decap_8 FILLER_39_188 ();
 sg13g2_decap_8 FILLER_39_195 ();
 sg13g2_fill_1 FILLER_39_202 ();
 sg13g2_decap_8 FILLER_39_230 ();
 sg13g2_decap_8 FILLER_39_237 ();
 sg13g2_fill_2 FILLER_39_244 ();
 sg13g2_decap_4 FILLER_39_267 ();
 sg13g2_fill_1 FILLER_39_271 ();
 sg13g2_decap_8 FILLER_39_281 ();
 sg13g2_decap_8 FILLER_39_288 ();
 sg13g2_decap_8 FILLER_39_295 ();
 sg13g2_decap_8 FILLER_39_302 ();
 sg13g2_fill_1 FILLER_39_309 ();
 sg13g2_decap_8 FILLER_39_337 ();
 sg13g2_decap_4 FILLER_39_344 ();
 sg13g2_fill_1 FILLER_39_348 ();
 sg13g2_fill_2 FILLER_39_362 ();
 sg13g2_fill_1 FILLER_39_364 ();
 sg13g2_decap_8 FILLER_39_395 ();
 sg13g2_fill_2 FILLER_39_402 ();
 sg13g2_decap_8 FILLER_39_431 ();
 sg13g2_decap_8 FILLER_39_438 ();
 sg13g2_decap_8 FILLER_39_445 ();
 sg13g2_decap_8 FILLER_39_452 ();
 sg13g2_fill_2 FILLER_39_459 ();
 sg13g2_fill_1 FILLER_39_461 ();
 sg13g2_decap_8 FILLER_39_470 ();
 sg13g2_decap_4 FILLER_39_481 ();
 sg13g2_fill_1 FILLER_39_485 ();
 sg13g2_decap_8 FILLER_39_490 ();
 sg13g2_fill_2 FILLER_39_497 ();
 sg13g2_decap_8 FILLER_39_508 ();
 sg13g2_decap_8 FILLER_39_515 ();
 sg13g2_decap_8 FILLER_39_522 ();
 sg13g2_decap_8 FILLER_39_529 ();
 sg13g2_decap_8 FILLER_39_536 ();
 sg13g2_decap_8 FILLER_39_543 ();
 sg13g2_decap_8 FILLER_39_550 ();
 sg13g2_decap_8 FILLER_39_557 ();
 sg13g2_decap_8 FILLER_39_564 ();
 sg13g2_decap_8 FILLER_39_571 ();
 sg13g2_decap_8 FILLER_39_578 ();
 sg13g2_decap_8 FILLER_39_585 ();
 sg13g2_decap_8 FILLER_39_592 ();
 sg13g2_decap_8 FILLER_39_599 ();
 sg13g2_decap_8 FILLER_39_606 ();
 sg13g2_decap_8 FILLER_39_613 ();
 sg13g2_decap_8 FILLER_39_620 ();
 sg13g2_decap_8 FILLER_39_627 ();
 sg13g2_decap_8 FILLER_39_634 ();
 sg13g2_decap_8 FILLER_39_641 ();
 sg13g2_decap_8 FILLER_39_648 ();
 sg13g2_decap_8 FILLER_39_655 ();
 sg13g2_decap_8 FILLER_39_662 ();
 sg13g2_decap_8 FILLER_39_669 ();
 sg13g2_decap_8 FILLER_39_676 ();
 sg13g2_decap_8 FILLER_39_683 ();
 sg13g2_decap_8 FILLER_39_690 ();
 sg13g2_decap_8 FILLER_39_697 ();
 sg13g2_decap_8 FILLER_39_704 ();
 sg13g2_decap_8 FILLER_39_711 ();
 sg13g2_decap_8 FILLER_39_718 ();
 sg13g2_decap_8 FILLER_39_725 ();
 sg13g2_decap_8 FILLER_39_732 ();
 sg13g2_decap_8 FILLER_39_739 ();
 sg13g2_decap_8 FILLER_39_746 ();
 sg13g2_decap_8 FILLER_39_753 ();
 sg13g2_decap_8 FILLER_39_760 ();
 sg13g2_decap_8 FILLER_39_767 ();
 sg13g2_decap_8 FILLER_39_774 ();
 sg13g2_decap_8 FILLER_39_781 ();
 sg13g2_decap_8 FILLER_39_788 ();
 sg13g2_decap_8 FILLER_39_795 ();
 sg13g2_decap_8 FILLER_39_802 ();
 sg13g2_decap_8 FILLER_39_809 ();
 sg13g2_decap_8 FILLER_39_816 ();
 sg13g2_decap_8 FILLER_39_823 ();
 sg13g2_decap_8 FILLER_39_830 ();
 sg13g2_decap_8 FILLER_39_837 ();
 sg13g2_decap_8 FILLER_39_844 ();
 sg13g2_decap_8 FILLER_39_851 ();
 sg13g2_decap_8 FILLER_39_858 ();
 sg13g2_decap_8 FILLER_39_865 ();
 sg13g2_decap_8 FILLER_39_872 ();
 sg13g2_decap_8 FILLER_39_879 ();
 sg13g2_decap_8 FILLER_39_886 ();
 sg13g2_decap_8 FILLER_39_893 ();
 sg13g2_decap_8 FILLER_39_900 ();
 sg13g2_decap_8 FILLER_39_907 ();
 sg13g2_decap_8 FILLER_39_914 ();
 sg13g2_decap_8 FILLER_39_921 ();
 sg13g2_decap_8 FILLER_39_928 ();
 sg13g2_decap_8 FILLER_39_935 ();
 sg13g2_decap_8 FILLER_39_942 ();
 sg13g2_decap_8 FILLER_39_949 ();
 sg13g2_decap_8 FILLER_39_956 ();
 sg13g2_decap_8 FILLER_39_963 ();
 sg13g2_decap_8 FILLER_39_970 ();
 sg13g2_decap_8 FILLER_39_977 ();
 sg13g2_decap_8 FILLER_39_984 ();
 sg13g2_decap_8 FILLER_39_991 ();
 sg13g2_decap_8 FILLER_39_998 ();
 sg13g2_decap_8 FILLER_39_1005 ();
 sg13g2_decap_8 FILLER_39_1012 ();
 sg13g2_decap_8 FILLER_39_1019 ();
 sg13g2_fill_2 FILLER_39_1026 ();
 sg13g2_fill_1 FILLER_39_1028 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_4 FILLER_40_28 ();
 sg13g2_fill_1 FILLER_40_32 ();
 sg13g2_decap_8 FILLER_40_46 ();
 sg13g2_decap_8 FILLER_40_53 ();
 sg13g2_decap_8 FILLER_40_60 ();
 sg13g2_decap_8 FILLER_40_67 ();
 sg13g2_decap_8 FILLER_40_74 ();
 sg13g2_decap_8 FILLER_40_81 ();
 sg13g2_decap_8 FILLER_40_88 ();
 sg13g2_decap_8 FILLER_40_95 ();
 sg13g2_decap_8 FILLER_40_102 ();
 sg13g2_decap_8 FILLER_40_118 ();
 sg13g2_decap_8 FILLER_40_125 ();
 sg13g2_decap_8 FILLER_40_132 ();
 sg13g2_decap_8 FILLER_40_139 ();
 sg13g2_decap_8 FILLER_40_146 ();
 sg13g2_decap_8 FILLER_40_153 ();
 sg13g2_decap_8 FILLER_40_160 ();
 sg13g2_decap_8 FILLER_40_167 ();
 sg13g2_decap_8 FILLER_40_174 ();
 sg13g2_decap_8 FILLER_40_181 ();
 sg13g2_decap_8 FILLER_40_188 ();
 sg13g2_decap_8 FILLER_40_195 ();
 sg13g2_decap_8 FILLER_40_202 ();
 sg13g2_decap_8 FILLER_40_209 ();
 sg13g2_fill_2 FILLER_40_216 ();
 sg13g2_fill_1 FILLER_40_218 ();
 sg13g2_decap_8 FILLER_40_232 ();
 sg13g2_fill_2 FILLER_40_239 ();
 sg13g2_fill_1 FILLER_40_241 ();
 sg13g2_decap_8 FILLER_40_250 ();
 sg13g2_decap_8 FILLER_40_257 ();
 sg13g2_decap_8 FILLER_40_264 ();
 sg13g2_fill_2 FILLER_40_271 ();
 sg13g2_fill_1 FILLER_40_273 ();
 sg13g2_decap_8 FILLER_40_283 ();
 sg13g2_decap_8 FILLER_40_290 ();
 sg13g2_decap_8 FILLER_40_297 ();
 sg13g2_decap_8 FILLER_40_304 ();
 sg13g2_decap_8 FILLER_40_320 ();
 sg13g2_decap_8 FILLER_40_327 ();
 sg13g2_decap_4 FILLER_40_334 ();
 sg13g2_decap_8 FILLER_40_351 ();
 sg13g2_decap_4 FILLER_40_358 ();
 sg13g2_fill_1 FILLER_40_362 ();
 sg13g2_decap_8 FILLER_40_402 ();
 sg13g2_decap_8 FILLER_40_409 ();
 sg13g2_decap_8 FILLER_40_416 ();
 sg13g2_decap_8 FILLER_40_423 ();
 sg13g2_decap_8 FILLER_40_430 ();
 sg13g2_decap_8 FILLER_40_437 ();
 sg13g2_decap_8 FILLER_40_444 ();
 sg13g2_decap_4 FILLER_40_451 ();
 sg13g2_decap_8 FILLER_40_460 ();
 sg13g2_decap_8 FILLER_40_467 ();
 sg13g2_decap_8 FILLER_40_474 ();
 sg13g2_decap_8 FILLER_40_481 ();
 sg13g2_decap_8 FILLER_40_488 ();
 sg13g2_decap_8 FILLER_40_495 ();
 sg13g2_decap_8 FILLER_40_502 ();
 sg13g2_decap_8 FILLER_40_509 ();
 sg13g2_decap_8 FILLER_40_516 ();
 sg13g2_decap_8 FILLER_40_523 ();
 sg13g2_decap_8 FILLER_40_530 ();
 sg13g2_decap_8 FILLER_40_537 ();
 sg13g2_decap_8 FILLER_40_544 ();
 sg13g2_decap_8 FILLER_40_551 ();
 sg13g2_decap_8 FILLER_40_558 ();
 sg13g2_decap_8 FILLER_40_565 ();
 sg13g2_decap_8 FILLER_40_572 ();
 sg13g2_decap_8 FILLER_40_579 ();
 sg13g2_decap_8 FILLER_40_586 ();
 sg13g2_decap_8 FILLER_40_593 ();
 sg13g2_decap_8 FILLER_40_600 ();
 sg13g2_decap_8 FILLER_40_607 ();
 sg13g2_decap_8 FILLER_40_614 ();
 sg13g2_decap_8 FILLER_40_621 ();
 sg13g2_decap_8 FILLER_40_628 ();
 sg13g2_decap_8 FILLER_40_635 ();
 sg13g2_decap_8 FILLER_40_642 ();
 sg13g2_decap_8 FILLER_40_649 ();
 sg13g2_decap_8 FILLER_40_656 ();
 sg13g2_decap_8 FILLER_40_663 ();
 sg13g2_decap_8 FILLER_40_670 ();
 sg13g2_decap_8 FILLER_40_677 ();
 sg13g2_decap_8 FILLER_40_684 ();
 sg13g2_decap_8 FILLER_40_691 ();
 sg13g2_decap_8 FILLER_40_698 ();
 sg13g2_decap_8 FILLER_40_705 ();
 sg13g2_decap_8 FILLER_40_712 ();
 sg13g2_decap_8 FILLER_40_719 ();
 sg13g2_decap_8 FILLER_40_726 ();
 sg13g2_decap_8 FILLER_40_733 ();
 sg13g2_decap_8 FILLER_40_740 ();
 sg13g2_decap_8 FILLER_40_747 ();
 sg13g2_decap_8 FILLER_40_754 ();
 sg13g2_decap_8 FILLER_40_761 ();
 sg13g2_decap_8 FILLER_40_768 ();
 sg13g2_decap_8 FILLER_40_775 ();
 sg13g2_decap_8 FILLER_40_782 ();
 sg13g2_decap_8 FILLER_40_789 ();
 sg13g2_decap_8 FILLER_40_796 ();
 sg13g2_decap_8 FILLER_40_803 ();
 sg13g2_decap_8 FILLER_40_810 ();
 sg13g2_decap_8 FILLER_40_817 ();
 sg13g2_decap_8 FILLER_40_824 ();
 sg13g2_decap_8 FILLER_40_831 ();
 sg13g2_decap_8 FILLER_40_838 ();
 sg13g2_decap_8 FILLER_40_845 ();
 sg13g2_decap_8 FILLER_40_852 ();
 sg13g2_decap_8 FILLER_40_859 ();
 sg13g2_decap_8 FILLER_40_866 ();
 sg13g2_decap_8 FILLER_40_873 ();
 sg13g2_decap_8 FILLER_40_880 ();
 sg13g2_decap_8 FILLER_40_887 ();
 sg13g2_decap_8 FILLER_40_894 ();
 sg13g2_decap_8 FILLER_40_901 ();
 sg13g2_decap_8 FILLER_40_908 ();
 sg13g2_decap_8 FILLER_40_915 ();
 sg13g2_decap_8 FILLER_40_922 ();
 sg13g2_decap_8 FILLER_40_929 ();
 sg13g2_decap_8 FILLER_40_936 ();
 sg13g2_decap_8 FILLER_40_943 ();
 sg13g2_decap_8 FILLER_40_950 ();
 sg13g2_decap_8 FILLER_40_957 ();
 sg13g2_decap_8 FILLER_40_964 ();
 sg13g2_decap_8 FILLER_40_971 ();
 sg13g2_decap_8 FILLER_40_978 ();
 sg13g2_decap_8 FILLER_40_985 ();
 sg13g2_decap_8 FILLER_40_992 ();
 sg13g2_decap_8 FILLER_40_999 ();
 sg13g2_decap_8 FILLER_40_1006 ();
 sg13g2_decap_8 FILLER_40_1013 ();
 sg13g2_decap_8 FILLER_40_1020 ();
 sg13g2_fill_2 FILLER_40_1027 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_fill_1 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_fill_2 FILLER_41_168 ();
 sg13g2_decap_8 FILLER_41_174 ();
 sg13g2_decap_8 FILLER_41_181 ();
 sg13g2_decap_8 FILLER_41_188 ();
 sg13g2_decap_8 FILLER_41_195 ();
 sg13g2_decap_8 FILLER_41_202 ();
 sg13g2_decap_8 FILLER_41_209 ();
 sg13g2_decap_8 FILLER_41_216 ();
 sg13g2_decap_8 FILLER_41_223 ();
 sg13g2_decap_8 FILLER_41_230 ();
 sg13g2_decap_8 FILLER_41_237 ();
 sg13g2_decap_8 FILLER_41_244 ();
 sg13g2_decap_8 FILLER_41_251 ();
 sg13g2_decap_8 FILLER_41_258 ();
 sg13g2_decap_8 FILLER_41_265 ();
 sg13g2_decap_8 FILLER_41_272 ();
 sg13g2_decap_8 FILLER_41_279 ();
 sg13g2_decap_8 FILLER_41_286 ();
 sg13g2_decap_8 FILLER_41_293 ();
 sg13g2_decap_8 FILLER_41_300 ();
 sg13g2_decap_8 FILLER_41_307 ();
 sg13g2_decap_8 FILLER_41_314 ();
 sg13g2_decap_8 FILLER_41_321 ();
 sg13g2_decap_8 FILLER_41_328 ();
 sg13g2_decap_8 FILLER_41_335 ();
 sg13g2_decap_4 FILLER_41_342 ();
 sg13g2_decap_8 FILLER_41_373 ();
 sg13g2_fill_1 FILLER_41_380 ();
 sg13g2_decap_8 FILLER_41_393 ();
 sg13g2_decap_8 FILLER_41_400 ();
 sg13g2_fill_1 FILLER_41_407 ();
 sg13g2_decap_8 FILLER_41_416 ();
 sg13g2_decap_8 FILLER_41_423 ();
 sg13g2_decap_4 FILLER_41_430 ();
 sg13g2_fill_2 FILLER_41_434 ();
 sg13g2_decap_4 FILLER_41_463 ();
 sg13g2_decap_8 FILLER_41_471 ();
 sg13g2_decap_8 FILLER_41_478 ();
 sg13g2_decap_8 FILLER_41_485 ();
 sg13g2_decap_8 FILLER_41_492 ();
 sg13g2_decap_8 FILLER_41_499 ();
 sg13g2_decap_8 FILLER_41_506 ();
 sg13g2_decap_8 FILLER_41_513 ();
 sg13g2_decap_8 FILLER_41_520 ();
 sg13g2_decap_8 FILLER_41_527 ();
 sg13g2_decap_8 FILLER_41_534 ();
 sg13g2_decap_8 FILLER_41_541 ();
 sg13g2_decap_8 FILLER_41_548 ();
 sg13g2_decap_8 FILLER_41_555 ();
 sg13g2_decap_8 FILLER_41_562 ();
 sg13g2_decap_8 FILLER_41_569 ();
 sg13g2_decap_8 FILLER_41_576 ();
 sg13g2_decap_8 FILLER_41_583 ();
 sg13g2_decap_8 FILLER_41_590 ();
 sg13g2_decap_8 FILLER_41_597 ();
 sg13g2_decap_8 FILLER_41_604 ();
 sg13g2_decap_8 FILLER_41_611 ();
 sg13g2_decap_8 FILLER_41_618 ();
 sg13g2_decap_8 FILLER_41_625 ();
 sg13g2_decap_8 FILLER_41_632 ();
 sg13g2_decap_8 FILLER_41_639 ();
 sg13g2_decap_8 FILLER_41_646 ();
 sg13g2_decap_8 FILLER_41_653 ();
 sg13g2_decap_8 FILLER_41_660 ();
 sg13g2_decap_8 FILLER_41_667 ();
 sg13g2_decap_8 FILLER_41_674 ();
 sg13g2_decap_8 FILLER_41_681 ();
 sg13g2_decap_8 FILLER_41_688 ();
 sg13g2_decap_8 FILLER_41_695 ();
 sg13g2_decap_8 FILLER_41_702 ();
 sg13g2_decap_8 FILLER_41_709 ();
 sg13g2_decap_8 FILLER_41_716 ();
 sg13g2_decap_8 FILLER_41_723 ();
 sg13g2_decap_8 FILLER_41_730 ();
 sg13g2_decap_8 FILLER_41_737 ();
 sg13g2_decap_8 FILLER_41_744 ();
 sg13g2_decap_8 FILLER_41_751 ();
 sg13g2_decap_8 FILLER_41_758 ();
 sg13g2_decap_8 FILLER_41_765 ();
 sg13g2_decap_8 FILLER_41_772 ();
 sg13g2_decap_8 FILLER_41_779 ();
 sg13g2_decap_8 FILLER_41_786 ();
 sg13g2_decap_8 FILLER_41_793 ();
 sg13g2_decap_8 FILLER_41_800 ();
 sg13g2_decap_8 FILLER_41_807 ();
 sg13g2_decap_8 FILLER_41_814 ();
 sg13g2_decap_8 FILLER_41_821 ();
 sg13g2_decap_8 FILLER_41_828 ();
 sg13g2_decap_8 FILLER_41_835 ();
 sg13g2_decap_8 FILLER_41_842 ();
 sg13g2_decap_8 FILLER_41_849 ();
 sg13g2_decap_8 FILLER_41_856 ();
 sg13g2_decap_8 FILLER_41_863 ();
 sg13g2_decap_8 FILLER_41_870 ();
 sg13g2_decap_8 FILLER_41_877 ();
 sg13g2_decap_8 FILLER_41_884 ();
 sg13g2_decap_8 FILLER_41_891 ();
 sg13g2_decap_8 FILLER_41_898 ();
 sg13g2_decap_8 FILLER_41_905 ();
 sg13g2_decap_8 FILLER_41_912 ();
 sg13g2_decap_8 FILLER_41_919 ();
 sg13g2_decap_8 FILLER_41_926 ();
 sg13g2_decap_8 FILLER_41_933 ();
 sg13g2_decap_8 FILLER_41_940 ();
 sg13g2_decap_8 FILLER_41_947 ();
 sg13g2_decap_8 FILLER_41_954 ();
 sg13g2_decap_8 FILLER_41_961 ();
 sg13g2_decap_8 FILLER_41_968 ();
 sg13g2_decap_8 FILLER_41_975 ();
 sg13g2_decap_8 FILLER_41_982 ();
 sg13g2_decap_8 FILLER_41_989 ();
 sg13g2_decap_8 FILLER_41_996 ();
 sg13g2_decap_8 FILLER_41_1003 ();
 sg13g2_decap_8 FILLER_41_1010 ();
 sg13g2_decap_8 FILLER_41_1017 ();
 sg13g2_decap_4 FILLER_41_1024 ();
 sg13g2_fill_1 FILLER_41_1028 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_4 FILLER_42_56 ();
 sg13g2_fill_1 FILLER_42_60 ();
 sg13g2_decap_8 FILLER_42_74 ();
 sg13g2_decap_4 FILLER_42_81 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_fill_1 FILLER_42_158 ();
 sg13g2_decap_8 FILLER_42_163 ();
 sg13g2_decap_8 FILLER_42_170 ();
 sg13g2_decap_8 FILLER_42_177 ();
 sg13g2_decap_8 FILLER_42_184 ();
 sg13g2_decap_8 FILLER_42_191 ();
 sg13g2_decap_8 FILLER_42_198 ();
 sg13g2_decap_8 FILLER_42_205 ();
 sg13g2_decap_8 FILLER_42_212 ();
 sg13g2_fill_1 FILLER_42_219 ();
 sg13g2_decap_8 FILLER_42_247 ();
 sg13g2_decap_4 FILLER_42_254 ();
 sg13g2_fill_2 FILLER_42_258 ();
 sg13g2_decap_8 FILLER_42_287 ();
 sg13g2_decap_8 FILLER_42_294 ();
 sg13g2_decap_8 FILLER_42_301 ();
 sg13g2_decap_8 FILLER_42_308 ();
 sg13g2_decap_8 FILLER_42_315 ();
 sg13g2_decap_8 FILLER_42_322 ();
 sg13g2_decap_8 FILLER_42_329 ();
 sg13g2_decap_8 FILLER_42_336 ();
 sg13g2_decap_8 FILLER_42_343 ();
 sg13g2_decap_8 FILLER_42_350 ();
 sg13g2_decap_8 FILLER_42_357 ();
 sg13g2_decap_8 FILLER_42_364 ();
 sg13g2_decap_8 FILLER_42_371 ();
 sg13g2_decap_8 FILLER_42_387 ();
 sg13g2_decap_8 FILLER_42_394 ();
 sg13g2_decap_8 FILLER_42_401 ();
 sg13g2_decap_8 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_42_415 ();
 sg13g2_decap_8 FILLER_42_422 ();
 sg13g2_decap_8 FILLER_42_429 ();
 sg13g2_decap_8 FILLER_42_436 ();
 sg13g2_fill_2 FILLER_42_443 ();
 sg13g2_decap_4 FILLER_42_449 ();
 sg13g2_fill_2 FILLER_42_453 ();
 sg13g2_fill_2 FILLER_42_464 ();
 sg13g2_decap_8 FILLER_42_493 ();
 sg13g2_decap_8 FILLER_42_500 ();
 sg13g2_decap_8 FILLER_42_507 ();
 sg13g2_decap_8 FILLER_42_514 ();
 sg13g2_decap_8 FILLER_42_521 ();
 sg13g2_decap_8 FILLER_42_528 ();
 sg13g2_decap_8 FILLER_42_535 ();
 sg13g2_decap_8 FILLER_42_542 ();
 sg13g2_decap_8 FILLER_42_549 ();
 sg13g2_decap_8 FILLER_42_556 ();
 sg13g2_decap_8 FILLER_42_563 ();
 sg13g2_decap_8 FILLER_42_570 ();
 sg13g2_decap_8 FILLER_42_577 ();
 sg13g2_decap_8 FILLER_42_584 ();
 sg13g2_decap_8 FILLER_42_591 ();
 sg13g2_decap_8 FILLER_42_598 ();
 sg13g2_decap_8 FILLER_42_605 ();
 sg13g2_decap_8 FILLER_42_612 ();
 sg13g2_decap_8 FILLER_42_619 ();
 sg13g2_decap_8 FILLER_42_626 ();
 sg13g2_decap_8 FILLER_42_633 ();
 sg13g2_decap_8 FILLER_42_640 ();
 sg13g2_decap_8 FILLER_42_647 ();
 sg13g2_decap_8 FILLER_42_654 ();
 sg13g2_decap_8 FILLER_42_661 ();
 sg13g2_decap_8 FILLER_42_668 ();
 sg13g2_decap_8 FILLER_42_675 ();
 sg13g2_decap_8 FILLER_42_682 ();
 sg13g2_decap_8 FILLER_42_689 ();
 sg13g2_decap_8 FILLER_42_696 ();
 sg13g2_decap_8 FILLER_42_703 ();
 sg13g2_decap_8 FILLER_42_710 ();
 sg13g2_decap_8 FILLER_42_717 ();
 sg13g2_decap_8 FILLER_42_724 ();
 sg13g2_decap_8 FILLER_42_731 ();
 sg13g2_decap_8 FILLER_42_738 ();
 sg13g2_decap_8 FILLER_42_745 ();
 sg13g2_decap_8 FILLER_42_752 ();
 sg13g2_decap_8 FILLER_42_759 ();
 sg13g2_decap_8 FILLER_42_766 ();
 sg13g2_decap_8 FILLER_42_773 ();
 sg13g2_decap_8 FILLER_42_780 ();
 sg13g2_decap_8 FILLER_42_787 ();
 sg13g2_decap_8 FILLER_42_794 ();
 sg13g2_decap_8 FILLER_42_801 ();
 sg13g2_decap_8 FILLER_42_808 ();
 sg13g2_decap_8 FILLER_42_815 ();
 sg13g2_decap_8 FILLER_42_822 ();
 sg13g2_decap_8 FILLER_42_829 ();
 sg13g2_decap_8 FILLER_42_836 ();
 sg13g2_decap_8 FILLER_42_843 ();
 sg13g2_decap_8 FILLER_42_850 ();
 sg13g2_decap_8 FILLER_42_857 ();
 sg13g2_decap_8 FILLER_42_864 ();
 sg13g2_decap_8 FILLER_42_871 ();
 sg13g2_decap_8 FILLER_42_878 ();
 sg13g2_decap_8 FILLER_42_885 ();
 sg13g2_decap_8 FILLER_42_892 ();
 sg13g2_decap_8 FILLER_42_899 ();
 sg13g2_decap_8 FILLER_42_906 ();
 sg13g2_decap_8 FILLER_42_913 ();
 sg13g2_decap_8 FILLER_42_920 ();
 sg13g2_decap_8 FILLER_42_927 ();
 sg13g2_decap_8 FILLER_42_934 ();
 sg13g2_decap_8 FILLER_42_941 ();
 sg13g2_decap_8 FILLER_42_948 ();
 sg13g2_decap_8 FILLER_42_955 ();
 sg13g2_decap_8 FILLER_42_962 ();
 sg13g2_decap_8 FILLER_42_969 ();
 sg13g2_decap_8 FILLER_42_976 ();
 sg13g2_decap_8 FILLER_42_983 ();
 sg13g2_decap_8 FILLER_42_990 ();
 sg13g2_decap_8 FILLER_42_997 ();
 sg13g2_decap_8 FILLER_42_1004 ();
 sg13g2_decap_8 FILLER_42_1011 ();
 sg13g2_decap_8 FILLER_42_1018 ();
 sg13g2_decap_4 FILLER_42_1025 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_121 ();
 sg13g2_decap_8 FILLER_43_128 ();
 sg13g2_decap_8 FILLER_43_135 ();
 sg13g2_decap_8 FILLER_43_142 ();
 sg13g2_decap_8 FILLER_43_185 ();
 sg13g2_decap_8 FILLER_43_192 ();
 sg13g2_decap_8 FILLER_43_199 ();
 sg13g2_decap_8 FILLER_43_206 ();
 sg13g2_decap_8 FILLER_43_213 ();
 sg13g2_decap_8 FILLER_43_220 ();
 sg13g2_decap_8 FILLER_43_227 ();
 sg13g2_decap_8 FILLER_43_234 ();
 sg13g2_decap_4 FILLER_43_241 ();
 sg13g2_decap_8 FILLER_43_261 ();
 sg13g2_decap_8 FILLER_43_268 ();
 sg13g2_decap_8 FILLER_43_275 ();
 sg13g2_decap_8 FILLER_43_282 ();
 sg13g2_decap_8 FILLER_43_289 ();
 sg13g2_decap_8 FILLER_43_296 ();
 sg13g2_decap_8 FILLER_43_303 ();
 sg13g2_decap_8 FILLER_43_310 ();
 sg13g2_decap_8 FILLER_43_317 ();
 sg13g2_decap_8 FILLER_43_324 ();
 sg13g2_decap_8 FILLER_43_331 ();
 sg13g2_decap_8 FILLER_43_338 ();
 sg13g2_decap_8 FILLER_43_345 ();
 sg13g2_decap_8 FILLER_43_352 ();
 sg13g2_decap_8 FILLER_43_359 ();
 sg13g2_decap_8 FILLER_43_366 ();
 sg13g2_decap_8 FILLER_43_373 ();
 sg13g2_decap_8 FILLER_43_380 ();
 sg13g2_decap_8 FILLER_43_387 ();
 sg13g2_decap_8 FILLER_43_394 ();
 sg13g2_decap_8 FILLER_43_401 ();
 sg13g2_decap_8 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_43_415 ();
 sg13g2_decap_8 FILLER_43_422 ();
 sg13g2_decap_8 FILLER_43_429 ();
 sg13g2_decap_8 FILLER_43_436 ();
 sg13g2_decap_8 FILLER_43_443 ();
 sg13g2_decap_8 FILLER_43_450 ();
 sg13g2_decap_8 FILLER_43_457 ();
 sg13g2_decap_8 FILLER_43_464 ();
 sg13g2_decap_8 FILLER_43_471 ();
 sg13g2_fill_2 FILLER_43_478 ();
 sg13g2_fill_1 FILLER_43_480 ();
 sg13g2_decap_8 FILLER_43_490 ();
 sg13g2_decap_8 FILLER_43_497 ();
 sg13g2_decap_8 FILLER_43_504 ();
 sg13g2_decap_8 FILLER_43_511 ();
 sg13g2_decap_8 FILLER_43_518 ();
 sg13g2_decap_8 FILLER_43_525 ();
 sg13g2_decap_8 FILLER_43_532 ();
 sg13g2_decap_8 FILLER_43_539 ();
 sg13g2_decap_8 FILLER_43_546 ();
 sg13g2_decap_8 FILLER_43_553 ();
 sg13g2_decap_8 FILLER_43_560 ();
 sg13g2_decap_8 FILLER_43_567 ();
 sg13g2_decap_8 FILLER_43_574 ();
 sg13g2_decap_8 FILLER_43_581 ();
 sg13g2_decap_8 FILLER_43_588 ();
 sg13g2_decap_8 FILLER_43_595 ();
 sg13g2_decap_8 FILLER_43_602 ();
 sg13g2_decap_8 FILLER_43_609 ();
 sg13g2_decap_8 FILLER_43_616 ();
 sg13g2_decap_8 FILLER_43_623 ();
 sg13g2_decap_8 FILLER_43_630 ();
 sg13g2_decap_8 FILLER_43_637 ();
 sg13g2_decap_8 FILLER_43_644 ();
 sg13g2_decap_8 FILLER_43_651 ();
 sg13g2_decap_8 FILLER_43_658 ();
 sg13g2_decap_8 FILLER_43_665 ();
 sg13g2_decap_8 FILLER_43_672 ();
 sg13g2_decap_8 FILLER_43_679 ();
 sg13g2_decap_8 FILLER_43_686 ();
 sg13g2_decap_8 FILLER_43_693 ();
 sg13g2_decap_8 FILLER_43_700 ();
 sg13g2_decap_8 FILLER_43_707 ();
 sg13g2_decap_8 FILLER_43_714 ();
 sg13g2_decap_8 FILLER_43_721 ();
 sg13g2_decap_8 FILLER_43_728 ();
 sg13g2_decap_8 FILLER_43_735 ();
 sg13g2_decap_8 FILLER_43_742 ();
 sg13g2_decap_8 FILLER_43_749 ();
 sg13g2_decap_8 FILLER_43_756 ();
 sg13g2_decap_8 FILLER_43_763 ();
 sg13g2_decap_8 FILLER_43_770 ();
 sg13g2_decap_8 FILLER_43_777 ();
 sg13g2_decap_8 FILLER_43_784 ();
 sg13g2_decap_8 FILLER_43_791 ();
 sg13g2_decap_8 FILLER_43_798 ();
 sg13g2_decap_8 FILLER_43_805 ();
 sg13g2_decap_8 FILLER_43_812 ();
 sg13g2_decap_8 FILLER_43_819 ();
 sg13g2_decap_8 FILLER_43_826 ();
 sg13g2_decap_8 FILLER_43_833 ();
 sg13g2_decap_8 FILLER_43_840 ();
 sg13g2_decap_8 FILLER_43_847 ();
 sg13g2_decap_8 FILLER_43_854 ();
 sg13g2_decap_8 FILLER_43_861 ();
 sg13g2_decap_8 FILLER_43_868 ();
 sg13g2_decap_8 FILLER_43_875 ();
 sg13g2_decap_8 FILLER_43_882 ();
 sg13g2_decap_8 FILLER_43_889 ();
 sg13g2_decap_8 FILLER_43_896 ();
 sg13g2_decap_8 FILLER_43_903 ();
 sg13g2_decap_8 FILLER_43_910 ();
 sg13g2_decap_8 FILLER_43_917 ();
 sg13g2_decap_8 FILLER_43_924 ();
 sg13g2_decap_8 FILLER_43_931 ();
 sg13g2_decap_8 FILLER_43_938 ();
 sg13g2_decap_8 FILLER_43_945 ();
 sg13g2_decap_8 FILLER_43_952 ();
 sg13g2_decap_8 FILLER_43_959 ();
 sg13g2_decap_8 FILLER_43_966 ();
 sg13g2_decap_8 FILLER_43_973 ();
 sg13g2_decap_8 FILLER_43_980 ();
 sg13g2_decap_8 FILLER_43_987 ();
 sg13g2_decap_8 FILLER_43_994 ();
 sg13g2_decap_8 FILLER_43_1001 ();
 sg13g2_decap_8 FILLER_43_1008 ();
 sg13g2_decap_8 FILLER_43_1015 ();
 sg13g2_decap_8 FILLER_43_1022 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_4 FILLER_44_28 ();
 sg13g2_fill_2 FILLER_44_32 ();
 sg13g2_decap_8 FILLER_44_61 ();
 sg13g2_decap_8 FILLER_44_68 ();
 sg13g2_fill_1 FILLER_44_75 ();
 sg13g2_decap_8 FILLER_44_89 ();
 sg13g2_decap_8 FILLER_44_96 ();
 sg13g2_decap_8 FILLER_44_103 ();
 sg13g2_decap_8 FILLER_44_110 ();
 sg13g2_decap_8 FILLER_44_117 ();
 sg13g2_decap_8 FILLER_44_124 ();
 sg13g2_decap_8 FILLER_44_131 ();
 sg13g2_decap_4 FILLER_44_138 ();
 sg13g2_fill_2 FILLER_44_142 ();
 sg13g2_decap_8 FILLER_44_180 ();
 sg13g2_decap_8 FILLER_44_187 ();
 sg13g2_decap_4 FILLER_44_194 ();
 sg13g2_fill_2 FILLER_44_198 ();
 sg13g2_decap_8 FILLER_44_213 ();
 sg13g2_decap_8 FILLER_44_220 ();
 sg13g2_decap_8 FILLER_44_227 ();
 sg13g2_decap_8 FILLER_44_234 ();
 sg13g2_decap_8 FILLER_44_241 ();
 sg13g2_decap_8 FILLER_44_248 ();
 sg13g2_decap_8 FILLER_44_255 ();
 sg13g2_decap_8 FILLER_44_262 ();
 sg13g2_decap_8 FILLER_44_269 ();
 sg13g2_decap_8 FILLER_44_276 ();
 sg13g2_decap_8 FILLER_44_283 ();
 sg13g2_decap_8 FILLER_44_290 ();
 sg13g2_decap_8 FILLER_44_297 ();
 sg13g2_decap_4 FILLER_44_304 ();
 sg13g2_fill_1 FILLER_44_308 ();
 sg13g2_decap_8 FILLER_44_336 ();
 sg13g2_fill_2 FILLER_44_343 ();
 sg13g2_decap_8 FILLER_44_350 ();
 sg13g2_decap_8 FILLER_44_357 ();
 sg13g2_decap_8 FILLER_44_364 ();
 sg13g2_decap_8 FILLER_44_371 ();
 sg13g2_decap_4 FILLER_44_378 ();
 sg13g2_decap_8 FILLER_44_409 ();
 sg13g2_decap_8 FILLER_44_416 ();
 sg13g2_decap_8 FILLER_44_423 ();
 sg13g2_decap_8 FILLER_44_430 ();
 sg13g2_decap_8 FILLER_44_437 ();
 sg13g2_decap_8 FILLER_44_444 ();
 sg13g2_decap_8 FILLER_44_451 ();
 sg13g2_decap_8 FILLER_44_458 ();
 sg13g2_decap_8 FILLER_44_465 ();
 sg13g2_decap_8 FILLER_44_472 ();
 sg13g2_decap_8 FILLER_44_479 ();
 sg13g2_decap_8 FILLER_44_486 ();
 sg13g2_decap_8 FILLER_44_493 ();
 sg13g2_decap_8 FILLER_44_500 ();
 sg13g2_decap_8 FILLER_44_507 ();
 sg13g2_decap_8 FILLER_44_514 ();
 sg13g2_decap_8 FILLER_44_521 ();
 sg13g2_decap_8 FILLER_44_528 ();
 sg13g2_decap_8 FILLER_44_535 ();
 sg13g2_decap_8 FILLER_44_542 ();
 sg13g2_decap_8 FILLER_44_549 ();
 sg13g2_decap_8 FILLER_44_556 ();
 sg13g2_decap_8 FILLER_44_563 ();
 sg13g2_decap_8 FILLER_44_570 ();
 sg13g2_decap_8 FILLER_44_577 ();
 sg13g2_decap_8 FILLER_44_584 ();
 sg13g2_decap_8 FILLER_44_591 ();
 sg13g2_decap_8 FILLER_44_598 ();
 sg13g2_decap_8 FILLER_44_605 ();
 sg13g2_decap_8 FILLER_44_612 ();
 sg13g2_decap_8 FILLER_44_619 ();
 sg13g2_decap_8 FILLER_44_626 ();
 sg13g2_decap_8 FILLER_44_633 ();
 sg13g2_decap_8 FILLER_44_640 ();
 sg13g2_decap_8 FILLER_44_647 ();
 sg13g2_decap_8 FILLER_44_654 ();
 sg13g2_decap_8 FILLER_44_661 ();
 sg13g2_decap_8 FILLER_44_668 ();
 sg13g2_decap_8 FILLER_44_675 ();
 sg13g2_decap_8 FILLER_44_682 ();
 sg13g2_decap_8 FILLER_44_689 ();
 sg13g2_decap_8 FILLER_44_696 ();
 sg13g2_decap_8 FILLER_44_703 ();
 sg13g2_decap_8 FILLER_44_710 ();
 sg13g2_decap_8 FILLER_44_717 ();
 sg13g2_decap_8 FILLER_44_724 ();
 sg13g2_decap_8 FILLER_44_731 ();
 sg13g2_decap_8 FILLER_44_738 ();
 sg13g2_decap_8 FILLER_44_745 ();
 sg13g2_decap_8 FILLER_44_752 ();
 sg13g2_decap_8 FILLER_44_759 ();
 sg13g2_decap_8 FILLER_44_766 ();
 sg13g2_decap_8 FILLER_44_773 ();
 sg13g2_decap_8 FILLER_44_780 ();
 sg13g2_decap_8 FILLER_44_787 ();
 sg13g2_decap_8 FILLER_44_794 ();
 sg13g2_decap_8 FILLER_44_801 ();
 sg13g2_decap_8 FILLER_44_808 ();
 sg13g2_decap_8 FILLER_44_815 ();
 sg13g2_decap_8 FILLER_44_822 ();
 sg13g2_decap_8 FILLER_44_829 ();
 sg13g2_decap_8 FILLER_44_836 ();
 sg13g2_decap_8 FILLER_44_843 ();
 sg13g2_decap_8 FILLER_44_850 ();
 sg13g2_decap_8 FILLER_44_857 ();
 sg13g2_decap_8 FILLER_44_864 ();
 sg13g2_decap_8 FILLER_44_871 ();
 sg13g2_decap_8 FILLER_44_878 ();
 sg13g2_decap_8 FILLER_44_885 ();
 sg13g2_decap_8 FILLER_44_892 ();
 sg13g2_decap_8 FILLER_44_899 ();
 sg13g2_decap_8 FILLER_44_906 ();
 sg13g2_decap_8 FILLER_44_913 ();
 sg13g2_decap_8 FILLER_44_920 ();
 sg13g2_decap_8 FILLER_44_927 ();
 sg13g2_decap_8 FILLER_44_934 ();
 sg13g2_decap_8 FILLER_44_941 ();
 sg13g2_decap_8 FILLER_44_948 ();
 sg13g2_decap_8 FILLER_44_955 ();
 sg13g2_decap_8 FILLER_44_962 ();
 sg13g2_decap_8 FILLER_44_969 ();
 sg13g2_decap_8 FILLER_44_976 ();
 sg13g2_decap_8 FILLER_44_983 ();
 sg13g2_decap_8 FILLER_44_990 ();
 sg13g2_decap_8 FILLER_44_997 ();
 sg13g2_decap_8 FILLER_44_1004 ();
 sg13g2_decap_8 FILLER_44_1011 ();
 sg13g2_decap_8 FILLER_44_1018 ();
 sg13g2_decap_4 FILLER_44_1025 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_fill_2 FILLER_45_42 ();
 sg13g2_decap_4 FILLER_45_48 ();
 sg13g2_fill_2 FILLER_45_52 ();
 sg13g2_decap_4 FILLER_45_63 ();
 sg13g2_fill_2 FILLER_45_67 ();
 sg13g2_decap_8 FILLER_45_73 ();
 sg13g2_decap_8 FILLER_45_80 ();
 sg13g2_fill_2 FILLER_45_87 ();
 sg13g2_fill_1 FILLER_45_89 ();
 sg13g2_decap_8 FILLER_45_103 ();
 sg13g2_decap_8 FILLER_45_110 ();
 sg13g2_decap_8 FILLER_45_117 ();
 sg13g2_decap_8 FILLER_45_124 ();
 sg13g2_decap_8 FILLER_45_131 ();
 sg13g2_decap_8 FILLER_45_138 ();
 sg13g2_decap_8 FILLER_45_145 ();
 sg13g2_decap_8 FILLER_45_152 ();
 sg13g2_decap_8 FILLER_45_159 ();
 sg13g2_decap_8 FILLER_45_166 ();
 sg13g2_decap_8 FILLER_45_173 ();
 sg13g2_decap_8 FILLER_45_180 ();
 sg13g2_decap_8 FILLER_45_187 ();
 sg13g2_decap_8 FILLER_45_194 ();
 sg13g2_decap_8 FILLER_45_201 ();
 sg13g2_decap_8 FILLER_45_208 ();
 sg13g2_decap_8 FILLER_45_227 ();
 sg13g2_decap_8 FILLER_45_234 ();
 sg13g2_decap_8 FILLER_45_241 ();
 sg13g2_fill_2 FILLER_45_248 ();
 sg13g2_fill_2 FILLER_45_254 ();
 sg13g2_decap_8 FILLER_45_261 ();
 sg13g2_decap_8 FILLER_45_268 ();
 sg13g2_decap_8 FILLER_45_275 ();
 sg13g2_decap_8 FILLER_45_282 ();
 sg13g2_decap_8 FILLER_45_289 ();
 sg13g2_decap_8 FILLER_45_296 ();
 sg13g2_decap_8 FILLER_45_303 ();
 sg13g2_decap_8 FILLER_45_310 ();
 sg13g2_fill_2 FILLER_45_317 ();
 sg13g2_decap_4 FILLER_45_323 ();
 sg13g2_fill_2 FILLER_45_327 ();
 sg13g2_decap_8 FILLER_45_342 ();
 sg13g2_decap_8 FILLER_45_349 ();
 sg13g2_decap_8 FILLER_45_356 ();
 sg13g2_fill_2 FILLER_45_363 ();
 sg13g2_fill_1 FILLER_45_365 ();
 sg13g2_decap_8 FILLER_45_374 ();
 sg13g2_decap_8 FILLER_45_381 ();
 sg13g2_decap_8 FILLER_45_388 ();
 sg13g2_decap_8 FILLER_45_395 ();
 sg13g2_decap_8 FILLER_45_402 ();
 sg13g2_decap_8 FILLER_45_409 ();
 sg13g2_decap_8 FILLER_45_416 ();
 sg13g2_decap_8 FILLER_45_423 ();
 sg13g2_decap_8 FILLER_45_430 ();
 sg13g2_decap_8 FILLER_45_437 ();
 sg13g2_decap_8 FILLER_45_444 ();
 sg13g2_decap_8 FILLER_45_451 ();
 sg13g2_decap_8 FILLER_45_458 ();
 sg13g2_decap_8 FILLER_45_465 ();
 sg13g2_decap_8 FILLER_45_472 ();
 sg13g2_decap_8 FILLER_45_479 ();
 sg13g2_decap_8 FILLER_45_486 ();
 sg13g2_decap_8 FILLER_45_493 ();
 sg13g2_decap_8 FILLER_45_500 ();
 sg13g2_decap_8 FILLER_45_507 ();
 sg13g2_decap_8 FILLER_45_514 ();
 sg13g2_decap_8 FILLER_45_521 ();
 sg13g2_decap_8 FILLER_45_528 ();
 sg13g2_decap_8 FILLER_45_535 ();
 sg13g2_decap_8 FILLER_45_542 ();
 sg13g2_decap_8 FILLER_45_549 ();
 sg13g2_decap_8 FILLER_45_556 ();
 sg13g2_decap_8 FILLER_45_563 ();
 sg13g2_decap_8 FILLER_45_570 ();
 sg13g2_decap_8 FILLER_45_577 ();
 sg13g2_decap_8 FILLER_45_584 ();
 sg13g2_decap_8 FILLER_45_591 ();
 sg13g2_decap_8 FILLER_45_598 ();
 sg13g2_decap_8 FILLER_45_605 ();
 sg13g2_decap_8 FILLER_45_612 ();
 sg13g2_decap_8 FILLER_45_619 ();
 sg13g2_decap_8 FILLER_45_626 ();
 sg13g2_decap_8 FILLER_45_633 ();
 sg13g2_decap_8 FILLER_45_640 ();
 sg13g2_decap_8 FILLER_45_647 ();
 sg13g2_decap_8 FILLER_45_654 ();
 sg13g2_decap_8 FILLER_45_661 ();
 sg13g2_decap_8 FILLER_45_668 ();
 sg13g2_decap_8 FILLER_45_675 ();
 sg13g2_decap_8 FILLER_45_682 ();
 sg13g2_decap_8 FILLER_45_689 ();
 sg13g2_decap_8 FILLER_45_696 ();
 sg13g2_decap_8 FILLER_45_703 ();
 sg13g2_decap_8 FILLER_45_710 ();
 sg13g2_decap_8 FILLER_45_717 ();
 sg13g2_decap_8 FILLER_45_724 ();
 sg13g2_decap_8 FILLER_45_731 ();
 sg13g2_decap_8 FILLER_45_738 ();
 sg13g2_decap_8 FILLER_45_745 ();
 sg13g2_decap_8 FILLER_45_752 ();
 sg13g2_decap_8 FILLER_45_759 ();
 sg13g2_decap_8 FILLER_45_766 ();
 sg13g2_decap_8 FILLER_45_773 ();
 sg13g2_decap_8 FILLER_45_780 ();
 sg13g2_decap_8 FILLER_45_787 ();
 sg13g2_decap_8 FILLER_45_794 ();
 sg13g2_decap_8 FILLER_45_801 ();
 sg13g2_decap_8 FILLER_45_808 ();
 sg13g2_decap_8 FILLER_45_815 ();
 sg13g2_decap_8 FILLER_45_822 ();
 sg13g2_decap_8 FILLER_45_829 ();
 sg13g2_decap_8 FILLER_45_836 ();
 sg13g2_decap_8 FILLER_45_843 ();
 sg13g2_decap_8 FILLER_45_850 ();
 sg13g2_decap_8 FILLER_45_857 ();
 sg13g2_decap_8 FILLER_45_864 ();
 sg13g2_decap_8 FILLER_45_871 ();
 sg13g2_decap_8 FILLER_45_878 ();
 sg13g2_decap_8 FILLER_45_885 ();
 sg13g2_decap_8 FILLER_45_892 ();
 sg13g2_decap_8 FILLER_45_899 ();
 sg13g2_decap_8 FILLER_45_906 ();
 sg13g2_decap_8 FILLER_45_913 ();
 sg13g2_decap_8 FILLER_45_920 ();
 sg13g2_decap_8 FILLER_45_927 ();
 sg13g2_decap_8 FILLER_45_934 ();
 sg13g2_decap_8 FILLER_45_941 ();
 sg13g2_decap_8 FILLER_45_948 ();
 sg13g2_decap_8 FILLER_45_955 ();
 sg13g2_decap_8 FILLER_45_962 ();
 sg13g2_decap_8 FILLER_45_969 ();
 sg13g2_decap_8 FILLER_45_976 ();
 sg13g2_decap_8 FILLER_45_983 ();
 sg13g2_decap_8 FILLER_45_990 ();
 sg13g2_decap_8 FILLER_45_997 ();
 sg13g2_decap_8 FILLER_45_1004 ();
 sg13g2_decap_8 FILLER_45_1011 ();
 sg13g2_decap_8 FILLER_45_1018 ();
 sg13g2_decap_4 FILLER_45_1025 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_69 ();
 sg13g2_decap_8 FILLER_46_76 ();
 sg13g2_decap_4 FILLER_46_83 ();
 sg13g2_fill_2 FILLER_46_87 ();
 sg13g2_decap_8 FILLER_46_120 ();
 sg13g2_decap_8 FILLER_46_127 ();
 sg13g2_decap_8 FILLER_46_134 ();
 sg13g2_decap_8 FILLER_46_141 ();
 sg13g2_decap_8 FILLER_46_148 ();
 sg13g2_decap_8 FILLER_46_155 ();
 sg13g2_decap_8 FILLER_46_162 ();
 sg13g2_decap_8 FILLER_46_169 ();
 sg13g2_decap_8 FILLER_46_176 ();
 sg13g2_decap_8 FILLER_46_183 ();
 sg13g2_decap_4 FILLER_46_190 ();
 sg13g2_fill_2 FILLER_46_198 ();
 sg13g2_decap_8 FILLER_46_204 ();
 sg13g2_decap_8 FILLER_46_211 ();
 sg13g2_decap_4 FILLER_46_218 ();
 sg13g2_fill_2 FILLER_46_222 ();
 sg13g2_decap_8 FILLER_46_228 ();
 sg13g2_decap_8 FILLER_46_275 ();
 sg13g2_decap_8 FILLER_46_282 ();
 sg13g2_decap_8 FILLER_46_289 ();
 sg13g2_decap_8 FILLER_46_296 ();
 sg13g2_decap_4 FILLER_46_303 ();
 sg13g2_fill_1 FILLER_46_307 ();
 sg13g2_decap_8 FILLER_46_335 ();
 sg13g2_decap_8 FILLER_46_342 ();
 sg13g2_decap_8 FILLER_46_349 ();
 sg13g2_decap_4 FILLER_46_356 ();
 sg13g2_decap_4 FILLER_46_364 ();
 sg13g2_fill_1 FILLER_46_368 ();
 sg13g2_decap_8 FILLER_46_386 ();
 sg13g2_decap_8 FILLER_46_393 ();
 sg13g2_decap_8 FILLER_46_400 ();
 sg13g2_decap_8 FILLER_46_407 ();
 sg13g2_decap_8 FILLER_46_414 ();
 sg13g2_decap_8 FILLER_46_421 ();
 sg13g2_decap_8 FILLER_46_428 ();
 sg13g2_decap_8 FILLER_46_435 ();
 sg13g2_decap_8 FILLER_46_442 ();
 sg13g2_decap_8 FILLER_46_449 ();
 sg13g2_decap_8 FILLER_46_456 ();
 sg13g2_decap_8 FILLER_46_463 ();
 sg13g2_decap_8 FILLER_46_470 ();
 sg13g2_decap_8 FILLER_46_477 ();
 sg13g2_decap_8 FILLER_46_484 ();
 sg13g2_decap_8 FILLER_46_491 ();
 sg13g2_decap_8 FILLER_46_498 ();
 sg13g2_decap_8 FILLER_46_505 ();
 sg13g2_decap_8 FILLER_46_512 ();
 sg13g2_decap_8 FILLER_46_519 ();
 sg13g2_decap_8 FILLER_46_526 ();
 sg13g2_decap_8 FILLER_46_533 ();
 sg13g2_decap_8 FILLER_46_540 ();
 sg13g2_decap_8 FILLER_46_547 ();
 sg13g2_decap_8 FILLER_46_554 ();
 sg13g2_decap_8 FILLER_46_561 ();
 sg13g2_decap_8 FILLER_46_568 ();
 sg13g2_decap_8 FILLER_46_575 ();
 sg13g2_decap_8 FILLER_46_582 ();
 sg13g2_decap_8 FILLER_46_589 ();
 sg13g2_decap_8 FILLER_46_596 ();
 sg13g2_decap_8 FILLER_46_603 ();
 sg13g2_decap_8 FILLER_46_610 ();
 sg13g2_decap_8 FILLER_46_617 ();
 sg13g2_decap_8 FILLER_46_624 ();
 sg13g2_decap_8 FILLER_46_631 ();
 sg13g2_decap_8 FILLER_46_638 ();
 sg13g2_decap_8 FILLER_46_645 ();
 sg13g2_decap_8 FILLER_46_652 ();
 sg13g2_decap_8 FILLER_46_659 ();
 sg13g2_decap_8 FILLER_46_666 ();
 sg13g2_decap_8 FILLER_46_673 ();
 sg13g2_decap_8 FILLER_46_680 ();
 sg13g2_decap_8 FILLER_46_687 ();
 sg13g2_decap_8 FILLER_46_694 ();
 sg13g2_decap_8 FILLER_46_701 ();
 sg13g2_decap_8 FILLER_46_708 ();
 sg13g2_decap_8 FILLER_46_715 ();
 sg13g2_decap_8 FILLER_46_722 ();
 sg13g2_decap_8 FILLER_46_729 ();
 sg13g2_decap_8 FILLER_46_736 ();
 sg13g2_decap_8 FILLER_46_743 ();
 sg13g2_decap_8 FILLER_46_750 ();
 sg13g2_decap_8 FILLER_46_757 ();
 sg13g2_decap_8 FILLER_46_764 ();
 sg13g2_decap_8 FILLER_46_771 ();
 sg13g2_decap_8 FILLER_46_778 ();
 sg13g2_decap_8 FILLER_46_785 ();
 sg13g2_decap_8 FILLER_46_792 ();
 sg13g2_decap_8 FILLER_46_799 ();
 sg13g2_decap_8 FILLER_46_806 ();
 sg13g2_decap_8 FILLER_46_813 ();
 sg13g2_decap_8 FILLER_46_820 ();
 sg13g2_decap_8 FILLER_46_827 ();
 sg13g2_decap_8 FILLER_46_834 ();
 sg13g2_decap_8 FILLER_46_841 ();
 sg13g2_decap_8 FILLER_46_848 ();
 sg13g2_decap_8 FILLER_46_855 ();
 sg13g2_decap_8 FILLER_46_862 ();
 sg13g2_decap_8 FILLER_46_869 ();
 sg13g2_decap_8 FILLER_46_876 ();
 sg13g2_decap_8 FILLER_46_883 ();
 sg13g2_decap_8 FILLER_46_890 ();
 sg13g2_decap_8 FILLER_46_897 ();
 sg13g2_decap_8 FILLER_46_904 ();
 sg13g2_decap_8 FILLER_46_911 ();
 sg13g2_decap_8 FILLER_46_918 ();
 sg13g2_decap_8 FILLER_46_925 ();
 sg13g2_decap_8 FILLER_46_932 ();
 sg13g2_decap_8 FILLER_46_939 ();
 sg13g2_decap_8 FILLER_46_946 ();
 sg13g2_decap_8 FILLER_46_953 ();
 sg13g2_decap_8 FILLER_46_960 ();
 sg13g2_decap_8 FILLER_46_967 ();
 sg13g2_decap_8 FILLER_46_974 ();
 sg13g2_decap_8 FILLER_46_981 ();
 sg13g2_decap_8 FILLER_46_988 ();
 sg13g2_decap_8 FILLER_46_995 ();
 sg13g2_decap_8 FILLER_46_1002 ();
 sg13g2_decap_8 FILLER_46_1009 ();
 sg13g2_decap_8 FILLER_46_1016 ();
 sg13g2_decap_4 FILLER_46_1023 ();
 sg13g2_fill_2 FILLER_46_1027 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_fill_2 FILLER_47_49 ();
 sg13g2_fill_1 FILLER_47_51 ();
 sg13g2_decap_4 FILLER_47_56 ();
 sg13g2_fill_2 FILLER_47_60 ();
 sg13g2_decap_8 FILLER_47_71 ();
 sg13g2_decap_8 FILLER_47_78 ();
 sg13g2_decap_4 FILLER_47_85 ();
 sg13g2_fill_2 FILLER_47_89 ();
 sg13g2_decap_8 FILLER_47_118 ();
 sg13g2_decap_8 FILLER_47_125 ();
 sg13g2_decap_8 FILLER_47_132 ();
 sg13g2_decap_8 FILLER_47_139 ();
 sg13g2_decap_8 FILLER_47_146 ();
 sg13g2_decap_8 FILLER_47_153 ();
 sg13g2_decap_8 FILLER_47_160 ();
 sg13g2_decap_8 FILLER_47_167 ();
 sg13g2_decap_8 FILLER_47_174 ();
 sg13g2_decap_8 FILLER_47_181 ();
 sg13g2_fill_1 FILLER_47_188 ();
 sg13g2_decap_8 FILLER_47_225 ();
 sg13g2_decap_8 FILLER_47_232 ();
 sg13g2_decap_8 FILLER_47_239 ();
 sg13g2_fill_2 FILLER_47_246 ();
 sg13g2_fill_1 FILLER_47_248 ();
 sg13g2_decap_8 FILLER_47_276 ();
 sg13g2_decap_8 FILLER_47_283 ();
 sg13g2_decap_8 FILLER_47_290 ();
 sg13g2_decap_8 FILLER_47_297 ();
 sg13g2_decap_8 FILLER_47_304 ();
 sg13g2_decap_8 FILLER_47_311 ();
 sg13g2_decap_4 FILLER_47_322 ();
 sg13g2_fill_2 FILLER_47_326 ();
 sg13g2_decap_8 FILLER_47_337 ();
 sg13g2_decap_8 FILLER_47_344 ();
 sg13g2_decap_8 FILLER_47_351 ();
 sg13g2_decap_8 FILLER_47_358 ();
 sg13g2_decap_8 FILLER_47_365 ();
 sg13g2_fill_2 FILLER_47_372 ();
 sg13g2_decap_8 FILLER_47_401 ();
 sg13g2_decap_8 FILLER_47_408 ();
 sg13g2_decap_8 FILLER_47_415 ();
 sg13g2_decap_8 FILLER_47_422 ();
 sg13g2_decap_8 FILLER_47_429 ();
 sg13g2_decap_8 FILLER_47_436 ();
 sg13g2_decap_8 FILLER_47_443 ();
 sg13g2_decap_8 FILLER_47_450 ();
 sg13g2_decap_8 FILLER_47_457 ();
 sg13g2_decap_8 FILLER_47_464 ();
 sg13g2_decap_8 FILLER_47_471 ();
 sg13g2_decap_8 FILLER_47_478 ();
 sg13g2_decap_8 FILLER_47_485 ();
 sg13g2_decap_8 FILLER_47_492 ();
 sg13g2_decap_8 FILLER_47_499 ();
 sg13g2_decap_8 FILLER_47_506 ();
 sg13g2_decap_8 FILLER_47_513 ();
 sg13g2_decap_8 FILLER_47_520 ();
 sg13g2_decap_8 FILLER_47_527 ();
 sg13g2_decap_8 FILLER_47_534 ();
 sg13g2_decap_8 FILLER_47_541 ();
 sg13g2_decap_8 FILLER_47_548 ();
 sg13g2_decap_8 FILLER_47_555 ();
 sg13g2_decap_8 FILLER_47_562 ();
 sg13g2_decap_8 FILLER_47_569 ();
 sg13g2_decap_8 FILLER_47_576 ();
 sg13g2_decap_8 FILLER_47_583 ();
 sg13g2_decap_8 FILLER_47_590 ();
 sg13g2_decap_8 FILLER_47_597 ();
 sg13g2_decap_8 FILLER_47_604 ();
 sg13g2_decap_8 FILLER_47_611 ();
 sg13g2_decap_8 FILLER_47_618 ();
 sg13g2_decap_8 FILLER_47_625 ();
 sg13g2_decap_8 FILLER_47_632 ();
 sg13g2_decap_8 FILLER_47_639 ();
 sg13g2_decap_8 FILLER_47_646 ();
 sg13g2_decap_8 FILLER_47_653 ();
 sg13g2_decap_8 FILLER_47_660 ();
 sg13g2_decap_8 FILLER_47_667 ();
 sg13g2_decap_8 FILLER_47_674 ();
 sg13g2_decap_8 FILLER_47_681 ();
 sg13g2_decap_8 FILLER_47_688 ();
 sg13g2_decap_8 FILLER_47_695 ();
 sg13g2_decap_8 FILLER_47_702 ();
 sg13g2_decap_8 FILLER_47_709 ();
 sg13g2_decap_8 FILLER_47_716 ();
 sg13g2_decap_8 FILLER_47_723 ();
 sg13g2_decap_8 FILLER_47_730 ();
 sg13g2_decap_8 FILLER_47_737 ();
 sg13g2_decap_8 FILLER_47_744 ();
 sg13g2_decap_8 FILLER_47_751 ();
 sg13g2_decap_8 FILLER_47_758 ();
 sg13g2_decap_8 FILLER_47_765 ();
 sg13g2_decap_8 FILLER_47_772 ();
 sg13g2_decap_8 FILLER_47_779 ();
 sg13g2_decap_8 FILLER_47_786 ();
 sg13g2_decap_8 FILLER_47_793 ();
 sg13g2_decap_8 FILLER_47_800 ();
 sg13g2_decap_8 FILLER_47_807 ();
 sg13g2_decap_8 FILLER_47_814 ();
 sg13g2_decap_8 FILLER_47_821 ();
 sg13g2_decap_8 FILLER_47_828 ();
 sg13g2_decap_8 FILLER_47_835 ();
 sg13g2_decap_8 FILLER_47_842 ();
 sg13g2_decap_8 FILLER_47_849 ();
 sg13g2_decap_8 FILLER_47_856 ();
 sg13g2_decap_8 FILLER_47_863 ();
 sg13g2_decap_8 FILLER_47_870 ();
 sg13g2_decap_8 FILLER_47_877 ();
 sg13g2_decap_8 FILLER_47_884 ();
 sg13g2_decap_8 FILLER_47_891 ();
 sg13g2_decap_8 FILLER_47_898 ();
 sg13g2_decap_8 FILLER_47_905 ();
 sg13g2_decap_8 FILLER_47_912 ();
 sg13g2_decap_8 FILLER_47_919 ();
 sg13g2_decap_8 FILLER_47_926 ();
 sg13g2_decap_8 FILLER_47_933 ();
 sg13g2_decap_8 FILLER_47_940 ();
 sg13g2_decap_8 FILLER_47_947 ();
 sg13g2_decap_8 FILLER_47_954 ();
 sg13g2_decap_8 FILLER_47_961 ();
 sg13g2_decap_8 FILLER_47_968 ();
 sg13g2_decap_8 FILLER_47_975 ();
 sg13g2_decap_8 FILLER_47_982 ();
 sg13g2_decap_8 FILLER_47_989 ();
 sg13g2_decap_8 FILLER_47_996 ();
 sg13g2_decap_8 FILLER_47_1003 ();
 sg13g2_decap_8 FILLER_47_1010 ();
 sg13g2_decap_8 FILLER_47_1017 ();
 sg13g2_decap_4 FILLER_47_1024 ();
 sg13g2_fill_1 FILLER_47_1028 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_4 FILLER_48_84 ();
 sg13g2_fill_2 FILLER_48_88 ();
 sg13g2_decap_8 FILLER_48_103 ();
 sg13g2_decap_8 FILLER_48_110 ();
 sg13g2_decap_8 FILLER_48_117 ();
 sg13g2_decap_8 FILLER_48_124 ();
 sg13g2_decap_8 FILLER_48_131 ();
 sg13g2_decap_8 FILLER_48_138 ();
 sg13g2_decap_8 FILLER_48_145 ();
 sg13g2_decap_8 FILLER_48_152 ();
 sg13g2_decap_8 FILLER_48_159 ();
 sg13g2_decap_8 FILLER_48_166 ();
 sg13g2_decap_8 FILLER_48_173 ();
 sg13g2_decap_4 FILLER_48_180 ();
 sg13g2_decap_8 FILLER_48_220 ();
 sg13g2_decap_8 FILLER_48_227 ();
 sg13g2_decap_8 FILLER_48_234 ();
 sg13g2_decap_8 FILLER_48_241 ();
 sg13g2_fill_2 FILLER_48_248 ();
 sg13g2_fill_1 FILLER_48_250 ();
 sg13g2_decap_8 FILLER_48_260 ();
 sg13g2_decap_8 FILLER_48_267 ();
 sg13g2_decap_8 FILLER_48_274 ();
 sg13g2_decap_8 FILLER_48_281 ();
 sg13g2_decap_8 FILLER_48_288 ();
 sg13g2_decap_8 FILLER_48_295 ();
 sg13g2_decap_8 FILLER_48_302 ();
 sg13g2_decap_8 FILLER_48_309 ();
 sg13g2_decap_8 FILLER_48_316 ();
 sg13g2_decap_8 FILLER_48_323 ();
 sg13g2_decap_8 FILLER_48_330 ();
 sg13g2_decap_8 FILLER_48_337 ();
 sg13g2_decap_8 FILLER_48_344 ();
 sg13g2_decap_8 FILLER_48_351 ();
 sg13g2_fill_2 FILLER_48_358 ();
 sg13g2_decap_8 FILLER_48_387 ();
 sg13g2_decap_8 FILLER_48_394 ();
 sg13g2_decap_8 FILLER_48_401 ();
 sg13g2_decap_8 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_48_415 ();
 sg13g2_decap_8 FILLER_48_422 ();
 sg13g2_decap_8 FILLER_48_429 ();
 sg13g2_decap_8 FILLER_48_436 ();
 sg13g2_decap_8 FILLER_48_443 ();
 sg13g2_decap_8 FILLER_48_450 ();
 sg13g2_decap_8 FILLER_48_457 ();
 sg13g2_decap_8 FILLER_48_464 ();
 sg13g2_decap_8 FILLER_48_471 ();
 sg13g2_decap_8 FILLER_48_478 ();
 sg13g2_decap_8 FILLER_48_485 ();
 sg13g2_decap_8 FILLER_48_492 ();
 sg13g2_decap_8 FILLER_48_499 ();
 sg13g2_decap_8 FILLER_48_506 ();
 sg13g2_decap_8 FILLER_48_513 ();
 sg13g2_decap_8 FILLER_48_520 ();
 sg13g2_decap_8 FILLER_48_527 ();
 sg13g2_decap_8 FILLER_48_534 ();
 sg13g2_decap_8 FILLER_48_541 ();
 sg13g2_decap_8 FILLER_48_548 ();
 sg13g2_decap_8 FILLER_48_555 ();
 sg13g2_decap_8 FILLER_48_562 ();
 sg13g2_decap_8 FILLER_48_569 ();
 sg13g2_decap_8 FILLER_48_576 ();
 sg13g2_decap_8 FILLER_48_583 ();
 sg13g2_decap_8 FILLER_48_590 ();
 sg13g2_decap_8 FILLER_48_597 ();
 sg13g2_decap_8 FILLER_48_604 ();
 sg13g2_decap_8 FILLER_48_611 ();
 sg13g2_decap_8 FILLER_48_618 ();
 sg13g2_decap_8 FILLER_48_625 ();
 sg13g2_decap_8 FILLER_48_632 ();
 sg13g2_decap_8 FILLER_48_639 ();
 sg13g2_decap_8 FILLER_48_646 ();
 sg13g2_decap_8 FILLER_48_653 ();
 sg13g2_decap_8 FILLER_48_660 ();
 sg13g2_decap_8 FILLER_48_667 ();
 sg13g2_decap_8 FILLER_48_674 ();
 sg13g2_decap_8 FILLER_48_681 ();
 sg13g2_decap_8 FILLER_48_688 ();
 sg13g2_decap_8 FILLER_48_695 ();
 sg13g2_decap_8 FILLER_48_702 ();
 sg13g2_decap_8 FILLER_48_709 ();
 sg13g2_decap_8 FILLER_48_716 ();
 sg13g2_decap_8 FILLER_48_723 ();
 sg13g2_decap_8 FILLER_48_730 ();
 sg13g2_decap_8 FILLER_48_737 ();
 sg13g2_decap_8 FILLER_48_744 ();
 sg13g2_decap_8 FILLER_48_751 ();
 sg13g2_decap_8 FILLER_48_758 ();
 sg13g2_decap_8 FILLER_48_765 ();
 sg13g2_decap_8 FILLER_48_772 ();
 sg13g2_decap_8 FILLER_48_779 ();
 sg13g2_decap_8 FILLER_48_786 ();
 sg13g2_decap_8 FILLER_48_793 ();
 sg13g2_decap_8 FILLER_48_800 ();
 sg13g2_decap_8 FILLER_48_807 ();
 sg13g2_decap_8 FILLER_48_814 ();
 sg13g2_decap_8 FILLER_48_821 ();
 sg13g2_decap_8 FILLER_48_828 ();
 sg13g2_decap_8 FILLER_48_835 ();
 sg13g2_decap_8 FILLER_48_842 ();
 sg13g2_decap_8 FILLER_48_849 ();
 sg13g2_decap_8 FILLER_48_856 ();
 sg13g2_decap_8 FILLER_48_863 ();
 sg13g2_decap_8 FILLER_48_870 ();
 sg13g2_decap_8 FILLER_48_877 ();
 sg13g2_decap_8 FILLER_48_884 ();
 sg13g2_decap_8 FILLER_48_891 ();
 sg13g2_decap_8 FILLER_48_898 ();
 sg13g2_decap_8 FILLER_48_905 ();
 sg13g2_decap_8 FILLER_48_912 ();
 sg13g2_decap_8 FILLER_48_919 ();
 sg13g2_decap_8 FILLER_48_926 ();
 sg13g2_decap_8 FILLER_48_933 ();
 sg13g2_decap_8 FILLER_48_940 ();
 sg13g2_decap_8 FILLER_48_947 ();
 sg13g2_decap_8 FILLER_48_954 ();
 sg13g2_decap_8 FILLER_48_961 ();
 sg13g2_decap_8 FILLER_48_968 ();
 sg13g2_decap_8 FILLER_48_975 ();
 sg13g2_decap_8 FILLER_48_982 ();
 sg13g2_decap_8 FILLER_48_989 ();
 sg13g2_decap_8 FILLER_48_996 ();
 sg13g2_decap_8 FILLER_48_1003 ();
 sg13g2_decap_8 FILLER_48_1010 ();
 sg13g2_decap_8 FILLER_48_1017 ();
 sg13g2_decap_4 FILLER_48_1024 ();
 sg13g2_fill_1 FILLER_48_1028 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_decap_8 FILLER_49_140 ();
 sg13g2_decap_8 FILLER_49_147 ();
 sg13g2_decap_8 FILLER_49_154 ();
 sg13g2_decap_8 FILLER_49_161 ();
 sg13g2_decap_8 FILLER_49_168 ();
 sg13g2_decap_8 FILLER_49_175 ();
 sg13g2_decap_8 FILLER_49_182 ();
 sg13g2_decap_8 FILLER_49_189 ();
 sg13g2_decap_8 FILLER_49_196 ();
 sg13g2_decap_8 FILLER_49_203 ();
 sg13g2_decap_8 FILLER_49_210 ();
 sg13g2_decap_8 FILLER_49_217 ();
 sg13g2_decap_8 FILLER_49_224 ();
 sg13g2_decap_8 FILLER_49_231 ();
 sg13g2_decap_8 FILLER_49_238 ();
 sg13g2_decap_8 FILLER_49_245 ();
 sg13g2_decap_8 FILLER_49_252 ();
 sg13g2_decap_8 FILLER_49_259 ();
 sg13g2_decap_8 FILLER_49_266 ();
 sg13g2_decap_8 FILLER_49_273 ();
 sg13g2_decap_8 FILLER_49_280 ();
 sg13g2_decap_8 FILLER_49_287 ();
 sg13g2_decap_8 FILLER_49_294 ();
 sg13g2_decap_8 FILLER_49_301 ();
 sg13g2_decap_8 FILLER_49_308 ();
 sg13g2_decap_8 FILLER_49_315 ();
 sg13g2_decap_8 FILLER_49_322 ();
 sg13g2_decap_8 FILLER_49_329 ();
 sg13g2_decap_8 FILLER_49_336 ();
 sg13g2_decap_8 FILLER_49_343 ();
 sg13g2_decap_8 FILLER_49_350 ();
 sg13g2_decap_8 FILLER_49_357 ();
 sg13g2_decap_8 FILLER_49_364 ();
 sg13g2_decap_4 FILLER_49_371 ();
 sg13g2_decap_8 FILLER_49_384 ();
 sg13g2_decap_8 FILLER_49_391 ();
 sg13g2_decap_8 FILLER_49_398 ();
 sg13g2_decap_8 FILLER_49_405 ();
 sg13g2_decap_8 FILLER_49_412 ();
 sg13g2_decap_8 FILLER_49_419 ();
 sg13g2_decap_8 FILLER_49_426 ();
 sg13g2_decap_8 FILLER_49_433 ();
 sg13g2_decap_8 FILLER_49_440 ();
 sg13g2_decap_8 FILLER_49_447 ();
 sg13g2_decap_8 FILLER_49_454 ();
 sg13g2_decap_8 FILLER_49_461 ();
 sg13g2_decap_8 FILLER_49_468 ();
 sg13g2_decap_8 FILLER_49_475 ();
 sg13g2_decap_8 FILLER_49_482 ();
 sg13g2_decap_8 FILLER_49_489 ();
 sg13g2_decap_8 FILLER_49_496 ();
 sg13g2_decap_8 FILLER_49_503 ();
 sg13g2_decap_8 FILLER_49_510 ();
 sg13g2_decap_8 FILLER_49_517 ();
 sg13g2_decap_8 FILLER_49_524 ();
 sg13g2_decap_8 FILLER_49_531 ();
 sg13g2_decap_8 FILLER_49_538 ();
 sg13g2_decap_8 FILLER_49_545 ();
 sg13g2_decap_8 FILLER_49_552 ();
 sg13g2_decap_8 FILLER_49_559 ();
 sg13g2_decap_8 FILLER_49_566 ();
 sg13g2_decap_8 FILLER_49_573 ();
 sg13g2_decap_8 FILLER_49_580 ();
 sg13g2_decap_8 FILLER_49_587 ();
 sg13g2_decap_8 FILLER_49_594 ();
 sg13g2_decap_8 FILLER_49_601 ();
 sg13g2_decap_8 FILLER_49_608 ();
 sg13g2_decap_8 FILLER_49_615 ();
 sg13g2_decap_8 FILLER_49_622 ();
 sg13g2_decap_8 FILLER_49_629 ();
 sg13g2_decap_8 FILLER_49_636 ();
 sg13g2_decap_8 FILLER_49_643 ();
 sg13g2_decap_8 FILLER_49_650 ();
 sg13g2_decap_8 FILLER_49_657 ();
 sg13g2_decap_8 FILLER_49_664 ();
 sg13g2_decap_8 FILLER_49_671 ();
 sg13g2_decap_8 FILLER_49_678 ();
 sg13g2_decap_8 FILLER_49_685 ();
 sg13g2_decap_8 FILLER_49_692 ();
 sg13g2_decap_8 FILLER_49_699 ();
 sg13g2_decap_8 FILLER_49_706 ();
 sg13g2_decap_8 FILLER_49_713 ();
 sg13g2_decap_8 FILLER_49_720 ();
 sg13g2_decap_8 FILLER_49_727 ();
 sg13g2_decap_8 FILLER_49_734 ();
 sg13g2_decap_8 FILLER_49_741 ();
 sg13g2_decap_8 FILLER_49_748 ();
 sg13g2_decap_8 FILLER_49_755 ();
 sg13g2_decap_8 FILLER_49_762 ();
 sg13g2_decap_8 FILLER_49_769 ();
 sg13g2_decap_8 FILLER_49_776 ();
 sg13g2_decap_8 FILLER_49_783 ();
 sg13g2_decap_8 FILLER_49_790 ();
 sg13g2_decap_8 FILLER_49_797 ();
 sg13g2_decap_8 FILLER_49_804 ();
 sg13g2_decap_8 FILLER_49_811 ();
 sg13g2_decap_8 FILLER_49_818 ();
 sg13g2_decap_8 FILLER_49_825 ();
 sg13g2_decap_8 FILLER_49_832 ();
 sg13g2_decap_8 FILLER_49_839 ();
 sg13g2_decap_8 FILLER_49_846 ();
 sg13g2_decap_8 FILLER_49_853 ();
 sg13g2_decap_8 FILLER_49_860 ();
 sg13g2_decap_8 FILLER_49_867 ();
 sg13g2_decap_8 FILLER_49_874 ();
 sg13g2_decap_8 FILLER_49_881 ();
 sg13g2_decap_8 FILLER_49_888 ();
 sg13g2_decap_8 FILLER_49_895 ();
 sg13g2_decap_8 FILLER_49_902 ();
 sg13g2_decap_8 FILLER_49_909 ();
 sg13g2_decap_8 FILLER_49_916 ();
 sg13g2_decap_8 FILLER_49_923 ();
 sg13g2_decap_8 FILLER_49_930 ();
 sg13g2_decap_8 FILLER_49_937 ();
 sg13g2_decap_8 FILLER_49_944 ();
 sg13g2_decap_8 FILLER_49_951 ();
 sg13g2_decap_8 FILLER_49_958 ();
 sg13g2_decap_8 FILLER_49_965 ();
 sg13g2_decap_8 FILLER_49_972 ();
 sg13g2_decap_8 FILLER_49_979 ();
 sg13g2_decap_8 FILLER_49_986 ();
 sg13g2_decap_8 FILLER_49_993 ();
 sg13g2_decap_8 FILLER_49_1000 ();
 sg13g2_decap_8 FILLER_49_1007 ();
 sg13g2_decap_8 FILLER_49_1014 ();
 sg13g2_decap_8 FILLER_49_1021 ();
 sg13g2_fill_1 FILLER_49_1028 ();
 assign uio_oe[0] = net17;
 assign uio_oe[1] = net18;
 assign uio_oe[2] = net19;
 assign uio_oe[3] = net20;
 assign uio_oe[4] = net21;
 assign uio_oe[5] = net22;
 assign uio_oe[6] = net23;
 assign uio_oe[7] = net24;
 assign uio_out[0] = net5;
 assign uio_out[1] = net6;
 assign uio_out[2] = net7;
 assign uio_out[3] = net8;
 assign uio_out[4] = net9;
 assign uio_out[5] = net10;
 assign uio_out[6] = net11;
 assign uio_out[7] = net12;
 assign uo_out[4] = net13;
 assign uo_out[5] = net14;
 assign uo_out[6] = net15;
 assign uo_out[7] = net16;
endmodule
