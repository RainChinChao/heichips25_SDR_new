* NGSPICE file created from heichips25_template.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

.subckt heichips25_template VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
XFILLER_27_417 VPWR VGND sg13g2_decap_8
XFILLER_36_940 VPWR VGND sg13g2_decap_8
XFILLER_39_288 VPWR VGND sg13g2_decap_8
XFILLER_35_494 VPWR VGND sg13g2_decap_8
XFILLER_10_317 VPWR VGND sg13g2_decap_8
XFILLER_22_155 VPWR VGND sg13g2_decap_8
XFILLER_23_667 VPWR VGND sg13g2_decap_8
XFILLER_7_7 VPWR VGND sg13g2_decap_8
XFILLER_46_704 VPWR VGND sg13g2_decap_8
XFILLER_33_409 VPWR VGND sg13g2_decap_8
X_501_ net82 VGND VPWR _062_ mac2.products_ff\[102\] clknet_5_30__leaf_clk sg13g2_dfrbpq_1
XFILLER_42_932 VPWR VGND sg13g2_decap_8
XFILLER_14_623 VPWR VGND sg13g2_decap_8
X_432_ net152 _126_ VPWR VGND sg13g2_buf_1
XFILLER_26_74 VPWR VGND sg13g2_decap_8
XFILLER_27_995 VPWR VGND sg13g2_decap_8
XFILLER_26_494 VPWR VGND sg13g2_decap_8
XFILLER_13_144 VPWR VGND sg13g2_decap_8
X_363_ net171 VPWR _019_ VGND _172_ _174_ sg13g2_o21ai_1
XFILLER_41_475 VPWR VGND sg13g2_decap_8
XFILLER_9_137 VPWR VGND sg13g2_decap_8
X_294_ _173_ net170 mac2.sum_lvl3_ff\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_42_73 VPWR VGND sg13g2_decap_8
XFILLER_10_851 VPWR VGND sg13g2_decap_8
XFILLER_6_844 VPWR VGND sg13g2_decap_8
XFILLER_5_310 VPWR VGND sg13g2_decap_8
XFILLER_5_387 VPWR VGND sg13g2_decap_8
XFILLER_49_520 VPWR VGND sg13g2_decap_8
XFILLER_1_593 VPWR VGND sg13g2_decap_8
XFILLER_3_1007 VPWR VGND sg13g2_decap_8
XFILLER_49_597 VPWR VGND sg13g2_decap_8
XFILLER_37_737 VPWR VGND sg13g2_decap_8
XFILLER_17_483 VPWR VGND sg13g2_decap_8
XFILLER_18_984 VPWR VGND sg13g2_decap_8
XFILLER_32_431 VPWR VGND sg13g2_decap_8
XFILLER_33_965 VPWR VGND sg13g2_decap_8
XFILLER_20_626 VPWR VGND sg13g2_decap_8
XFILLER_9_682 VPWR VGND sg13g2_decap_8
XFILLER_41_1002 VPWR VGND sg13g2_decap_8
XFILLER_27_203 VPWR VGND sg13g2_decap_8
XFILLER_27_247 VPWR VGND sg13g2_decap_8
XFILLER_42_206 VPWR VGND sg13g2_decap_8
XFILLER_24_965 VPWR VGND sg13g2_decap_8
XFILLER_35_280 VPWR VGND sg13g2_decap_8
XFILLER_11_648 VPWR VGND sg13g2_decap_8
XFILLER_12_76 VPWR VGND sg13g2_decap_8
XFILLER_3_825 VPWR VGND sg13g2_decap_8
XFILLER_5_4 VPWR VGND sg13g2_decap_8
XFILLER_2_335 VPWR VGND sg13g2_decap_8
XFILLER_46_501 VPWR VGND sg13g2_decap_8
XFILLER_19_748 VPWR VGND sg13g2_decap_8
XFILLER_46_578 VPWR VGND sg13g2_decap_8
XFILLER_15_932 VPWR VGND sg13g2_decap_8
XFILLER_27_792 VPWR VGND sg13g2_decap_8
XFILLER_18_1026 VPWR VGND sg13g2_fill_2
X_415_ net57 _109_ VPWR VGND sg13g2_buf_1
XFILLER_30_913 VPWR VGND sg13g2_decap_8
XFILLER_14_475 VPWR VGND sg13g2_decap_4
XFILLER_14_497 VPWR VGND sg13g2_decap_8
X_346_ _203_ net134 net98 VPWR VGND sg13g2_nand2_1
XFILLER_41_272 VPWR VGND sg13g2_decap_8
X_277_ _164_ net187 net113 VPWR VGND sg13g2_nand2_1
XFILLER_6_641 VPWR VGND sg13g2_decap_8
XFILLER_5_140 VPWR VGND sg13g2_decap_8
XFILLER_2_880 VPWR VGND sg13g2_decap_8
XFILLER_25_1019 VPWR VGND sg13g2_decap_8
XFILLER_1_390 VPWR VGND sg13g2_decap_8
XFILLER_37_534 VPWR VGND sg13g2_decap_8
XFILLER_49_394 VPWR VGND sg13g2_decap_8
XFILLER_18_781 VPWR VGND sg13g2_decap_8
XFILLER_25_718 VPWR VGND sg13g2_decap_8
XFILLER_33_762 VPWR VGND sg13g2_decap_8
XFILLER_20_423 VPWR VGND sg13g2_decap_8
XFILLER_21_946 VPWR VGND sg13g2_decap_8
Xclkbuf_4_12_0_clk clknet_0_clk clknet_4_12_0_clk VPWR VGND sg13g2_buf_8
XFILLER_28_567 VPWR VGND sg13g2_decap_8
XFILLER_16_718 VPWR VGND sg13g2_decap_8
XFILLER_43_559 VPWR VGND sg13g2_decap_8
XFILLER_24_762 VPWR VGND sg13g2_decap_8
XFILLER_12_935 VPWR VGND sg13g2_decap_8
XFILLER_11_456 VPWR VGND sg13g2_decap_8
XFILLER_20_990 VPWR VGND sg13g2_decap_8
XFILLER_3_622 VPWR VGND sg13g2_decap_8
XFILLER_3_699 VPWR VGND sg13g2_decap_8
XFILLER_47_854 VPWR VGND sg13g2_decap_8
XFILLER_46_331 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_19_545 VPWR VGND sg13g2_decap_8
XFILLER_34_559 VPWR VGND sg13g2_decap_8
XFILLER_9_11 VPWR VGND sg13g2_decap_4
XFILLER_14_272 VPWR VGND sg13g2_decap_8
XFILLER_30_710 VPWR VGND sg13g2_decap_8
XFILLER_9_55 VPWR VGND sg13g2_decap_8
X_329_ _192_ net131 net58 VPWR VGND sg13g2_nand2_1
XFILLER_30_787 VPWR VGND sg13g2_decap_8
XFILLER_29_0 VPWR VGND sg13g2_decap_8
XFILLER_38_810 VPWR VGND sg13g2_decap_8
XFILLER_49_191 VPWR VGND sg13g2_decap_8
XFILLER_25_504 VPWR VGND sg13g2_fill_2
XFILLER_25_515 VPWR VGND sg13g2_decap_8
XFILLER_38_887 VPWR VGND sg13g2_decap_8
XFILLER_37_397 VPWR VGND sg13g2_decap_8
XFILLER_20_242 VPWR VGND sg13g2_decap_8
XFILLER_21_743 VPWR VGND sg13g2_decap_8
XFILLER_4_419 VPWR VGND sg13g2_fill_2
XFILLER_4_408 VPWR VGND sg13g2_fill_2
XFILLER_0_658 VPWR VGND sg13g2_decap_8
XFILLER_48_629 VPWR VGND sg13g2_decap_8
XFILLER_18_53 VPWR VGND sg13g2_decap_8
XFILLER_29_876 VPWR VGND sg13g2_decap_8
XFILLER_44_857 VPWR VGND sg13g2_decap_8
XFILLER_43_323 VPWR VGND sg13g2_decap_8
XFILLER_28_397 VPWR VGND sg13g2_decap_8
XFILLER_12_732 VPWR VGND sg13g2_decap_8
XFILLER_8_769 VPWR VGND sg13g2_decap_8
XFILLER_11_297 VPWR VGND sg13g2_decap_8
XFILLER_7_279 VPWR VGND sg13g2_decap_8
XFILLER_4_920 VPWR VGND sg13g2_decap_8
XFILLER_4_997 VPWR VGND sg13g2_decap_8
XFILLER_3_496 VPWR VGND sg13g2_decap_8
XFILLER_3_485 VPWR VGND sg13g2_fill_2
XFILLER_38_117 VPWR VGND sg13g2_decap_8
XFILLER_47_651 VPWR VGND sg13g2_decap_8
XFILLER_19_353 VPWR VGND sg13g2_decap_8
XFILLER_19_364 VPWR VGND sg13g2_fill_1
XFILLER_35_802 VPWR VGND sg13g2_decap_8
XFILLER_46_194 VPWR VGND sg13g2_decap_8
XFILLER_35_879 VPWR VGND sg13g2_decap_8
XFILLER_15_570 VPWR VGND sg13g2_decap_8
XFILLER_22_529 VPWR VGND sg13g2_decap_8
XFILLER_30_584 VPWR VGND sg13g2_decap_8
XFILLER_6_290 VPWR VGND sg13g2_decap_8
XFILLER_29_106 VPWR VGND sg13g2_decap_8
XFILLER_26_802 VPWR VGND sg13g2_decap_8
XFILLER_25_323 VPWR VGND sg13g2_decap_8
XFILLER_38_684 VPWR VGND sg13g2_decap_8
XFILLER_26_879 VPWR VGND sg13g2_decap_8
XFILLER_40_326 VPWR VGND sg13g2_decap_4
XFILLER_41_827 VPWR VGND sg13g2_decap_8
XFILLER_5_717 VPWR VGND sg13g2_decap_8
XFILLER_20_32 VPWR VGND sg13g2_decap_8
XFILLER_1_901 VPWR VGND sg13g2_decap_8
XFILLER_49_905 VPWR VGND sg13g2_decap_8
XFILLER_0_455 VPWR VGND sg13g2_decap_8
XFILLER_1_978 VPWR VGND sg13g2_decap_8
XFILLER_48_426 VPWR VGND sg13g2_decap_8
Xhold30 DP_1.matrix\[55\] VPWR VGND net54 sg13g2_dlygate4sd3_1
Xhold41 DP_1.matrix\[73\] VPWR VGND net91 sg13g2_dlygate4sd3_1
Xhold52 DP_3.matrix\[46\] VPWR VGND net102 sg13g2_dlygate4sd3_1
Xhold63 mac1.products_ff\[68\] VPWR VGND net113 sg13g2_dlygate4sd3_1
Xhold74 _028_ VPWR VGND net124 sg13g2_dlygate4sd3_1
Xhold85 DP_2.matrix\[63\] VPWR VGND net135 sg13g2_dlygate4sd3_1
Xhold96 _010_ VPWR VGND net146 sg13g2_dlygate4sd3_1
XFILLER_29_673 VPWR VGND sg13g2_decap_8
XFILLER_17_824 VPWR VGND sg13g2_decap_8
XFILLER_44_654 VPWR VGND sg13g2_decap_8
XFILLER_43_120 VPWR VGND sg13g2_decap_8
XFILLER_16_334 VPWR VGND sg13g2_decap_8
X_594_ net72 VGND VPWR _134_ DP_4.matrix\[45\] clknet_5_13__leaf_clk sg13g2_dfrbpq_2
XFILLER_32_816 VPWR VGND sg13g2_decap_8
XFILLER_31_315 VPWR VGND sg13g2_decap_8
XFILLER_8_566 VPWR VGND sg13g2_decap_8
XFILLER_6_67 VPWR VGND sg13g2_decap_8
XFILLER_4_794 VPWR VGND sg13g2_decap_8
XFILLER_6_1005 VPWR VGND sg13g2_decap_8
XFILLER_20_4 VPWR VGND sg13g2_decap_8
XFILLER_48_993 VPWR VGND sg13g2_decap_8
XFILLER_19_172 VPWR VGND sg13g2_decap_8
XFILLER_22_304 VPWR VGND sg13g2_fill_1
XFILLER_23_849 VPWR VGND sg13g2_decap_8
XFILLER_35_676 VPWR VGND sg13g2_decap_8
XFILLER_31_860 VPWR VGND sg13g2_decap_8
XFILLER_1_208 VPWR VGND sg13g2_decap_8
XFILLER_44_1011 VPWR VGND sg13g2_decap_8
Xheichips25_template_10 VPWR VGND uio_out[5] sg13g2_tielo
Xheichips25_template_21 VPWR VGND uio_oe[4] sg13g2_tiehi
XFILLER_17_109 VPWR VGND sg13g2_decap_8
XFILLER_45_429 VPWR VGND sg13g2_decap_8
XFILLER_14_805 VPWR VGND sg13g2_decap_8
XFILLER_26_676 VPWR VGND sg13g2_decap_8
XFILLER_41_624 VPWR VGND sg13g2_decap_8
XFILLER_15_54 VPWR VGND sg13g2_decap_4
XFILLER_9_308 VPWR VGND sg13g2_fill_1
XFILLER_40_145 VPWR VGND sg13g2_decap_8
XFILLER_22_893 VPWR VGND sg13g2_decap_8
XFILLER_31_42 VPWR VGND sg13g2_decap_8
XFILLER_49_702 VPWR VGND sg13g2_decap_8
XFILLER_0_252 VPWR VGND sg13g2_decap_8
XFILLER_1_775 VPWR VGND sg13g2_decap_8
XFILLER_48_212 VPWR VGND sg13g2_decap_8
XFILLER_48_223 VPWR VGND sg13g2_fill_1
XFILLER_49_779 VPWR VGND sg13g2_decap_8
XFILLER_37_919 VPWR VGND sg13g2_decap_8
XFILLER_17_621 VPWR VGND sg13g2_decap_8
XFILLER_29_481 VPWR VGND sg13g2_decap_8
XFILLER_16_120 VPWR VGND sg13g2_fill_1
X_577_ net70 VGND VPWR _117_ DP_3.matrix\[46\] clknet_5_14__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_996 VPWR VGND sg13g2_decap_8
XFILLER_44_451 VPWR VGND sg13g2_decap_8
XFILLER_17_698 VPWR VGND sg13g2_decap_8
XFILLER_32_613 VPWR VGND sg13g2_decap_8
XFILLER_31_112 VPWR VGND sg13g2_decap_8
XFILLER_20_808 VPWR VGND sg13g2_decap_8
XFILLER_13_893 VPWR VGND sg13g2_decap_8
XFILLER_31_189 VPWR VGND sg13g2_decap_8
XFILLER_8_341 VPWR VGND sg13g2_fill_1
Xclkbuf_5_17__f_clk clknet_4_8_0_clk clknet_5_17__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_9_864 VPWR VGND sg13g2_decap_8
XFILLER_4_591 VPWR VGND sg13g2_decap_8
XFILLER_48_790 VPWR VGND sg13g2_decap_8
XFILLER_36_996 VPWR VGND sg13g2_decap_8
XFILLER_22_134 VPWR VGND sg13g2_decap_8
XFILLER_23_646 VPWR VGND sg13g2_decap_8
X_500_ net80 VGND VPWR _061_ mac2.products_ff\[86\] clknet_5_14__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_248 VPWR VGND sg13g2_decap_8
XFILLER_42_911 VPWR VGND sg13g2_decap_8
XFILLER_14_602 VPWR VGND sg13g2_decap_8
X_431_ net101 _125_ VPWR VGND sg13g2_buf_1
XFILLER_26_53 VPWR VGND sg13g2_decap_8
XFILLER_26_473 VPWR VGND sg13g2_decap_8
XFILLER_27_974 VPWR VGND sg13g2_decap_8
X_362_ _213_ _212_ _057_ VPWR VGND sg13g2_xor2_1
XFILLER_13_123 VPWR VGND sg13g2_decap_8
XFILLER_42_988 VPWR VGND sg13g2_decap_8
XFILLER_9_116 VPWR VGND sg13g2_decap_8
XFILLER_14_679 VPWR VGND sg13g2_decap_8
XFILLER_41_454 VPWR VGND sg13g2_decap_8
XFILLER_42_52 VPWR VGND sg13g2_decap_8
XFILLER_10_830 VPWR VGND sg13g2_decap_8
XFILLER_13_189 VPWR VGND sg13g2_decap_8
X_293_ _172_ net201 net115 VPWR VGND sg13g2_nand2_1
XFILLER_22_690 VPWR VGND sg13g2_decap_8
XFILLER_6_823 VPWR VGND sg13g2_decap_8
XFILLER_5_366 VPWR VGND sg13g2_decap_8
XFILLER_3_46 VPWR VGND sg13g2_decap_8
XFILLER_1_572 VPWR VGND sg13g2_decap_8
XFILLER_49_576 VPWR VGND sg13g2_decap_8
XFILLER_37_716 VPWR VGND sg13g2_decap_8
XFILLER_18_963 VPWR VGND sg13g2_decap_8
XFILLER_36_237 VPWR VGND sg13g2_decap_8
XFILLER_17_462 VPWR VGND sg13g2_decap_8
XFILLER_45_793 VPWR VGND sg13g2_decap_8
XFILLER_32_421 VPWR VGND sg13g2_fill_2
XFILLER_33_944 VPWR VGND sg13g2_decap_8
XFILLER_20_605 VPWR VGND sg13g2_decap_8
XFILLER_32_487 VPWR VGND sg13g2_decap_8
XFILLER_34_1021 VPWR VGND sg13g2_decap_8
XFILLER_9_661 VPWR VGND sg13g2_decap_8
XFILLER_13_690 VPWR VGND sg13g2_decap_8
XFILLER_28_749 VPWR VGND sg13g2_decap_8
XFILLER_24_944 VPWR VGND sg13g2_decap_8
XFILLER_36_793 VPWR VGND sg13g2_decap_8
XFILLER_11_627 VPWR VGND sg13g2_decap_8
XFILLER_23_476 VPWR VGND sg13g2_decap_4
XFILLER_10_159 VPWR VGND sg13g2_decap_8
XFILLER_12_11 VPWR VGND sg13g2_decap_8
XFILLER_3_804 VPWR VGND sg13g2_decap_8
XFILLER_12_55 VPWR VGND sg13g2_decap_8
XFILLER_2_314 VPWR VGND sg13g2_decap_8
XFILLER_19_727 VPWR VGND sg13g2_decap_8
XFILLER_46_557 VPWR VGND sg13g2_decap_8
XFILLER_15_911 VPWR VGND sg13g2_decap_8
XFILLER_27_771 VPWR VGND sg13g2_decap_8
X_414_ net157 _108_ VPWR VGND sg13g2_buf_1
XFILLER_14_454 VPWR VGND sg13g2_decap_8
XFILLER_15_988 VPWR VGND sg13g2_decap_8
XFILLER_18_1005 VPWR VGND sg13g2_decap_8
XFILLER_41_251 VPWR VGND sg13g2_decap_8
XFILLER_42_785 VPWR VGND sg13g2_decap_8
X_345_ _202_ net129 net55 VPWR VGND sg13g2_nand2_1
XFILLER_41_262 VPWR VGND sg13g2_fill_2
X_276_ net111 mac1.products_ff\[34\] _004_ VPWR VGND sg13g2_xor2_1
XFILLER_30_969 VPWR VGND sg13g2_decap_8
XFILLER_6_620 VPWR VGND sg13g2_decap_8
XFILLER_6_697 VPWR VGND sg13g2_decap_8
XFILLER_5_196 VPWR VGND sg13g2_decap_8
XFILLER_49_373 VPWR VGND sg13g2_decap_8
XFILLER_37_513 VPWR VGND sg13g2_decap_8
XFILLER_18_760 VPWR VGND sg13g2_decap_8
XFILLER_45_590 VPWR VGND sg13g2_decap_8
XFILLER_24_229 VPWR VGND sg13g2_decap_8
XFILLER_33_741 VPWR VGND sg13g2_decap_8
XFILLER_20_402 VPWR VGND sg13g2_decap_8
XFILLER_21_925 VPWR VGND sg13g2_decap_8
XFILLER_32_295 VPWR VGND sg13g2_decap_8
XFILLER_20_479 VPWR VGND sg13g2_decap_8
XFILLER_9_491 VPWR VGND sg13g2_decap_8
XFILLER_28_546 VPWR VGND sg13g2_decap_8
XFILLER_43_538 VPWR VGND sg13g2_decap_8
XFILLER_36_590 VPWR VGND sg13g2_decap_8
XFILLER_12_914 VPWR VGND sg13g2_decap_8
XFILLER_23_240 VPWR VGND sg13g2_decap_8
XFILLER_24_741 VPWR VGND sg13g2_decap_8
XFILLER_11_435 VPWR VGND sg13g2_decap_8
XFILLER_23_87 VPWR VGND sg13g2_decap_8
XFILLER_3_601 VPWR VGND sg13g2_decap_8
XFILLER_3_678 VPWR VGND sg13g2_decap_8
XFILLER_47_833 VPWR VGND sg13g2_decap_8
XFILLER_48_84 VPWR VGND sg13g2_decap_8
XFILLER_46_310 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_19_535 VPWR VGND sg13g2_fill_1
XFILLER_46_387 VPWR VGND sg13g2_decap_8
XFILLER_34_538 VPWR VGND sg13g2_decap_8
XFILLER_42_582 VPWR VGND sg13g2_decap_8
XFILLER_14_251 VPWR VGND sg13g2_decap_8
XFILLER_15_785 VPWR VGND sg13g2_decap_8
XFILLER_30_766 VPWR VGND sg13g2_decap_8
X_328_ _191_ _190_ _035_ VPWR VGND sg13g2_xor2_1
X_259_ _153_ mac1.total_sum\[1\] mac2.total_sum\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_11_991 VPWR VGND sg13g2_decap_8
XFILLER_7_995 VPWR VGND sg13g2_decap_8
XFILLER_9_1025 VPWR VGND sg13g2_decap_4
XFILLER_49_170 VPWR VGND sg13g2_decap_8
XFILLER_38_866 VPWR VGND sg13g2_decap_8
XFILLER_37_376 VPWR VGND sg13g2_decap_8
XFILLER_21_722 VPWR VGND sg13g2_decap_8
XFILLER_20_221 VPWR VGND sg13g2_decap_8
XFILLER_21_799 VPWR VGND sg13g2_decap_8
XFILLER_20_298 VPWR VGND sg13g2_decap_8
XFILLER_0_637 VPWR VGND sg13g2_decap_8
XFILLER_48_608 VPWR VGND sg13g2_decap_8
XFILLER_18_32 VPWR VGND sg13g2_decap_8
XFILLER_29_855 VPWR VGND sg13g2_decap_8
XFILLER_44_836 VPWR VGND sg13g2_decap_8
XFILLER_43_302 VPWR VGND sg13g2_decap_8
XFILLER_16_527 VPWR VGND sg13g2_decap_4
XFILLER_18_98 VPWR VGND sg13g2_decap_8
XFILLER_28_376 VPWR VGND sg13g2_decap_8
XFILLER_43_379 VPWR VGND sg13g2_decap_8
XFILLER_12_711 VPWR VGND sg13g2_decap_8
XFILLER_34_75 VPWR VGND sg13g2_decap_8
XFILLER_7_203 VPWR VGND sg13g2_decap_8
XFILLER_12_788 VPWR VGND sg13g2_decap_8
XFILLER_8_748 VPWR VGND sg13g2_decap_8
XFILLER_11_276 VPWR VGND sg13g2_decap_8
XFILLER_7_258 VPWR VGND sg13g2_decap_8
XFILLER_4_976 VPWR VGND sg13g2_decap_8
XFILLER_3_464 VPWR VGND sg13g2_decap_8
XFILLER_47_630 VPWR VGND sg13g2_decap_8
XFILLER_46_140 VPWR VGND sg13g2_decap_8
Xclkbuf_4_11_0_clk clknet_0_clk clknet_4_11_0_clk VPWR VGND sg13g2_buf_8
XFILLER_35_858 VPWR VGND sg13g2_decap_8
XFILLER_22_508 VPWR VGND sg13g2_decap_8
XFILLER_34_379 VPWR VGND sg13g2_fill_1
XFILLER_30_563 VPWR VGND sg13g2_decap_8
XFILLER_7_792 VPWR VGND sg13g2_decap_8
XFILLER_41_0 VPWR VGND sg13g2_decap_8
XFILLER_38_663 VPWR VGND sg13g2_decap_8
XFILLER_37_184 VPWR VGND sg13g2_decap_8
XFILLER_26_858 VPWR VGND sg13g2_decap_8
XFILLER_41_806 VPWR VGND sg13g2_decap_8
XFILLER_40_305 VPWR VGND sg13g2_decap_8
XFILLER_21_596 VPWR VGND sg13g2_decap_8
XFILLER_20_11 VPWR VGND sg13g2_decap_8
XFILLER_20_88 VPWR VGND sg13g2_decap_8
XFILLER_0_434 VPWR VGND sg13g2_decap_8
XFILLER_1_957 VPWR VGND sg13g2_decap_8
XFILLER_48_405 VPWR VGND sg13g2_fill_1
Xhold20 DP_2.matrix\[37\] VPWR VGND net44 sg13g2_dlygate4sd3_1
Xhold31 DP_1.matrix\[19\] VPWR VGND net55 sg13g2_dlygate4sd3_1
Xhold53 mac2.products_ff\[85\] VPWR VGND net103 sg13g2_dlygate4sd3_1
Xhold42 DP_1.matrix\[64\] VPWR VGND net92 sg13g2_dlygate4sd3_1
Xhold64 _006_ VPWR VGND net114 sg13g2_dlygate4sd3_1
Xhold75 DP_3.matrix\[45\] VPWR VGND net125 sg13g2_dlygate4sd3_1
XFILLER_17_803 VPWR VGND sg13g2_decap_8
XFILLER_21_1023 VPWR VGND sg13g2_decap_4
Xhold97 DP_1.matrix\[9\] VPWR VGND net147 sg13g2_dlygate4sd3_1
XFILLER_29_652 VPWR VGND sg13g2_decap_8
Xhold86 mac2.sum_lvl1_ff\[24\] VPWR VGND net136 sg13g2_dlygate4sd3_1
XFILLER_44_633 VPWR VGND sg13g2_decap_8
XFILLER_16_324 VPWR VGND sg13g2_decap_4
X_593_ net70 VGND VPWR _133_ DP_4.matrix\[37\] clknet_5_11__leaf_clk sg13g2_dfrbpq_1
XFILLER_28_195 VPWR VGND sg13g2_decap_4
XFILLER_24_390 VPWR VGND sg13g2_decap_8
XFILLER_8_545 VPWR VGND sg13g2_decap_8
XFILLER_40_883 VPWR VGND sg13g2_decap_8
XFILLER_6_46 VPWR VGND sg13g2_decap_8
XFILLER_4_773 VPWR VGND sg13g2_decap_8
XFILLER_6_1028 VPWR VGND sg13g2_fill_1
XFILLER_13_4 VPWR VGND sg13g2_decap_8
XFILLER_48_972 VPWR VGND sg13g2_decap_8
XFILLER_19_151 VPWR VGND sg13g2_decap_8
XFILLER_35_655 VPWR VGND sg13g2_decap_8
XFILLER_23_828 VPWR VGND sg13g2_decap_8
XFILLER_34_187 VPWR VGND sg13g2_decap_8
Xheichips25_template_11 VPWR VGND uio_out[6] sg13g2_tielo
XFILLER_45_408 VPWR VGND sg13g2_decap_8
Xheichips25_template_22 VPWR VGND uio_oe[5] sg13g2_tiehi
XFILLER_39_994 VPWR VGND sg13g2_decap_8
XFILLER_26_655 VPWR VGND sg13g2_decap_8
XFILLER_13_316 VPWR VGND sg13g2_decap_8
XFILLER_15_11 VPWR VGND sg13g2_decap_4
XFILLER_41_603 VPWR VGND sg13g2_decap_8
XFILLER_13_327 VPWR VGND sg13g2_decap_8
XFILLER_25_198 VPWR VGND sg13g2_decap_8
XFILLER_40_124 VPWR VGND sg13g2_decap_8
XFILLER_22_872 VPWR VGND sg13g2_decap_8
XFILLER_31_21 VPWR VGND sg13g2_decap_8
XFILLER_31_98 VPWR VGND sg13g2_decap_8
XFILLER_1_754 VPWR VGND sg13g2_decap_8
XFILLER_0_231 VPWR VGND sg13g2_decap_8
XFILLER_49_758 VPWR VGND sg13g2_decap_8
XFILLER_48_257 VPWR VGND sg13g2_fill_2
XFILLER_48_246 VPWR VGND sg13g2_decap_8
XFILLER_44_430 VPWR VGND sg13g2_decap_8
X_576_ net80 VGND VPWR _116_ DP_3.matrix\[45\] clknet_5_15__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_975 VPWR VGND sg13g2_decap_8
XFILLER_17_677 VPWR VGND sg13g2_decap_8
XFILLER_16_176 VPWR VGND sg13g2_decap_8
XFILLER_13_872 VPWR VGND sg13g2_decap_8
XFILLER_31_168 VPWR VGND sg13g2_decap_8
XFILLER_32_669 VPWR VGND sg13g2_decap_8
XFILLER_9_843 VPWR VGND sg13g2_decap_8
XFILLER_40_680 VPWR VGND sg13g2_decap_8
XFILLER_36_975 VPWR VGND sg13g2_decap_8
XFILLER_23_625 VPWR VGND sg13g2_decap_8
XFILLER_11_809 VPWR VGND sg13g2_decap_8
XFILLER_2_518 VPWR VGND sg13g2_fill_1
XFILLER_19_909 VPWR VGND sg13g2_decap_8
XFILLER_46_739 VPWR VGND sg13g2_decap_8
XFILLER_45_227 VPWR VGND sg13g2_decap_8
XFILLER_45_205 VPWR VGND sg13g2_fill_2
Xclkbuf_5_23__f_clk clknet_4_11_0_clk clknet_5_23__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_26_32 VPWR VGND sg13g2_decap_8
XFILLER_27_953 VPWR VGND sg13g2_decap_8
XFILLER_39_791 VPWR VGND sg13g2_decap_8
XFILLER_26_452 VPWR VGND sg13g2_decap_8
X_430_ net119 _124_ VPWR VGND sg13g2_buf_1
X_361_ _213_ net126 net40 VPWR VGND sg13g2_nand2_1
XFILLER_13_102 VPWR VGND sg13g2_decap_8
XFILLER_41_433 VPWR VGND sg13g2_decap_4
XFILLER_42_967 VPWR VGND sg13g2_decap_8
XFILLER_14_658 VPWR VGND sg13g2_decap_8
X_292_ net161 mac1.sum_lvl1_ff\[24\] _012_ VPWR VGND sg13g2_xor2_1
XFILLER_13_168 VPWR VGND sg13g2_decap_8
XFILLER_6_802 VPWR VGND sg13g2_decap_8
XFILLER_10_886 VPWR VGND sg13g2_decap_8
XFILLER_6_879 VPWR VGND sg13g2_decap_8
XFILLER_5_345 VPWR VGND sg13g2_decap_8
XFILLER_3_25 VPWR VGND sg13g2_decap_8
XFILLER_1_551 VPWR VGND sg13g2_decap_8
XFILLER_49_555 VPWR VGND sg13g2_decap_8
XFILLER_36_216 VPWR VGND sg13g2_decap_8
XFILLER_18_942 VPWR VGND sg13g2_decap_8
XFILLER_45_772 VPWR VGND sg13g2_decap_8
XFILLER_17_441 VPWR VGND sg13g2_decap_8
XFILLER_33_923 VPWR VGND sg13g2_decap_8
X_559_ net83 VGND VPWR _099_ DP_2.matrix\[46\] clknet_5_29__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_466 VPWR VGND sg13g2_decap_8
XFILLER_34_1000 VPWR VGND sg13g2_decap_8
XFILLER_9_640 VPWR VGND sg13g2_decap_8
XFILLER_28_728 VPWR VGND sg13g2_decap_8
XFILLER_36_772 VPWR VGND sg13g2_decap_8
XFILLER_24_923 VPWR VGND sg13g2_decap_8
XFILLER_11_606 VPWR VGND sg13g2_decap_8
XFILLER_23_455 VPWR VGND sg13g2_decap_8
XFILLER_10_138 VPWR VGND sg13g2_decap_8
XFILLER_6_109 VPWR VGND sg13g2_decap_8
Xhold150 _001_ VPWR VGND net200 sg13g2_dlygate4sd3_1
XFILLER_19_706 VPWR VGND sg13g2_decap_8
XFILLER_18_216 VPWR VGND sg13g2_fill_1
XFILLER_46_536 VPWR VGND sg13g2_decap_8
XFILLER_2_1020 VPWR VGND sg13g2_decap_8
XFILLER_37_64 VPWR VGND sg13g2_decap_8
XFILLER_27_750 VPWR VGND sg13g2_decap_8
XFILLER_26_271 VPWR VGND sg13g2_fill_2
XFILLER_26_282 VPWR VGND sg13g2_decap_8
X_413_ net88 _107_ VPWR VGND sg13g2_buf_1
XFILLER_42_764 VPWR VGND sg13g2_decap_8
XFILLER_14_433 VPWR VGND sg13g2_decap_8
XFILLER_15_967 VPWR VGND sg13g2_decap_8
XFILLER_18_1028 VPWR VGND sg13g2_fill_1
XFILLER_41_230 VPWR VGND sg13g2_decap_8
XFILLER_30_948 VPWR VGND sg13g2_decap_8
X_344_ _201_ _200_ _045_ VPWR VGND sg13g2_xor2_1
X_275_ _005_ _162_ _163_ VPWR VGND sg13g2_xnor2_1
XFILLER_10_683 VPWR VGND sg13g2_decap_8
XFILLER_6_676 VPWR VGND sg13g2_decap_8
XFILLER_45_7 VPWR VGND sg13g2_decap_8
XFILLER_5_175 VPWR VGND sg13g2_decap_8
XFILLER_49_352 VPWR VGND sg13g2_decap_8
XFILLER_24_208 VPWR VGND sg13g2_decap_8
XFILLER_37_569 VPWR VGND sg13g2_decap_8
XFILLER_33_720 VPWR VGND sg13g2_decap_8
XFILLER_17_293 VPWR VGND sg13g2_decap_8
XFILLER_21_904 VPWR VGND sg13g2_decap_8
XFILLER_32_230 VPWR VGND sg13g2_fill_1
XFILLER_32_274 VPWR VGND sg13g2_decap_8
XFILLER_33_797 VPWR VGND sg13g2_decap_8
XFILLER_20_458 VPWR VGND sg13g2_decap_8
XFILLER_0_819 VPWR VGND sg13g2_decap_8
XFILLER_28_525 VPWR VGND sg13g2_decap_8
XFILLER_43_517 VPWR VGND sg13g2_decap_8
XFILLER_24_720 VPWR VGND sg13g2_decap_8
XFILLER_24_797 VPWR VGND sg13g2_decap_8
XFILLER_23_296 VPWR VGND sg13g2_decap_8
XFILLER_7_429 VPWR VGND sg13g2_decap_8
XFILLER_2_112 VPWR VGND sg13g2_fill_2
XFILLER_3_657 VPWR VGND sg13g2_decap_8
XFILLER_2_123 VPWR VGND sg13g2_decap_8
XFILLER_2_167 VPWR VGND sg13g2_decap_8
XFILLER_24_1021 VPWR VGND sg13g2_decap_8
XFILLER_47_812 VPWR VGND sg13g2_decap_8
XFILLER_48_63 VPWR VGND sg13g2_decap_8
XFILLER_47_889 VPWR VGND sg13g2_decap_8
XFILLER_46_366 VPWR VGND sg13g2_decap_8
XFILLER_34_517 VPWR VGND sg13g2_decap_8
XFILLER_14_230 VPWR VGND sg13g2_decap_8
XFILLER_15_764 VPWR VGND sg13g2_decap_8
XFILLER_42_561 VPWR VGND sg13g2_decap_8
X_327_ _191_ net141 net51 VPWR VGND sg13g2_nand2_1
XFILLER_30_745 VPWR VGND sg13g2_decap_8
XFILLER_11_970 VPWR VGND sg13g2_decap_8
XFILLER_31_1014 VPWR VGND sg13g2_decap_8
X_258_ _152_ mac1.total_sum\[0\] mac2.total_sum\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_7_974 VPWR VGND sg13g2_decap_8
XFILLER_6_462 VPWR VGND sg13g2_fill_2
XFILLER_9_1004 VPWR VGND sg13g2_decap_8
XFILLER_38_845 VPWR VGND sg13g2_decap_8
XFILLER_25_506 VPWR VGND sg13g2_fill_1
XFILLER_37_355 VPWR VGND sg13g2_decap_8
XFILLER_21_701 VPWR VGND sg13g2_decap_8
XFILLER_20_200 VPWR VGND sg13g2_decap_8
XFILLER_33_594 VPWR VGND sg13g2_decap_8
XFILLER_21_778 VPWR VGND sg13g2_decap_8
XFILLER_20_277 VPWR VGND sg13g2_decap_8
XFILLER_0_616 VPWR VGND sg13g2_decap_8
XFILLER_18_11 VPWR VGND sg13g2_decap_8
XFILLER_29_834 VPWR VGND sg13g2_decap_8
XFILLER_44_815 VPWR VGND sg13g2_decap_8
XFILLER_16_506 VPWR VGND sg13g2_fill_1
XFILLER_28_355 VPWR VGND sg13g2_decap_8
XFILLER_43_358 VPWR VGND sg13g2_decap_8
XFILLER_34_21 VPWR VGND sg13g2_decap_8
XFILLER_15_1009 VPWR VGND sg13g2_decap_8
XFILLER_24_594 VPWR VGND sg13g2_decap_8
XFILLER_8_727 VPWR VGND sg13g2_decap_8
XFILLER_11_244 VPWR VGND sg13g2_decap_8
XFILLER_12_767 VPWR VGND sg13g2_decap_8
XFILLER_7_237 VPWR VGND sg13g2_decap_8
XFILLER_4_955 VPWR VGND sg13g2_decap_8
XFILLER_3_443 VPWR VGND sg13g2_decap_8
XFILLER_3_487 VPWR VGND sg13g2_fill_1
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_39_609 VPWR VGND sg13g2_decap_8
XFILLER_38_108 VPWR VGND sg13g2_fill_1
XFILLER_47_686 VPWR VGND sg13g2_decap_8
XFILLER_19_399 VPWR VGND sg13g2_decap_8
XFILLER_35_837 VPWR VGND sg13g2_decap_8
XFILLER_34_358 VPWR VGND sg13g2_decap_8
XFILLER_43_881 VPWR VGND sg13g2_decap_8
XFILLER_15_550 VPWR VGND sg13g2_decap_8
XFILLER_30_542 VPWR VGND sg13g2_decap_8
XFILLER_7_771 VPWR VGND sg13g2_decap_8
XFILLER_34_0 VPWR VGND sg13g2_decap_8
Xclkbuf_5_4__f_clk clknet_4_2_0_clk clknet_5_4__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_38_642 VPWR VGND sg13g2_decap_8
XFILLER_26_837 VPWR VGND sg13g2_decap_8
XFILLER_37_163 VPWR VGND sg13g2_decap_8
XFILLER_25_358 VPWR VGND sg13g2_decap_8
XFILLER_34_881 VPWR VGND sg13g2_decap_8
XFILLER_33_380 VPWR VGND sg13g2_decap_8
XFILLER_21_542 VPWR VGND sg13g2_decap_8
XFILLER_20_67 VPWR VGND sg13g2_decap_8
XFILLER_0_413 VPWR VGND sg13g2_decap_8
XFILLER_1_936 VPWR VGND sg13g2_decap_8
Xhold32 DP_3.matrix\[19\] VPWR VGND net56 sg13g2_dlygate4sd3_1
Xhold21 DP_4.matrix\[19\] VPWR VGND net45 sg13g2_dlygate4sd3_1
Xhold10 mac2.sum_lvl2_ff\[9\] VPWR VGND net34 sg13g2_dlygate4sd3_1
Xhold65 mac2.sum_lvl3_ff\[0\] VPWR VGND net115 sg13g2_dlygate4sd3_1
XFILLER_21_1002 VPWR VGND sg13g2_decap_8
Xhold43 mac1.products_ff\[0\] VPWR VGND net93 sg13g2_dlygate4sd3_1
XFILLER_29_631 VPWR VGND sg13g2_decap_8
Xhold54 _026_ VPWR VGND net104 sg13g2_dlygate4sd3_1
Xhold98 DP_3.matrix\[18\] VPWR VGND net148 sg13g2_dlygate4sd3_1
Xhold76 DP_1.matrix\[63\] VPWR VGND net126 sg13g2_dlygate4sd3_1
Xhold87 _032_ VPWR VGND net137 sg13g2_dlygate4sd3_1
XFILLER_44_612 VPWR VGND sg13g2_decap_8
X_592_ net71 VGND VPWR _132_ DP_4.matrix\[36\] clknet_5_14__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_53 VPWR VGND sg13g2_fill_2
XFILLER_45_42 VPWR VGND sg13g2_decap_8
XFILLER_17_859 VPWR VGND sg13g2_decap_8
XFILLER_45_97 VPWR VGND sg13g2_decap_8
XFILLER_44_689 VPWR VGND sg13g2_decap_8
XFILLER_16_369 VPWR VGND sg13g2_decap_8
XFILLER_40_862 VPWR VGND sg13g2_decap_8
XFILLER_8_524 VPWR VGND sg13g2_decap_8
XFILLER_6_25 VPWR VGND sg13g2_decap_8
XFILLER_4_752 VPWR VGND sg13g2_decap_8
XFILLER_39_406 VPWR VGND sg13g2_decap_8
XFILLER_0_980 VPWR VGND sg13g2_decap_8
XFILLER_48_951 VPWR VGND sg13g2_decap_8
XFILLER_19_130 VPWR VGND sg13g2_decap_8
XFILLER_47_483 VPWR VGND sg13g2_decap_8
XFILLER_35_634 VPWR VGND sg13g2_decap_8
XFILLER_23_807 VPWR VGND sg13g2_decap_8
XFILLER_22_339 VPWR VGND sg13g2_decap_8
XFILLER_30_372 VPWR VGND sg13g2_decap_4
XFILLER_31_895 VPWR VGND sg13g2_decap_8
Xheichips25_template_12 VPWR VGND uio_out[7] sg13g2_tielo
Xheichips25_template_23 VPWR VGND uio_oe[6] sg13g2_tiehi
XFILLER_39_973 VPWR VGND sg13g2_decap_8
XFILLER_25_111 VPWR VGND sg13g2_decap_8
XFILLER_26_634 VPWR VGND sg13g2_decap_8
XFILLER_25_177 VPWR VGND sg13g2_decap_8
XFILLER_22_851 VPWR VGND sg13g2_decap_8
XFILLER_41_659 VPWR VGND sg13g2_decap_8
Xclkbuf_4_10_0_clk clknet_0_clk clknet_4_10_0_clk VPWR VGND sg13g2_buf_8
XFILLER_5_527 VPWR VGND sg13g2_decap_8
XFILLER_31_77 VPWR VGND sg13g2_decap_8
XFILLER_0_210 VPWR VGND sg13g2_decap_8
XFILLER_1_733 VPWR VGND sg13g2_decap_8
XFILLER_49_737 VPWR VGND sg13g2_decap_8
XFILLER_0_287 VPWR VGND sg13g2_decap_8
XFILLER_45_954 VPWR VGND sg13g2_decap_8
XFILLER_17_656 VPWR VGND sg13g2_decap_8
X_575_ net70 VGND VPWR _115_ DP_3.matrix\[37\] clknet_5_14__leaf_clk sg13g2_dfrbpq_1
XFILLER_16_155 VPWR VGND sg13g2_decap_8
XFILLER_44_486 VPWR VGND sg13g2_decap_8
XFILLER_32_648 VPWR VGND sg13g2_decap_8
XFILLER_13_851 VPWR VGND sg13g2_decap_8
XFILLER_31_147 VPWR VGND sg13g2_decap_8
XFILLER_9_822 VPWR VGND sg13g2_decap_8
XFILLER_12_372 VPWR VGND sg13g2_decap_8
XFILLER_8_332 VPWR VGND sg13g2_decap_8
XFILLER_8_387 VPWR VGND sg13g2_fill_2
XFILLER_8_376 VPWR VGND sg13g2_decap_8
XFILLER_9_899 VPWR VGND sg13g2_decap_8
XFILLER_8_398 VPWR VGND sg13g2_decap_8
XFILLER_4_560 VPWR VGND sg13g2_decap_8
XFILLER_28_1008 VPWR VGND sg13g2_decap_8
XFILLER_39_203 VPWR VGND sg13g2_decap_8
XFILLER_35_431 VPWR VGND sg13g2_decap_4
XFILLER_36_954 VPWR VGND sg13g2_decap_8
XFILLER_23_604 VPWR VGND sg13g2_decap_8
XFILLER_22_103 VPWR VGND sg13g2_decap_4
XFILLER_22_169 VPWR VGND sg13g2_decap_8
XFILLER_31_692 VPWR VGND sg13g2_decap_8
XFILLER_11_1012 VPWR VGND sg13g2_decap_8
XFILLER_46_718 VPWR VGND sg13g2_decap_8
XFILLER_39_770 VPWR VGND sg13g2_decap_8
XFILLER_26_11 VPWR VGND sg13g2_decap_8
XFILLER_26_431 VPWR VGND sg13g2_decap_8
XFILLER_27_932 VPWR VGND sg13g2_decap_8
XFILLER_42_946 VPWR VGND sg13g2_decap_8
X_360_ _212_ net135 net92 VPWR VGND sg13g2_nand2_1
XFILLER_14_637 VPWR VGND sg13g2_decap_8
XFILLER_26_88 VPWR VGND sg13g2_decap_8
XFILLER_41_412 VPWR VGND sg13g2_decap_8
XFILLER_13_158 VPWR VGND sg13g2_fill_1
X_291_ _013_ _170_ _171_ VPWR VGND sg13g2_xnor2_1
XFILLER_41_489 VPWR VGND sg13g2_decap_8
XFILLER_42_21 VPWR VGND sg13g2_decap_8
XFILLER_42_87 VPWR VGND sg13g2_decap_8
XFILLER_10_865 VPWR VGND sg13g2_decap_8
XFILLER_6_858 VPWR VGND sg13g2_decap_8
XFILLER_5_324 VPWR VGND sg13g2_decap_8
XFILLER_1_530 VPWR VGND sg13g2_decap_8
XFILLER_49_534 VPWR VGND sg13g2_decap_8
XFILLER_18_921 VPWR VGND sg13g2_decap_8
XFILLER_45_751 VPWR VGND sg13g2_decap_8
XFILLER_33_902 VPWR VGND sg13g2_decap_8
XFILLER_44_283 VPWR VGND sg13g2_decap_8
XFILLER_18_998 VPWR VGND sg13g2_decap_8
X_558_ net77 VGND VPWR _098_ DP_2.matrix\[45\] clknet_5_29__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_445 VPWR VGND sg13g2_decap_8
XFILLER_33_979 VPWR VGND sg13g2_decap_8
X_489_ net69 VGND VPWR _064_ mac2.products_ff\[0\] clknet_5_9__leaf_clk sg13g2_dfrbpq_1
XFILLER_9_696 VPWR VGND sg13g2_decap_8
XFILLER_28_707 VPWR VGND sg13g2_decap_8
XFILLER_41_1016 VPWR VGND sg13g2_decap_8
XFILLER_41_1027 VPWR VGND sg13g2_fill_2
XFILLER_24_902 VPWR VGND sg13g2_decap_8
XFILLER_36_751 VPWR VGND sg13g2_decap_8
XFILLER_23_401 VPWR VGND sg13g2_decap_8
XFILLER_24_979 VPWR VGND sg13g2_decap_8
XFILLER_35_294 VPWR VGND sg13g2_decap_8
XFILLER_3_839 VPWR VGND sg13g2_decap_8
Xhold151 mac2.sum_lvl3_ff\[2\] VPWR VGND net201 sg13g2_dlygate4sd3_1
Xhold140 _033_ VPWR VGND net190 sg13g2_dlygate4sd3_1
XFILLER_2_349 VPWR VGND sg13g2_decap_8
XFILLER_46_515 VPWR VGND sg13g2_decap_8
XFILLER_37_21 VPWR VGND sg13g2_decap_8
XFILLER_37_98 VPWR VGND sg13g2_decap_8
XFILLER_14_412 VPWR VGND sg13g2_decap_4
XFILLER_15_946 VPWR VGND sg13g2_decap_8
XFILLER_26_261 VPWR VGND sg13g2_fill_2
X_412_ net132 _106_ VPWR VGND sg13g2_buf_1
XFILLER_42_743 VPWR VGND sg13g2_decap_8
XFILLER_30_927 VPWR VGND sg13g2_decap_8
X_343_ _201_ net147 net48 VPWR VGND sg13g2_nand2_1
X_274_ mac1.products_ff\[52\] mac1.products_ff\[35\] _163_ VPWR VGND sg13g2_xor2_1
XFILLER_10_662 VPWR VGND sg13g2_decap_8
XFILLER_6_655 VPWR VGND sg13g2_decap_8
XFILLER_5_154 VPWR VGND sg13g2_decap_8
XFILLER_2_894 VPWR VGND sg13g2_decap_8
XFILLER_38_7 VPWR VGND sg13g2_decap_8
XFILLER_49_331 VPWR VGND sg13g2_decap_8
XFILLER_37_548 VPWR VGND sg13g2_decap_8
XFILLER_17_272 VPWR VGND sg13g2_decap_8
XFILLER_18_795 VPWR VGND sg13g2_decap_8
XFILLER_33_776 VPWR VGND sg13g2_decap_8
XFILLER_20_437 VPWR VGND sg13g2_decap_8
XFILLER_24_776 VPWR VGND sg13g2_decap_8
XFILLER_8_909 VPWR VGND sg13g2_decap_8
XFILLER_12_949 VPWR VGND sg13g2_decap_8
XFILLER_23_45 VPWR VGND sg13g2_decap_8
XFILLER_3_636 VPWR VGND sg13g2_decap_8
XFILLER_3_4 VPWR VGND sg13g2_decap_8
XFILLER_48_42 VPWR VGND sg13g2_decap_8
XFILLER_24_1000 VPWR VGND sg13g2_decap_8
XFILLER_19_504 VPWR VGND sg13g2_fill_2
XFILLER_47_868 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_19_559 VPWR VGND sg13g2_decap_8
XFILLER_42_540 VPWR VGND sg13g2_decap_8
XFILLER_15_743 VPWR VGND sg13g2_decap_8
X_326_ _190_ net121 net86 VPWR VGND sg13g2_nand2_1
XFILLER_9_69 VPWR VGND sg13g2_decap_8
XFILLER_14_286 VPWR VGND sg13g2_decap_8
XFILLER_30_724 VPWR VGND sg13g2_decap_8
XFILLER_7_953 VPWR VGND sg13g2_decap_8
X_257_ mac2.sum_lvl2_ff\[4\] net163 _000_ VPWR VGND sg13g2_xor2_1
XFILLER_6_441 VPWR VGND sg13g2_decap_8
XFILLER_6_474 VPWR VGND sg13g2_fill_2
XFILLER_2_691 VPWR VGND sg13g2_decap_8
XFILLER_38_824 VPWR VGND sg13g2_decap_8
XFILLER_18_570 VPWR VGND sg13g2_decap_8
XFILLER_25_529 VPWR VGND sg13g2_decap_8
XFILLER_33_573 VPWR VGND sg13g2_decap_8
XFILLER_20_256 VPWR VGND sg13g2_decap_8
XFILLER_21_757 VPWR VGND sg13g2_decap_8
XFILLER_47_1022 VPWR VGND sg13g2_decap_8
XFILLER_29_813 VPWR VGND sg13g2_decap_8
XFILLER_18_67 VPWR VGND sg13g2_decap_8
XFILLER_43_337 VPWR VGND sg13g2_decap_8
XFILLER_24_573 VPWR VGND sg13g2_decap_8
XFILLER_34_44 VPWR VGND sg13g2_decap_8
XFILLER_11_223 VPWR VGND sg13g2_decap_8
XFILLER_12_746 VPWR VGND sg13g2_decap_8
XFILLER_8_706 VPWR VGND sg13g2_decap_8
XFILLER_4_934 VPWR VGND sg13g2_decap_8
XFILLER_47_665 VPWR VGND sg13g2_decap_8
XFILLER_19_378 VPWR VGND sg13g2_decap_8
XFILLER_35_816 VPWR VGND sg13g2_decap_8
XFILLER_34_337 VPWR VGND sg13g2_decap_8
XFILLER_43_860 VPWR VGND sg13g2_decap_8
XFILLER_30_521 VPWR VGND sg13g2_decap_8
XFILLER_30_598 VPWR VGND sg13g2_decap_8
X_309_ _029_ _180_ _181_ VPWR VGND sg13g2_xnor2_1
XFILLER_7_750 VPWR VGND sg13g2_decap_8
XFILLER_27_0 VPWR VGND sg13g2_decap_8
XFILLER_38_621 VPWR VGND sg13g2_decap_8
XFILLER_37_142 VPWR VGND sg13g2_decap_8
XFILLER_1_70 VPWR VGND sg13g2_decap_4
XFILLER_26_816 VPWR VGND sg13g2_decap_8
XFILLER_38_698 VPWR VGND sg13g2_decap_8
XFILLER_25_337 VPWR VGND sg13g2_decap_8
XFILLER_34_860 VPWR VGND sg13g2_decap_8
XFILLER_21_521 VPWR VGND sg13g2_decap_8
XFILLER_20_46 VPWR VGND sg13g2_decap_8
XFILLER_1_915 VPWR VGND sg13g2_decap_8
XFILLER_49_919 VPWR VGND sg13g2_decap_8
Xhold11 mac1.sum_lvl1_ff\[32\] VPWR VGND net35 sg13g2_dlygate4sd3_1
XFILLER_0_469 VPWR VGND sg13g2_decap_8
Xhold22 DP_1.matrix\[1\] VPWR VGND net46 sg13g2_dlygate4sd3_1
Xhold33 DP_3.matrix\[10\] VPWR VGND net57 sg13g2_dlygate4sd3_1
Xhold44 _002_ VPWR VGND net94 sg13g2_dlygate4sd3_1
Xhold55 DP_1.matrix\[46\] VPWR VGND net105 sg13g2_dlygate4sd3_1
XFILLER_29_610 VPWR VGND sg13g2_decap_8
Xhold77 DP_3.matrix\[72\] VPWR VGND net127 sg13g2_dlygate4sd3_1
Xhold66 _020_ VPWR VGND net116 sg13g2_dlygate4sd3_1
Xhold88 DP_1.matrix\[45\] VPWR VGND net138 sg13g2_dlygate4sd3_1
XFILLER_29_99 VPWR VGND sg13g2_decap_8
XFILLER_28_131 VPWR VGND sg13g2_decap_8
Xhold99 DP_3.matrix\[27\] VPWR VGND net149 sg13g2_dlygate4sd3_1
XFILLER_45_21 VPWR VGND sg13g2_decap_8
XFILLER_17_838 VPWR VGND sg13g2_decap_8
XFILLER_28_142 VPWR VGND sg13g2_fill_2
XFILLER_29_687 VPWR VGND sg13g2_decap_8
X_591_ net68 VGND VPWR _131_ DP_4.matrix\[28\] clknet_5_8__leaf_clk sg13g2_dfrbpq_1
XFILLER_43_134 VPWR VGND sg13g2_decap_8
XFILLER_16_348 VPWR VGND sg13g2_decap_8
XFILLER_44_668 VPWR VGND sg13g2_decap_8
XFILLER_12_510 VPWR VGND sg13g2_fill_1
XFILLER_25_893 VPWR VGND sg13g2_decap_8
XFILLER_40_841 VPWR VGND sg13g2_decap_8
XFILLER_12_576 VPWR VGND sg13g2_decap_8
XFILLER_4_731 VPWR VGND sg13g2_decap_8
XFILLER_3_285 VPWR VGND sg13g2_decap_8
XFILLER_6_1019 VPWR VGND sg13g2_decap_8
XFILLER_48_930 VPWR VGND sg13g2_decap_8
XFILLER_47_462 VPWR VGND sg13g2_decap_8
XFILLER_35_613 VPWR VGND sg13g2_decap_8
XFILLER_19_186 VPWR VGND sg13g2_decap_8
XFILLER_34_123 VPWR VGND sg13g2_fill_2
XFILLER_37_1010 VPWR VGND sg13g2_decap_8
XFILLER_16_893 VPWR VGND sg13g2_decap_8
XFILLER_30_351 VPWR VGND sg13g2_decap_8
XFILLER_31_874 VPWR VGND sg13g2_decap_8
XFILLER_44_1025 VPWR VGND sg13g2_decap_4
Xheichips25_template_13 VPWR VGND uo_out[4] sg13g2_tielo
Xheichips25_template_24 VPWR VGND uio_oe[7] sg13g2_tiehi
XFILLER_39_952 VPWR VGND sg13g2_decap_8
XFILLER_26_613 VPWR VGND sg13g2_decap_8
XFILLER_38_451 VPWR VGND sg13g2_decap_8
XFILLER_38_495 VPWR VGND sg13g2_decap_8
XFILLER_14_819 VPWR VGND sg13g2_decap_8
XFILLER_25_156 VPWR VGND sg13g2_decap_8
XFILLER_41_638 VPWR VGND sg13g2_decap_8
XFILLER_22_830 VPWR VGND sg13g2_decap_8
XFILLER_40_159 VPWR VGND sg13g2_decap_8
XFILLER_21_351 VPWR VGND sg13g2_decap_8
XFILLER_5_506 VPWR VGND sg13g2_decap_8
XFILLER_31_56 VPWR VGND sg13g2_decap_8
XFILLER_5_539 VPWR VGND sg13g2_decap_8
XFILLER_1_712 VPWR VGND sg13g2_decap_8
XFILLER_49_716 VPWR VGND sg13g2_decap_8
XFILLER_0_266 VPWR VGND sg13g2_decap_8
XFILLER_1_789 VPWR VGND sg13g2_decap_8
XFILLER_45_933 VPWR VGND sg13g2_decap_8
XFILLER_17_635 VPWR VGND sg13g2_decap_8
XFILLER_44_465 VPWR VGND sg13g2_decap_8
X_574_ net71 VGND VPWR _114_ DP_3.matrix\[36\] clknet_5_12__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_627 VPWR VGND sg13g2_decap_8
XFILLER_9_801 VPWR VGND sg13g2_decap_8
XFILLER_13_830 VPWR VGND sg13g2_decap_8
XFILLER_25_690 VPWR VGND sg13g2_decap_8
XFILLER_31_126 VPWR VGND sg13g2_decap_8
XFILLER_12_351 VPWR VGND sg13g2_decap_8
XFILLER_9_878 VPWR VGND sg13g2_decap_8
XFILLER_35_410 VPWR VGND sg13g2_decap_8
XFILLER_36_933 VPWR VGND sg13g2_decap_8
XFILLER_35_476 VPWR VGND sg13g2_decap_4
XFILLER_16_690 VPWR VGND sg13g2_decap_8
XFILLER_22_148 VPWR VGND sg13g2_decap_8
XFILLER_31_671 VPWR VGND sg13g2_decap_8
XFILLER_30_170 VPWR VGND sg13g2_decap_8
XFILLER_7_91 VPWR VGND sg13g2_decap_8
XFILLER_27_911 VPWR VGND sg13g2_decap_8
XFILLER_27_988 VPWR VGND sg13g2_decap_8
XFILLER_42_925 VPWR VGND sg13g2_decap_8
XFILLER_14_616 VPWR VGND sg13g2_decap_8
XFILLER_26_67 VPWR VGND sg13g2_decap_8
XFILLER_26_487 VPWR VGND sg13g2_decap_8
X_290_ mac1.sum_lvl1_ff\[17\] mac1.sum_lvl1_ff\[25\] _171_ VPWR VGND sg13g2_xor2_1
XFILLER_13_137 VPWR VGND sg13g2_decap_8
XFILLER_41_468 VPWR VGND sg13g2_decap_8
XFILLER_42_66 VPWR VGND sg13g2_decap_8
XFILLER_10_844 VPWR VGND sg13g2_decap_8
XFILLER_6_837 VPWR VGND sg13g2_decap_8
XFILLER_5_303 VPWR VGND sg13g2_decap_8
XFILLER_49_513 VPWR VGND sg13g2_decap_8
XFILLER_1_586 VPWR VGND sg13g2_decap_8
XFILLER_18_900 VPWR VGND sg13g2_decap_8
XFILLER_45_730 VPWR VGND sg13g2_decap_8
XFILLER_18_977 VPWR VGND sg13g2_decap_8
XFILLER_29_292 VPWR VGND sg13g2_fill_1
X_557_ net76 VGND VPWR _097_ DP_2.matrix\[37\] clknet_5_23__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_476 VPWR VGND sg13g2_decap_8
XFILLER_33_958 VPWR VGND sg13g2_decap_8
X_488_ net60 VGND VPWR net169 mac1.total_sum\[2\] clknet_5_5__leaf_clk sg13g2_dfrbpq_1
XFILLER_20_619 VPWR VGND sg13g2_decap_8
XFILLER_9_675 VPWR VGND sg13g2_decap_8
XFILLER_8_141 VPWR VGND sg13g2_decap_8
XFILLER_8_196 VPWR VGND sg13g2_decap_8
XFILLER_5_892 VPWR VGND sg13g2_decap_8
XFILLER_4_391 VPWR VGND sg13g2_fill_1
XFILLER_36_730 VPWR VGND sg13g2_decap_8
XFILLER_35_273 VPWR VGND sg13g2_decap_8
XFILLER_24_958 VPWR VGND sg13g2_decap_8
XFILLER_32_991 VPWR VGND sg13g2_decap_8
XFILLER_12_25 VPWR VGND sg13g2_fill_2
XFILLER_12_69 VPWR VGND sg13g2_decap_8
XFILLER_3_818 VPWR VGND sg13g2_decap_8
XFILLER_2_328 VPWR VGND sg13g2_decap_8
Xhold152 _021_ VPWR VGND net202 sg13g2_dlygate4sd3_1
Xhold141 mac2.products_ff\[0\] VPWR VGND net191 sg13g2_dlygate4sd3_1
Xhold130 _025_ VPWR VGND net180 sg13g2_dlygate4sd3_1
XFILLER_26_240 VPWR VGND sg13g2_decap_8
XFILLER_42_722 VPWR VGND sg13g2_decap_8
X_411_ net106 _105_ VPWR VGND sg13g2_buf_1
XFILLER_15_925 VPWR VGND sg13g2_decap_8
XFILLER_27_785 VPWR VGND sg13g2_decap_8
XFILLER_18_1019 VPWR VGND sg13g2_decap_8
XFILLER_30_906 VPWR VGND sg13g2_decap_8
XFILLER_42_799 VPWR VGND sg13g2_decap_8
XFILLER_14_468 VPWR VGND sg13g2_decap_8
XFILLER_14_479 VPWR VGND sg13g2_fill_2
X_342_ _200_ net128 net97 VPWR VGND sg13g2_nand2_1
X_273_ _162_ net183 net111 VPWR VGND sg13g2_nand2_1
XFILLER_10_641 VPWR VGND sg13g2_decap_8
XFILLER_6_634 VPWR VGND sg13g2_decap_8
XFILLER_2_873 VPWR VGND sg13g2_decap_8
XFILLER_49_310 VPWR VGND sg13g2_decap_8
XFILLER_1_383 VPWR VGND sg13g2_decap_8
XFILLER_49_387 VPWR VGND sg13g2_decap_8
XFILLER_37_527 VPWR VGND sg13g2_decap_8
XFILLER_18_774 VPWR VGND sg13g2_decap_8
XFILLER_33_755 VPWR VGND sg13g2_decap_8
XFILLER_21_939 VPWR VGND sg13g2_decap_8
XFILLER_14_980 VPWR VGND sg13g2_decap_8
XFILLER_20_416 VPWR VGND sg13g2_decap_8
XFILLER_4_81 VPWR VGND sg13g2_decap_8
XFILLER_24_755 VPWR VGND sg13g2_decap_8
XFILLER_12_928 VPWR VGND sg13g2_decap_8
XFILLER_23_254 VPWR VGND sg13g2_fill_1
XFILLER_11_449 VPWR VGND sg13g2_decap_8
XFILLER_20_983 VPWR VGND sg13g2_decap_8
XFILLER_3_615 VPWR VGND sg13g2_decap_8
XFILLER_2_114 VPWR VGND sg13g2_fill_1
XFILLER_48_21 VPWR VGND sg13g2_decap_8
XFILLER_47_847 VPWR VGND sg13g2_decap_8
XFILLER_48_98 VPWR VGND sg13g2_decap_8
XFILLER_46_324 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_15_722 VPWR VGND sg13g2_decap_8
XFILLER_27_582 VPWR VGND sg13g2_decap_8
XFILLER_9_15 VPWR VGND sg13g2_fill_2
XFILLER_14_265 VPWR VGND sg13g2_decap_8
XFILLER_30_703 VPWR VGND sg13g2_decap_8
XFILLER_42_596 VPWR VGND sg13g2_decap_8
XFILLER_9_48 VPWR VGND sg13g2_decap_8
X_325_ _189_ _188_ _069_ VPWR VGND sg13g2_xor2_1
XFILLER_15_799 VPWR VGND sg13g2_decap_8
Xfanout80 net81 net80 VPWR VGND sg13g2_buf_8
XFILLER_7_932 VPWR VGND sg13g2_decap_8
XFILLER_6_420 VPWR VGND sg13g2_decap_8
X_256_ _001_ _150_ _151_ VPWR VGND sg13g2_xnor2_1
XFILLER_6_464 VPWR VGND sg13g2_fill_1
XFILLER_2_670 VPWR VGND sg13g2_decap_8
XFILLER_1_180 VPWR VGND sg13g2_decap_8
XFILLER_38_803 VPWR VGND sg13g2_decap_8
XFILLER_49_184 VPWR VGND sg13g2_decap_8
XFILLER_33_552 VPWR VGND sg13g2_decap_8
XFILLER_21_736 VPWR VGND sg13g2_decap_8
XFILLER_20_235 VPWR VGND sg13g2_decap_8
XFILLER_9_280 VPWR VGND sg13g2_decap_8
XFILLER_47_1001 VPWR VGND sg13g2_decap_8
XFILLER_18_46 VPWR VGND sg13g2_decap_8
XFILLER_29_869 VPWR VGND sg13g2_decap_8
XFILLER_43_316 VPWR VGND sg13g2_decap_8
XFILLER_37_891 VPWR VGND sg13g2_decap_8
XFILLER_24_552 VPWR VGND sg13g2_decap_8
XFILLER_11_202 VPWR VGND sg13g2_decap_8
XFILLER_12_725 VPWR VGND sg13g2_decap_8
Xclkload0 VPWR clkload0/Y clknet_5_7__leaf_clk VGND sg13g2_inv_1
XFILLER_20_780 VPWR VGND sg13g2_decap_8
XFILLER_4_913 VPWR VGND sg13g2_decap_8
XFILLER_3_478 VPWR VGND sg13g2_decap_8
Xclkbuf_5_29__f_clk clknet_4_14_0_clk clknet_5_29__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_47_644 VPWR VGND sg13g2_decap_8
XFILLER_19_346 VPWR VGND sg13g2_decap_8
XFILLER_46_154 VPWR VGND sg13g2_decap_4
XFILLER_30_500 VPWR VGND sg13g2_decap_8
XFILLER_42_393 VPWR VGND sg13g2_decap_8
XFILLER_30_577 VPWR VGND sg13g2_decap_8
X_308_ mac2.products_ff\[103\] mac2.products_ff\[120\] _181_ VPWR VGND sg13g2_xor2_1
X_239_ net150 net138 _052_ VPWR VGND sg13g2_and2_1
XFILLER_6_283 VPWR VGND sg13g2_decap_8
XFILLER_38_600 VPWR VGND sg13g2_decap_8
XFILLER_38_677 VPWR VGND sg13g2_decap_8
XFILLER_37_198 VPWR VGND sg13g2_decap_8
XFILLER_18_390 VPWR VGND sg13g2_decap_8
XFILLER_21_500 VPWR VGND sg13g2_decap_8
XFILLER_40_319 VPWR VGND sg13g2_decap_8
XFILLER_14_1022 VPWR VGND sg13g2_decap_8
XFILLER_20_25 VPWR VGND sg13g2_decap_8
Xhold12 mac1.sum_lvl2_ff\[8\] VPWR VGND net36 sg13g2_dlygate4sd3_1
XFILLER_0_448 VPWR VGND sg13g2_decap_8
Xhold23 DP_1.matrix\[28\] VPWR VGND net47 sg13g2_dlygate4sd3_1
XFILLER_48_419 VPWR VGND sg13g2_decap_8
Xhold34 DP_3.matrix\[37\] VPWR VGND net58 sg13g2_dlygate4sd3_1
Xhold56 DP_2.matrix\[73\] VPWR VGND net106 sg13g2_dlygate4sd3_1
Xhold45 mac2.products_ff\[17\] VPWR VGND net95 sg13g2_dlygate4sd3_1
Xhold89 DP_1.matrix\[36\] VPWR VGND net139 sg13g2_dlygate4sd3_1
Xhold67 DP_1.matrix\[27\] VPWR VGND net117 sg13g2_dlygate4sd3_1
Xhold78 DP_2.matrix\[9\] VPWR VGND net128 sg13g2_dlygate4sd3_1
XFILLER_17_817 VPWR VGND sg13g2_decap_8
XFILLER_29_666 VPWR VGND sg13g2_decap_8
X_590_ net68 VGND VPWR _130_ DP_4.matrix\[27\] clknet_5_10__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_647 VPWR VGND sg13g2_decap_8
XFILLER_43_113 VPWR VGND sg13g2_decap_8
XFILLER_31_308 VPWR VGND sg13g2_decap_8
XFILLER_32_809 VPWR VGND sg13g2_decap_8
XFILLER_25_872 VPWR VGND sg13g2_decap_8
XFILLER_40_820 VPWR VGND sg13g2_decap_8
XFILLER_40_897 VPWR VGND sg13g2_decap_8
XFILLER_8_559 VPWR VGND sg13g2_decap_8
XFILLER_12_599 VPWR VGND sg13g2_decap_8
XFILLER_4_710 VPWR VGND sg13g2_decap_8
XFILLER_4_787 VPWR VGND sg13g2_decap_8
XFILLER_47_441 VPWR VGND sg13g2_decap_8
XFILLER_48_986 VPWR VGND sg13g2_decap_8
XFILLER_19_165 VPWR VGND sg13g2_decap_8
XFILLER_34_102 VPWR VGND sg13g2_decap_8
XFILLER_35_669 VPWR VGND sg13g2_decap_8
XFILLER_16_872 VPWR VGND sg13g2_decap_8
XFILLER_15_382 VPWR VGND sg13g2_decap_8
XFILLER_30_330 VPWR VGND sg13g2_decap_8
XFILLER_31_853 VPWR VGND sg13g2_decap_8
XFILLER_44_1004 VPWR VGND sg13g2_decap_8
Xclkbuf_5_12__f_clk clknet_4_6_0_clk clknet_5_12__leaf_clk VPWR VGND sg13g2_buf_8
Xheichips25_template_14 VPWR VGND uo_out[5] sg13g2_tielo
XFILLER_39_931 VPWR VGND sg13g2_decap_8
XFILLER_26_669 VPWR VGND sg13g2_decap_8
XFILLER_15_47 VPWR VGND sg13g2_decap_8
XFILLER_41_617 VPWR VGND sg13g2_decap_8
XFILLER_33_190 VPWR VGND sg13g2_fill_1
XFILLER_40_138 VPWR VGND sg13g2_decap_8
XFILLER_22_886 VPWR VGND sg13g2_decap_8
XFILLER_31_35 VPWR VGND sg13g2_decap_8
XFILLER_0_245 VPWR VGND sg13g2_decap_8
XFILLER_1_768 VPWR VGND sg13g2_decap_8
XFILLER_48_205 VPWR VGND sg13g2_decap_8
XFILLER_29_430 VPWR VGND sg13g2_decap_8
XFILLER_45_912 VPWR VGND sg13g2_decap_8
XFILLER_17_614 VPWR VGND sg13g2_decap_8
XFILLER_29_474 VPWR VGND sg13g2_decap_8
XFILLER_45_989 VPWR VGND sg13g2_decap_8
XFILLER_44_444 VPWR VGND sg13g2_decap_8
XFILLER_32_606 VPWR VGND sg13g2_decap_8
X_573_ net68 VGND VPWR _113_ DP_3.matrix\[28\] clknet_5_10__leaf_clk sg13g2_dfrbpq_1
XFILLER_31_105 VPWR VGND sg13g2_decap_8
XFILLER_13_886 VPWR VGND sg13g2_decap_8
XFILLER_9_857 VPWR VGND sg13g2_decap_8
XFILLER_40_694 VPWR VGND sg13g2_decap_8
XFILLER_21_90 VPWR VGND sg13g2_decap_8
XFILLER_4_584 VPWR VGND sg13g2_decap_8
XFILLER_39_249 VPWR VGND sg13g2_decap_4
XFILLER_11_4 VPWR VGND sg13g2_decap_8
XFILLER_36_912 VPWR VGND sg13g2_decap_8
XFILLER_48_783 VPWR VGND sg13g2_decap_8
XFILLER_47_282 VPWR VGND sg13g2_decap_8
XFILLER_47_293 VPWR VGND sg13g2_fill_2
XFILLER_36_989 VPWR VGND sg13g2_decap_8
XFILLER_23_639 VPWR VGND sg13g2_decap_8
XFILLER_31_650 VPWR VGND sg13g2_decap_8
XFILLER_7_70 VPWR VGND sg13g2_decap_8
XFILLER_38_260 VPWR VGND sg13g2_fill_1
XFILLER_42_904 VPWR VGND sg13g2_decap_8
XFILLER_26_46 VPWR VGND sg13g2_decap_8
XFILLER_27_967 VPWR VGND sg13g2_decap_8
XFILLER_26_466 VPWR VGND sg13g2_decap_8
XFILLER_13_116 VPWR VGND sg13g2_decap_8
XFILLER_41_447 VPWR VGND sg13g2_decap_8
XFILLER_9_109 VPWR VGND sg13g2_decap_8
XFILLER_10_823 VPWR VGND sg13g2_decap_8
XFILLER_21_160 VPWR VGND sg13g2_decap_4
XFILLER_22_683 VPWR VGND sg13g2_decap_8
XFILLER_42_45 VPWR VGND sg13g2_decap_8
XFILLER_6_816 VPWR VGND sg13g2_decap_8
XFILLER_5_359 VPWR VGND sg13g2_decap_8
XFILLER_3_39 VPWR VGND sg13g2_decap_8
XFILLER_1_565 VPWR VGND sg13g2_decap_8
XFILLER_49_569 VPWR VGND sg13g2_decap_8
XFILLER_37_709 VPWR VGND sg13g2_decap_8
XFILLER_17_411 VPWR VGND sg13g2_fill_2
XFILLER_17_422 VPWR VGND sg13g2_fill_2
XFILLER_17_455 VPWR VGND sg13g2_decap_8
XFILLER_18_956 VPWR VGND sg13g2_decap_8
XFILLER_45_786 VPWR VGND sg13g2_decap_8
X_556_ net77 VGND VPWR _096_ DP_2.matrix\[36\] clknet_5_23__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_403 VPWR VGND sg13g2_fill_2
XFILLER_33_937 VPWR VGND sg13g2_decap_8
X_487_ net60 VGND VPWR net204 mac1.total_sum\[1\] clknet_5_5__leaf_clk sg13g2_dfrbpq_1
XFILLER_34_1014 VPWR VGND sg13g2_decap_8
XFILLER_8_120 VPWR VGND sg13g2_decap_8
XFILLER_13_683 VPWR VGND sg13g2_decap_8
XFILLER_41_981 VPWR VGND sg13g2_decap_8
XFILLER_9_654 VPWR VGND sg13g2_decap_8
XFILLER_12_182 VPWR VGND sg13g2_decap_8
XFILLER_5_871 VPWR VGND sg13g2_decap_8
XFILLER_48_580 VPWR VGND sg13g2_decap_8
XFILLER_24_937 VPWR VGND sg13g2_decap_8
XFILLER_35_252 VPWR VGND sg13g2_decap_8
XFILLER_36_786 VPWR VGND sg13g2_decap_8
XFILLER_23_469 VPWR VGND sg13g2_decap_8
XFILLER_32_970 VPWR VGND sg13g2_decap_8
XFILLER_12_48 VPWR VGND sg13g2_decap_8
Xhold153 mac1.sum_lvl3_ff\[0\] VPWR VGND net203 sg13g2_dlygate4sd3_1
XFILLER_2_307 VPWR VGND sg13g2_decap_8
Xhold120 mac2.sum_lvl3_ff\[3\] VPWR VGND net170 sg13g2_dlygate4sd3_1
Xhold142 _023_ VPWR VGND net192 sg13g2_dlygate4sd3_1
Xhold131 mac2.products_ff\[68\] VPWR VGND net181 sg13g2_dlygate4sd3_1
XFILLER_15_904 VPWR VGND sg13g2_decap_8
XFILLER_37_78 VPWR VGND sg13g2_decap_8
XFILLER_42_701 VPWR VGND sg13g2_decap_8
X_410_ net118 _104_ VPWR VGND sg13g2_buf_1
XFILLER_27_764 VPWR VGND sg13g2_decap_8
XFILLER_14_447 VPWR VGND sg13g2_decap_8
XFILLER_26_296 VPWR VGND sg13g2_decap_8
X_341_ _199_ _198_ _043_ VPWR VGND sg13g2_xor2_1
XFILLER_42_778 VPWR VGND sg13g2_decap_8
XFILLER_41_244 VPWR VGND sg13g2_decap_8
XFILLER_10_620 VPWR VGND sg13g2_decap_8
X_272_ net93 mac1.products_ff\[17\] _002_ VPWR VGND sg13g2_xor2_1
XFILLER_6_613 VPWR VGND sg13g2_decap_8
XFILLER_10_697 VPWR VGND sg13g2_decap_8
XFILLER_5_189 VPWR VGND sg13g2_decap_8
XFILLER_2_852 VPWR VGND sg13g2_decap_8
XFILLER_1_362 VPWR VGND sg13g2_decap_8
XFILLER_49_366 VPWR VGND sg13g2_decap_8
XFILLER_37_506 VPWR VGND sg13g2_decap_8
XFILLER_18_753 VPWR VGND sg13g2_decap_8
XFILLER_45_583 VPWR VGND sg13g2_decap_8
XFILLER_32_200 VPWR VGND sg13g2_decap_8
XFILLER_33_734 VPWR VGND sg13g2_decap_8
X_539_ net77 VGND VPWR _079_ DP_1.matrix\[37\] clknet_5_23__leaf_clk sg13g2_dfrbpq_1
XFILLER_21_918 VPWR VGND sg13g2_decap_8
XFILLER_32_288 VPWR VGND sg13g2_decap_8
XFILLER_9_451 VPWR VGND sg13g2_decap_8
XFILLER_9_484 VPWR VGND sg13g2_decap_8
XFILLER_4_60 VPWR VGND sg13g2_decap_8
XFILLER_28_539 VPWR VGND sg13g2_decap_8
XFILLER_23_222 VPWR VGND sg13g2_decap_8
XFILLER_24_734 VPWR VGND sg13g2_decap_8
XFILLER_36_583 VPWR VGND sg13g2_decap_8
XFILLER_12_907 VPWR VGND sg13g2_decap_8
XFILLER_11_428 VPWR VGND sg13g2_decap_8
XFILLER_17_1020 VPWR VGND sg13g2_decap_8
XFILLER_20_962 VPWR VGND sg13g2_decap_8
XFILLER_2_137 VPWR VGND sg13g2_fill_2
XFILLER_47_826 VPWR VGND sg13g2_decap_8
XFILLER_48_77 VPWR VGND sg13g2_decap_8
XFILLER_15_701 VPWR VGND sg13g2_decap_8
XFILLER_27_561 VPWR VGND sg13g2_decap_8
XFILLER_14_244 VPWR VGND sg13g2_decap_8
XFILLER_15_778 VPWR VGND sg13g2_decap_8
XFILLER_42_575 VPWR VGND sg13g2_decap_8
X_324_ _189_ net133 net106 VPWR VGND sg13g2_nand2_1
XFILLER_30_759 VPWR VGND sg13g2_decap_8
X_255_ mac2.sum_lvl2_ff\[5\] mac2.sum_lvl2_ff\[1\] _151_ VPWR VGND sg13g2_xor2_1
Xfanout81 net84 net81 VPWR VGND sg13g2_buf_8
Xfanout70 net71 net70 VPWR VGND sg13g2_buf_8
XFILLER_7_911 VPWR VGND sg13g2_decap_8
XFILLER_11_984 VPWR VGND sg13g2_decap_8
XFILLER_31_1028 VPWR VGND sg13g2_fill_1
XFILLER_10_494 VPWR VGND sg13g2_decap_8
XFILLER_7_988 VPWR VGND sg13g2_decap_8
XFILLER_6_476 VPWR VGND sg13g2_fill_1
XFILLER_43_7 VPWR VGND sg13g2_decap_8
XFILLER_9_1018 VPWR VGND sg13g2_decap_8
XFILLER_49_163 VPWR VGND sg13g2_decap_8
XFILLER_38_859 VPWR VGND sg13g2_decap_8
XFILLER_37_369 VPWR VGND sg13g2_decap_8
XFILLER_33_531 VPWR VGND sg13g2_decap_8
XFILLER_45_391 VPWR VGND sg13g2_decap_8
XFILLER_20_214 VPWR VGND sg13g2_decap_8
XFILLER_21_715 VPWR VGND sg13g2_decap_8
XFILLER_18_25 VPWR VGND sg13g2_decap_8
XFILLER_28_314 VPWR VGND sg13g2_fill_1
XFILLER_29_848 VPWR VGND sg13g2_decap_8
XFILLER_44_829 VPWR VGND sg13g2_decap_8
XFILLER_28_369 VPWR VGND sg13g2_decap_8
XFILLER_37_870 VPWR VGND sg13g2_decap_8
XFILLER_12_704 VPWR VGND sg13g2_decap_8
XFILLER_24_531 VPWR VGND sg13g2_decap_8
XFILLER_34_35 VPWR VGND sg13g2_decap_4
XFILLER_34_68 VPWR VGND sg13g2_decap_8
Xclkload1 VPWR clkload1/Y clknet_5_11__leaf_clk VGND sg13g2_inv_1
XFILLER_4_969 VPWR VGND sg13g2_decap_8
XFILLER_3_457 VPWR VGND sg13g2_decap_8
XFILLER_47_623 VPWR VGND sg13g2_decap_8
XFILLER_46_133 VPWR VGND sg13g2_decap_8
XFILLER_34_317 VPWR VGND sg13g2_decap_4
XFILLER_43_895 VPWR VGND sg13g2_decap_8
XFILLER_42_372 VPWR VGND sg13g2_decap_8
XFILLER_15_564 VPWR VGND sg13g2_fill_1
XFILLER_30_556 VPWR VGND sg13g2_decap_8
X_307_ _180_ net195 net123 VPWR VGND sg13g2_nand2_1
XFILLER_11_781 VPWR VGND sg13g2_decap_8
X_238_ net122 net139 _050_ VPWR VGND sg13g2_and2_1
XFILLER_7_785 VPWR VGND sg13g2_decap_8
XFILLER_6_262 VPWR VGND sg13g2_decap_8
XFILLER_38_656 VPWR VGND sg13g2_decap_8
XFILLER_1_83 VPWR VGND sg13g2_fill_2
XFILLER_19_881 VPWR VGND sg13g2_decap_8
XFILLER_37_177 VPWR VGND sg13g2_decap_8
XFILLER_34_895 VPWR VGND sg13g2_decap_8
XFILLER_21_556 VPWR VGND sg13g2_decap_4
XFILLER_14_1001 VPWR VGND sg13g2_decap_8
XFILLER_0_427 VPWR VGND sg13g2_decap_8
Xhold13 DP_4.matrix\[55\] VPWR VGND net37 sg13g2_dlygate4sd3_1
Xhold35 DP_2.matrix\[46\] VPWR VGND net59 sg13g2_dlygate4sd3_1
XFILLER_29_68 VPWR VGND sg13g2_decap_4
Xhold46 _022_ VPWR VGND net96 sg13g2_dlygate4sd3_1
Xhold24 DP_2.matrix\[10\] VPWR VGND net48 sg13g2_dlygate4sd3_1
Xhold68 DP_2.matrix\[72\] VPWR VGND net118 sg13g2_dlygate4sd3_1
Xhold79 DP_2.matrix\[18\] VPWR VGND net129 sg13g2_dlygate4sd3_1
XFILLER_21_1016 VPWR VGND sg13g2_decap_8
XFILLER_21_1027 VPWR VGND sg13g2_fill_2
XFILLER_29_645 VPWR VGND sg13g2_decap_8
Xhold57 mac2.sum_lvl1_ff\[8\] VPWR VGND net107 sg13g2_dlygate4sd3_1
XFILLER_44_626 VPWR VGND sg13g2_decap_8
XFILLER_16_317 VPWR VGND sg13g2_decap_8
XFILLER_16_328 VPWR VGND sg13g2_fill_1
XFILLER_28_188 VPWR VGND sg13g2_decap_8
XFILLER_25_851 VPWR VGND sg13g2_decap_8
XFILLER_24_383 VPWR VGND sg13g2_decap_8
XFILLER_40_876 VPWR VGND sg13g2_decap_8
XFILLER_8_538 VPWR VGND sg13g2_decap_8
XFILLER_6_39 VPWR VGND sg13g2_decap_8
XFILLER_4_766 VPWR VGND sg13g2_decap_8
XFILLER_0_994 VPWR VGND sg13g2_decap_8
XFILLER_48_965 VPWR VGND sg13g2_decap_8
XFILLER_19_144 VPWR VGND sg13g2_decap_8
XFILLER_47_497 VPWR VGND sg13g2_decap_8
XFILLER_35_648 VPWR VGND sg13g2_decap_8
XFILLER_16_851 VPWR VGND sg13g2_decap_8
XFILLER_34_125 VPWR VGND sg13g2_fill_1
XFILLER_15_361 VPWR VGND sg13g2_decap_8
XFILLER_43_692 VPWR VGND sg13g2_decap_8
XFILLER_42_180 VPWR VGND sg13g2_fill_1
XFILLER_31_832 VPWR VGND sg13g2_decap_8
XFILLER_7_582 VPWR VGND sg13g2_decap_8
XFILLER_32_0 VPWR VGND sg13g2_decap_8
XFILLER_39_910 VPWR VGND sg13g2_decap_8
Xheichips25_template_15 VPWR VGND uo_out[6] sg13g2_tielo
XFILLER_38_420 VPWR VGND sg13g2_decap_8
XFILLER_39_987 VPWR VGND sg13g2_decap_8
XFILLER_26_648 VPWR VGND sg13g2_decap_8
XFILLER_25_125 VPWR VGND sg13g2_decap_4
XFILLER_13_309 VPWR VGND sg13g2_decap_8
XFILLER_15_15 VPWR VGND sg13g2_fill_1
XFILLER_40_117 VPWR VGND sg13g2_decap_8
XFILLER_34_692 VPWR VGND sg13g2_decap_8
XFILLER_22_865 VPWR VGND sg13g2_decap_8
XFILLER_31_14 VPWR VGND sg13g2_decap_8
XFILLER_0_224 VPWR VGND sg13g2_decap_8
XFILLER_1_747 VPWR VGND sg13g2_decap_8
XFILLER_48_239 VPWR VGND sg13g2_decap_8
XFILLER_44_423 VPWR VGND sg13g2_decap_8
X_572_ net68 VGND VPWR _112_ DP_3.matrix\[27\] clknet_5_8__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_968 VPWR VGND sg13g2_decap_8
XFILLER_16_169 VPWR VGND sg13g2_decap_8
XFILLER_24_180 VPWR VGND sg13g2_decap_8
XFILLER_9_836 VPWR VGND sg13g2_decap_8
XFILLER_13_865 VPWR VGND sg13g2_decap_8
XFILLER_12_386 VPWR VGND sg13g2_decap_8
XFILLER_40_673 VPWR VGND sg13g2_decap_8
XFILLER_4_541 VPWR VGND sg13g2_decap_8
XFILLER_4_574 VPWR VGND sg13g2_fill_1
XFILLER_0_791 VPWR VGND sg13g2_decap_8
XFILLER_39_217 VPWR VGND sg13g2_decap_4
XFILLER_48_762 VPWR VGND sg13g2_decap_8
XFILLER_36_968 VPWR VGND sg13g2_decap_8
XFILLER_23_618 VPWR VGND sg13g2_decap_8
XFILLER_44_990 VPWR VGND sg13g2_decap_8
XFILLER_11_1026 VPWR VGND sg13g2_fill_2
XFILLER_7_390 VPWR VGND sg13g2_decap_4
XFILLER_27_946 VPWR VGND sg13g2_decap_8
XFILLER_39_784 VPWR VGND sg13g2_decap_8
XFILLER_26_25 VPWR VGND sg13g2_decap_8
XFILLER_26_445 VPWR VGND sg13g2_decap_8
XFILLER_41_426 VPWR VGND sg13g2_decap_8
XFILLER_41_437 VPWR VGND sg13g2_fill_2
XFILLER_10_802 VPWR VGND sg13g2_decap_8
XFILLER_22_662 VPWR VGND sg13g2_decap_8
XFILLER_10_879 VPWR VGND sg13g2_decap_8
XFILLER_5_338 VPWR VGND sg13g2_decap_8
XFILLER_3_18 VPWR VGND sg13g2_decap_8
XFILLER_1_544 VPWR VGND sg13g2_decap_8
XFILLER_49_548 VPWR VGND sg13g2_decap_8
XFILLER_18_935 VPWR VGND sg13g2_decap_8
XFILLER_36_209 VPWR VGND sg13g2_decap_8
XFILLER_17_434 VPWR VGND sg13g2_decap_8
XFILLER_45_765 VPWR VGND sg13g2_decap_8
XFILLER_44_253 VPWR VGND sg13g2_fill_2
X_555_ net66 VGND VPWR _095_ DP_2.matrix\[28\] clknet_5_24__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_916 VPWR VGND sg13g2_decap_8
XFILLER_44_297 VPWR VGND sg13g2_decap_8
X_486_ net60 VGND VPWR net166 mac1.total_sum\[0\] clknet_5_6__leaf_clk sg13g2_dfrbpq_1
XFILLER_16_80 VPWR VGND sg13g2_decap_8
XFILLER_13_662 VPWR VGND sg13g2_decap_8
XFILLER_32_459 VPWR VGND sg13g2_decap_8
XFILLER_41_960 VPWR VGND sg13g2_decap_8
XFILLER_9_633 VPWR VGND sg13g2_decap_8
XFILLER_5_850 VPWR VGND sg13g2_decap_8
XFILLER_4_382 VPWR VGND sg13g2_decap_8
XFILLER_24_916 VPWR VGND sg13g2_decap_8
XFILLER_36_765 VPWR VGND sg13g2_decap_8
XFILLER_23_448 VPWR VGND sg13g2_decap_8
XFILLER_12_27 VPWR VGND sg13g2_fill_1
Xhold110 DP_2.matrix\[27\] VPWR VGND net160 sg13g2_dlygate4sd3_1
Xhold132 _027_ VPWR VGND net182 sg13g2_dlygate4sd3_1
Xhold143 mac1.products_ff\[102\] VPWR VGND net193 sg13g2_dlygate4sd3_1
Xhold121 _173_ VPWR VGND net171 sg13g2_dlygate4sd3_1
Xhold154 _018_ VPWR VGND net204 sg13g2_dlygate4sd3_1
XFILLER_46_529 VPWR VGND sg13g2_decap_8
XFILLER_2_1013 VPWR VGND sg13g2_decap_8
XFILLER_18_209 VPWR VGND sg13g2_decap_8
XFILLER_37_35 VPWR VGND sg13g2_fill_2
XFILLER_37_57 VPWR VGND sg13g2_decap_8
XFILLER_39_581 VPWR VGND sg13g2_decap_8
XFILLER_27_743 VPWR VGND sg13g2_decap_8
XFILLER_14_426 VPWR VGND sg13g2_decap_8
X_340_ _199_ net159 net38 VPWR VGND sg13g2_nand2_1
XFILLER_41_223 VPWR VGND sg13g2_decap_8
XFILLER_42_757 VPWR VGND sg13g2_decap_8
XFILLER_23_982 VPWR VGND sg13g2_decap_8
X_271_ _003_ _160_ _161_ VPWR VGND sg13g2_xnor2_1
XFILLER_10_676 VPWR VGND sg13g2_decap_8
XFILLER_5_102 VPWR VGND sg13g2_decap_8
XFILLER_6_669 VPWR VGND sg13g2_decap_8
XFILLER_5_168 VPWR VGND sg13g2_decap_8
XFILLER_2_831 VPWR VGND sg13g2_decap_8
XFILLER_1_341 VPWR VGND sg13g2_decap_8
XFILLER_49_345 VPWR VGND sg13g2_decap_8
XFILLER_18_732 VPWR VGND sg13g2_decap_8
XFILLER_45_562 VPWR VGND sg13g2_decap_8
XFILLER_17_242 VPWR VGND sg13g2_decap_8
XFILLER_17_253 VPWR VGND sg13g2_fill_2
XFILLER_27_90 VPWR VGND sg13g2_decap_8
XFILLER_33_713 VPWR VGND sg13g2_decap_8
XFILLER_17_286 VPWR VGND sg13g2_decap_8
X_538_ net75 VGND VPWR _078_ DP_1.matrix\[36\] clknet_5_21__leaf_clk sg13g2_dfrbpq_1
X_469_ net74 VGND VPWR net184 mac1.sum_lvl1_ff\[9\] clknet_5_25__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_267 VPWR VGND sg13g2_decap_8
XFILLER_9_430 VPWR VGND sg13g2_decap_8
XFILLER_13_492 VPWR VGND sg13g2_decap_8
XFILLER_24_713 VPWR VGND sg13g2_decap_8
XFILLER_36_562 VPWR VGND sg13g2_decap_8
XFILLER_23_201 VPWR VGND sg13g2_decap_8
XFILLER_23_289 VPWR VGND sg13g2_decap_8
XFILLER_20_941 VPWR VGND sg13g2_decap_8
XFILLER_23_59 VPWR VGND sg13g2_fill_2
XFILLER_2_105 VPWR VGND sg13g2_decap_8
XFILLER_47_805 VPWR VGND sg13g2_decap_8
XFILLER_48_56 VPWR VGND sg13g2_decap_8
XFILLER_24_1014 VPWR VGND sg13g2_decap_8
XFILLER_27_540 VPWR VGND sg13g2_decap_8
XFILLER_42_554 VPWR VGND sg13g2_decap_8
XFILLER_14_223 VPWR VGND sg13g2_decap_8
XFILLER_15_757 VPWR VGND sg13g2_decap_8
X_323_ _188_ net118 net91 VPWR VGND sg13g2_nand2_1
XFILLER_30_738 VPWR VGND sg13g2_decap_8
Xfanout60 net61 net60 VPWR VGND sg13g2_buf_8
X_254_ _150_ net163 net199 VPWR VGND sg13g2_nand2_1
Xfanout71 net72 net71 VPWR VGND sg13g2_buf_8
Xfanout82 net83 net82 VPWR VGND sg13g2_buf_8
XFILLER_11_963 VPWR VGND sg13g2_decap_8
XFILLER_31_1007 VPWR VGND sg13g2_decap_8
XFILLER_7_967 VPWR VGND sg13g2_decap_8
XFILLER_13_81 VPWR VGND sg13g2_decap_8
XFILLER_6_455 VPWR VGND sg13g2_decap_8
XFILLER_36_7 VPWR VGND sg13g2_decap_8
XFILLER_49_142 VPWR VGND sg13g2_decap_8
XFILLER_38_838 VPWR VGND sg13g2_decap_8
XFILLER_37_326 VPWR VGND sg13g2_fill_2
XFILLER_18_540 VPWR VGND sg13g2_fill_1
XFILLER_46_893 VPWR VGND sg13g2_decap_8
XFILLER_18_584 VPWR VGND sg13g2_fill_1
XFILLER_33_510 VPWR VGND sg13g2_decap_8
XFILLER_33_587 VPWR VGND sg13g2_decap_8
XFILLER_0_609 VPWR VGND sg13g2_decap_8
XFILLER_29_827 VPWR VGND sg13g2_decap_8
XFILLER_44_808 VPWR VGND sg13g2_decap_8
XFILLER_24_510 VPWR VGND sg13g2_decap_4
XFILLER_34_14 VPWR VGND sg13g2_decap_8
XFILLER_24_587 VPWR VGND sg13g2_decap_8
XFILLER_11_237 VPWR VGND sg13g2_decap_8
Xclkload2 clknet_5_12__leaf_clk clkload2/X VPWR VGND sg13g2_buf_1
XFILLER_4_948 VPWR VGND sg13g2_decap_8
XFILLER_3_436 VPWR VGND sg13g2_decap_8
XFILLER_47_602 VPWR VGND sg13g2_decap_8
XFILLER_46_101 VPWR VGND sg13g2_fill_1
XFILLER_47_679 VPWR VGND sg13g2_decap_8
XFILLER_28_882 VPWR VGND sg13g2_decap_8
XFILLER_15_543 VPWR VGND sg13g2_decap_8
XFILLER_43_874 VPWR VGND sg13g2_decap_8
XFILLER_42_351 VPWR VGND sg13g2_decap_8
XFILLER_15_587 VPWR VGND sg13g2_decap_8
XFILLER_30_535 VPWR VGND sg13g2_decap_8
X_306_ net103 mac2.products_ff\[68\] _026_ VPWR VGND sg13g2_xor2_1
XFILLER_11_760 VPWR VGND sg13g2_decap_8
X_237_ net160 net117 _048_ VPWR VGND sg13g2_and2_1
XFILLER_10_281 VPWR VGND sg13g2_decap_8
XFILLER_7_764 VPWR VGND sg13g2_decap_8
XFILLER_6_241 VPWR VGND sg13g2_decap_8
XFILLER_37_112 VPWR VGND sg13g2_decap_8
XFILLER_38_635 VPWR VGND sg13g2_decap_8
XFILLER_19_860 VPWR VGND sg13g2_decap_8
XFILLER_37_156 VPWR VGND sg13g2_decap_8
XFILLER_1_95 VPWR VGND sg13g2_decap_8
XFILLER_46_690 VPWR VGND sg13g2_decap_8
XFILLER_34_874 VPWR VGND sg13g2_decap_8
XFILLER_21_535 VPWR VGND sg13g2_decap_8
XFILLER_33_395 VPWR VGND sg13g2_decap_8
XFILLER_0_406 VPWR VGND sg13g2_decap_8
XFILLER_1_929 VPWR VGND sg13g2_decap_8
XFILLER_29_14 VPWR VGND sg13g2_decap_8
Xhold14 DP_2.matrix\[1\] VPWR VGND net38 sg13g2_dlygate4sd3_1
Xhold36 DP_3.matrix\[64\] VPWR VGND net86 sg13g2_dlygate4sd3_1
Xhold47 DP_1.matrix\[10\] VPWR VGND net97 sg13g2_dlygate4sd3_1
Xhold25 DP_4.matrix\[28\] VPWR VGND net49 sg13g2_dlygate4sd3_1
Xhold58 _030_ VPWR VGND net108 sg13g2_dlygate4sd3_1
XFILLER_29_624 VPWR VGND sg13g2_decap_8
Xhold69 DP_4.matrix\[0\] VPWR VGND net119 sg13g2_dlygate4sd3_1
XFILLER_44_605 VPWR VGND sg13g2_decap_8
XFILLER_45_35 VPWR VGND sg13g2_decap_8
XFILLER_43_159 VPWR VGND sg13g2_decap_4
XFILLER_43_148 VPWR VGND sg13g2_decap_8
XFILLER_25_830 VPWR VGND sg13g2_decap_8
XFILLER_40_855 VPWR VGND sg13g2_decap_8
XFILLER_6_18 VPWR VGND sg13g2_decap_8
XFILLER_3_211 VPWR VGND sg13g2_fill_2
XFILLER_4_745 VPWR VGND sg13g2_decap_8
XFILLER_3_222 VPWR VGND sg13g2_fill_2
XFILLER_3_299 VPWR VGND sg13g2_decap_8
XFILLER_0_973 VPWR VGND sg13g2_decap_8
XFILLER_48_944 VPWR VGND sg13g2_decap_8
XFILLER_19_123 VPWR VGND sg13g2_decap_8
XFILLER_47_476 VPWR VGND sg13g2_decap_8
XFILLER_35_627 VPWR VGND sg13g2_decap_8
XFILLER_16_830 VPWR VGND sg13g2_decap_8
XFILLER_43_671 VPWR VGND sg13g2_decap_8
XFILLER_31_811 VPWR VGND sg13g2_decap_8
XFILLER_37_1024 VPWR VGND sg13g2_decap_4
XFILLER_42_192 VPWR VGND sg13g2_decap_8
XFILLER_31_888 VPWR VGND sg13g2_decap_8
XFILLER_30_365 VPWR VGND sg13g2_decap_8
XFILLER_30_376 VPWR VGND sg13g2_fill_1
Xheichips25_template_16 VPWR VGND uo_out[7] sg13g2_tielo
XFILLER_38_465 VPWR VGND sg13g2_decap_4
XFILLER_39_966 VPWR VGND sg13g2_decap_8
XFILLER_26_627 VPWR VGND sg13g2_decap_8
XFILLER_34_671 VPWR VGND sg13g2_decap_8
XFILLER_22_844 VPWR VGND sg13g2_decap_8
XFILLER_21_365 VPWR VGND sg13g2_decap_8
XFILLER_0_203 VPWR VGND sg13g2_decap_8
XFILLER_1_726 VPWR VGND sg13g2_decap_8
XFILLER_5_1011 VPWR VGND sg13g2_decap_8
X_571_ net70 VGND VPWR _111_ DP_3.matrix\[19\] clknet_5_11__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_947 VPWR VGND sg13g2_decap_8
XFILLER_44_402 VPWR VGND sg13g2_decap_8
XFILLER_16_148 VPWR VGND sg13g2_decap_8
XFILLER_17_649 VPWR VGND sg13g2_decap_8
XFILLER_44_479 VPWR VGND sg13g2_decap_8
XFILLER_13_844 VPWR VGND sg13g2_decap_8
XFILLER_9_815 VPWR VGND sg13g2_decap_8
XFILLER_40_652 VPWR VGND sg13g2_decap_8
XFILLER_12_365 VPWR VGND sg13g2_decap_8
XFILLER_8_369 VPWR VGND sg13g2_decap_8
XFILLER_4_520 VPWR VGND sg13g2_decap_8
XFILLER_0_770 VPWR VGND sg13g2_decap_8
XFILLER_48_741 VPWR VGND sg13g2_decap_8
XFILLER_36_947 VPWR VGND sg13g2_decap_8
XFILLER_35_424 VPWR VGND sg13g2_decap_8
XFILLER_35_435 VPWR VGND sg13g2_fill_1
XFILLER_31_685 VPWR VGND sg13g2_decap_8
XFILLER_11_1005 VPWR VGND sg13g2_decap_8
XFILLER_30_184 VPWR VGND sg13g2_decap_4
XFILLER_8_881 VPWR VGND sg13g2_decap_8
XFILLER_39_763 VPWR VGND sg13g2_decap_8
XFILLER_27_925 VPWR VGND sg13g2_decap_8
XFILLER_38_251 VPWR VGND sg13g2_decap_8
XFILLER_26_424 VPWR VGND sg13g2_decap_8
XFILLER_42_939 VPWR VGND sg13g2_decap_8
XFILLER_41_405 VPWR VGND sg13g2_decap_8
XFILLER_35_991 VPWR VGND sg13g2_decap_8
XFILLER_22_641 VPWR VGND sg13g2_decap_8
XFILLER_42_14 VPWR VGND sg13g2_decap_8
XFILLER_10_858 VPWR VGND sg13g2_decap_8
XFILLER_5_317 VPWR VGND sg13g2_decap_8
XFILLER_1_523 VPWR VGND sg13g2_decap_8
XFILLER_27_1023 VPWR VGND sg13g2_decap_4
XFILLER_49_527 VPWR VGND sg13g2_decap_8
XFILLER_18_914 VPWR VGND sg13g2_decap_8
XFILLER_29_251 VPWR VGND sg13g2_fill_1
XFILLER_45_744 VPWR VGND sg13g2_decap_8
XFILLER_17_424 VPWR VGND sg13g2_fill_1
X_554_ net66 VGND VPWR _094_ DP_2.matrix\[27\] clknet_5_7__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_276 VPWR VGND sg13g2_decap_8
X_485_ net64 VGND VPWR net30 mac1.sum_lvl3_ff\[3\] clknet_5_16__leaf_clk sg13g2_dfrbpq_1
XFILLER_26_991 VPWR VGND sg13g2_decap_8
XFILLER_32_438 VPWR VGND sg13g2_decap_8
XFILLER_13_641 VPWR VGND sg13g2_decap_8
XFILLER_9_612 VPWR VGND sg13g2_decap_8
XFILLER_12_151 VPWR VGND sg13g2_decap_8
XFILLER_9_689 VPWR VGND sg13g2_decap_8
XFILLER_8_155 VPWR VGND sg13g2_decap_8
XFILLER_32_80 VPWR VGND sg13g2_decap_8
XFILLER_4_361 VPWR VGND sg13g2_decap_8
XFILLER_41_1009 VPWR VGND sg13g2_decap_8
XFILLER_35_210 VPWR VGND sg13g2_fill_1
XFILLER_36_744 VPWR VGND sg13g2_decap_8
XFILLER_35_287 VPWR VGND sg13g2_decap_8
XFILLER_31_482 VPWR VGND sg13g2_decap_8
Xhold100 DP_2.matrix\[45\] VPWR VGND net150 sg13g2_dlygate4sd3_1
Xhold144 _009_ VPWR VGND net194 sg13g2_dlygate4sd3_1
Xhold111 mac1.sum_lvl1_ff\[16\] VPWR VGND net161 sg13g2_dlygate4sd3_1
Xhold122 _019_ VPWR VGND net172 sg13g2_dlygate4sd3_1
Xhold133 mac1.products_ff\[34\] VPWR VGND net183 sg13g2_dlygate4sd3_1
XFILLER_37_14 VPWR VGND sg13g2_decap_8
XFILLER_46_508 VPWR VGND sg13g2_decap_8
XFILLER_39_560 VPWR VGND sg13g2_decap_8
XFILLER_27_722 VPWR VGND sg13g2_decap_8
XFILLER_14_405 VPWR VGND sg13g2_decap_8
XFILLER_26_254 VPWR VGND sg13g2_decap_8
XFILLER_42_736 VPWR VGND sg13g2_decap_8
XFILLER_14_416 VPWR VGND sg13g2_fill_1
XFILLER_15_939 VPWR VGND sg13g2_decap_8
XFILLER_27_799 VPWR VGND sg13g2_decap_8
XFILLER_41_202 VPWR VGND sg13g2_decap_8
XFILLER_23_961 VPWR VGND sg13g2_decap_8
X_270_ mac1.products_ff\[1\] mac1.products_ff\[18\] _161_ VPWR VGND sg13g2_xor2_1
XFILLER_41_279 VPWR VGND sg13g2_decap_8
XFILLER_22_482 VPWR VGND sg13g2_fill_2
XFILLER_22_493 VPWR VGND sg13g2_fill_1
XFILLER_10_655 VPWR VGND sg13g2_decap_8
XFILLER_6_648 VPWR VGND sg13g2_decap_8
XFILLER_5_147 VPWR VGND sg13g2_decap_8
XFILLER_2_810 VPWR VGND sg13g2_decap_8
XFILLER_1_320 VPWR VGND sg13g2_decap_8
XFILLER_49_324 VPWR VGND sg13g2_decap_8
XFILLER_2_887 VPWR VGND sg13g2_decap_8
XFILLER_1_397 VPWR VGND sg13g2_decap_8
XFILLER_18_711 VPWR VGND sg13g2_decap_8
XFILLER_17_221 VPWR VGND sg13g2_decap_8
XFILLER_45_541 VPWR VGND sg13g2_decap_8
XFILLER_18_788 VPWR VGND sg13g2_decap_8
X_537_ net65 VGND VPWR _077_ DP_1.matrix\[28\] clknet_5_24__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_769 VPWR VGND sg13g2_decap_8
XFILLER_14_994 VPWR VGND sg13g2_decap_8
X_468_ net74 VGND VPWR net112 mac1.sum_lvl1_ff\[8\] clknet_5_19__leaf_clk sg13g2_dfrbpq_1
XFILLER_13_471 VPWR VGND sg13g2_decap_8
X_399_ net98 _093_ VPWR VGND sg13g2_buf_1
XFILLER_4_95 VPWR VGND sg13g2_decap_8
XFILLER_49_891 VPWR VGND sg13g2_decap_8
XFILLER_36_541 VPWR VGND sg13g2_decap_8
XFILLER_24_769 VPWR VGND sg13g2_decap_8
Xclkbuf_5_18__f_clk clknet_4_9_0_clk clknet_5_18__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_20_920 VPWR VGND sg13g2_decap_8
XFILLER_23_38 VPWR VGND sg13g2_decap_8
XFILLER_20_997 VPWR VGND sg13g2_decap_8
XFILLER_3_629 VPWR VGND sg13g2_decap_8
XFILLER_2_139 VPWR VGND sg13g2_fill_1
XFILLER_48_35 VPWR VGND sg13g2_decap_8
XFILLER_46_338 VPWR VGND sg13g2_fill_1
XFILLER_14_202 VPWR VGND sg13g2_decap_8
XFILLER_15_736 VPWR VGND sg13g2_decap_8
XFILLER_27_596 VPWR VGND sg13g2_decap_8
XFILLER_42_533 VPWR VGND sg13g2_decap_8
X_322_ _187_ _186_ _067_ VPWR VGND sg13g2_xor2_1
XFILLER_14_279 VPWR VGND sg13g2_decap_8
XFILLER_30_717 VPWR VGND sg13g2_decap_8
Xfanout61 net63 net61 VPWR VGND sg13g2_buf_8
XFILLER_11_942 VPWR VGND sg13g2_decap_8
X_253_ net107 mac2.sum_lvl1_ff\[0\] _030_ VPWR VGND sg13g2_xor2_1
Xfanout72 rst_n net72 VPWR VGND sg13g2_buf_8
Xfanout83 net84 net83 VPWR VGND sg13g2_buf_8
XFILLER_10_452 VPWR VGND sg13g2_decap_8
XFILLER_13_60 VPWR VGND sg13g2_decap_8
XFILLER_7_946 VPWR VGND sg13g2_decap_8
XFILLER_6_434 VPWR VGND sg13g2_decap_8
XFILLER_2_684 VPWR VGND sg13g2_decap_8
XFILLER_1_194 VPWR VGND sg13g2_decap_8
XFILLER_29_7 VPWR VGND sg13g2_decap_8
XFILLER_38_817 VPWR VGND sg13g2_decap_8
XFILLER_49_198 VPWR VGND sg13g2_decap_8
XFILLER_38_90 VPWR VGND sg13g2_decap_8
XFILLER_46_872 VPWR VGND sg13g2_decap_8
XFILLER_18_563 VPWR VGND sg13g2_decap_8
XFILLER_18_596 VPWR VGND sg13g2_fill_1
XFILLER_33_566 VPWR VGND sg13g2_decap_8
XFILLER_14_791 VPWR VGND sg13g2_decap_8
XFILLER_20_249 VPWR VGND sg13g2_decap_8
XFILLER_9_294 VPWR VGND sg13g2_decap_8
XFILLER_47_1015 VPWR VGND sg13g2_decap_8
XFILLER_29_806 VPWR VGND sg13g2_decap_8
XFILLER_36_382 VPWR VGND sg13g2_decap_8
XFILLER_24_566 VPWR VGND sg13g2_decap_8
XFILLER_11_216 VPWR VGND sg13g2_decap_8
XFILLER_12_739 VPWR VGND sg13g2_decap_8
Xclkload3 VPWR clkload3/Y clknet_5_15__leaf_clk VGND sg13g2_inv_1
XFILLER_20_794 VPWR VGND sg13g2_decap_8
XFILLER_4_927 VPWR VGND sg13g2_decap_8
XFILLER_19_305 VPWR VGND sg13g2_decap_8
XFILLER_47_658 VPWR VGND sg13g2_decap_8
XFILLER_28_861 VPWR VGND sg13g2_decap_8
XFILLER_35_809 VPWR VGND sg13g2_decap_8
XFILLER_27_371 VPWR VGND sg13g2_decap_8
XFILLER_43_853 VPWR VGND sg13g2_decap_8
XFILLER_42_330 VPWR VGND sg13g2_decap_8
XFILLER_15_522 VPWR VGND sg13g2_decap_8
XFILLER_27_382 VPWR VGND sg13g2_fill_1
XFILLER_15_577 VPWR VGND sg13g2_fill_2
XFILLER_30_514 VPWR VGND sg13g2_decap_8
X_305_ _027_ _178_ _179_ VPWR VGND sg13g2_xnor2_1
XFILLER_7_743 VPWR VGND sg13g2_decap_8
X_236_ net129 net134 _046_ VPWR VGND sg13g2_and2_1
XFILLER_6_220 VPWR VGND sg13g2_decap_8
XFILLER_6_297 VPWR VGND sg13g2_decap_8
XFILLER_3_993 VPWR VGND sg13g2_decap_8
XFILLER_38_614 VPWR VGND sg13g2_decap_8
XFILLER_1_74 VPWR VGND sg13g2_fill_1
XFILLER_1_63 VPWR VGND sg13g2_decap_8
XFILLER_26_809 VPWR VGND sg13g2_decap_8
XFILLER_37_135 VPWR VGND sg13g2_decap_8
XFILLER_1_85 VPWR VGND sg13g2_fill_1
XFILLER_34_853 VPWR VGND sg13g2_decap_8
XFILLER_21_514 VPWR VGND sg13g2_decap_8
XFILLER_20_39 VPWR VGND sg13g2_decap_8
XFILLER_1_908 VPWR VGND sg13g2_decap_8
Xhold15 DP_4.matrix\[46\] VPWR VGND net39 sg13g2_dlygate4sd3_1
Xhold26 DP_3.matrix\[28\] VPWR VGND net50 sg13g2_dlygate4sd3_1
Xhold37 DP_1.matrix\[37\] VPWR VGND net87 sg13g2_dlygate4sd3_1
XFILLER_29_603 VPWR VGND sg13g2_decap_8
Xhold48 DP_2.matrix\[19\] VPWR VGND net98 sg13g2_dlygate4sd3_1
Xhold59 mac2.products_ff\[34\] VPWR VGND net109 sg13g2_dlygate4sd3_1
XFILLER_28_124 VPWR VGND sg13g2_decap_8
XFILLER_45_14 VPWR VGND sg13g2_decap_8
XFILLER_43_127 VPWR VGND sg13g2_decap_8
XFILLER_12_503 VPWR VGND sg13g2_decap_8
XFILLER_25_886 VPWR VGND sg13g2_decap_8
XFILLER_40_834 VPWR VGND sg13g2_decap_8
XFILLER_20_591 VPWR VGND sg13g2_decap_8
XFILLER_4_724 VPWR VGND sg13g2_decap_8
XFILLER_3_278 VPWR VGND sg13g2_decap_8
XFILLER_0_952 VPWR VGND sg13g2_decap_8
XFILLER_48_923 VPWR VGND sg13g2_decap_8
XFILLER_19_102 VPWR VGND sg13g2_decap_8
XFILLER_47_455 VPWR VGND sg13g2_decap_8
XFILLER_19_81 VPWR VGND sg13g2_decap_8
XFILLER_19_179 VPWR VGND sg13g2_decap_8
XFILLER_35_606 VPWR VGND sg13g2_decap_8
XFILLER_34_116 VPWR VGND sg13g2_decap_8
XFILLER_43_650 VPWR VGND sg13g2_decap_8
XFILLER_16_886 VPWR VGND sg13g2_decap_8
XFILLER_37_1003 VPWR VGND sg13g2_decap_8
XFILLER_42_171 VPWR VGND sg13g2_decap_8
XFILLER_15_396 VPWR VGND sg13g2_decap_8
XFILLER_30_344 VPWR VGND sg13g2_decap_8
XFILLER_31_867 VPWR VGND sg13g2_decap_8
XFILLER_44_1018 VPWR VGND sg13g2_decap_8
XFILLER_3_790 VPWR VGND sg13g2_decap_8
Xheichips25_template_17 VPWR VGND uio_oe[0] sg13g2_tiehi
XFILLER_39_945 VPWR VGND sg13g2_decap_8
XFILLER_26_606 VPWR VGND sg13g2_decap_8
XFILLER_34_650 VPWR VGND sg13g2_decap_8
XFILLER_22_823 VPWR VGND sg13g2_decap_8
XFILLER_31_49 VPWR VGND sg13g2_decap_8
XFILLER_1_705 VPWR VGND sg13g2_decap_8
XFILLER_49_709 VPWR VGND sg13g2_decap_8
XFILLER_0_259 VPWR VGND sg13g2_decap_8
XFILLER_48_219 VPWR VGND sg13g2_decap_4
XFILLER_45_926 VPWR VGND sg13g2_decap_8
X_570_ net69 VGND VPWR _110_ DP_3.matrix\[18\] clknet_5_10__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_628 VPWR VGND sg13g2_decap_8
XFILLER_29_488 VPWR VGND sg13g2_decap_4
XFILLER_44_458 VPWR VGND sg13g2_decap_8
XFILLER_13_823 VPWR VGND sg13g2_decap_8
XFILLER_25_683 VPWR VGND sg13g2_decap_8
XFILLER_31_119 VPWR VGND sg13g2_decap_8
XFILLER_12_344 VPWR VGND sg13g2_decap_8
XFILLER_40_631 VPWR VGND sg13g2_decap_8
XFILLER_4_598 VPWR VGND sg13g2_decap_8
XFILLER_48_720 VPWR VGND sg13g2_decap_8
XFILLER_48_797 VPWR VGND sg13g2_decap_8
XFILLER_35_403 VPWR VGND sg13g2_decap_8
XFILLER_36_926 VPWR VGND sg13g2_decap_8
XFILLER_16_683 VPWR VGND sg13g2_decap_8
XFILLER_15_182 VPWR VGND sg13g2_fill_1
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
XFILLER_31_664 VPWR VGND sg13g2_decap_8
XFILLER_8_860 VPWR VGND sg13g2_decap_8
XFILLER_11_1028 VPWR VGND sg13g2_fill_1
XFILLER_7_84 VPWR VGND sg13g2_decap_8
XFILLER_38_230 VPWR VGND sg13g2_decap_8
XFILLER_39_742 VPWR VGND sg13g2_decap_8
XFILLER_27_904 VPWR VGND sg13g2_decap_8
XFILLER_42_918 VPWR VGND sg13g2_decap_8
XFILLER_14_609 VPWR VGND sg13g2_decap_8
XFILLER_35_970 VPWR VGND sg13g2_decap_8
XFILLER_22_620 VPWR VGND sg13g2_decap_8
XFILLER_42_59 VPWR VGND sg13g2_decap_8
XFILLER_10_837 VPWR VGND sg13g2_decap_8
XFILLER_22_697 VPWR VGND sg13g2_decap_8
XFILLER_1_502 VPWR VGND sg13g2_decap_8
XFILLER_27_1002 VPWR VGND sg13g2_decap_8
XFILLER_49_506 VPWR VGND sg13g2_decap_8
XFILLER_1_579 VPWR VGND sg13g2_decap_8
XFILLER_45_723 VPWR VGND sg13g2_decap_8
XFILLER_29_285 VPWR VGND sg13g2_decap_8
XFILLER_44_255 VPWR VGND sg13g2_fill_1
X_553_ net66 VGND VPWR _093_ DP_2.matrix\[19\] clknet_5_18__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_469 VPWR VGND sg13g2_decap_8
X_484_ net64 VGND VPWR net36 mac1.sum_lvl3_ff\[2\] clknet_5_16__leaf_clk sg13g2_dfrbpq_1
XFILLER_26_970 VPWR VGND sg13g2_decap_8
XFILLER_13_620 VPWR VGND sg13g2_decap_8
XFILLER_12_130 VPWR VGND sg13g2_decap_8
XFILLER_34_1028 VPWR VGND sg13g2_fill_1
XFILLER_41_995 VPWR VGND sg13g2_decap_8
XFILLER_9_668 VPWR VGND sg13g2_decap_8
XFILLER_8_134 VPWR VGND sg13g2_decap_8
XFILLER_13_697 VPWR VGND sg13g2_decap_8
XFILLER_8_189 VPWR VGND sg13g2_decap_8
XFILLER_5_885 VPWR VGND sg13g2_decap_8
XFILLER_48_594 VPWR VGND sg13g2_decap_8
XFILLER_36_723 VPWR VGND sg13g2_decap_8
XFILLER_17_992 VPWR VGND sg13g2_decap_8
XFILLER_35_266 VPWR VGND sg13g2_decap_8
XFILLER_31_461 VPWR VGND sg13g2_decap_8
XFILLER_32_984 VPWR VGND sg13g2_decap_8
XFILLER_12_18 VPWR VGND sg13g2_decap_8
Xhold101 DP_1.matrix\[54\] VPWR VGND net151 sg13g2_dlygate4sd3_1
Xhold123 mac1.sum_lvl1_ff\[24\] VPWR VGND net173 sg13g2_dlygate4sd3_1
Xhold112 _012_ VPWR VGND net162 sg13g2_dlygate4sd3_1
Xhold134 _005_ VPWR VGND net184 sg13g2_dlygate4sd3_1
Xhold145 mac2.products_ff\[119\] VPWR VGND net195 sg13g2_dlygate4sd3_1
XFILLER_27_701 VPWR VGND sg13g2_decap_8
XFILLER_15_918 VPWR VGND sg13g2_decap_8
XFILLER_26_233 VPWR VGND sg13g2_decap_8
XFILLER_27_778 VPWR VGND sg13g2_decap_8
XFILLER_42_715 VPWR VGND sg13g2_decap_8
XFILLER_23_940 VPWR VGND sg13g2_decap_8
XFILLER_22_461 VPWR VGND sg13g2_decap_8
XFILLER_41_258 VPWR VGND sg13g2_decap_4
XFILLER_10_634 VPWR VGND sg13g2_decap_8
XFILLER_6_627 VPWR VGND sg13g2_decap_8
XFILLER_2_866 VPWR VGND sg13g2_decap_8
XFILLER_49_303 VPWR VGND sg13g2_decap_8
XFILLER_1_376 VPWR VGND sg13g2_decap_8
XFILLER_45_520 VPWR VGND sg13g2_decap_8
XFILLER_17_200 VPWR VGND sg13g2_decap_8
XFILLER_18_767 VPWR VGND sg13g2_decap_8
XFILLER_45_597 VPWR VGND sg13g2_decap_8
X_536_ net65 VGND VPWR _076_ DP_1.matrix\[27\] clknet_5_24__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_214 VPWR VGND sg13g2_decap_8
XFILLER_33_748 VPWR VGND sg13g2_decap_8
XFILLER_14_973 VPWR VGND sg13g2_decap_8
XFILLER_20_409 VPWR VGND sg13g2_decap_8
X_467_ net74 VGND VPWR net178 mac1.sum_lvl1_ff\[1\] clknet_5_19__leaf_clk sg13g2_dfrbpq_1
X_398_ net129 _092_ VPWR VGND sg13g2_buf_1
XFILLER_41_792 VPWR VGND sg13g2_decap_8
XFILLER_9_465 VPWR VGND sg13g2_fill_2
XFILLER_40_291 VPWR VGND sg13g2_decap_8
XFILLER_9_498 VPWR VGND sg13g2_decap_8
XFILLER_5_682 VPWR VGND sg13g2_decap_8
XFILLER_4_74 VPWR VGND sg13g2_decap_8
XFILLER_49_870 VPWR VGND sg13g2_decap_8
XFILLER_36_520 VPWR VGND sg13g2_decap_8
XFILLER_36_597 VPWR VGND sg13g2_decap_8
XFILLER_23_247 VPWR VGND sg13g2_decap_8
XFILLER_24_748 VPWR VGND sg13g2_decap_8
XFILLER_31_280 VPWR VGND sg13g2_decap_8
XFILLER_32_781 VPWR VGND sg13g2_decap_8
XFILLER_20_976 VPWR VGND sg13g2_decap_8
XFILLER_3_608 VPWR VGND sg13g2_decap_8
XFILLER_48_14 VPWR VGND sg13g2_decap_8
XFILLER_46_317 VPWR VGND sg13g2_decap_8
XFILLER_42_512 VPWR VGND sg13g2_decap_8
XFILLER_15_715 VPWR VGND sg13g2_decap_8
XFILLER_27_575 VPWR VGND sg13g2_decap_8
X_321_ _187_ net130 net56 VPWR VGND sg13g2_nand2_1
XFILLER_42_589 VPWR VGND sg13g2_decap_8
XFILLER_14_258 VPWR VGND sg13g2_decap_8
Xfanout73 net74 net73 VPWR VGND sg13g2_buf_8
XFILLER_11_921 VPWR VGND sg13g2_decap_8
Xfanout62 net63 net62 VPWR VGND sg13g2_buf_8
X_252_ _031_ _148_ _149_ VPWR VGND sg13g2_xnor2_1
XFILLER_10_431 VPWR VGND sg13g2_decap_8
XFILLER_7_925 VPWR VGND sg13g2_decap_8
Xfanout84 net85 net84 VPWR VGND sg13g2_buf_8
XFILLER_6_413 VPWR VGND sg13g2_decap_8
XFILLER_11_998 VPWR VGND sg13g2_decap_8
XFILLER_1_151 VPWR VGND sg13g2_decap_8
XFILLER_2_663 VPWR VGND sg13g2_decap_8
XFILLER_49_177 VPWR VGND sg13g2_decap_8
XFILLER_46_851 VPWR VGND sg13g2_decap_8
Xclkbuf_5_24__f_clk clknet_4_12_0_clk clknet_5_24__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_33_545 VPWR VGND sg13g2_decap_8
XFILLER_21_729 VPWR VGND sg13g2_decap_8
X_519_ net71 VGND VPWR net137 mac2.sum_lvl2_ff\[4\] clknet_5_13__leaf_clk sg13g2_dfrbpq_1
XFILLER_14_770 VPWR VGND sg13g2_decap_8
XFILLER_20_228 VPWR VGND sg13g2_decap_8
XFILLER_9_251 VPWR VGND sg13g2_fill_2
XFILLER_6_991 VPWR VGND sg13g2_decap_8
XFILLER_48_0 VPWR VGND sg13g2_decap_8
XFILLER_18_39 VPWR VGND sg13g2_decap_8
XFILLER_43_309 VPWR VGND sg13g2_decap_8
XFILLER_36_361 VPWR VGND sg13g2_decap_8
XFILLER_37_884 VPWR VGND sg13g2_decap_8
XFILLER_24_545 VPWR VGND sg13g2_decap_8
XFILLER_12_718 VPWR VGND sg13g2_decap_8
Xclkload4 clknet_5_17__leaf_clk clkload4/X VPWR VGND sg13g2_buf_1
XFILLER_20_773 VPWR VGND sg13g2_decap_8
XFILLER_4_906 VPWR VGND sg13g2_decap_8
XFILLER_3_416 VPWR VGND sg13g2_decap_4
XFILLER_8_1021 VPWR VGND sg13g2_decap_8
XFILLER_47_637 VPWR VGND sg13g2_decap_8
XFILLER_19_339 VPWR VGND sg13g2_decap_8
XFILLER_46_147 VPWR VGND sg13g2_decap_8
XFILLER_28_840 VPWR VGND sg13g2_decap_8
XFILLER_15_501 VPWR VGND sg13g2_decap_8
XFILLER_27_350 VPWR VGND sg13g2_decap_8
XFILLER_43_832 VPWR VGND sg13g2_decap_8
X_304_ mac2.products_ff\[86\] mac2.products_ff\[69\] _179_ VPWR VGND sg13g2_xor2_1
XFILLER_42_386 VPWR VGND sg13g2_decap_8
XFILLER_24_82 VPWR VGND sg13g2_decap_8
X_235_ net128 net147 _044_ VPWR VGND sg13g2_and2_1
XFILLER_7_722 VPWR VGND sg13g2_decap_8
XFILLER_11_795 VPWR VGND sg13g2_decap_8
XFILLER_7_799 VPWR VGND sg13g2_decap_8
XFILLER_6_276 VPWR VGND sg13g2_decap_8
XFILLER_3_972 VPWR VGND sg13g2_decap_8
XFILLER_41_7 VPWR VGND sg13g2_decap_4
XFILLER_1_42 VPWR VGND sg13g2_decap_8
XFILLER_45_180 VPWR VGND sg13g2_decap_8
XFILLER_18_383 VPWR VGND sg13g2_decap_8
XFILLER_19_895 VPWR VGND sg13g2_decap_8
XFILLER_34_832 VPWR VGND sg13g2_decap_8
XFILLER_33_342 VPWR VGND sg13g2_decap_8
XFILLER_14_1015 VPWR VGND sg13g2_decap_8
XFILLER_20_18 VPWR VGND sg13g2_decap_8
Xhold27 DP_4.matrix\[64\] VPWR VGND net51 sg13g2_dlygate4sd3_1
Xhold16 DP_2.matrix\[64\] VPWR VGND net40 sg13g2_dlygate4sd3_1
Xhold38 DP_3.matrix\[1\] VPWR VGND net88 sg13g2_dlygate4sd3_1
Xhold49 mac1.products_ff\[119\] VPWR VGND net99 sg13g2_dlygate4sd3_1
XFILLER_29_659 VPWR VGND sg13g2_decap_8
XFILLER_43_106 VPWR VGND sg13g2_decap_8
XFILLER_37_681 VPWR VGND sg13g2_decap_8
XFILLER_24_353 VPWR VGND sg13g2_fill_2
XFILLER_25_865 VPWR VGND sg13g2_decap_8
XFILLER_12_526 VPWR VGND sg13g2_decap_4
XFILLER_24_397 VPWR VGND sg13g2_decap_4
XFILLER_40_813 VPWR VGND sg13g2_decap_8
XFILLER_20_570 VPWR VGND sg13g2_decap_8
XFILLER_4_703 VPWR VGND sg13g2_decap_8
XFILLER_0_931 VPWR VGND sg13g2_decap_8
XFILLER_48_902 VPWR VGND sg13g2_decap_8
XFILLER_48_979 VPWR VGND sg13g2_decap_8
XFILLER_47_434 VPWR VGND sg13g2_decap_8
XFILLER_19_60 VPWR VGND sg13g2_decap_8
XFILLER_19_158 VPWR VGND sg13g2_decap_8
XFILLER_15_331 VPWR VGND sg13g2_fill_1
XFILLER_16_865 VPWR VGND sg13g2_decap_8
XFILLER_15_375 VPWR VGND sg13g2_decap_8
XFILLER_30_323 VPWR VGND sg13g2_decap_8
XFILLER_31_846 VPWR VGND sg13g2_decap_8
XFILLER_7_530 VPWR VGND sg13g2_decap_8
XFILLER_11_592 VPWR VGND sg13g2_decap_8
XFILLER_7_596 VPWR VGND sg13g2_decap_8
Xheichips25_template_18 VPWR VGND uio_oe[1] sg13g2_tiehi
XFILLER_39_924 VPWR VGND sg13g2_decap_8
XFILLER_38_434 VPWR VGND sg13g2_decap_4
XFILLER_19_692 VPWR VGND sg13g2_decap_8
XFILLER_22_802 VPWR VGND sg13g2_decap_8
XFILLER_33_172 VPWR VGND sg13g2_decap_8
XFILLER_22_879 VPWR VGND sg13g2_decap_8
XFILLER_31_28 VPWR VGND sg13g2_decap_8
XFILLER_0_238 VPWR VGND sg13g2_decap_8
XFILLER_29_423 VPWR VGND sg13g2_decap_8
XFILLER_45_905 VPWR VGND sg13g2_decap_8
XFILLER_17_607 VPWR VGND sg13g2_decap_8
XFILLER_44_437 VPWR VGND sg13g2_decap_8
XFILLER_13_802 VPWR VGND sg13g2_decap_8
XFILLER_25_662 VPWR VGND sg13g2_decap_8
XFILLER_12_301 VPWR VGND sg13g2_decap_8
XFILLER_40_610 VPWR VGND sg13g2_decap_8
XFILLER_24_194 VPWR VGND sg13g2_decap_8
XFILLER_8_316 VPWR VGND sg13g2_decap_8
XFILLER_13_879 VPWR VGND sg13g2_decap_8
XFILLER_40_687 VPWR VGND sg13g2_decap_8
XFILLER_21_890 VPWR VGND sg13g2_decap_8
XFILLER_4_555 VPWR VGND sg13g2_fill_1
XFILLER_21_83 VPWR VGND sg13g2_decap_8
XFILLER_47_220 VPWR VGND sg13g2_fill_1
XFILLER_48_776 VPWR VGND sg13g2_decap_8
XFILLER_36_905 VPWR VGND sg13g2_decap_8
XFILLER_46_80 VPWR VGND sg13g2_decap_8
XFILLER_15_161 VPWR VGND sg13g2_decap_8
XFILLER_16_662 VPWR VGND sg13g2_decap_8
XFILLER_31_643 VPWR VGND sg13g2_decap_8
XFILLER_30_197 VPWR VGND sg13g2_decap_8
XFILLER_7_63 VPWR VGND sg13g2_decap_8
XFILLER_30_0 VPWR VGND sg13g2_decap_8
XFILLER_39_721 VPWR VGND sg13g2_decap_8
XFILLER_26_39 VPWR VGND sg13g2_decap_8
XFILLER_39_798 VPWR VGND sg13g2_decap_8
XFILLER_26_459 VPWR VGND sg13g2_decap_8
XFILLER_13_109 VPWR VGND sg13g2_decap_8
XFILLER_34_481 VPWR VGND sg13g2_fill_2
XFILLER_10_816 VPWR VGND sg13g2_decap_8
XFILLER_21_153 VPWR VGND sg13g2_decap_8
XFILLER_22_676 VPWR VGND sg13g2_decap_8
XFILLER_42_38 VPWR VGND sg13g2_decap_8
XFILLER_6_809 VPWR VGND sg13g2_decap_8
XFILLER_21_164 VPWR VGND sg13g2_fill_1
XFILLER_1_558 VPWR VGND sg13g2_decap_8
Xclkbuf_5_5__f_clk clknet_4_2_0_clk clknet_5_5__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_45_702 VPWR VGND sg13g2_decap_8
XFILLER_29_242 VPWR VGND sg13g2_decap_8
XFILLER_18_949 VPWR VGND sg13g2_decap_8
XFILLER_45_779 VPWR VGND sg13g2_decap_8
X_552_ net64 VGND VPWR _092_ DP_2.matrix\[18\] clknet_5_18__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_448 VPWR VGND sg13g2_decap_8
X_483_ net73 VGND VPWR net198 mac1.sum_lvl3_ff\[1\] clknet_5_16__leaf_clk sg13g2_dfrbpq_2
XFILLER_12_120 VPWR VGND sg13g2_fill_1
XFILLER_8_102 VPWR VGND sg13g2_decap_4
XFILLER_13_676 VPWR VGND sg13g2_decap_8
XFILLER_34_1007 VPWR VGND sg13g2_decap_8
XFILLER_41_974 VPWR VGND sg13g2_decap_8
XFILLER_9_647 VPWR VGND sg13g2_decap_8
XFILLER_12_175 VPWR VGND sg13g2_decap_8
XFILLER_40_473 VPWR VGND sg13g2_decap_8
XFILLER_5_864 VPWR VGND sg13g2_decap_8
XFILLER_36_702 VPWR VGND sg13g2_decap_8
XFILLER_48_573 VPWR VGND sg13g2_decap_8
XFILLER_35_245 VPWR VGND sg13g2_decap_8
XFILLER_36_779 VPWR VGND sg13g2_decap_8
XFILLER_17_971 VPWR VGND sg13g2_decap_8
XFILLER_16_470 VPWR VGND sg13g2_fill_2
XFILLER_32_963 VPWR VGND sg13g2_decap_8
Xhold124 _013_ VPWR VGND net174 sg13g2_dlygate4sd3_1
Xhold102 DP_4.matrix\[9\] VPWR VGND net152 sg13g2_dlygate4sd3_1
Xhold113 mac2.sum_lvl2_ff\[0\] VPWR VGND net163 sg13g2_dlygate4sd3_1
Xhold135 mac2.sum_lvl1_ff\[0\] VPWR VGND net185 sg13g2_dlygate4sd3_1
Xhold146 _029_ VPWR VGND net196 sg13g2_dlygate4sd3_1
XFILLER_2_1027 VPWR VGND sg13g2_fill_2
XFILLER_26_212 VPWR VGND sg13g2_decap_8
XFILLER_39_595 VPWR VGND sg13g2_decap_8
XFILLER_27_757 VPWR VGND sg13g2_decap_8
XFILLER_26_267 VPWR VGND sg13g2_decap_4
XFILLER_26_289 VPWR VGND sg13g2_decap_8
XFILLER_41_237 VPWR VGND sg13g2_decap_8
XFILLER_22_440 VPWR VGND sg13g2_decap_8
XFILLER_10_613 VPWR VGND sg13g2_decap_8
XFILLER_22_484 VPWR VGND sg13g2_fill_1
XFILLER_23_996 VPWR VGND sg13g2_decap_8
XFILLER_6_606 VPWR VGND sg13g2_decap_8
XFILLER_2_845 VPWR VGND sg13g2_decap_8
XFILLER_1_355 VPWR VGND sg13g2_decap_8
XFILLER_49_359 VPWR VGND sg13g2_decap_8
XFILLER_18_746 VPWR VGND sg13g2_decap_8
XFILLER_45_576 VPWR VGND sg13g2_decap_8
X_535_ net64 VGND VPWR _075_ DP_1.matrix\[19\] clknet_5_18__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_727 VPWR VGND sg13g2_decap_8
XFILLER_14_952 VPWR VGND sg13g2_decap_8
X_466_ net74 VGND VPWR net94 mac1.sum_lvl1_ff\[0\] clknet_5_19__leaf_clk sg13g2_dfrbpq_1
XFILLER_43_92 VPWR VGND sg13g2_decap_8
XFILLER_9_444 VPWR VGND sg13g2_decap_8
X_397_ net48 _091_ VPWR VGND sg13g2_buf_1
XFILLER_40_270 VPWR VGND sg13g2_decap_8
XFILLER_41_771 VPWR VGND sg13g2_decap_8
XFILLER_9_477 VPWR VGND sg13g2_decap_8
Xheichips25_template_5 VPWR VGND uio_out[0] sg13g2_tielo
XFILLER_5_661 VPWR VGND sg13g2_decap_8
XFILLER_4_193 VPWR VGND sg13g2_decap_8
XFILLER_4_53 VPWR VGND sg13g2_decap_8
XFILLER_24_727 VPWR VGND sg13g2_decap_8
XFILLER_36_576 VPWR VGND sg13g2_decap_8
XFILLER_23_215 VPWR VGND sg13g2_decap_8
XFILLER_17_1013 VPWR VGND sg13g2_decap_8
XFILLER_32_760 VPWR VGND sg13g2_decap_8
XFILLER_20_955 VPWR VGND sg13g2_decap_8
XFILLER_47_819 VPWR VGND sg13g2_decap_8
XFILLER_24_1028 VPWR VGND sg13g2_fill_1
XFILLER_27_554 VPWR VGND sg13g2_decap_8
X_320_ _186_ net148 net45 VPWR VGND sg13g2_nand2_1
XFILLER_14_237 VPWR VGND sg13g2_decap_8
XFILLER_42_568 VPWR VGND sg13g2_decap_8
XFILLER_11_900 VPWR VGND sg13g2_decap_8
Xfanout63 net72 net63 VPWR VGND sg13g2_buf_8
Xfanout74 net85 net74 VPWR VGND sg13g2_buf_8
XFILLER_23_793 VPWR VGND sg13g2_decap_8
X_251_ mac2.sum_lvl1_ff\[9\] mac2.sum_lvl1_ff\[1\] _149_ VPWR VGND sg13g2_xor2_1
XFILLER_7_904 VPWR VGND sg13g2_decap_8
XFILLER_11_977 VPWR VGND sg13g2_decap_8
Xfanout85 rst_n net85 VPWR VGND sg13g2_buf_8
XFILLER_13_95 VPWR VGND sg13g2_decap_8
XFILLER_2_642 VPWR VGND sg13g2_decap_8
XFILLER_1_130 VPWR VGND sg13g2_decap_8
XFILLER_49_112 VPWR VGND sg13g2_decap_8
XFILLER_49_156 VPWR VGND sg13g2_decap_8
XFILLER_46_830 VPWR VGND sg13g2_decap_8
XFILLER_45_384 VPWR VGND sg13g2_decap_8
XFILLER_33_524 VPWR VGND sg13g2_decap_8
XFILLER_21_708 VPWR VGND sg13g2_decap_8
X_518_ net71 VGND VPWR net186 mac2.sum_lvl2_ff\[1\] clknet_5_12__leaf_clk sg13g2_dfrbpq_1
XFILLER_20_207 VPWR VGND sg13g2_decap_8
X_449_ net81 VGND VPWR _043_ mac1.products_ff\[1\] clknet_5_31__leaf_clk sg13g2_dfrbpq_1
XFILLER_13_281 VPWR VGND sg13g2_decap_8
XFILLER_6_970 VPWR VGND sg13g2_decap_8
XFILLER_18_18 VPWR VGND sg13g2_decap_8
XFILLER_36_340 VPWR VGND sg13g2_decap_8
XFILLER_37_863 VPWR VGND sg13g2_decap_8
XFILLER_24_524 VPWR VGND sg13g2_decap_8
XFILLER_34_28 VPWR VGND sg13g2_decap_8
XFILLER_34_39 VPWR VGND sg13g2_fill_1
Xclkload5 VPWR clkload5/Y clknet_5_23__leaf_clk VGND sg13g2_inv_1
XFILLER_20_752 VPWR VGND sg13g2_decap_8
Xclkbuf_5_30__f_clk clknet_4_15_0_clk clknet_5_30__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_8_1000 VPWR VGND sg13g2_decap_8
XFILLER_47_616 VPWR VGND sg13g2_decap_8
XFILLER_46_126 VPWR VGND sg13g2_decap_8
XFILLER_43_811 VPWR VGND sg13g2_decap_8
XFILLER_28_896 VPWR VGND sg13g2_decap_8
XFILLER_43_888 VPWR VGND sg13g2_decap_8
XFILLER_15_557 VPWR VGND sg13g2_decap_8
XFILLER_42_365 VPWR VGND sg13g2_decap_8
X_303_ _178_ net181 net103 VPWR VGND sg13g2_nand2_1
XFILLER_23_590 VPWR VGND sg13g2_decap_8
XFILLER_24_61 VPWR VGND sg13g2_decap_8
X_234_ net159 net142 _042_ VPWR VGND sg13g2_and2_1
XFILLER_30_549 VPWR VGND sg13g2_decap_8
XFILLER_7_701 VPWR VGND sg13g2_decap_8
XFILLER_11_774 VPWR VGND sg13g2_decap_8
XFILLER_7_778 VPWR VGND sg13g2_decap_8
XFILLER_6_255 VPWR VGND sg13g2_decap_8
XFILLER_40_82 VPWR VGND sg13g2_decap_8
XFILLER_3_951 VPWR VGND sg13g2_decap_8
XFILLER_2_483 VPWR VGND sg13g2_fill_1
XFILLER_34_7 VPWR VGND sg13g2_decap_8
XFILLER_49_91 VPWR VGND sg13g2_decap_8
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_38_649 VPWR VGND sg13g2_decap_8
XFILLER_18_362 VPWR VGND sg13g2_decap_4
XFILLER_19_874 VPWR VGND sg13g2_decap_8
XFILLER_34_811 VPWR VGND sg13g2_decap_8
XFILLER_33_387 VPWR VGND sg13g2_decap_4
XFILLER_34_888 VPWR VGND sg13g2_decap_8
XFILLER_21_549 VPWR VGND sg13g2_decap_8
Xhold28 DP_4.matrix\[37\] VPWR VGND net52 sg13g2_dlygate4sd3_1
Xhold17 DP_3.matrix\[73\] VPWR VGND net41 sg13g2_dlygate4sd3_1
XFILLER_21_1009 VPWR VGND sg13g2_decap_8
XFILLER_29_638 VPWR VGND sg13g2_decap_8
Xhold39 DP_3.matrix\[55\] VPWR VGND net89 sg13g2_dlygate4sd3_1
XFILLER_44_619 VPWR VGND sg13g2_decap_8
XFILLER_37_660 VPWR VGND sg13g2_decap_8
XFILLER_45_49 VPWR VGND sg13g2_decap_4
XFILLER_25_844 VPWR VGND sg13g2_decap_8
XFILLER_24_332 VPWR VGND sg13g2_decap_8
XFILLER_36_181 VPWR VGND sg13g2_decap_8
XFILLER_24_376 VPWR VGND sg13g2_decap_8
XFILLER_40_869 VPWR VGND sg13g2_decap_8
XFILLER_4_759 VPWR VGND sg13g2_decap_8
XFILLER_10_41 VPWR VGND sg13g2_fill_2
XFILLER_0_910 VPWR VGND sg13g2_decap_8
XFILLER_0_987 VPWR VGND sg13g2_decap_8
XFILLER_48_958 VPWR VGND sg13g2_decap_8
XFILLER_19_137 VPWR VGND sg13g2_decap_8
XFILLER_16_844 VPWR VGND sg13g2_decap_8
XFILLER_28_693 VPWR VGND sg13g2_decap_8
XFILLER_15_354 VPWR VGND sg13g2_decap_8
XFILLER_43_685 VPWR VGND sg13g2_decap_8
XFILLER_30_302 VPWR VGND sg13g2_decap_8
XFILLER_31_825 VPWR VGND sg13g2_decap_8
XFILLER_35_82 VPWR VGND sg13g2_fill_1
XFILLER_7_575 VPWR VGND sg13g2_decap_8
XFILLER_39_903 VPWR VGND sg13g2_decap_8
Xheichips25_template_19 VPWR VGND uio_oe[2] sg13g2_tiehi
XFILLER_38_413 VPWR VGND sg13g2_decap_8
XFILLER_47_980 VPWR VGND sg13g2_decap_8
XFILLER_19_671 VPWR VGND sg13g2_decap_8
XFILLER_25_118 VPWR VGND sg13g2_decap_8
XFILLER_18_181 VPWR VGND sg13g2_decap_8
XFILLER_33_151 VPWR VGND sg13g2_decap_8
XFILLER_34_685 VPWR VGND sg13g2_decap_8
XFILLER_21_313 VPWR VGND sg13g2_fill_2
XFILLER_22_858 VPWR VGND sg13g2_decap_8
XFILLER_0_217 VPWR VGND sg13g2_decap_8
XFILLER_29_402 VPWR VGND sg13g2_decap_8
XFILLER_5_1025 VPWR VGND sg13g2_decap_4
XFILLER_44_416 VPWR VGND sg13g2_decap_8
XFILLER_16_118 VPWR VGND sg13g2_fill_2
XFILLER_25_641 VPWR VGND sg13g2_decap_8
XFILLER_13_858 VPWR VGND sg13g2_decap_8
XFILLER_24_173 VPWR VGND sg13g2_decap_8
XFILLER_9_829 VPWR VGND sg13g2_decap_8
XFILLER_12_379 VPWR VGND sg13g2_decap_8
XFILLER_40_666 VPWR VGND sg13g2_decap_8
XFILLER_8_339 VPWR VGND sg13g2_fill_2
XFILLER_4_534 VPWR VGND sg13g2_decap_8
XFILLER_4_567 VPWR VGND sg13g2_decap_8
XFILLER_48_755 VPWR VGND sg13g2_decap_8
XFILLER_0_784 VPWR VGND sg13g2_decap_8
XFILLER_16_641 VPWR VGND sg13g2_decap_8
XFILLER_44_983 VPWR VGND sg13g2_decap_8
XFILLER_15_140 VPWR VGND sg13g2_decap_8
XFILLER_43_482 VPWR VGND sg13g2_decap_8
XFILLER_31_622 VPWR VGND sg13g2_decap_8
XFILLER_31_699 VPWR VGND sg13g2_decap_8
XFILLER_7_42 VPWR VGND sg13g2_decap_8
XFILLER_11_1019 VPWR VGND sg13g2_decap_8
XFILLER_8_895 VPWR VGND sg13g2_decap_8
XFILLER_7_383 VPWR VGND sg13g2_decap_8
XFILLER_7_394 VPWR VGND sg13g2_fill_1
XFILLER_39_700 VPWR VGND sg13g2_decap_8
XFILLER_39_777 VPWR VGND sg13g2_decap_8
XFILLER_26_18 VPWR VGND sg13g2_decap_8
XFILLER_26_438 VPWR VGND sg13g2_decap_8
XFILLER_27_939 VPWR VGND sg13g2_decap_8
XFILLER_38_298 VPWR VGND sg13g2_decap_8
XFILLER_19_490 VPWR VGND sg13g2_decap_8
XFILLER_34_460 VPWR VGND sg13g2_decap_8
XFILLER_41_419 VPWR VGND sg13g2_decap_8
XFILLER_21_132 VPWR VGND sg13g2_decap_8
XFILLER_22_655 VPWR VGND sg13g2_decap_8
XFILLER_42_28 VPWR VGND sg13g2_fill_1
XFILLER_1_537 VPWR VGND sg13g2_decap_8
XFILLER_44_202 VPWR VGND sg13g2_decap_8
XFILLER_18_928 VPWR VGND sg13g2_decap_8
X_551_ net79 VGND VPWR _091_ DP_2.matrix\[10\] clknet_5_26__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_758 VPWR VGND sg13g2_decap_8
XFILLER_33_909 VPWR VGND sg13g2_decap_8
X_482_ net73 VGND VPWR net154 mac1.sum_lvl3_ff\[0\] clknet_5_16__leaf_clk sg13g2_dfrbpq_1
XFILLER_25_493 VPWR VGND sg13g2_fill_2
XFILLER_41_953 VPWR VGND sg13g2_decap_8
XFILLER_9_626 VPWR VGND sg13g2_decap_8
XFILLER_13_655 VPWR VGND sg13g2_decap_8
XFILLER_40_452 VPWR VGND sg13g2_decap_8
XFILLER_32_94 VPWR VGND sg13g2_decap_8
XFILLER_5_843 VPWR VGND sg13g2_decap_8
XFILLER_4_375 VPWR VGND sg13g2_decap_8
XFILLER_0_581 VPWR VGND sg13g2_decap_8
XFILLER_48_552 VPWR VGND sg13g2_decap_8
XFILLER_17_950 VPWR VGND sg13g2_decap_8
XFILLER_24_909 VPWR VGND sg13g2_decap_8
XFILLER_36_758 VPWR VGND sg13g2_decap_8
XFILLER_23_408 VPWR VGND sg13g2_fill_2
XFILLER_23_419 VPWR VGND sg13g2_fill_2
XFILLER_44_780 VPWR VGND sg13g2_decap_8
XFILLER_32_942 VPWR VGND sg13g2_decap_8
XFILLER_31_496 VPWR VGND sg13g2_decap_8
XFILLER_8_692 VPWR VGND sg13g2_decap_8
Xhold103 mac1.sum_lvl2_ff\[4\] VPWR VGND net153 sg13g2_dlygate4sd3_1
Xhold125 mac1.sum_lvl1_ff\[8\] VPWR VGND net175 sg13g2_dlygate4sd3_1
Xhold114 _000_ VPWR VGND net164 sg13g2_dlygate4sd3_1
Xhold147 mac1.sum_lvl2_ff\[0\] VPWR VGND net197 sg13g2_dlygate4sd3_1
Xhold136 _031_ VPWR VGND net186 sg13g2_dlygate4sd3_1
XFILLER_37_28 VPWR VGND sg13g2_decap_8
XFILLER_2_1006 VPWR VGND sg13g2_decap_8
XFILLER_27_736 VPWR VGND sg13g2_decap_8
XFILLER_39_574 VPWR VGND sg13g2_decap_8
XFILLER_41_216 VPWR VGND sg13g2_decap_8
XFILLER_23_975 VPWR VGND sg13g2_decap_8
XFILLER_10_669 VPWR VGND sg13g2_decap_8
XFILLER_2_824 VPWR VGND sg13g2_decap_8
XFILLER_1_334 VPWR VGND sg13g2_decap_8
XFILLER_49_338 VPWR VGND sg13g2_decap_8
XFILLER_40_1023 VPWR VGND sg13g2_decap_4
XFILLER_18_725 VPWR VGND sg13g2_decap_8
XFILLER_45_555 VPWR VGND sg13g2_decap_8
XFILLER_17_235 VPWR VGND sg13g2_decap_8
X_534_ net64 VGND VPWR _074_ DP_1.matrix\[18\] clknet_5_18__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_279 VPWR VGND sg13g2_decap_8
XFILLER_27_83 VPWR VGND sg13g2_decap_8
XFILLER_33_706 VPWR VGND sg13g2_decap_8
X_465_ net61 VGND VPWR _069_ mac1.products_ff\[137\] clknet_5_4__leaf_clk sg13g2_dfrbpq_1
XFILLER_14_931 VPWR VGND sg13g2_decap_8
XFILLER_41_750 VPWR VGND sg13g2_decap_8
XFILLER_43_71 VPWR VGND sg13g2_decap_8
XFILLER_9_423 VPWR VGND sg13g2_decap_8
XFILLER_13_485 VPWR VGND sg13g2_decap_8
X_396_ net128 _090_ VPWR VGND sg13g2_buf_1
XFILLER_9_467 VPWR VGND sg13g2_fill_1
Xheichips25_template_6 VPWR VGND uio_out[1] sg13g2_tielo
XFILLER_5_640 VPWR VGND sg13g2_decap_8
XFILLER_4_172 VPWR VGND sg13g2_decap_8
XFILLER_4_32 VPWR VGND sg13g2_decap_8
XFILLER_48_393 VPWR VGND sg13g2_fill_2
XFILLER_24_706 VPWR VGND sg13g2_decap_8
XFILLER_36_555 VPWR VGND sg13g2_decap_8
XFILLER_20_934 VPWR VGND sg13g2_decap_8
XFILLER_9_990 VPWR VGND sg13g2_decap_8
XFILLER_48_49 VPWR VGND sg13g2_decap_8
XFILLER_24_1007 VPWR VGND sg13g2_decap_8
XFILLER_27_533 VPWR VGND sg13g2_decap_8
XFILLER_42_547 VPWR VGND sg13g2_decap_8
XFILLER_14_216 VPWR VGND sg13g2_decap_8
Xfanout64 net66 net64 VPWR VGND sg13g2_buf_8
XFILLER_23_772 VPWR VGND sg13g2_decap_8
X_250_ _148_ net185 net107 VPWR VGND sg13g2_nand2_1
Xfanout75 net78 net75 VPWR VGND sg13g2_buf_8
XFILLER_11_956 VPWR VGND sg13g2_decap_8
XFILLER_10_466 VPWR VGND sg13g2_fill_1
XFILLER_13_74 VPWR VGND sg13g2_decap_8
XFILLER_6_448 VPWR VGND sg13g2_decap_8
XFILLER_2_621 VPWR VGND sg13g2_decap_8
XFILLER_2_698 VPWR VGND sg13g2_decap_8
XFILLER_49_135 VPWR VGND sg13g2_decap_8
XFILLER_37_319 VPWR VGND sg13g2_decap_8
XFILLER_46_886 VPWR VGND sg13g2_decap_8
XFILLER_18_577 VPWR VGND sg13g2_decap_8
XFILLER_33_503 VPWR VGND sg13g2_decap_8
X_517_ net71 VGND VPWR net108 mac2.sum_lvl2_ff\[0\] clknet_5_12__leaf_clk sg13g2_dfrbpq_1
XFILLER_13_260 VPWR VGND sg13g2_decap_8
X_448_ net79 VGND VPWR _042_ mac1.products_ff\[0\] clknet_5_25__leaf_clk sg13g2_dfrbpq_1
X_379_ net97 _073_ VPWR VGND sg13g2_buf_1
XFILLER_5_492 VPWR VGND sg13g2_decap_8
XFILLER_37_842 VPWR VGND sg13g2_decap_8
XFILLER_24_503 VPWR VGND sg13g2_decap_8
XFILLER_24_514 VPWR VGND sg13g2_fill_2
XFILLER_36_396 VPWR VGND sg13g2_decap_8
XFILLER_20_731 VPWR VGND sg13g2_decap_8
Xclkload6 VPWR clkload6/Y clknet_5_27__leaf_clk VGND sg13g2_inv_1
XFILLER_30_1011 VPWR VGND sg13g2_decap_8
XFILLER_3_407 VPWR VGND sg13g2_fill_1
XFILLER_3_429 VPWR VGND sg13g2_decap_8
XFILLER_28_875 VPWR VGND sg13g2_decap_8
XFILLER_15_536 VPWR VGND sg13g2_decap_8
XFILLER_43_867 VPWR VGND sg13g2_decap_8
XFILLER_42_344 VPWR VGND sg13g2_decap_8
XFILLER_24_40 VPWR VGND sg13g2_decap_8
XFILLER_30_528 VPWR VGND sg13g2_decap_8
X_302_ net109 mac2.products_ff\[51\] _024_ VPWR VGND sg13g2_xor2_1
X_233_ net157 net152 _040_ VPWR VGND sg13g2_and2_1
XFILLER_10_241 VPWR VGND sg13g2_decap_8
XFILLER_11_753 VPWR VGND sg13g2_decap_8
XFILLER_10_274 VPWR VGND sg13g2_decap_8
XFILLER_7_757 VPWR VGND sg13g2_decap_8
XFILLER_6_234 VPWR VGND sg13g2_decap_8
XFILLER_40_61 VPWR VGND sg13g2_decap_8
XFILLER_3_930 VPWR VGND sg13g2_decap_8
XFILLER_2_451 VPWR VGND sg13g2_fill_1
XFILLER_49_70 VPWR VGND sg13g2_decap_8
XFILLER_27_7 VPWR VGND sg13g2_decap_8
XFILLER_37_105 VPWR VGND sg13g2_decap_8
XFILLER_38_628 VPWR VGND sg13g2_decap_8
XFILLER_18_341 VPWR VGND sg13g2_decap_8
XFILLER_19_853 VPWR VGND sg13g2_decap_8
XFILLER_37_149 VPWR VGND sg13g2_decap_8
XFILLER_46_683 VPWR VGND sg13g2_decap_8
XFILLER_45_160 VPWR VGND sg13g2_decap_8
XFILLER_34_867 VPWR VGND sg13g2_decap_8
XFILLER_21_528 VPWR VGND sg13g2_decap_8
Xhold18 DP_4.matrix\[10\] VPWR VGND net42 sg13g2_dlygate4sd3_1
Xhold29 DP_2.matrix\[28\] VPWR VGND net53 sg13g2_dlygate4sd3_1
XFILLER_28_105 VPWR VGND sg13g2_decap_4
XFILLER_29_617 VPWR VGND sg13g2_decap_8
XFILLER_45_28 VPWR VGND sg13g2_decap_8
XFILLER_24_311 VPWR VGND sg13g2_decap_8
XFILLER_25_823 VPWR VGND sg13g2_decap_8
XFILLER_36_160 VPWR VGND sg13g2_decap_8
XFILLER_24_355 VPWR VGND sg13g2_fill_1
XFILLER_40_848 VPWR VGND sg13g2_decap_8
XFILLER_4_738 VPWR VGND sg13g2_decap_8
XFILLER_3_204 VPWR VGND sg13g2_decap_8
XFILLER_0_966 VPWR VGND sg13g2_decap_8
XFILLER_48_937 VPWR VGND sg13g2_decap_8
XFILLER_19_116 VPWR VGND sg13g2_decap_8
XFILLER_47_469 VPWR VGND sg13g2_decap_8
XFILLER_19_95 VPWR VGND sg13g2_decap_8
XFILLER_16_823 VPWR VGND sg13g2_decap_8
XFILLER_28_672 VPWR VGND sg13g2_decap_8
XFILLER_15_322 VPWR VGND sg13g2_decap_4
XFILLER_27_182 VPWR VGND sg13g2_decap_8
XFILLER_35_61 VPWR VGND sg13g2_decap_8
XFILLER_43_664 VPWR VGND sg13g2_decap_8
XFILLER_31_804 VPWR VGND sg13g2_decap_8
XFILLER_37_1017 VPWR VGND sg13g2_decap_8
XFILLER_37_1028 VPWR VGND sg13g2_fill_1
XFILLER_42_185 VPWR VGND sg13g2_decap_8
XFILLER_30_358 VPWR VGND sg13g2_decap_8
XFILLER_25_4 VPWR VGND sg13g2_decap_8
XFILLER_39_959 VPWR VGND sg13g2_decap_8
XFILLER_19_650 VPWR VGND sg13g2_decap_8
XFILLER_38_458 VPWR VGND sg13g2_decap_8
XFILLER_46_480 VPWR VGND sg13g2_decap_8
XFILLER_33_130 VPWR VGND sg13g2_decap_8
XFILLER_34_664 VPWR VGND sg13g2_decap_8
XFILLER_22_837 VPWR VGND sg13g2_decap_8
XFILLER_21_358 VPWR VGND sg13g2_decap_8
XFILLER_30_892 VPWR VGND sg13g2_decap_8
XFILLER_1_719 VPWR VGND sg13g2_decap_8
XFILLER_5_1004 VPWR VGND sg13g2_decap_8
XFILLER_38_992 VPWR VGND sg13g2_decap_8
XFILLER_25_620 VPWR VGND sg13g2_decap_8
XFILLER_24_152 VPWR VGND sg13g2_decap_8
XFILLER_9_808 VPWR VGND sg13g2_decap_8
XFILLER_13_837 VPWR VGND sg13g2_decap_8
XFILLER_25_697 VPWR VGND sg13g2_decap_8
XFILLER_40_645 VPWR VGND sg13g2_decap_8
XFILLER_12_358 VPWR VGND sg13g2_decap_8
XFILLER_4_513 VPWR VGND sg13g2_decap_8
XFILLER_43_1021 VPWR VGND sg13g2_decap_8
XFILLER_0_763 VPWR VGND sg13g2_decap_8
XFILLER_48_734 VPWR VGND sg13g2_decap_8
XFILLER_29_981 VPWR VGND sg13g2_decap_8
XFILLER_35_417 VPWR VGND sg13g2_decap_8
XFILLER_16_620 VPWR VGND sg13g2_decap_8
XFILLER_44_962 VPWR VGND sg13g2_decap_8
XFILLER_43_461 VPWR VGND sg13g2_decap_8
XFILLER_31_601 VPWR VGND sg13g2_decap_8
XFILLER_16_697 VPWR VGND sg13g2_decap_8
XFILLER_30_122 VPWR VGND sg13g2_decap_8
XFILLER_30_133 VPWR VGND sg13g2_fill_1
XFILLER_31_678 VPWR VGND sg13g2_decap_8
XFILLER_7_21 VPWR VGND sg13g2_decap_8
XFILLER_30_177 VPWR VGND sg13g2_decap_8
XFILLER_8_874 VPWR VGND sg13g2_decap_8
XFILLER_7_362 VPWR VGND sg13g2_decap_8
XFILLER_7_98 VPWR VGND sg13g2_decap_8
XFILLER_27_918 VPWR VGND sg13g2_decap_8
XFILLER_38_244 VPWR VGND sg13g2_decap_8
XFILLER_39_756 VPWR VGND sg13g2_decap_8
XFILLER_26_417 VPWR VGND sg13g2_decap_8
XFILLER_38_288 VPWR VGND sg13g2_fill_1
XFILLER_35_984 VPWR VGND sg13g2_decap_8
XFILLER_22_634 VPWR VGND sg13g2_decap_8
XFILLER_1_516 VPWR VGND sg13g2_decap_8
XFILLER_27_1016 VPWR VGND sg13g2_decap_8
XFILLER_27_1027 VPWR VGND sg13g2_fill_2
XFILLER_18_907 VPWR VGND sg13g2_decap_8
XFILLER_45_737 VPWR VGND sg13g2_decap_8
X_550_ net79 VGND VPWR _090_ DP_2.matrix\[9\] clknet_5_26__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_269 VPWR VGND sg13g2_decap_8
X_481_ net64 VGND VPWR net31 mac1.sum_lvl2_ff\[9\] clknet_5_5__leaf_clk sg13g2_dfrbpq_1
XFILLER_26_984 VPWR VGND sg13g2_decap_8
XFILLER_32_409 VPWR VGND sg13g2_decap_4
XFILLER_12_111 VPWR VGND sg13g2_decap_8
XFILLER_13_634 VPWR VGND sg13g2_decap_8
XFILLER_16_63 VPWR VGND sg13g2_decap_4
XFILLER_25_472 VPWR VGND sg13g2_decap_8
XFILLER_41_932 VPWR VGND sg13g2_decap_8
XFILLER_9_605 VPWR VGND sg13g2_decap_8
XFILLER_12_144 VPWR VGND sg13g2_decap_8
XFILLER_8_148 VPWR VGND sg13g2_decap_8
XFILLER_32_73 VPWR VGND sg13g2_decap_8
XFILLER_5_822 VPWR VGND sg13g2_decap_8
XFILLER_4_332 VPWR VGND sg13g2_decap_8
XFILLER_5_899 VPWR VGND sg13g2_decap_8
XFILLER_4_354 VPWR VGND sg13g2_decap_8
XFILLER_0_560 VPWR VGND sg13g2_decap_8
XFILLER_48_531 VPWR VGND sg13g2_decap_8
XFILLER_35_203 VPWR VGND sg13g2_decap_8
XFILLER_36_737 VPWR VGND sg13g2_decap_8
XFILLER_32_921 VPWR VGND sg13g2_decap_8
XFILLER_31_475 VPWR VGND sg13g2_decap_8
XFILLER_32_998 VPWR VGND sg13g2_decap_8
XFILLER_8_671 VPWR VGND sg13g2_decap_8
Xhold104 _014_ VPWR VGND net154 sg13g2_dlygate4sd3_1
Xhold115 mac1.sum_lvl3_ff\[2\] VPWR VGND net165 sg13g2_dlygate4sd3_1
Xhold126 _011_ VPWR VGND net176 sg13g2_dlygate4sd3_1
Xhold148 _015_ VPWR VGND net198 sg13g2_dlygate4sd3_1
Xhold137 mac1.products_ff\[85\] VPWR VGND net187 sg13g2_dlygate4sd3_1
XFILLER_39_553 VPWR VGND sg13g2_decap_8
XFILLER_27_715 VPWR VGND sg13g2_decap_8
XFILLER_42_729 VPWR VGND sg13g2_decap_8
XFILLER_26_247 VPWR VGND sg13g2_decap_8
XFILLER_35_781 VPWR VGND sg13g2_decap_8
XFILLER_23_954 VPWR VGND sg13g2_decap_8
XFILLER_34_280 VPWR VGND sg13g2_fill_2
XFILLER_22_475 VPWR VGND sg13g2_decap_8
XFILLER_10_648 VPWR VGND sg13g2_decap_8
XFILLER_2_803 VPWR VGND sg13g2_decap_8
XFILLER_1_313 VPWR VGND sg13g2_decap_8
Xclkbuf_5_13__f_clk clknet_4_6_0_clk clknet_5_13__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_49_317 VPWR VGND sg13g2_decap_8
XFILLER_40_1002 VPWR VGND sg13g2_decap_8
XFILLER_18_704 VPWR VGND sg13g2_decap_8
XFILLER_45_534 VPWR VGND sg13g2_decap_8
XFILLER_17_214 VPWR VGND sg13g2_decap_8
XFILLER_27_62 VPWR VGND sg13g2_decap_8
X_533_ net79 VGND VPWR _073_ DP_1.matrix\[10\] clknet_5_24__leaf_clk sg13g2_dfrbpq_1
X_464_ net61 VGND VPWR _068_ mac1.products_ff\[136\] clknet_5_4__leaf_clk sg13g2_dfrbpq_1
XFILLER_14_910 VPWR VGND sg13g2_decap_8
XFILLER_26_781 VPWR VGND sg13g2_decap_8
XFILLER_25_280 VPWR VGND sg13g2_decap_8
XFILLER_13_464 VPWR VGND sg13g2_decap_8
XFILLER_14_987 VPWR VGND sg13g2_decap_8
X_395_ net38 _089_ VPWR VGND sg13g2_buf_1
Xheichips25_template_7 VPWR VGND uio_out[2] sg13g2_tielo
XFILLER_4_151 VPWR VGND sg13g2_decap_8
XFILLER_5_696 VPWR VGND sg13g2_decap_8
XFILLER_4_11 VPWR VGND sg13g2_decap_8
XFILLER_4_88 VPWR VGND sg13g2_decap_8
XFILLER_1_880 VPWR VGND sg13g2_decap_8
XFILLER_49_884 VPWR VGND sg13g2_decap_8
XFILLER_48_372 VPWR VGND sg13g2_decap_8
XFILLER_36_534 VPWR VGND sg13g2_decap_8
XFILLER_20_913 VPWR VGND sg13g2_decap_8
XFILLER_31_294 VPWR VGND sg13g2_decap_8
XFILLER_32_795 VPWR VGND sg13g2_decap_8
XFILLER_48_28 VPWR VGND sg13g2_decap_8
XFILLER_42_526 VPWR VGND sg13g2_decap_8
XFILLER_15_729 VPWR VGND sg13g2_decap_8
XFILLER_27_589 VPWR VGND sg13g2_decap_8
XFILLER_23_751 VPWR VGND sg13g2_decap_8
Xfanout65 net66 net65 VPWR VGND sg13g2_buf_8
Xfanout76 net78 net76 VPWR VGND sg13g2_buf_2
XFILLER_11_935 VPWR VGND sg13g2_decap_8
XFILLER_10_445 VPWR VGND sg13g2_decap_8
XFILLER_7_939 VPWR VGND sg13g2_decap_8
XFILLER_6_427 VPWR VGND sg13g2_decap_8
XFILLER_13_53 VPWR VGND sg13g2_decap_8
XFILLER_2_600 VPWR VGND sg13g2_decap_8
XFILLER_1_165 VPWR VGND sg13g2_decap_4
XFILLER_2_677 VPWR VGND sg13g2_decap_8
XFILLER_1_187 VPWR VGND sg13g2_decap_8
XFILLER_45_320 VPWR VGND sg13g2_decap_8
XFILLER_18_512 VPWR VGND sg13g2_decap_8
XFILLER_38_83 VPWR VGND sg13g2_decap_8
XFILLER_46_865 VPWR VGND sg13g2_decap_8
XFILLER_18_556 VPWR VGND sg13g2_decap_8
X_516_ net63 VGND VPWR net29 mac2.sum_lvl1_ff\[33\] clknet_5_3__leaf_clk sg13g2_dfrbpq_1
XFILLER_18_589 VPWR VGND sg13g2_decap_8
XFILLER_33_559 VPWR VGND sg13g2_decap_8
X_447_ net43 _141_ VPWR VGND sg13g2_buf_1
XFILLER_14_784 VPWR VGND sg13g2_decap_8
X_378_ net147 _072_ VPWR VGND sg13g2_buf_1
XFILLER_9_287 VPWR VGND sg13g2_decap_8
XFILLER_47_1008 VPWR VGND sg13g2_decap_8
XFILLER_49_681 VPWR VGND sg13g2_decap_8
XFILLER_37_821 VPWR VGND sg13g2_decap_8
XFILLER_36_375 VPWR VGND sg13g2_decap_8
XFILLER_37_898 VPWR VGND sg13g2_decap_8
XFILLER_24_559 VPWR VGND sg13g2_decap_8
XFILLER_11_209 VPWR VGND sg13g2_decap_8
XFILLER_20_710 VPWR VGND sg13g2_decap_8
XFILLER_32_592 VPWR VGND sg13g2_decap_8
Xclkload7 VPWR clkload7/Y clknet_5_31__leaf_clk VGND sg13g2_inv_1
XFILLER_20_787 VPWR VGND sg13g2_decap_8
XFILLER_28_854 VPWR VGND sg13g2_decap_8
XFILLER_15_515 VPWR VGND sg13g2_decap_8
XFILLER_27_364 VPWR VGND sg13g2_decap_8
XFILLER_43_846 VPWR VGND sg13g2_decap_8
XFILLER_42_323 VPWR VGND sg13g2_decap_8
XFILLER_30_507 VPWR VGND sg13g2_decap_8
X_301_ _025_ _176_ _177_ VPWR VGND sg13g2_xnor2_1
X_232_ _018_ _142_ _145_ VPWR VGND sg13g2_xnor2_1
XFILLER_11_732 VPWR VGND sg13g2_decap_8
XFILLER_24_96 VPWR VGND sg13g2_decap_8
XFILLER_7_736 VPWR VGND sg13g2_decap_8
XFILLER_6_213 VPWR VGND sg13g2_decap_8
XFILLER_2_430 VPWR VGND sg13g2_decap_8
XFILLER_3_986 VPWR VGND sg13g2_decap_8
XFILLER_38_607 VPWR VGND sg13g2_decap_8
XFILLER_1_56 VPWR VGND sg13g2_decap_8
XFILLER_19_832 VPWR VGND sg13g2_decap_8
XFILLER_37_128 VPWR VGND sg13g2_decap_8
XFILLER_46_662 VPWR VGND sg13g2_decap_8
XFILLER_18_320 VPWR VGND sg13g2_decap_8
XFILLER_33_301 VPWR VGND sg13g2_fill_1
XFILLER_45_194 VPWR VGND sg13g2_decap_8
XFILLER_18_397 VPWR VGND sg13g2_decap_8
XFILLER_34_846 VPWR VGND sg13g2_decap_8
XFILLER_21_507 VPWR VGND sg13g2_decap_8
XFILLER_42_890 VPWR VGND sg13g2_decap_8
XFILLER_14_581 VPWR VGND sg13g2_decap_8
XFILLER_46_0 VPWR VGND sg13g2_decap_8
Xhold19 DP_4.matrix\[73\] VPWR VGND net43 sg13g2_dlygate4sd3_1
XFILLER_28_117 VPWR VGND sg13g2_decap_8
XFILLER_25_802 VPWR VGND sg13g2_decap_8
XFILLER_37_695 VPWR VGND sg13g2_decap_8
XFILLER_25_879 VPWR VGND sg13g2_decap_8
XFILLER_40_827 VPWR VGND sg13g2_decap_8
XFILLER_20_584 VPWR VGND sg13g2_decap_8
XFILLER_4_717 VPWR VGND sg13g2_decap_8
XFILLER_0_945 VPWR VGND sg13g2_decap_8
XFILLER_48_916 VPWR VGND sg13g2_decap_8
XFILLER_19_74 VPWR VGND sg13g2_decap_8
XFILLER_47_448 VPWR VGND sg13g2_decap_8
XFILLER_28_651 VPWR VGND sg13g2_decap_8
XFILLER_16_802 VPWR VGND sg13g2_decap_8
XFILLER_27_150 VPWR VGND sg13g2_fill_2
XFILLER_27_161 VPWR VGND sg13g2_decap_8
XFILLER_34_109 VPWR VGND sg13g2_decap_8
XFILLER_43_643 VPWR VGND sg13g2_decap_8
XFILLER_16_879 VPWR VGND sg13g2_decap_8
XFILLER_15_389 VPWR VGND sg13g2_decap_8
XFILLER_30_337 VPWR VGND sg13g2_decap_8
XFILLER_7_544 VPWR VGND sg13g2_fill_2
XFILLER_3_783 VPWR VGND sg13g2_decap_8
XFILLER_2_293 VPWR VGND sg13g2_decap_8
XFILLER_18_4 VPWR VGND sg13g2_decap_8
XFILLER_39_938 VPWR VGND sg13g2_decap_8
XFILLER_20_1011 VPWR VGND sg13g2_decap_8
XFILLER_18_161 VPWR VGND sg13g2_decap_4
XFILLER_34_643 VPWR VGND sg13g2_decap_8
XFILLER_22_816 VPWR VGND sg13g2_decap_8
XFILLER_15_890 VPWR VGND sg13g2_decap_8
XFILLER_21_315 VPWR VGND sg13g2_fill_1
XFILLER_33_186 VPWR VGND sg13g2_decap_4
XFILLER_30_871 VPWR VGND sg13g2_decap_8
XFILLER_29_437 VPWR VGND sg13g2_fill_1
XFILLER_45_919 VPWR VGND sg13g2_decap_8
XFILLER_38_971 VPWR VGND sg13g2_decap_8
XFILLER_37_492 VPWR VGND sg13g2_decap_8
XFILLER_13_816 VPWR VGND sg13g2_decap_8
XFILLER_24_131 VPWR VGND sg13g2_decap_8
XFILLER_25_676 VPWR VGND sg13g2_decap_8
XFILLER_12_315 VPWR VGND sg13g2_fill_2
XFILLER_40_624 VPWR VGND sg13g2_decap_8
XFILLER_20_381 VPWR VGND sg13g2_decap_8
XFILLER_21_97 VPWR VGND sg13g2_decap_4
XFILLER_43_1000 VPWR VGND sg13g2_decap_8
XFILLER_0_742 VPWR VGND sg13g2_decap_8
XFILLER_48_713 VPWR VGND sg13g2_decap_8
XFILLER_36_919 VPWR VGND sg13g2_decap_8
XFILLER_47_289 VPWR VGND sg13g2_decap_4
XFILLER_29_960 VPWR VGND sg13g2_decap_8
XFILLER_46_94 VPWR VGND sg13g2_decap_8
XFILLER_44_941 VPWR VGND sg13g2_decap_8
XFILLER_43_440 VPWR VGND sg13g2_decap_8
XFILLER_16_676 VPWR VGND sg13g2_decap_8
XFILLER_15_175 VPWR VGND sg13g2_decap_8
XFILLER_31_657 VPWR VGND sg13g2_decap_8
XFILLER_8_853 VPWR VGND sg13g2_decap_8
XFILLER_7_341 VPWR VGND sg13g2_decap_8
XFILLER_11_381 VPWR VGND sg13g2_decap_8
XFILLER_12_893 VPWR VGND sg13g2_decap_8
XFILLER_7_77 VPWR VGND sg13g2_decap_8
XFILLER_39_735 VPWR VGND sg13g2_decap_8
XFILLER_38_223 VPWR VGND sg13g2_decap_8
XFILLER_35_963 VPWR VGND sg13g2_decap_8
XFILLER_22_613 VPWR VGND sg13g2_decap_8
XFILLER_45_716 VPWR VGND sg13g2_decap_8
XFILLER_29_278 VPWR VGND sg13g2_decap_8
X_480_ net64 VGND VPWR net35 mac1.sum_lvl2_ff\[8\] clknet_5_5__leaf_clk sg13g2_dfrbpq_1
XFILLER_16_42 VPWR VGND sg13g2_decap_8
XFILLER_25_451 VPWR VGND sg13g2_decap_8
XFILLER_26_963 VPWR VGND sg13g2_decap_8
XFILLER_13_613 VPWR VGND sg13g2_decap_8
XFILLER_41_911 VPWR VGND sg13g2_decap_8
XFILLER_8_127 VPWR VGND sg13g2_decap_8
XFILLER_41_988 VPWR VGND sg13g2_decap_8
XFILLER_12_189 VPWR VGND sg13g2_fill_2
XFILLER_32_52 VPWR VGND sg13g2_decap_8
XFILLER_5_801 VPWR VGND sg13g2_decap_8
XFILLER_4_311 VPWR VGND sg13g2_decap_8
XFILLER_5_878 VPWR VGND sg13g2_decap_8
XFILLER_48_510 VPWR VGND sg13g2_decap_8
XFILLER_48_587 VPWR VGND sg13g2_decap_8
XFILLER_36_716 VPWR VGND sg13g2_decap_8
XFILLER_32_900 VPWR VGND sg13g2_decap_8
XFILLER_35_259 VPWR VGND sg13g2_decap_8
XFILLER_17_985 VPWR VGND sg13g2_decap_8
XFILLER_32_977 VPWR VGND sg13g2_decap_8
XFILLER_31_454 VPWR VGND sg13g2_decap_8
XFILLER_12_690 VPWR VGND sg13g2_decap_8
XFILLER_8_650 VPWR VGND sg13g2_decap_8
Xhold116 _017_ VPWR VGND net166 sg13g2_dlygate4sd3_1
XFILLER_7_182 VPWR VGND sg13g2_decap_8
Xhold105 DP_4.matrix\[27\] VPWR VGND net155 sg13g2_dlygate4sd3_1
Xhold138 _007_ VPWR VGND net188 sg13g2_dlygate4sd3_1
Xhold127 mac1.products_ff\[17\] VPWR VGND net177 sg13g2_dlygate4sd3_1
Xhold149 mac2.sum_lvl2_ff\[4\] VPWR VGND net199 sg13g2_dlygate4sd3_1
XFILLER_39_532 VPWR VGND sg13g2_decap_8
XFILLER_26_226 VPWR VGND sg13g2_decap_8
XFILLER_42_708 VPWR VGND sg13g2_decap_8
XFILLER_35_760 VPWR VGND sg13g2_decap_8
XFILLER_23_933 VPWR VGND sg13g2_decap_8
XFILLER_10_627 VPWR VGND sg13g2_decap_8
XFILLER_22_454 VPWR VGND sg13g2_decap_8
XFILLER_33_1021 VPWR VGND sg13g2_decap_8
XFILLER_2_859 VPWR VGND sg13g2_decap_8
XFILLER_1_369 VPWR VGND sg13g2_decap_8
X_601_ net62 VGND VPWR _141_ DP_4.matrix\[73\] clknet_5_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_513 VPWR VGND sg13g2_decap_8
XFILLER_17_259 VPWR VGND sg13g2_decap_4
X_532_ net79 VGND VPWR _072_ DP_1.matrix\[9\] clknet_5_26__leaf_clk sg13g2_dfrbpq_1
X_463_ net75 VGND VPWR _057_ mac1.products_ff\[120\] clknet_5_20__leaf_clk sg13g2_dfrbpq_1
XFILLER_26_760 VPWR VGND sg13g2_decap_8
XFILLER_32_207 VPWR VGND sg13g2_decap_8
XFILLER_13_432 VPWR VGND sg13g2_decap_8
XFILLER_14_966 VPWR VGND sg13g2_decap_8
X_394_ net142 _088_ VPWR VGND sg13g2_buf_1
XFILLER_40_240 VPWR VGND sg13g2_decap_8
XFILLER_41_785 VPWR VGND sg13g2_decap_8
XFILLER_9_458 VPWR VGND sg13g2_decap_8
XFILLER_40_284 VPWR VGND sg13g2_decap_8
Xheichips25_template_8 VPWR VGND uio_out[3] sg13g2_tielo
XFILLER_5_675 VPWR VGND sg13g2_decap_8
XFILLER_4_67 VPWR VGND sg13g2_decap_8
XFILLER_49_863 VPWR VGND sg13g2_decap_8
XFILLER_48_351 VPWR VGND sg13g2_decap_8
XFILLER_48_395 VPWR VGND sg13g2_fill_1
XFILLER_36_513 VPWR VGND sg13g2_decap_8
XFILLER_17_782 VPWR VGND sg13g2_decap_8
XFILLER_23_229 VPWR VGND sg13g2_fill_2
XFILLER_17_1027 VPWR VGND sg13g2_fill_2
XFILLER_32_774 VPWR VGND sg13g2_decap_8
XFILLER_31_273 VPWR VGND sg13g2_decap_8
XFILLER_20_969 VPWR VGND sg13g2_decap_8
XFILLER_8_491 VPWR VGND sg13g2_decap_4
XFILLER_27_502 VPWR VGND sg13g2_fill_2
XFILLER_15_708 VPWR VGND sg13g2_decap_8
XFILLER_27_568 VPWR VGND sg13g2_decap_8
XFILLER_42_505 VPWR VGND sg13g2_decap_8
XFILLER_23_730 VPWR VGND sg13g2_decap_8
XFILLER_10_402 VPWR VGND sg13g2_fill_2
XFILLER_11_914 VPWR VGND sg13g2_decap_8
XFILLER_10_424 VPWR VGND sg13g2_decap_8
XFILLER_13_32 VPWR VGND sg13g2_decap_8
Xfanout66 net72 net66 VPWR VGND sg13g2_buf_8
Xfanout77 net78 net77 VPWR VGND sg13g2_buf_8
XFILLER_22_273 VPWR VGND sg13g2_fill_2
XFILLER_22_295 VPWR VGND sg13g2_decap_8
XFILLER_7_918 VPWR VGND sg13g2_decap_8
XFILLER_2_656 VPWR VGND sg13g2_decap_8
XFILLER_1_144 VPWR VGND sg13g2_decap_8
XFILLER_38_62 VPWR VGND sg13g2_decap_8
XFILLER_46_844 VPWR VGND sg13g2_decap_8
X_515_ net62 VGND VPWR net25 mac2.sum_lvl1_ff\[32\] clknet_5_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_398 VPWR VGND sg13g2_fill_2
XFILLER_33_538 VPWR VGND sg13g2_decap_8
X_446_ net140 _140_ VPWR VGND sg13g2_buf_1
XFILLER_14_763 VPWR VGND sg13g2_decap_8
X_377_ net46 _071_ VPWR VGND sg13g2_buf_1
XFILLER_41_582 VPWR VGND sg13g2_decap_8
XFILLER_9_244 VPWR VGND sg13g2_decap_8
XFILLER_13_295 VPWR VGND sg13g2_decap_8
XFILLER_10_991 VPWR VGND sg13g2_decap_8
XFILLER_5_450 VPWR VGND sg13g2_decap_8
XFILLER_6_984 VPWR VGND sg13g2_decap_8
XFILLER_49_660 VPWR VGND sg13g2_decap_8
XFILLER_37_800 VPWR VGND sg13g2_decap_8
XFILLER_36_354 VPWR VGND sg13g2_decap_8
XFILLER_37_877 VPWR VGND sg13g2_decap_8
XFILLER_24_538 VPWR VGND sg13g2_decap_8
XFILLER_32_571 VPWR VGND sg13g2_decap_8
XFILLER_20_766 VPWR VGND sg13g2_decap_8
XFILLER_8_1014 VPWR VGND sg13g2_decap_8
XFILLER_28_833 VPWR VGND sg13g2_decap_8
XFILLER_27_343 VPWR VGND sg13g2_fill_2
XFILLER_43_825 VPWR VGND sg13g2_decap_8
XFILLER_42_302 VPWR VGND sg13g2_decap_8
X_300_ mac2.products_ff\[35\] mac2.products_ff\[52\] _177_ VPWR VGND sg13g2_xor2_1
XFILLER_42_379 VPWR VGND sg13g2_decap_8
XFILLER_24_20 VPWR VGND sg13g2_fill_1
XFILLER_10_210 VPWR VGND sg13g2_fill_1
X_231_ mac1.sum_lvl3_ff\[3\] net167 _145_ VPWR VGND sg13g2_xor2_1
XFILLER_11_711 VPWR VGND sg13g2_decap_8
XFILLER_24_75 VPWR VGND sg13g2_decap_8
XFILLER_7_715 VPWR VGND sg13g2_decap_8
XFILLER_11_788 VPWR VGND sg13g2_decap_8
XFILLER_6_269 VPWR VGND sg13g2_decap_8
XFILLER_3_965 VPWR VGND sg13g2_decap_8
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_19_811 VPWR VGND sg13g2_decap_8
XFILLER_46_641 VPWR VGND sg13g2_decap_8
XFILLER_18_376 VPWR VGND sg13g2_decap_8
XFILLER_19_888 VPWR VGND sg13g2_decap_8
XFILLER_34_825 VPWR VGND sg13g2_decap_8
XFILLER_45_173 VPWR VGND sg13g2_decap_8
XFILLER_14_560 VPWR VGND sg13g2_decap_8
X_429_ net41 _123_ VPWR VGND sg13g2_buf_1
XFILLER_14_1008 VPWR VGND sg13g2_decap_8
XFILLER_6_781 VPWR VGND sg13g2_decap_8
XFILLER_39_0 VPWR VGND sg13g2_decap_8
XFILLER_37_674 VPWR VGND sg13g2_decap_8
XFILLER_25_858 VPWR VGND sg13g2_decap_8
XFILLER_36_195 VPWR VGND sg13g2_decap_8
XFILLER_12_519 VPWR VGND sg13g2_decap_8
XFILLER_24_346 VPWR VGND sg13g2_decap_8
XFILLER_40_806 VPWR VGND sg13g2_decap_8
XFILLER_20_563 VPWR VGND sg13g2_decap_8
XFILLER_10_11 VPWR VGND sg13g2_fill_2
XFILLER_0_924 VPWR VGND sg13g2_decap_8
XFILLER_19_53 VPWR VGND sg13g2_decap_8
XFILLER_28_630 VPWR VGND sg13g2_decap_8
XFILLER_43_622 VPWR VGND sg13g2_decap_8
XFILLER_16_858 VPWR VGND sg13g2_decap_8
XFILLER_42_143 VPWR VGND sg13g2_fill_1
XFILLER_15_368 VPWR VGND sg13g2_decap_8
XFILLER_43_699 VPWR VGND sg13g2_decap_8
XFILLER_30_316 VPWR VGND sg13g2_decap_8
XFILLER_31_839 VPWR VGND sg13g2_decap_8
XFILLER_11_541 VPWR VGND sg13g2_fill_2
XFILLER_7_523 VPWR VGND sg13g2_decap_8
XFILLER_11_563 VPWR VGND sg13g2_fill_2
XFILLER_7_589 VPWR VGND sg13g2_decap_8
XFILLER_3_762 VPWR VGND sg13g2_decap_8
XFILLER_2_272 VPWR VGND sg13g2_decap_8
XFILLER_32_7 VPWR VGND sg13g2_decap_8
XFILLER_39_917 VPWR VGND sg13g2_decap_8
XFILLER_38_427 VPWR VGND sg13g2_decap_8
XFILLER_47_994 VPWR VGND sg13g2_decap_8
XFILLER_18_140 VPWR VGND sg13g2_decap_8
XFILLER_19_685 VPWR VGND sg13g2_decap_8
XFILLER_18_195 VPWR VGND sg13g2_decap_8
XFILLER_34_622 VPWR VGND sg13g2_decap_8
XFILLER_33_165 VPWR VGND sg13g2_decap_8
XFILLER_34_699 VPWR VGND sg13g2_decap_8
XFILLER_30_850 VPWR VGND sg13g2_decap_8
XFILLER_29_416 VPWR VGND sg13g2_decap_8
XFILLER_38_950 VPWR VGND sg13g2_decap_8
XFILLER_37_460 VPWR VGND sg13g2_decap_8
XFILLER_24_110 VPWR VGND sg13g2_decap_8
XFILLER_25_655 VPWR VGND sg13g2_decap_8
XFILLER_40_603 VPWR VGND sg13g2_decap_8
XFILLER_24_187 VPWR VGND sg13g2_decap_8
XFILLER_21_883 VPWR VGND sg13g2_decap_8
XFILLER_21_32 VPWR VGND sg13g2_decap_8
XFILLER_4_548 VPWR VGND sg13g2_decap_8
XFILLER_0_721 VPWR VGND sg13g2_decap_8
XFILLER_47_202 VPWR VGND sg13g2_decap_8
XFILLER_0_798 VPWR VGND sg13g2_decap_8
XFILLER_48_769 VPWR VGND sg13g2_decap_8
XFILLER_44_920 VPWR VGND sg13g2_decap_8
XFILLER_28_471 VPWR VGND sg13g2_decap_8
XFILLER_16_655 VPWR VGND sg13g2_decap_8
XFILLER_44_997 VPWR VGND sg13g2_decap_8
XFILLER_43_496 VPWR VGND sg13g2_decap_8
Xclkbuf_5_0__f_clk clknet_4_0_0_clk clknet_5_0__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_15_154 VPWR VGND sg13g2_decap_8
XFILLER_31_636 VPWR VGND sg13g2_decap_8
XFILLER_8_832 VPWR VGND sg13g2_decap_8
XFILLER_12_872 VPWR VGND sg13g2_decap_8
XFILLER_7_320 VPWR VGND sg13g2_decap_8
XFILLER_11_360 VPWR VGND sg13g2_decap_8
XFILLER_7_56 VPWR VGND sg13g2_decap_8
XFILLER_38_202 VPWR VGND sg13g2_decap_8
XFILLER_39_714 VPWR VGND sg13g2_decap_8
XFILLER_47_791 VPWR VGND sg13g2_decap_8
XFILLER_35_942 VPWR VGND sg13g2_decap_8
XFILLER_34_430 VPWR VGND sg13g2_decap_8
XFILLER_34_474 VPWR VGND sg13g2_decap_8
XFILLER_10_809 VPWR VGND sg13g2_decap_8
XFILLER_22_669 VPWR VGND sg13g2_decap_8
XFILLER_21_146 VPWR VGND sg13g2_decap_8
XFILLER_29_213 VPWR VGND sg13g2_decap_4
XFILLER_29_235 VPWR VGND sg13g2_decap_8
XFILLER_44_238 VPWR VGND sg13g2_decap_8
XFILLER_26_942 VPWR VGND sg13g2_decap_8
XFILLER_25_430 VPWR VGND sg13g2_decap_8
XFILLER_16_87 VPWR VGND sg13g2_fill_2
XFILLER_16_98 VPWR VGND sg13g2_decap_8
XFILLER_41_967 VPWR VGND sg13g2_decap_8
XFILLER_8_106 VPWR VGND sg13g2_fill_1
XFILLER_12_168 VPWR VGND sg13g2_decap_8
XFILLER_13_669 VPWR VGND sg13g2_decap_8
XFILLER_40_466 VPWR VGND sg13g2_decap_8
XFILLER_21_680 VPWR VGND sg13g2_decap_8
XFILLER_5_857 VPWR VGND sg13g2_decap_8
XFILLER_4_389 VPWR VGND sg13g2_fill_2
XFILLER_0_595 VPWR VGND sg13g2_decap_8
XFILLER_48_566 VPWR VGND sg13g2_decap_8
XFILLER_35_238 VPWR VGND sg13g2_decap_8
XFILLER_17_964 VPWR VGND sg13g2_decap_8
XFILLER_44_794 VPWR VGND sg13g2_decap_8
XFILLER_16_452 VPWR VGND sg13g2_decap_8
XFILLER_31_433 VPWR VGND sg13g2_fill_1
XFILLER_32_956 VPWR VGND sg13g2_decap_8
Xhold117 mac1.sum_lvl3_ff\[1\] VPWR VGND net167 sg13g2_dlygate4sd3_1
XFILLER_7_161 VPWR VGND sg13g2_decap_8
Xhold106 DP_3.matrix\[36\] VPWR VGND net156 sg13g2_dlygate4sd3_1
Xhold128 _003_ VPWR VGND net178 sg13g2_dlygate4sd3_1
Xhold139 mac2.sum_lvl1_ff\[16\] VPWR VGND net189 sg13g2_dlygate4sd3_1
XFILLER_26_205 VPWR VGND sg13g2_decap_8
XFILLER_39_588 VPWR VGND sg13g2_decap_8
XFILLER_23_912 VPWR VGND sg13g2_decap_8
XFILLER_22_433 VPWR VGND sg13g2_decap_8
XFILLER_34_282 VPWR VGND sg13g2_fill_1
XFILLER_10_606 VPWR VGND sg13g2_decap_8
XFILLER_23_989 VPWR VGND sg13g2_decap_8
XFILLER_33_1000 VPWR VGND sg13g2_decap_8
XFILLER_5_109 VPWR VGND sg13g2_decap_4
XFILLER_2_838 VPWR VGND sg13g2_decap_8
XFILLER_1_348 VPWR VGND sg13g2_decap_8
X_600_ net62 VGND VPWR _140_ DP_4.matrix\[72\] clknet_5_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_18_739 VPWR VGND sg13g2_decap_8
X_531_ net79 VGND VPWR _071_ DP_1.matrix\[1\] clknet_5_30__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_569 VPWR VGND sg13g2_decap_8
XFILLER_17_249 VPWR VGND sg13g2_decap_4
X_462_ net75 VGND VPWR _056_ mac1.products_ff\[119\] clknet_5_20__leaf_clk sg13g2_dfrbpq_1
XFILLER_27_97 VPWR VGND sg13g2_decap_8
X_393_ net91 _087_ VPWR VGND sg13g2_buf_1
XFILLER_14_945 VPWR VGND sg13g2_decap_8
XFILLER_41_764 VPWR VGND sg13g2_decap_8
XFILLER_43_85 VPWR VGND sg13g2_decap_8
XFILLER_9_437 VPWR VGND sg13g2_decap_8
XFILLER_13_499 VPWR VGND sg13g2_decap_8
Xheichips25_template_9 VPWR VGND uio_out[4] sg13g2_tielo
XFILLER_5_654 VPWR VGND sg13g2_decap_8
XFILLER_4_186 VPWR VGND sg13g2_decap_8
XFILLER_4_46 VPWR VGND sg13g2_decap_8
XFILLER_49_842 VPWR VGND sg13g2_decap_8
XFILLER_48_330 VPWR VGND sg13g2_decap_8
XFILLER_0_392 VPWR VGND sg13g2_decap_8
XFILLER_1_1020 VPWR VGND sg13g2_decap_8
XFILLER_36_569 VPWR VGND sg13g2_decap_8
XFILLER_17_761 VPWR VGND sg13g2_decap_8
XFILLER_23_208 VPWR VGND sg13g2_decap_8
XFILLER_44_591 VPWR VGND sg13g2_decap_8
XFILLER_16_293 VPWR VGND sg13g2_fill_1
XFILLER_17_1006 VPWR VGND sg13g2_decap_8
XFILLER_31_252 VPWR VGND sg13g2_decap_8
XFILLER_32_753 VPWR VGND sg13g2_decap_8
XFILLER_20_948 VPWR VGND sg13g2_decap_8
XFILLER_8_470 VPWR VGND sg13g2_decap_8
XFILLER_39_341 VPWR VGND sg13g2_decap_8
XFILLER_27_547 VPWR VGND sg13g2_decap_8
XFILLER_10_414 VPWR VGND sg13g2_fill_2
XFILLER_13_11 VPWR VGND sg13g2_decap_8
Xfanout78 net85 net78 VPWR VGND sg13g2_buf_8
XFILLER_23_786 VPWR VGND sg13g2_decap_8
Xfanout67 net69 net67 VPWR VGND sg13g2_buf_8
XFILLER_13_88 VPWR VGND sg13g2_decap_8
XFILLER_8_4 VPWR VGND sg13g2_decap_8
XFILLER_1_123 VPWR VGND sg13g2_decap_8
XFILLER_2_635 VPWR VGND sg13g2_decap_8
XFILLER_49_105 VPWR VGND sg13g2_decap_8
XFILLER_49_149 VPWR VGND sg13g2_decap_8
XFILLER_46_823 VPWR VGND sg13g2_decap_8
XFILLER_33_517 VPWR VGND sg13g2_decap_8
X_514_ net82 VGND VPWR net196 mac2.sum_lvl1_ff\[25\] clknet_5_27__leaf_clk sg13g2_dfrbpq_1
XFILLER_14_742 VPWR VGND sg13g2_decap_8
X_445_ net51 _139_ VPWR VGND sg13g2_buf_1
XFILLER_41_561 VPWR VGND sg13g2_decap_8
XFILLER_13_274 VPWR VGND sg13g2_decap_8
X_376_ net159 _070_ VPWR VGND sg13g2_buf_1
XFILLER_10_970 VPWR VGND sg13g2_decap_8
XFILLER_6_963 VPWR VGND sg13g2_decap_8
XFILLER_23_1010 VPWR VGND sg13g2_decap_8
XFILLER_36_333 VPWR VGND sg13g2_decap_8
XFILLER_37_856 VPWR VGND sg13g2_decap_8
XFILLER_32_550 VPWR VGND sg13g2_decap_8
XFILLER_20_745 VPWR VGND sg13g2_decap_8
XFILLER_30_1025 VPWR VGND sg13g2_decap_4
XFILLER_47_609 VPWR VGND sg13g2_decap_8
XFILLER_46_119 VPWR VGND sg13g2_decap_8
XFILLER_28_812 VPWR VGND sg13g2_decap_8
XFILLER_39_171 VPWR VGND sg13g2_decap_4
XFILLER_43_804 VPWR VGND sg13g2_decap_8
XFILLER_28_889 VPWR VGND sg13g2_decap_8
XFILLER_42_358 VPWR VGND sg13g2_decap_8
X_230_ net167 mac1.sum_lvl3_ff\[3\] _144_ VPWR VGND sg13g2_nor2_1
XFILLER_23_583 VPWR VGND sg13g2_decap_8
XFILLER_24_54 VPWR VGND sg13g2_decap_8
XFILLER_11_767 VPWR VGND sg13g2_decap_8
XFILLER_10_255 VPWR VGND sg13g2_decap_8
XFILLER_10_288 VPWR VGND sg13g2_decap_4
XFILLER_6_248 VPWR VGND sg13g2_decap_8
XFILLER_40_75 VPWR VGND sg13g2_decap_8
XFILLER_3_944 VPWR VGND sg13g2_decap_8
XFILLER_49_84 VPWR VGND sg13g2_decap_8
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_37_119 VPWR VGND sg13g2_fill_1
XFILLER_46_620 VPWR VGND sg13g2_decap_8
XFILLER_19_867 VPWR VGND sg13g2_decap_8
XFILLER_18_355 VPWR VGND sg13g2_decap_8
XFILLER_18_366 VPWR VGND sg13g2_fill_2
XFILLER_34_804 VPWR VGND sg13g2_decap_8
XFILLER_46_697 VPWR VGND sg13g2_decap_8
X_428_ net127 _122_ VPWR VGND sg13g2_buf_1
X_359_ _211_ _210_ _055_ VPWR VGND sg13g2_xor2_1
XFILLER_6_760 VPWR VGND sg13g2_decap_8
XFILLER_37_653 VPWR VGND sg13g2_decap_8
XFILLER_24_325 VPWR VGND sg13g2_decap_8
XFILLER_25_837 VPWR VGND sg13g2_decap_8
XFILLER_36_174 VPWR VGND sg13g2_decap_8
XFILLER_24_369 VPWR VGND sg13g2_decap_8
XFILLER_33_881 VPWR VGND sg13g2_decap_8
XFILLER_20_542 VPWR VGND sg13g2_decap_8
XFILLER_0_903 VPWR VGND sg13g2_decap_8
XFILLER_19_32 VPWR VGND sg13g2_decap_8
XFILLER_43_601 VPWR VGND sg13g2_decap_8
XFILLER_16_837 VPWR VGND sg13g2_decap_8
XFILLER_28_686 VPWR VGND sg13g2_decap_8
XFILLER_35_31 VPWR VGND sg13g2_fill_2
XFILLER_43_678 VPWR VGND sg13g2_decap_8
XFILLER_42_122 VPWR VGND sg13g2_decap_8
XFILLER_27_196 VPWR VGND sg13g2_decap_8
XFILLER_31_818 VPWR VGND sg13g2_decap_8
XFILLER_35_75 VPWR VGND sg13g2_decap_8
XFILLER_24_881 VPWR VGND sg13g2_decap_8
XFILLER_42_199 VPWR VGND sg13g2_decap_8
Xclkbuf_5_19__f_clk clknet_4_9_0_clk clknet_5_19__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_23_380 VPWR VGND sg13g2_decap_8
XFILLER_7_502 VPWR VGND sg13g2_decap_8
XFILLER_7_568 VPWR VGND sg13g2_decap_8
XFILLER_3_741 VPWR VGND sg13g2_decap_8
XFILLER_2_251 VPWR VGND sg13g2_decap_8
XFILLER_38_406 VPWR VGND sg13g2_decap_8
XFILLER_47_973 VPWR VGND sg13g2_decap_8
XFILLER_19_664 VPWR VGND sg13g2_decap_8
XFILLER_34_601 VPWR VGND sg13g2_decap_8
XFILLER_46_494 VPWR VGND sg13g2_decap_8
XFILLER_18_174 VPWR VGND sg13g2_decap_8
XFILLER_33_144 VPWR VGND sg13g2_decap_8
XFILLER_34_678 VPWR VGND sg13g2_decap_8
XFILLER_21_306 VPWR VGND sg13g2_decap_8
XFILLER_14_391 VPWR VGND sg13g2_decap_8
XFILLER_5_1018 VPWR VGND sg13g2_decap_8
XFILLER_44_409 VPWR VGND sg13g2_decap_8
XFILLER_25_634 VPWR VGND sg13g2_decap_8
XFILLER_24_166 VPWR VGND sg13g2_decap_8
XFILLER_40_659 VPWR VGND sg13g2_decap_8
XFILLER_21_862 VPWR VGND sg13g2_decap_8
XFILLER_21_11 VPWR VGND sg13g2_decap_8
XFILLER_4_527 VPWR VGND sg13g2_decap_8
XFILLER_0_700 VPWR VGND sg13g2_decap_8
XFILLER_0_777 VPWR VGND sg13g2_decap_8
XFILLER_48_748 VPWR VGND sg13g2_decap_8
XFILLER_16_634 VPWR VGND sg13g2_decap_8
XFILLER_29_995 VPWR VGND sg13g2_decap_8
XFILLER_44_976 VPWR VGND sg13g2_decap_8
XFILLER_15_133 VPWR VGND sg13g2_decap_8
XFILLER_43_475 VPWR VGND sg13g2_decap_8
XFILLER_31_615 VPWR VGND sg13g2_decap_8
XFILLER_8_811 VPWR VGND sg13g2_decap_8
XFILLER_12_851 VPWR VGND sg13g2_decap_8
XFILLER_7_35 VPWR VGND sg13g2_decap_8
XFILLER_8_888 VPWR VGND sg13g2_decap_8
XFILLER_7_376 VPWR VGND sg13g2_decap_8
XFILLER_23_4 VPWR VGND sg13g2_decap_8
XFILLER_38_258 VPWR VGND sg13g2_fill_2
XFILLER_47_770 VPWR VGND sg13g2_decap_8
XFILLER_19_483 VPWR VGND sg13g2_decap_8
XFILLER_35_921 VPWR VGND sg13g2_decap_8
XFILLER_35_998 VPWR VGND sg13g2_decap_8
XFILLER_22_648 VPWR VGND sg13g2_decap_8
XFILLER_16_11 VPWR VGND sg13g2_decap_4
XFILLER_26_921 VPWR VGND sg13g2_decap_8
XFILLER_25_486 VPWR VGND sg13g2_decap_8
XFILLER_26_998 VPWR VGND sg13g2_decap_8
XFILLER_13_648 VPWR VGND sg13g2_decap_8
XFILLER_40_412 VPWR VGND sg13g2_decap_8
XFILLER_40_423 VPWR VGND sg13g2_fill_2
XFILLER_40_445 VPWR VGND sg13g2_decap_8
XFILLER_41_946 VPWR VGND sg13g2_decap_8
XFILLER_9_619 VPWR VGND sg13g2_decap_8
XFILLER_12_158 VPWR VGND sg13g2_fill_2
XFILLER_32_87 VPWR VGND sg13g2_decap_8
XFILLER_5_836 VPWR VGND sg13g2_decap_8
XFILLER_10_1012 VPWR VGND sg13g2_decap_8
XFILLER_4_346 VPWR VGND sg13g2_decap_4
XFILLER_4_368 VPWR VGND sg13g2_decap_8
XFILLER_0_574 VPWR VGND sg13g2_decap_8
XFILLER_48_545 VPWR VGND sg13g2_decap_8
XFILLER_29_792 VPWR VGND sg13g2_decap_8
XFILLER_17_943 VPWR VGND sg13g2_decap_8
XFILLER_44_773 VPWR VGND sg13g2_decap_8
XFILLER_31_412 VPWR VGND sg13g2_decap_8
XFILLER_32_935 VPWR VGND sg13g2_decap_8
XFILLER_31_489 VPWR VGND sg13g2_decap_8
XFILLER_7_140 VPWR VGND sg13g2_decap_8
XFILLER_8_685 VPWR VGND sg13g2_decap_8
Xhold107 DP_3.matrix\[9\] VPWR VGND net157 sg13g2_dlygate4sd3_1
Xhold118 _143_ VPWR VGND net168 sg13g2_dlygate4sd3_1
Xhold129 mac2.products_ff\[51\] VPWR VGND net179 sg13g2_dlygate4sd3_1
XFILLER_39_567 VPWR VGND sg13g2_decap_8
XFILLER_27_729 VPWR VGND sg13g2_decap_8
XFILLER_19_291 VPWR VGND sg13g2_decap_8
XFILLER_41_209 VPWR VGND sg13g2_decap_8
XFILLER_22_423 VPWR VGND sg13g2_fill_2
XFILLER_35_795 VPWR VGND sg13g2_decap_8
XFILLER_23_968 VPWR VGND sg13g2_decap_8
XFILLER_2_817 VPWR VGND sg13g2_decap_8
XFILLER_1_327 VPWR VGND sg13g2_decap_8
XFILLER_18_718 VPWR VGND sg13g2_decap_8
XFILLER_40_1016 VPWR VGND sg13g2_decap_8
XFILLER_40_1027 VPWR VGND sg13g2_fill_2
XFILLER_17_228 VPWR VGND sg13g2_decap_8
X_530_ net83 VGND VPWR _070_ DP_1.matrix\[0\] clknet_5_28__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_548 VPWR VGND sg13g2_decap_8
XFILLER_27_76 VPWR VGND sg13g2_decap_8
X_461_ net75 VGND VPWR _055_ mac1.products_ff\[103\] clknet_5_20__leaf_clk sg13g2_dfrbpq_1
XFILLER_14_924 VPWR VGND sg13g2_decap_8
XFILLER_25_250 VPWR VGND sg13g2_fill_2
X_392_ net133 _086_ VPWR VGND sg13g2_buf_1
XFILLER_25_294 VPWR VGND sg13g2_fill_2
XFILLER_26_795 VPWR VGND sg13g2_decap_8
XFILLER_41_743 VPWR VGND sg13g2_decap_8
XFILLER_43_42 VPWR VGND sg13g2_decap_8
XFILLER_9_416 VPWR VGND sg13g2_decap_8
XFILLER_13_478 VPWR VGND sg13g2_decap_8
XFILLER_5_633 VPWR VGND sg13g2_decap_8
XFILLER_4_165 VPWR VGND sg13g2_decap_8
XFILLER_4_25 VPWR VGND sg13g2_decap_8
XFILLER_49_821 VPWR VGND sg13g2_decap_8
XFILLER_0_371 VPWR VGND sg13g2_decap_8
XFILLER_1_894 VPWR VGND sg13g2_decap_8
XFILLER_49_898 VPWR VGND sg13g2_decap_8
XFILLER_48_386 VPWR VGND sg13g2_decap_8
XFILLER_17_740 VPWR VGND sg13g2_decap_8
XFILLER_36_548 VPWR VGND sg13g2_decap_8
XFILLER_44_570 VPWR VGND sg13g2_decap_8
XFILLER_16_283 VPWR VGND sg13g2_decap_4
XFILLER_32_732 VPWR VGND sg13g2_decap_8
XFILLER_31_231 VPWR VGND sg13g2_decap_8
XFILLER_20_927 VPWR VGND sg13g2_decap_8
XFILLER_9_983 VPWR VGND sg13g2_decap_8
XFILLER_39_320 VPWR VGND sg13g2_decap_8
XFILLER_27_526 VPWR VGND sg13g2_decap_8
XFILLER_14_209 VPWR VGND sg13g2_decap_8
XFILLER_35_592 VPWR VGND sg13g2_decap_8
XFILLER_23_765 VPWR VGND sg13g2_decap_8
XFILLER_10_404 VPWR VGND sg13g2_fill_1
XFILLER_11_949 VPWR VGND sg13g2_decap_8
Xfanout79 net81 net79 VPWR VGND sg13g2_buf_8
Xfanout68 net69 net68 VPWR VGND sg13g2_buf_8
XFILLER_10_459 VPWR VGND sg13g2_decap_8
XFILLER_13_67 VPWR VGND sg13g2_decap_8
XFILLER_2_614 VPWR VGND sg13g2_decap_8
XFILLER_1_102 VPWR VGND sg13g2_decap_8
XFILLER_49_128 VPWR VGND sg13g2_decap_8
XFILLER_46_802 VPWR VGND sg13g2_decap_8
XFILLER_38_42 VPWR VGND sg13g2_decap_4
XFILLER_18_526 VPWR VGND sg13g2_fill_1
XFILLER_38_97 VPWR VGND sg13g2_decap_8
XFILLER_45_334 VPWR VGND sg13g2_decap_4
XFILLER_46_879 VPWR VGND sg13g2_decap_8
X_513_ net81 VGND VPWR net124 mac2.sum_lvl1_ff\[24\] clknet_5_26__leaf_clk sg13g2_dfrbpq_1
X_444_ net121 _138_ VPWR VGND sg13g2_buf_1
XFILLER_14_721 VPWR VGND sg13g2_decap_8
XFILLER_26_592 VPWR VGND sg13g2_decap_8
XFILLER_13_231 VPWR VGND sg13g2_fill_2
XFILLER_41_540 VPWR VGND sg13g2_decap_8
XFILLER_9_202 VPWR VGND sg13g2_decap_8
XFILLER_14_798 VPWR VGND sg13g2_decap_8
X_375_ _221_ _220_ _065_ VPWR VGND sg13g2_xor2_1
XFILLER_6_942 VPWR VGND sg13g2_decap_8
XFILLER_1_691 VPWR VGND sg13g2_decap_8
XFILLER_37_835 VPWR VGND sg13g2_decap_8
XFILLER_49_695 VPWR VGND sg13g2_decap_8
XFILLER_36_312 VPWR VGND sg13g2_decap_8
XFILLER_36_389 VPWR VGND sg13g2_decap_8
XFILLER_20_724 VPWR VGND sg13g2_decap_8
XFILLER_9_780 VPWR VGND sg13g2_decap_8
XFILLER_30_1004 VPWR VGND sg13g2_decap_8
XFILLER_39_150 VPWR VGND sg13g2_decap_8
XFILLER_28_868 VPWR VGND sg13g2_decap_8
XFILLER_27_378 VPWR VGND sg13g2_decap_4
XFILLER_42_337 VPWR VGND sg13g2_decap_8
XFILLER_15_529 VPWR VGND sg13g2_decap_8
XFILLER_24_11 VPWR VGND sg13g2_decap_8
XFILLER_23_562 VPWR VGND sg13g2_decap_8
XFILLER_10_234 VPWR VGND sg13g2_decap_8
XFILLER_11_746 VPWR VGND sg13g2_decap_8
XFILLER_10_267 VPWR VGND sg13g2_decap_8
XFILLER_6_227 VPWR VGND sg13g2_decap_8
XFILLER_40_54 VPWR VGND sg13g2_decap_8
XFILLER_3_923 VPWR VGND sg13g2_decap_8
XFILLER_2_444 VPWR VGND sg13g2_decap_8
XFILLER_49_63 VPWR VGND sg13g2_decap_8
XFILLER_18_334 VPWR VGND sg13g2_decap_8
XFILLER_19_846 VPWR VGND sg13g2_decap_8
XFILLER_46_676 VPWR VGND sg13g2_decap_8
XFILLER_45_153 VPWR VGND sg13g2_decap_8
XFILLER_27_890 VPWR VGND sg13g2_decap_8
X_427_ net86 _121_ VPWR VGND sg13g2_buf_1
X_358_ _211_ net151 net90 VPWR VGND sg13g2_nand2_1
XFILLER_14_595 VPWR VGND sg13g2_decap_8
X_289_ _170_ net173 net161 VPWR VGND sg13g2_nand2_1
XFILLER_49_492 VPWR VGND sg13g2_decap_8
XFILLER_37_632 VPWR VGND sg13g2_decap_8
XFILLER_25_816 VPWR VGND sg13g2_decap_8
XFILLER_36_153 VPWR VGND sg13g2_decap_8
XFILLER_24_304 VPWR VGND sg13g2_decap_8
XFILLER_33_860 VPWR VGND sg13g2_decap_8
XFILLER_20_521 VPWR VGND sg13g2_decap_8
XFILLER_20_598 VPWR VGND sg13g2_decap_8
XFILLER_10_13 VPWR VGND sg13g2_fill_1
XFILLER_0_959 VPWR VGND sg13g2_decap_8
XFILLER_19_11 VPWR VGND sg13g2_decap_8
XFILLER_19_109 VPWR VGND sg13g2_decap_8
XFILLER_19_88 VPWR VGND sg13g2_decap_8
XFILLER_16_816 VPWR VGND sg13g2_decap_8
XFILLER_28_665 VPWR VGND sg13g2_decap_8
XFILLER_42_101 VPWR VGND sg13g2_decap_8
XFILLER_15_315 VPWR VGND sg13g2_decap_8
XFILLER_15_326 VPWR VGND sg13g2_fill_1
XFILLER_27_175 VPWR VGND sg13g2_decap_8
XFILLER_35_21 VPWR VGND sg13g2_decap_4
XFILLER_43_657 VPWR VGND sg13g2_decap_8
XFILLER_42_178 VPWR VGND sg13g2_fill_2
XFILLER_24_860 VPWR VGND sg13g2_decap_8
XFILLER_11_543 VPWR VGND sg13g2_fill_1
XFILLER_3_720 VPWR VGND sg13g2_decap_8
XFILLER_2_230 VPWR VGND sg13g2_decap_8
XFILLER_3_797 VPWR VGND sg13g2_decap_8
XFILLER_47_952 VPWR VGND sg13g2_decap_8
XFILLER_19_643 VPWR VGND sg13g2_decap_8
XFILLER_20_1025 VPWR VGND sg13g2_decap_4
XFILLER_46_473 VPWR VGND sg13g2_decap_8
XFILLER_33_123 VPWR VGND sg13g2_decap_8
XFILLER_34_657 VPWR VGND sg13g2_decap_8
XFILLER_14_370 VPWR VGND sg13g2_decap_8
XFILLER_30_885 VPWR VGND sg13g2_decap_8
XFILLER_44_0 VPWR VGND sg13g2_decap_8
Xclkbuf_5_25__f_clk clknet_4_12_0_clk clknet_5_25__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_25_613 VPWR VGND sg13g2_decap_8
XFILLER_38_985 VPWR VGND sg13g2_decap_8
XFILLER_24_145 VPWR VGND sg13g2_decap_8
XFILLER_36_1010 VPWR VGND sg13g2_decap_8
XFILLER_21_841 VPWR VGND sg13g2_decap_8
XFILLER_40_638 VPWR VGND sg13g2_decap_8
XFILLER_20_340 VPWR VGND sg13g2_decap_8
XFILLER_4_506 VPWR VGND sg13g2_decap_8
XFILLER_20_395 VPWR VGND sg13g2_decap_8
XFILLER_43_1014 VPWR VGND sg13g2_decap_8
XFILLER_0_756 VPWR VGND sg13g2_decap_8
XFILLER_48_727 VPWR VGND sg13g2_decap_8
XFILLER_47_248 VPWR VGND sg13g2_decap_8
XFILLER_46_42 VPWR VGND sg13g2_decap_8
XFILLER_29_974 VPWR VGND sg13g2_decap_8
XFILLER_16_613 VPWR VGND sg13g2_decap_8
XFILLER_44_955 VPWR VGND sg13g2_decap_8
XFILLER_43_454 VPWR VGND sg13g2_decap_8
XFILLER_12_830 VPWR VGND sg13g2_decap_8
XFILLER_30_115 VPWR VGND sg13g2_decap_8
XFILLER_7_14 VPWR VGND sg13g2_decap_8
XFILLER_8_867 VPWR VGND sg13g2_decap_8
XFILLER_7_355 VPWR VGND sg13g2_decap_8
XFILLER_11_395 VPWR VGND sg13g2_fill_2
XFILLER_7_399 VPWR VGND sg13g2_fill_2
XFILLER_3_594 VPWR VGND sg13g2_decap_8
XFILLER_16_4 VPWR VGND sg13g2_decap_8
XFILLER_38_237 VPWR VGND sg13g2_decap_8
XFILLER_39_749 VPWR VGND sg13g2_decap_8
XFILLER_35_900 VPWR VGND sg13g2_decap_8
XFILLER_19_462 VPWR VGND sg13g2_decap_8
XFILLER_46_270 VPWR VGND sg13g2_decap_8
XFILLER_35_977 VPWR VGND sg13g2_decap_8
XFILLER_22_627 VPWR VGND sg13g2_decap_8
XFILLER_30_682 VPWR VGND sg13g2_decap_8
XFILLER_1_509 VPWR VGND sg13g2_decap_8
XFILLER_27_1009 VPWR VGND sg13g2_decap_8
XFILLER_26_900 VPWR VGND sg13g2_decap_8
XFILLER_38_782 VPWR VGND sg13g2_decap_8
XFILLER_16_56 VPWR VGND sg13g2_decap_8
XFILLER_25_465 VPWR VGND sg13g2_decap_8
XFILLER_26_977 VPWR VGND sg13g2_decap_8
XFILLER_41_925 VPWR VGND sg13g2_decap_8
XFILLER_12_104 VPWR VGND sg13g2_decap_8
XFILLER_13_627 VPWR VGND sg13g2_decap_8
XFILLER_12_137 VPWR VGND sg13g2_decap_8
XFILLER_5_815 VPWR VGND sg13g2_decap_8
XFILLER_32_66 VPWR VGND sg13g2_decap_8
XFILLER_4_325 VPWR VGND sg13g2_decap_8
XFILLER_0_553 VPWR VGND sg13g2_decap_8
XFILLER_48_524 VPWR VGND sg13g2_decap_8
XFILLER_17_922 VPWR VGND sg13g2_decap_8
XFILLER_29_771 VPWR VGND sg13g2_decap_8
XFILLER_28_281 VPWR VGND sg13g2_decap_4
XFILLER_44_752 VPWR VGND sg13g2_decap_8
XFILLER_17_999 VPWR VGND sg13g2_decap_8
XFILLER_32_914 VPWR VGND sg13g2_decap_8
XFILLER_43_295 VPWR VGND sg13g2_decap_8
XFILLER_31_468 VPWR VGND sg13g2_decap_8
XFILLER_8_664 VPWR VGND sg13g2_decap_8
Xhold108 DP_4.matrix\[45\] VPWR VGND net158 sg13g2_dlygate4sd3_1
Xhold119 _016_ VPWR VGND net169 sg13g2_dlygate4sd3_1
XFILLER_7_196 VPWR VGND sg13g2_decap_8
XFILLER_4_892 VPWR VGND sg13g2_decap_8
XFILLER_27_708 VPWR VGND sg13g2_decap_8
XFILLER_39_546 VPWR VGND sg13g2_decap_8
XFILLER_19_270 VPWR VGND sg13g2_decap_8
XFILLER_35_774 VPWR VGND sg13g2_decap_8
XFILLER_22_402 VPWR VGND sg13g2_decap_8
XFILLER_23_947 VPWR VGND sg13g2_decap_8
XFILLER_34_273 VPWR VGND sg13g2_decap_8
XFILLER_22_468 VPWR VGND sg13g2_decap_8
XFILLER_1_306 VPWR VGND sg13g2_decap_8
XFILLER_45_527 VPWR VGND sg13g2_decap_8
XFILLER_17_207 VPWR VGND sg13g2_decap_8
XFILLER_27_55 VPWR VGND sg13g2_decap_8
X_460_ net73 VGND VPWR _054_ mac1.products_ff\[102\] clknet_5_17__leaf_clk sg13g2_dfrbpq_1
XFILLER_14_903 VPWR VGND sg13g2_decap_8
XFILLER_26_774 VPWR VGND sg13g2_decap_8
XFILLER_43_21 VPWR VGND sg13g2_decap_8
X_391_ net92 _085_ VPWR VGND sg13g2_buf_1
XFILLER_41_722 VPWR VGND sg13g2_decap_8
XFILLER_9_406 VPWR VGND sg13g2_fill_2
XFILLER_13_446 VPWR VGND sg13g2_fill_1
XFILLER_40_221 VPWR VGND sg13g2_decap_4
XFILLER_40_254 VPWR VGND sg13g2_fill_2
XFILLER_41_799 VPWR VGND sg13g2_decap_8
XFILLER_22_991 VPWR VGND sg13g2_decap_8
XFILLER_40_298 VPWR VGND sg13g2_decap_8
XFILLER_5_612 VPWR VGND sg13g2_decap_8
XFILLER_5_689 VPWR VGND sg13g2_decap_8
XFILLER_4_144 VPWR VGND sg13g2_decap_8
XFILLER_49_800 VPWR VGND sg13g2_decap_8
XFILLER_0_350 VPWR VGND sg13g2_decap_8
XFILLER_1_873 VPWR VGND sg13g2_decap_8
XFILLER_49_877 VPWR VGND sg13g2_decap_8
XFILLER_48_365 VPWR VGND sg13g2_decap_8
XFILLER_36_527 VPWR VGND sg13g2_decap_8
X_589_ net69 VGND VPWR _129_ DP_4.matrix\[19\] clknet_5_10__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_796 VPWR VGND sg13g2_decap_8
XFILLER_31_210 VPWR VGND sg13g2_decap_8
XFILLER_32_711 VPWR VGND sg13g2_decap_8
XFILLER_20_906 VPWR VGND sg13g2_decap_8
XFILLER_32_788 VPWR VGND sg13g2_decap_8
XFILLER_9_962 VPWR VGND sg13g2_decap_8
XFILLER_13_991 VPWR VGND sg13g2_decap_8
XFILLER_31_287 VPWR VGND sg13g2_decap_8
XFILLER_39_365 VPWR VGND sg13g2_fill_2
XFILLER_42_519 VPWR VGND sg13g2_decap_8
XFILLER_35_571 VPWR VGND sg13g2_decap_8
XFILLER_23_744 VPWR VGND sg13g2_decap_8
XFILLER_11_928 VPWR VGND sg13g2_decap_8
Xfanout69 net72 net69 VPWR VGND sg13g2_buf_8
XFILLER_10_438 VPWR VGND sg13g2_decap_8
XFILLER_13_46 VPWR VGND sg13g2_decap_8
XFILLER_1_158 VPWR VGND sg13g2_decap_8
XFILLER_1_169 VPWR VGND sg13g2_fill_2
XFILLER_38_21 VPWR VGND sg13g2_decap_8
XFILLER_18_505 VPWR VGND sg13g2_decap_8
XFILLER_38_76 VPWR VGND sg13g2_decap_8
XFILLER_46_858 VPWR VGND sg13g2_decap_8
XFILLER_45_313 VPWR VGND sg13g2_decap_8
XFILLER_18_549 VPWR VGND sg13g2_decap_8
X_512_ net80 VGND VPWR net182 mac2.sum_lvl1_ff\[17\] clknet_5_15__leaf_clk sg13g2_dfrbpq_1
XFILLER_14_700 VPWR VGND sg13g2_decap_8
XFILLER_26_571 VPWR VGND sg13g2_decap_8
X_443_ net37 _137_ VPWR VGND sg13g2_buf_1
XFILLER_13_210 VPWR VGND sg13g2_decap_8
XFILLER_14_777 VPWR VGND sg13g2_decap_8
X_374_ _221_ net132 net101 VPWR VGND sg13g2_nand2_1
XFILLER_41_596 VPWR VGND sg13g2_decap_8
XFILLER_6_921 VPWR VGND sg13g2_decap_8
XFILLER_5_420 VPWR VGND sg13g2_fill_2
XFILLER_6_998 VPWR VGND sg13g2_decap_8
XFILLER_5_464 VPWR VGND sg13g2_fill_1
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_1_670 VPWR VGND sg13g2_decap_8
Xclkbuf_5_6__f_clk clknet_4_3_0_clk clknet_5_6__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_49_674 VPWR VGND sg13g2_decap_8
XFILLER_48_162 VPWR VGND sg13g2_decap_8
XFILLER_37_814 VPWR VGND sg13g2_decap_8
XFILLER_48_184 VPWR VGND sg13g2_decap_4
XFILLER_36_368 VPWR VGND sg13g2_decap_8
XFILLER_45_891 VPWR VGND sg13g2_decap_8
XFILLER_20_703 VPWR VGND sg13g2_decap_8
XFILLER_32_585 VPWR VGND sg13g2_decap_8
XFILLER_8_280 VPWR VGND sg13g2_decap_8
XFILLER_8_1028 VPWR VGND sg13g2_fill_1
XFILLER_28_847 VPWR VGND sg13g2_decap_8
XFILLER_15_508 VPWR VGND sg13g2_decap_8
XFILLER_27_357 VPWR VGND sg13g2_decap_8
XFILLER_43_839 VPWR VGND sg13g2_decap_8
XFILLER_42_316 VPWR VGND sg13g2_decap_8
XFILLER_36_891 VPWR VGND sg13g2_decap_8
XFILLER_11_725 VPWR VGND sg13g2_decap_8
XFILLER_24_89 VPWR VGND sg13g2_decap_8
XFILLER_7_729 VPWR VGND sg13g2_decap_8
XFILLER_6_206 VPWR VGND sg13g2_decap_8
XFILLER_3_902 VPWR VGND sg13g2_decap_8
XFILLER_46_1012 VPWR VGND sg13g2_decap_8
XFILLER_3_979 VPWR VGND sg13g2_decap_8
XFILLER_49_42 VPWR VGND sg13g2_decap_8
XFILLER_19_825 VPWR VGND sg13g2_decap_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_18_313 VPWR VGND sg13g2_decap_8
XFILLER_46_655 VPWR VGND sg13g2_decap_8
XFILLER_45_132 VPWR VGND sg13g2_decap_8
XFILLER_45_187 VPWR VGND sg13g2_decap_8
XFILLER_34_839 VPWR VGND sg13g2_decap_8
XFILLER_33_349 VPWR VGND sg13g2_decap_4
X_426_ net141 _120_ VPWR VGND sg13g2_buf_1
XFILLER_42_883 VPWR VGND sg13g2_decap_8
XFILLER_14_574 VPWR VGND sg13g2_decap_8
X_357_ _210_ net120 net54 VPWR VGND sg13g2_nand2_1
X_288_ net145 mac1.sum_lvl1_ff\[8\] _010_ VPWR VGND sg13g2_xor2_1
XFILLER_6_795 VPWR VGND sg13g2_decap_8
XFILLER_49_471 VPWR VGND sg13g2_decap_8
XFILLER_37_611 VPWR VGND sg13g2_decap_8
XFILLER_36_132 VPWR VGND sg13g2_decap_8
XFILLER_37_688 VPWR VGND sg13g2_decap_8
XFILLER_20_500 VPWR VGND sg13g2_decap_8
XFILLER_32_382 VPWR VGND sg13g2_decap_8
XFILLER_20_577 VPWR VGND sg13g2_decap_8
XFILLER_0_938 VPWR VGND sg13g2_decap_8
XFILLER_48_909 VPWR VGND sg13g2_decap_8
XFILLER_19_67 VPWR VGND sg13g2_decap_8
XFILLER_27_132 VPWR VGND sg13g2_decap_8
XFILLER_28_644 VPWR VGND sg13g2_decap_8
XFILLER_35_33 VPWR VGND sg13g2_fill_1
XFILLER_43_636 VPWR VGND sg13g2_decap_8
XFILLER_11_522 VPWR VGND sg13g2_decap_4
XFILLER_7_537 VPWR VGND sg13g2_decap_8
XFILLER_11_599 VPWR VGND sg13g2_decap_8
XFILLER_3_776 VPWR VGND sg13g2_decap_8
XFILLER_2_286 VPWR VGND sg13g2_decap_8
XFILLER_47_931 VPWR VGND sg13g2_decap_8
XFILLER_19_622 VPWR VGND sg13g2_decap_8
XFILLER_20_1004 VPWR VGND sg13g2_decap_8
XFILLER_46_452 VPWR VGND sg13g2_decap_8
XFILLER_18_154 VPWR VGND sg13g2_decap_8
XFILLER_19_699 VPWR VGND sg13g2_decap_8
XFILLER_33_102 VPWR VGND sg13g2_decap_8
XFILLER_22_809 VPWR VGND sg13g2_decap_8
XFILLER_34_636 VPWR VGND sg13g2_decap_8
XFILLER_33_179 VPWR VGND sg13g2_decap_8
XFILLER_42_680 VPWR VGND sg13g2_decap_8
X_409_ net40 _103_ VPWR VGND sg13g2_buf_1
XFILLER_15_883 VPWR VGND sg13g2_decap_8
XFILLER_30_864 VPWR VGND sg13g2_decap_8
XFILLER_6_592 VPWR VGND sg13g2_decap_8
XFILLER_37_0 VPWR VGND sg13g2_decap_8
XFILLER_38_964 VPWR VGND sg13g2_decap_8
XFILLER_37_474 VPWR VGND sg13g2_decap_8
XFILLER_37_485 VPWR VGND sg13g2_decap_8
XFILLER_24_124 VPWR VGND sg13g2_decap_8
XFILLER_12_308 VPWR VGND sg13g2_decap_8
XFILLER_13_809 VPWR VGND sg13g2_decap_8
XFILLER_25_669 VPWR VGND sg13g2_decap_8
XFILLER_40_617 VPWR VGND sg13g2_decap_8
XFILLER_21_820 VPWR VGND sg13g2_decap_8
XFILLER_20_374 VPWR VGND sg13g2_decap_8
XFILLER_21_897 VPWR VGND sg13g2_decap_8
XFILLER_21_46 VPWR VGND sg13g2_fill_2
XFILLER_0_735 VPWR VGND sg13g2_decap_8
XFILLER_48_706 VPWR VGND sg13g2_decap_8
XFILLER_47_216 VPWR VGND sg13g2_decap_4
XFILLER_46_21 VPWR VGND sg13g2_decap_8
XFILLER_29_953 VPWR VGND sg13g2_decap_8
XFILLER_44_934 VPWR VGND sg13g2_decap_8
XFILLER_43_400 VPWR VGND sg13g2_decap_8
XFILLER_46_87 VPWR VGND sg13g2_decap_8
XFILLER_43_411 VPWR VGND sg13g2_fill_2
XFILLER_15_168 VPWR VGND sg13g2_decap_8
XFILLER_16_669 VPWR VGND sg13g2_decap_8
XFILLER_8_846 VPWR VGND sg13g2_decap_8
XFILLER_11_374 VPWR VGND sg13g2_decap_8
XFILLER_12_886 VPWR VGND sg13g2_decap_8
XFILLER_7_334 VPWR VGND sg13g2_decap_8
Xclkbuf_5_31__f_clk clknet_4_15_0_clk clknet_5_31__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_30_7 VPWR VGND sg13g2_decap_8
XFILLER_38_216 VPWR VGND sg13g2_decap_8
XFILLER_39_728 VPWR VGND sg13g2_decap_8
XFILLER_19_441 VPWR VGND sg13g2_decap_8
XFILLER_35_956 VPWR VGND sg13g2_decap_8
XFILLER_22_606 VPWR VGND sg13g2_decap_8
XFILLER_34_444 VPWR VGND sg13g2_fill_2
XFILLER_15_680 VPWR VGND sg13g2_decap_8
XFILLER_30_661 VPWR VGND sg13g2_decap_8
XFILLER_7_890 VPWR VGND sg13g2_decap_8
XFILLER_45_709 VPWR VGND sg13g2_decap_8
XFILLER_29_249 VPWR VGND sg13g2_fill_2
XFILLER_38_761 VPWR VGND sg13g2_decap_8
XFILLER_25_411 VPWR VGND sg13g2_fill_2
XFILLER_26_956 VPWR VGND sg13g2_decap_8
XFILLER_13_606 VPWR VGND sg13g2_decap_8
XFILLER_25_444 VPWR VGND sg13g2_decap_8
XFILLER_41_904 VPWR VGND sg13g2_decap_8
XFILLER_32_45 VPWR VGND sg13g2_decap_8
XFILLER_20_193 VPWR VGND sg13g2_decap_8
XFILLER_21_694 VPWR VGND sg13g2_decap_8
XFILLER_0_532 VPWR VGND sg13g2_decap_8
XFILLER_48_503 VPWR VGND sg13g2_decap_8
XFILLER_29_750 VPWR VGND sg13g2_decap_8
XFILLER_36_709 VPWR VGND sg13g2_decap_8
XFILLER_17_901 VPWR VGND sg13g2_decap_8
XFILLER_44_731 VPWR VGND sg13g2_decap_8
XFILLER_28_260 VPWR VGND sg13g2_decap_8
XFILLER_43_252 VPWR VGND sg13g2_decap_4
XFILLER_16_466 VPWR VGND sg13g2_decap_4
XFILLER_17_978 VPWR VGND sg13g2_decap_8
XFILLER_16_499 VPWR VGND sg13g2_decap_8
XFILLER_31_447 VPWR VGND sg13g2_decap_8
XFILLER_40_981 VPWR VGND sg13g2_decap_8
XFILLER_8_643 VPWR VGND sg13g2_decap_8
XFILLER_12_683 VPWR VGND sg13g2_decap_8
XFILLER_7_175 VPWR VGND sg13g2_decap_8
Xhold109 DP_1.matrix\[0\] VPWR VGND net159 sg13g2_dlygate4sd3_1
XFILLER_4_871 VPWR VGND sg13g2_decap_8
XFILLER_26_219 VPWR VGND sg13g2_decap_8
XFILLER_34_252 VPWR VGND sg13g2_decap_8
XFILLER_35_753 VPWR VGND sg13g2_decap_8
XFILLER_23_926 VPWR VGND sg13g2_decap_8
XFILLER_22_447 VPWR VGND sg13g2_decap_8
XFILLER_33_1014 VPWR VGND sg13g2_decap_8
XFILLER_45_506 VPWR VGND sg13g2_decap_8
XFILLER_26_753 VPWR VGND sg13g2_decap_8
XFILLER_41_701 VPWR VGND sg13g2_decap_8
X_390_ net126 _084_ VPWR VGND sg13g2_buf_1
XFILLER_13_403 VPWR VGND sg13g2_decap_4
XFILLER_13_425 VPWR VGND sg13g2_decap_8
XFILLER_25_252 VPWR VGND sg13g2_fill_1
XFILLER_14_959 VPWR VGND sg13g2_decap_8
XFILLER_25_296 VPWR VGND sg13g2_fill_1
XFILLER_43_99 VPWR VGND sg13g2_decap_8
XFILLER_22_970 VPWR VGND sg13g2_decap_8
XFILLER_40_277 VPWR VGND sg13g2_decap_8
XFILLER_41_778 VPWR VGND sg13g2_decap_8
XFILLER_49_1010 VPWR VGND sg13g2_decap_8
XFILLER_5_668 VPWR VGND sg13g2_decap_8
XFILLER_1_852 VPWR VGND sg13g2_decap_8
XFILLER_49_856 VPWR VGND sg13g2_decap_8
XFILLER_48_344 VPWR VGND sg13g2_decap_8
XFILLER_36_506 VPWR VGND sg13g2_decap_8
X_588_ net70 VGND VPWR _128_ DP_4.matrix\[18\] clknet_5_11__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_775 VPWR VGND sg13g2_decap_8
XFILLER_32_767 VPWR VGND sg13g2_decap_8
XFILLER_13_970 VPWR VGND sg13g2_decap_8
XFILLER_31_266 VPWR VGND sg13g2_decap_8
XFILLER_9_941 VPWR VGND sg13g2_decap_8
XFILLER_12_480 VPWR VGND sg13g2_fill_2
XFILLER_8_495 VPWR VGND sg13g2_fill_2
XFILLER_8_484 VPWR VGND sg13g2_decap_8
XFILLER_39_311 VPWR VGND sg13g2_fill_1
XFILLER_39_377 VPWR VGND sg13g2_fill_2
XFILLER_35_550 VPWR VGND sg13g2_decap_8
XFILLER_23_723 VPWR VGND sg13g2_decap_8
XFILLER_11_907 VPWR VGND sg13g2_decap_8
XFILLER_13_25 VPWR VGND sg13g2_decap_8
XFILLER_22_288 VPWR VGND sg13g2_decap_8
XFILLER_1_137 VPWR VGND sg13g2_decap_8
XFILLER_2_649 VPWR VGND sg13g2_decap_8
XFILLER_38_55 VPWR VGND sg13g2_decap_8
XFILLER_46_837 VPWR VGND sg13g2_decap_8
XFILLER_26_550 VPWR VGND sg13g2_decap_8
X_511_ net80 VGND VPWR net104 mac2.sum_lvl1_ff\[16\] clknet_5_13__leaf_clk sg13g2_dfrbpq_1
X_442_ net143 _136_ VPWR VGND sg13g2_buf_1
XFILLER_14_756 VPWR VGND sg13g2_decap_8
X_373_ _220_ net119 net88 VPWR VGND sg13g2_nand2_1
XFILLER_41_575 VPWR VGND sg13g2_decap_8
XFILLER_9_237 VPWR VGND sg13g2_decap_8
XFILLER_13_288 VPWR VGND sg13g2_decap_8
XFILLER_6_900 VPWR VGND sg13g2_decap_8
XFILLER_10_984 VPWR VGND sg13g2_decap_8
XFILLER_6_977 VPWR VGND sg13g2_decap_8
XFILLER_49_653 VPWR VGND sg13g2_decap_8
XFILLER_48_141 VPWR VGND sg13g2_decap_8
XFILLER_23_1024 VPWR VGND sg13g2_decap_4
XFILLER_36_347 VPWR VGND sg13g2_decap_8
XFILLER_45_870 VPWR VGND sg13g2_decap_8
XFILLER_32_564 VPWR VGND sg13g2_decap_8
XFILLER_20_759 VPWR VGND sg13g2_decap_8
XFILLER_5_81 VPWR VGND sg13g2_decap_8
XFILLER_8_1007 VPWR VGND sg13g2_decap_8
XFILLER_27_303 VPWR VGND sg13g2_decap_4
XFILLER_28_826 VPWR VGND sg13g2_decap_8
XFILLER_43_818 VPWR VGND sg13g2_decap_8
XFILLER_27_336 VPWR VGND sg13g2_decap_8
XFILLER_36_870 VPWR VGND sg13g2_decap_8
XFILLER_11_704 VPWR VGND sg13g2_decap_8
XFILLER_10_203 VPWR VGND sg13g2_decap_8
XFILLER_23_597 VPWR VGND sg13g2_decap_8
XFILLER_24_68 VPWR VGND sg13g2_decap_8
XFILLER_7_708 VPWR VGND sg13g2_decap_8
XFILLER_40_89 VPWR VGND sg13g2_fill_1
XFILLER_49_21 VPWR VGND sg13g2_decap_8
XFILLER_6_4 VPWR VGND sg13g2_decap_8
XFILLER_3_958 VPWR VGND sg13g2_decap_8
XFILLER_2_479 VPWR VGND sg13g2_decap_4
XFILLER_49_98 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_19_804 VPWR VGND sg13g2_decap_8
XFILLER_46_634 VPWR VGND sg13g2_decap_8
XFILLER_45_111 VPWR VGND sg13g2_decap_8
XFILLER_34_818 VPWR VGND sg13g2_decap_8
XFILLER_26_380 VPWR VGND sg13g2_decap_8
XFILLER_42_862 VPWR VGND sg13g2_decap_8
XFILLER_14_553 VPWR VGND sg13g2_decap_8
X_425_ net89 _119_ VPWR VGND sg13g2_buf_1
X_356_ _209_ _208_ _053_ VPWR VGND sg13g2_xor2_1
XFILLER_14_90 VPWR VGND sg13g2_decap_8
XFILLER_10_781 VPWR VGND sg13g2_decap_8
X_287_ _011_ _168_ _169_ VPWR VGND sg13g2_xnor2_1
XFILLER_6_774 VPWR VGND sg13g2_decap_8
XFILLER_49_450 VPWR VGND sg13g2_decap_8
XFILLER_36_100 VPWR VGND sg13g2_decap_8
XFILLER_37_667 VPWR VGND sg13g2_decap_8
XFILLER_24_339 VPWR VGND sg13g2_decap_8
XFILLER_36_188 VPWR VGND sg13g2_decap_8
XFILLER_32_361 VPWR VGND sg13g2_decap_8
XFILLER_33_895 VPWR VGND sg13g2_decap_8
XFILLER_20_556 VPWR VGND sg13g2_decap_8
XFILLER_0_917 VPWR VGND sg13g2_decap_8
XFILLER_19_46 VPWR VGND sg13g2_decap_8
XFILLER_28_623 VPWR VGND sg13g2_decap_8
XFILLER_27_111 VPWR VGND sg13g2_decap_8
XFILLER_43_615 VPWR VGND sg13g2_decap_8
XFILLER_42_136 VPWR VGND sg13g2_decap_8
XFILLER_30_309 VPWR VGND sg13g2_decap_8
XFILLER_11_501 VPWR VGND sg13g2_decap_8
XFILLER_24_895 VPWR VGND sg13g2_decap_8
XFILLER_11_556 VPWR VGND sg13g2_decap_8
XFILLER_23_394 VPWR VGND sg13g2_decap_8
XFILLER_7_516 VPWR VGND sg13g2_decap_8
XFILLER_13_1012 VPWR VGND sg13g2_decap_8
XFILLER_3_755 VPWR VGND sg13g2_decap_8
XFILLER_2_265 VPWR VGND sg13g2_decap_8
XFILLER_47_910 VPWR VGND sg13g2_decap_8
XFILLER_19_601 VPWR VGND sg13g2_decap_8
XFILLER_46_431 VPWR VGND sg13g2_decap_8
XFILLER_18_133 VPWR VGND sg13g2_decap_8
XFILLER_47_987 VPWR VGND sg13g2_decap_8
XFILLER_19_678 VPWR VGND sg13g2_decap_8
XFILLER_34_615 VPWR VGND sg13g2_decap_8
XFILLER_18_188 VPWR VGND sg13g2_decap_8
XFILLER_15_862 VPWR VGND sg13g2_decap_8
XFILLER_33_158 VPWR VGND sg13g2_decap_8
X_408_ net135 _102_ VPWR VGND sg13g2_buf_1
XFILLER_30_843 VPWR VGND sg13g2_decap_8
X_339_ _198_ net142 net46 VPWR VGND sg13g2_nand2_1
XFILLER_29_409 VPWR VGND sg13g2_decap_8
XFILLER_2_60 VPWR VGND sg13g2_decap_8
XFILLER_38_943 VPWR VGND sg13g2_decap_8
XFILLER_37_453 VPWR VGND sg13g2_decap_8
XFILLER_24_103 VPWR VGND sg13g2_decap_8
XFILLER_25_648 VPWR VGND sg13g2_decap_8
XFILLER_33_692 VPWR VGND sg13g2_decap_8
XFILLER_21_876 VPWR VGND sg13g2_decap_8
XFILLER_21_25 VPWR VGND sg13g2_decap_8
XFILLER_0_714 VPWR VGND sg13g2_decap_8
XFILLER_29_932 VPWR VGND sg13g2_decap_8
XFILLER_44_913 VPWR VGND sg13g2_decap_8
XFILLER_28_464 VPWR VGND sg13g2_decap_8
XFILLER_16_648 VPWR VGND sg13g2_decap_8
XFILLER_15_147 VPWR VGND sg13g2_decap_8
XFILLER_43_489 VPWR VGND sg13g2_decap_8
XFILLER_31_629 VPWR VGND sg13g2_decap_8
XFILLER_12_865 VPWR VGND sg13g2_decap_8
XFILLER_24_692 VPWR VGND sg13g2_decap_8
XFILLER_8_825 VPWR VGND sg13g2_decap_8
XFILLER_7_313 VPWR VGND sg13g2_decap_8
XFILLER_11_353 VPWR VGND sg13g2_decap_8
XFILLER_7_49 VPWR VGND sg13g2_decap_8
Xclkbuf_4_9_0_clk clknet_0_clk clknet_4_9_0_clk VPWR VGND sg13g2_buf_8
XFILLER_39_707 VPWR VGND sg13g2_decap_8
XFILLER_47_784 VPWR VGND sg13g2_decap_8
XFILLER_19_497 VPWR VGND sg13g2_decap_8
XFILLER_34_423 VPWR VGND sg13g2_decap_8
XFILLER_35_935 VPWR VGND sg13g2_decap_8
XFILLER_34_467 VPWR VGND sg13g2_decap_8
XFILLER_21_139 VPWR VGND sg13g2_decap_8
XFILLER_30_640 VPWR VGND sg13g2_decap_8
XFILLER_29_206 VPWR VGND sg13g2_decap_8
XFILLER_29_217 VPWR VGND sg13g2_fill_1
XFILLER_38_740 VPWR VGND sg13g2_decap_8
XFILLER_44_209 VPWR VGND sg13g2_fill_2
XFILLER_26_935 VPWR VGND sg13g2_decap_8
XFILLER_37_272 VPWR VGND sg13g2_decap_8
XFILLER_37_294 VPWR VGND sg13g2_fill_2
XFILLER_40_459 VPWR VGND sg13g2_decap_8
XFILLER_21_673 VPWR VGND sg13g2_decap_8
XFILLER_20_172 VPWR VGND sg13g2_decap_8
XFILLER_10_1026 VPWR VGND sg13g2_fill_2
XFILLER_0_511 VPWR VGND sg13g2_decap_8
XFILLER_0_588 VPWR VGND sg13g2_decap_8
XFILLER_48_559 VPWR VGND sg13g2_decap_8
XFILLER_44_710 VPWR VGND sg13g2_decap_8
XFILLER_16_423 VPWR VGND sg13g2_fill_2
XFILLER_17_957 VPWR VGND sg13g2_decap_8
XFILLER_43_231 VPWR VGND sg13g2_decap_8
XFILLER_44_787 VPWR VGND sg13g2_decap_8
XFILLER_31_426 VPWR VGND sg13g2_decap_8
XFILLER_32_949 VPWR VGND sg13g2_decap_8
XFILLER_8_622 VPWR VGND sg13g2_decap_8
XFILLER_12_662 VPWR VGND sg13g2_decap_8
XFILLER_40_960 VPWR VGND sg13g2_decap_8
XFILLER_7_154 VPWR VGND sg13g2_decap_8
XFILLER_8_699 VPWR VGND sg13g2_decap_8
XFILLER_4_850 VPWR VGND sg13g2_decap_8
XFILLER_3_382 VPWR VGND sg13g2_decap_8
XFILLER_21_4 VPWR VGND sg13g2_decap_8
XFILLER_47_581 VPWR VGND sg13g2_decap_8
XFILLER_35_732 VPWR VGND sg13g2_decap_8
XFILLER_23_905 VPWR VGND sg13g2_decap_8
XFILLER_34_231 VPWR VGND sg13g2_decap_8
XFILLER_31_993 VPWR VGND sg13g2_decap_8
XFILLER_8_81 VPWR VGND sg13g2_decap_8
XFILLER_26_732 VPWR VGND sg13g2_decap_8
XFILLER_14_938 VPWR VGND sg13g2_decap_8
XFILLER_43_56 VPWR VGND sg13g2_fill_2
XFILLER_41_757 VPWR VGND sg13g2_decap_8
XFILLER_43_78 VPWR VGND sg13g2_decap_8
XFILLER_40_256 VPWR VGND sg13g2_fill_1
XFILLER_5_647 VPWR VGND sg13g2_decap_8
XFILLER_4_102 VPWR VGND sg13g2_decap_4
XFILLER_4_179 VPWR VGND sg13g2_decap_8
XFILLER_4_39 VPWR VGND sg13g2_decap_8
XFILLER_1_831 VPWR VGND sg13g2_decap_8
XFILLER_49_835 VPWR VGND sg13g2_decap_8
XFILLER_48_323 VPWR VGND sg13g2_decap_8
XFILLER_0_385 VPWR VGND sg13g2_decap_8
XFILLER_1_1013 VPWR VGND sg13g2_decap_8
XFILLER_17_754 VPWR VGND sg13g2_decap_8
XFILLER_44_584 VPWR VGND sg13g2_decap_8
X_587_ net67 VGND VPWR _127_ DP_4.matrix\[10\] clknet_5_2__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_746 VPWR VGND sg13g2_decap_8
XFILLER_9_920 VPWR VGND sg13g2_decap_8
XFILLER_31_245 VPWR VGND sg13g2_decap_8
XFILLER_8_463 VPWR VGND sg13g2_decap_8
XFILLER_9_997 VPWR VGND sg13g2_decap_8
XFILLER_39_334 VPWR VGND sg13g2_decap_8
XFILLER_39_367 VPWR VGND sg13g2_fill_1
XFILLER_22_201 VPWR VGND sg13g2_decap_8
XFILLER_23_702 VPWR VGND sg13g2_decap_8
XFILLER_22_245 VPWR VGND sg13g2_decap_4
XFILLER_22_267 VPWR VGND sg13g2_fill_2
XFILLER_23_779 VPWR VGND sg13g2_decap_8
XFILLER_31_790 VPWR VGND sg13g2_decap_8
XFILLER_1_116 VPWR VGND sg13g2_decap_8
XFILLER_2_628 VPWR VGND sg13g2_decap_8
XFILLER_46_816 VPWR VGND sg13g2_decap_8
X_510_ net70 VGND VPWR net180 mac2.sum_lvl1_ff\[9\] clknet_5_9__leaf_clk sg13g2_dfrbpq_1
X_441_ net39 _135_ VPWR VGND sg13g2_buf_1
XFILLER_14_735 VPWR VGND sg13g2_decap_8
X_372_ _219_ _218_ _063_ VPWR VGND sg13g2_xor2_1
XFILLER_9_216 VPWR VGND sg13g2_decap_4
XFILLER_13_267 VPWR VGND sg13g2_decap_8
XFILLER_41_554 VPWR VGND sg13g2_decap_8
XFILLER_10_963 VPWR VGND sg13g2_decap_8
XFILLER_5_422 VPWR VGND sg13g2_fill_1
XFILLER_6_956 VPWR VGND sg13g2_decap_8
XFILLER_5_499 VPWR VGND sg13g2_decap_8
XFILLER_49_632 VPWR VGND sg13g2_decap_8
XFILLER_23_1003 VPWR VGND sg13g2_decap_8
XFILLER_0_182 VPWR VGND sg13g2_decap_8
XFILLER_36_326 VPWR VGND sg13g2_decap_8
XFILLER_37_849 VPWR VGND sg13g2_decap_8
XFILLER_44_381 VPWR VGND sg13g2_decap_8
XFILLER_32_543 VPWR VGND sg13g2_decap_8
XFILLER_20_738 VPWR VGND sg13g2_decap_8
XFILLER_9_794 VPWR VGND sg13g2_decap_8
XFILLER_30_1018 VPWR VGND sg13g2_decap_8
XFILLER_5_60 VPWR VGND sg13g2_decap_8
XFILLER_28_805 VPWR VGND sg13g2_decap_8
XFILLER_39_131 VPWR VGND sg13g2_fill_2
XFILLER_39_164 VPWR VGND sg13g2_decap_8
XFILLER_39_175 VPWR VGND sg13g2_fill_1
XFILLER_23_521 VPWR VGND sg13g2_decap_8
XFILLER_24_25 VPWR VGND sg13g2_decap_4
XFILLER_24_47 VPWR VGND sg13g2_decap_8
XFILLER_23_576 VPWR VGND sg13g2_decap_8
XFILLER_10_248 VPWR VGND sg13g2_decap_8
XFILLER_40_68 VPWR VGND sg13g2_decap_8
XFILLER_3_937 VPWR VGND sg13g2_decap_8
XFILLER_49_77 VPWR VGND sg13g2_decap_8
XFILLER_46_613 VPWR VGND sg13g2_decap_8
XFILLER_18_348 VPWR VGND sg13g2_decap_8
XFILLER_45_167 VPWR VGND sg13g2_fill_2
XFILLER_42_841 VPWR VGND sg13g2_decap_8
XFILLER_14_532 VPWR VGND sg13g2_decap_8
X_424_ net144 _118_ VPWR VGND sg13g2_buf_1
X_355_ _209_ net138 net59 VPWR VGND sg13g2_nand2_1
XFILLER_41_362 VPWR VGND sg13g2_fill_1
X_286_ mac1.sum_lvl1_ff\[1\] mac1.sum_lvl1_ff\[9\] _169_ VPWR VGND sg13g2_xor2_1
XFILLER_10_760 VPWR VGND sg13g2_decap_8
XFILLER_6_753 VPWR VGND sg13g2_decap_8
XFILLER_5_252 VPWR VGND sg13g2_decap_8
Xclkbuf_5_14__f_clk clknet_4_7_0_clk clknet_5_14__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_5_296 VPWR VGND sg13g2_decap_8
XFILLER_2_992 VPWR VGND sg13g2_decap_8
XFILLER_37_646 VPWR VGND sg13g2_decap_8
XFILLER_24_318 VPWR VGND sg13g2_decap_8
XFILLER_36_167 VPWR VGND sg13g2_decap_8
XFILLER_18_893 VPWR VGND sg13g2_decap_8
XFILLER_33_874 VPWR VGND sg13g2_decap_8
XFILLER_20_535 VPWR VGND sg13g2_decap_8
XFILLER_9_591 VPWR VGND sg13g2_decap_8
XFILLER_19_25 VPWR VGND sg13g2_decap_8
XFILLER_28_602 VPWR VGND sg13g2_decap_8
XFILLER_28_679 VPWR VGND sg13g2_decap_8
XFILLER_42_115 VPWR VGND sg13g2_decap_8
XFILLER_27_189 VPWR VGND sg13g2_decap_8
XFILLER_24_874 VPWR VGND sg13g2_decap_8
XFILLER_35_68 VPWR VGND sg13g2_decap_8
XFILLER_23_373 VPWR VGND sg13g2_decap_8
XFILLER_3_734 VPWR VGND sg13g2_decap_8
XFILLER_2_244 VPWR VGND sg13g2_decap_8
XFILLER_47_966 VPWR VGND sg13g2_decap_8
XFILLER_46_410 VPWR VGND sg13g2_decap_8
XFILLER_18_112 VPWR VGND sg13g2_decap_8
XFILLER_19_657 VPWR VGND sg13g2_decap_8
XFILLER_46_487 VPWR VGND sg13g2_decap_8
XFILLER_15_841 VPWR VGND sg13g2_decap_8
XFILLER_33_137 VPWR VGND sg13g2_decap_8
X_407_ net90 _101_ VPWR VGND sg13g2_buf_1
XFILLER_30_822 VPWR VGND sg13g2_decap_8
XFILLER_14_384 VPWR VGND sg13g2_decap_8
X_338_ _197_ _196_ _041_ VPWR VGND sg13g2_xor2_1
XFILLER_41_170 VPWR VGND sg13g2_decap_8
XFILLER_41_192 VPWR VGND sg13g2_fill_1
XFILLER_30_899 VPWR VGND sg13g2_decap_8
X_269_ _160_ net177 net93 VPWR VGND sg13g2_nand2_1
XFILLER_38_922 VPWR VGND sg13g2_decap_8
XFILLER_37_432 VPWR VGND sg13g2_decap_8
XFILLER_38_999 VPWR VGND sg13g2_decap_8
XFILLER_18_690 VPWR VGND sg13g2_decap_8
XFILLER_25_627 VPWR VGND sg13g2_decap_8
XFILLER_24_159 VPWR VGND sg13g2_decap_8
XFILLER_33_671 VPWR VGND sg13g2_decap_8
XFILLER_36_1024 VPWR VGND sg13g2_decap_4
XFILLER_21_855 VPWR VGND sg13g2_decap_8
XFILLER_20_354 VPWR VGND sg13g2_fill_2
XFILLER_43_1028 VPWR VGND sg13g2_fill_1
XFILLER_29_911 VPWR VGND sg13g2_decap_8
XFILLER_28_432 VPWR VGND sg13g2_fill_1
XFILLER_29_988 VPWR VGND sg13g2_decap_8
XFILLER_15_126 VPWR VGND sg13g2_decap_8
XFILLER_16_627 VPWR VGND sg13g2_decap_8
XFILLER_44_969 VPWR VGND sg13g2_decap_8
XFILLER_43_468 VPWR VGND sg13g2_decap_8
XFILLER_31_608 VPWR VGND sg13g2_decap_8
XFILLER_24_671 VPWR VGND sg13g2_decap_8
XFILLER_8_804 VPWR VGND sg13g2_decap_8
XFILLER_11_332 VPWR VGND sg13g2_decap_8
XFILLER_12_844 VPWR VGND sg13g2_decap_8
XFILLER_30_129 VPWR VGND sg13g2_decap_4
XFILLER_7_28 VPWR VGND sg13g2_decap_8
XFILLER_7_369 VPWR VGND sg13g2_decap_8
XFILLER_3_531 VPWR VGND sg13g2_fill_2
XFILLER_4_1011 VPWR VGND sg13g2_decap_8
XFILLER_47_763 VPWR VGND sg13g2_decap_8
XFILLER_35_914 VPWR VGND sg13g2_decap_8
XFILLER_19_476 VPWR VGND sg13g2_decap_8
XFILLER_34_446 VPWR VGND sg13g2_fill_1
XFILLER_30_696 VPWR VGND sg13g2_decap_8
XFILLER_42_0 VPWR VGND sg13g2_decap_8
XFILLER_26_914 VPWR VGND sg13g2_decap_8
XFILLER_37_251 VPWR VGND sg13g2_decap_8
XFILLER_38_796 VPWR VGND sg13g2_decap_8
XFILLER_12_118 VPWR VGND sg13g2_fill_2
XFILLER_25_479 VPWR VGND sg13g2_decap_8
XFILLER_40_405 VPWR VGND sg13g2_decap_8
XFILLER_41_939 VPWR VGND sg13g2_decap_8
XFILLER_40_438 VPWR VGND sg13g2_decap_8
XFILLER_21_652 VPWR VGND sg13g2_decap_8
XFILLER_32_14 VPWR VGND sg13g2_decap_4
XFILLER_20_151 VPWR VGND sg13g2_decap_8
XFILLER_5_829 VPWR VGND sg13g2_decap_8
XFILLER_10_1005 VPWR VGND sg13g2_decap_8
XFILLER_4_339 VPWR VGND sg13g2_decap_8
XFILLER_0_567 VPWR VGND sg13g2_decap_8
XFILLER_48_538 VPWR VGND sg13g2_decap_8
XFILLER_43_210 VPWR VGND sg13g2_decap_8
XFILLER_17_936 VPWR VGND sg13g2_decap_8
XFILLER_29_785 VPWR VGND sg13g2_decap_8
XFILLER_44_766 VPWR VGND sg13g2_decap_8
XFILLER_31_405 VPWR VGND sg13g2_decap_8
XFILLER_32_928 VPWR VGND sg13g2_decap_8
XFILLER_25_991 VPWR VGND sg13g2_decap_8
XFILLER_8_601 VPWR VGND sg13g2_decap_8
XFILLER_12_641 VPWR VGND sg13g2_decap_8
XFILLER_11_151 VPWR VGND sg13g2_decap_8
XFILLER_8_678 VPWR VGND sg13g2_decap_8
XFILLER_7_133 VPWR VGND sg13g2_decap_8
XFILLER_26_1012 VPWR VGND sg13g2_decap_8
XFILLER_14_4 VPWR VGND sg13g2_decap_8
XFILLER_47_560 VPWR VGND sg13g2_decap_8
XFILLER_19_284 VPWR VGND sg13g2_decap_8
XFILLER_35_711 VPWR VGND sg13g2_decap_8
XFILLER_34_210 VPWR VGND sg13g2_decap_8
XFILLER_22_416 VPWR VGND sg13g2_decap_8
XFILLER_35_788 VPWR VGND sg13g2_decap_8
XFILLER_16_991 VPWR VGND sg13g2_decap_8
XFILLER_31_972 VPWR VGND sg13g2_decap_8
XFILLER_8_60 VPWR VGND sg13g2_decap_8
XFILLER_30_493 VPWR VGND sg13g2_decap_8
XFILLER_40_1009 VPWR VGND sg13g2_decap_8
XFILLER_27_14 VPWR VGND sg13g2_decap_8
XFILLER_26_711 VPWR VGND sg13g2_decap_8
XFILLER_27_69 VPWR VGND sg13g2_decap_8
XFILLER_38_593 VPWR VGND sg13g2_decap_8
XFILLER_14_917 VPWR VGND sg13g2_decap_8
XFILLER_25_243 VPWR VGND sg13g2_decap_8
XFILLER_26_788 VPWR VGND sg13g2_decap_8
XFILLER_43_35 VPWR VGND sg13g2_decap_8
Xclkbuf_4_8_0_clk clknet_0_clk clknet_4_8_0_clk VPWR VGND sg13g2_buf_8
XFILLER_25_287 VPWR VGND sg13g2_decap_8
XFILLER_41_736 VPWR VGND sg13g2_decap_8
XFILLER_21_493 VPWR VGND sg13g2_decap_8
XFILLER_5_626 VPWR VGND sg13g2_decap_8
XFILLER_4_158 VPWR VGND sg13g2_decap_8
XFILLER_4_18 VPWR VGND sg13g2_decap_8
XFILLER_1_810 VPWR VGND sg13g2_decap_8
XFILLER_49_814 VPWR VGND sg13g2_decap_8
XFILLER_48_302 VPWR VGND sg13g2_decap_8
XFILLER_0_364 VPWR VGND sg13g2_decap_8
XFILLER_1_887 VPWR VGND sg13g2_decap_8
XFILLER_48_379 VPWR VGND sg13g2_decap_8
XFILLER_29_582 VPWR VGND sg13g2_decap_8
XFILLER_17_733 VPWR VGND sg13g2_decap_8
XFILLER_44_563 VPWR VGND sg13g2_decap_8
X_586_ net67 VGND VPWR _126_ DP_4.matrix\[9\] clknet_5_3__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_725 VPWR VGND sg13g2_decap_8
XFILLER_16_276 VPWR VGND sg13g2_decap_8
XFILLER_16_287 VPWR VGND sg13g2_fill_2
XFILLER_16_298 VPWR VGND sg13g2_fill_2
XFILLER_31_224 VPWR VGND sg13g2_decap_8
XFILLER_8_442 VPWR VGND sg13g2_decap_8
XFILLER_9_976 VPWR VGND sg13g2_decap_8
XFILLER_39_302 VPWR VGND sg13g2_decap_8
XFILLER_23_758 VPWR VGND sg13g2_decap_8
XFILLER_35_585 VPWR VGND sg13g2_decap_8
XFILLER_2_607 VPWR VGND sg13g2_decap_8
XFILLER_38_35 VPWR VGND sg13g2_decap_8
XFILLER_38_46 VPWR VGND sg13g2_fill_1
XFILLER_45_327 VPWR VGND sg13g2_decap_8
XFILLER_18_519 VPWR VGND sg13g2_decap_8
XFILLER_45_338 VPWR VGND sg13g2_fill_1
XFILLER_14_714 VPWR VGND sg13g2_decap_8
X_440_ net158 _134_ VPWR VGND sg13g2_buf_1
XFILLER_13_224 VPWR VGND sg13g2_decap_8
XFILLER_26_585 VPWR VGND sg13g2_decap_8
X_371_ _219_ net144 net37 VPWR VGND sg13g2_nand2_1
XFILLER_41_533 VPWR VGND sg13g2_decap_8
XFILLER_9_228 VPWR VGND sg13g2_decap_4
XFILLER_10_942 VPWR VGND sg13g2_decap_8
XFILLER_6_935 VPWR VGND sg13g2_decap_8
XFILLER_5_401 VPWR VGND sg13g2_fill_1
XFILLER_49_611 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_1_684 VPWR VGND sg13g2_decap_8
XFILLER_49_688 VPWR VGND sg13g2_decap_8
XFILLER_48_176 VPWR VGND sg13g2_decap_4
XFILLER_36_305 VPWR VGND sg13g2_decap_8
XFILLER_37_828 VPWR VGND sg13g2_decap_8
XFILLER_48_198 VPWR VGND sg13g2_decap_8
XFILLER_17_552 VPWR VGND sg13g2_decap_8
XFILLER_44_360 VPWR VGND sg13g2_decap_8
XFILLER_32_522 VPWR VGND sg13g2_decap_8
X_569_ net67 VGND VPWR _109_ DP_3.matrix\[10\] clknet_5_2__leaf_clk sg13g2_dfrbpq_1
XFILLER_20_717 VPWR VGND sg13g2_decap_8
XFILLER_32_599 VPWR VGND sg13g2_decap_8
XFILLER_9_773 VPWR VGND sg13g2_decap_8
XFILLER_5_990 VPWR VGND sg13g2_decap_8
XFILLER_39_110 VPWR VGND sg13g2_decap_8
XFILLER_39_143 VPWR VGND sg13g2_decap_8
XFILLER_35_382 VPWR VGND sg13g2_decap_8
XFILLER_39_1022 VPWR VGND sg13g2_decap_8
XFILLER_11_739 VPWR VGND sg13g2_decap_8
XFILLER_10_227 VPWR VGND sg13g2_decap_8
XFILLER_40_14 VPWR VGND sg13g2_fill_2
XFILLER_40_47 VPWR VGND sg13g2_decap_8
XFILLER_3_916 VPWR VGND sg13g2_decap_8
XFILLER_2_437 VPWR VGND sg13g2_decap_8
XFILLER_46_1026 VPWR VGND sg13g2_fill_2
XFILLER_49_56 VPWR VGND sg13g2_decap_8
XFILLER_19_839 VPWR VGND sg13g2_decap_8
XFILLER_18_327 VPWR VGND sg13g2_decap_8
XFILLER_46_669 VPWR VGND sg13g2_decap_8
XFILLER_45_146 VPWR VGND sg13g2_decap_8
X_423_ net102 _117_ VPWR VGND sg13g2_buf_1
XFILLER_42_820 VPWR VGND sg13g2_decap_8
XFILLER_14_511 VPWR VGND sg13g2_decap_8
XFILLER_27_883 VPWR VGND sg13g2_decap_8
XFILLER_41_341 VPWR VGND sg13g2_decap_8
XFILLER_42_897 VPWR VGND sg13g2_decap_8
XFILLER_14_588 VPWR VGND sg13g2_decap_8
X_354_ _208_ net150 net105 VPWR VGND sg13g2_nand2_1
X_285_ _168_ net175 net145 VPWR VGND sg13g2_nand2_1
XFILLER_6_732 VPWR VGND sg13g2_decap_8
XFILLER_5_231 VPWR VGND sg13g2_decap_8
XFILLER_46_7 VPWR VGND sg13g2_decap_8
XFILLER_2_971 VPWR VGND sg13g2_decap_8
XFILLER_1_481 VPWR VGND sg13g2_decap_8
XFILLER_49_485 VPWR VGND sg13g2_decap_8
XFILLER_37_625 VPWR VGND sg13g2_decap_8
XFILLER_18_872 VPWR VGND sg13g2_decap_8
XFILLER_25_809 VPWR VGND sg13g2_decap_8
XFILLER_36_146 VPWR VGND sg13g2_decap_8
XFILLER_17_371 VPWR VGND sg13g2_decap_8
XFILLER_33_853 VPWR VGND sg13g2_decap_8
XFILLER_20_514 VPWR VGND sg13g2_decap_8
XFILLER_32_396 VPWR VGND sg13g2_decap_8
XFILLER_9_570 VPWR VGND sg13g2_decap_8
XFILLER_28_658 VPWR VGND sg13g2_decap_8
XFILLER_15_308 VPWR VGND sg13g2_decap_8
XFILLER_16_809 VPWR VGND sg13g2_decap_8
XFILLER_27_146 VPWR VGND sg13g2_decap_4
XFILLER_27_168 VPWR VGND sg13g2_decap_8
XFILLER_35_14 VPWR VGND sg13g2_decap_8
XFILLER_35_25 VPWR VGND sg13g2_fill_2
XFILLER_24_853 VPWR VGND sg13g2_decap_8
Xclkbuf_5_20__f_clk clknet_4_10_0_clk clknet_5_20__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_23_352 VPWR VGND sg13g2_decap_8
XFILLER_3_713 VPWR VGND sg13g2_decap_8
XFILLER_2_223 VPWR VGND sg13g2_decap_8
XFILLER_47_945 VPWR VGND sg13g2_decap_8
XFILLER_19_636 VPWR VGND sg13g2_decap_8
XFILLER_20_1018 VPWR VGND sg13g2_decap_8
XFILLER_46_466 VPWR VGND sg13g2_decap_8
XFILLER_15_820 VPWR VGND sg13g2_decap_8
XFILLER_27_680 VPWR VGND sg13g2_decap_8
X_406_ net120 _100_ VPWR VGND sg13g2_buf_1
XFILLER_14_363 VPWR VGND sg13g2_decap_8
XFILLER_15_897 VPWR VGND sg13g2_decap_8
XFILLER_30_801 VPWR VGND sg13g2_decap_8
XFILLER_42_694 VPWR VGND sg13g2_decap_8
X_337_ _197_ net157 net42 VPWR VGND sg13g2_nand2_1
XFILLER_30_878 VPWR VGND sg13g2_decap_8
X_268_ mac2.total_sum\[0\] mac1.total_sum\[0\] net1 VPWR VGND sg13g2_xor2_1
XFILLER_38_901 VPWR VGND sg13g2_decap_8
XFILLER_49_282 VPWR VGND sg13g2_decap_8
XFILLER_37_411 VPWR VGND sg13g2_decap_8
XFILLER_25_606 VPWR VGND sg13g2_decap_8
XFILLER_38_978 VPWR VGND sg13g2_decap_8
XFILLER_37_499 VPWR VGND sg13g2_decap_8
XFILLER_24_138 VPWR VGND sg13g2_decap_8
XFILLER_36_1003 VPWR VGND sg13g2_decap_8
XFILLER_33_650 VPWR VGND sg13g2_decap_8
XFILLER_20_333 VPWR VGND sg13g2_decap_8
XFILLER_21_834 VPWR VGND sg13g2_decap_8
XFILLER_20_388 VPWR VGND sg13g2_decap_8
XFILLER_43_1007 VPWR VGND sg13g2_decap_8
XFILLER_0_749 VPWR VGND sg13g2_decap_8
XFILLER_28_411 VPWR VGND sg13g2_decap_8
XFILLER_46_35 VPWR VGND sg13g2_decap_8
XFILLER_16_606 VPWR VGND sg13g2_decap_8
XFILLER_29_967 VPWR VGND sg13g2_decap_8
XFILLER_44_948 VPWR VGND sg13g2_decap_8
XFILLER_43_447 VPWR VGND sg13g2_decap_8
XFILLER_24_650 VPWR VGND sg13g2_decap_8
XFILLER_11_311 VPWR VGND sg13g2_decap_8
XFILLER_12_823 VPWR VGND sg13g2_decap_8
XFILLER_7_348 VPWR VGND sg13g2_decap_8
XFILLER_11_388 VPWR VGND sg13g2_decap_8
XFILLER_3_510 VPWR VGND sg13g2_decap_8
XFILLER_11_60 VPWR VGND sg13g2_decap_8
XFILLER_11_93 VPWR VGND sg13g2_decap_4
XFILLER_3_587 VPWR VGND sg13g2_decap_8
XFILLER_47_742 VPWR VGND sg13g2_decap_8
XFILLER_19_455 VPWR VGND sg13g2_decap_8
XFILLER_46_252 VPWR VGND sg13g2_decap_8
XFILLER_42_491 VPWR VGND sg13g2_decap_8
XFILLER_14_171 VPWR VGND sg13g2_fill_1
XFILLER_15_694 VPWR VGND sg13g2_decap_8
XFILLER_30_675 VPWR VGND sg13g2_decap_8
XFILLER_6_370 VPWR VGND sg13g2_decap_8
XFILLER_35_0 VPWR VGND sg13g2_decap_8
XFILLER_38_775 VPWR VGND sg13g2_decap_8
XFILLER_25_403 VPWR VGND sg13g2_decap_4
XFILLER_16_49 VPWR VGND sg13g2_decap_8
XFILLER_25_458 VPWR VGND sg13g2_decap_8
XFILLER_37_296 VPWR VGND sg13g2_fill_1
XFILLER_41_918 VPWR VGND sg13g2_decap_8
XFILLER_21_631 VPWR VGND sg13g2_decap_8
XFILLER_32_59 VPWR VGND sg13g2_decap_8
XFILLER_5_808 VPWR VGND sg13g2_decap_8
XFILLER_4_318 VPWR VGND sg13g2_decap_8
XFILLER_10_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_546 VPWR VGND sg13g2_decap_8
XFILLER_48_517 VPWR VGND sg13g2_decap_8
XFILLER_29_764 VPWR VGND sg13g2_decap_8
XFILLER_17_915 VPWR VGND sg13g2_decap_8
XFILLER_28_274 VPWR VGND sg13g2_decap_8
XFILLER_44_745 VPWR VGND sg13g2_decap_8
XFILLER_28_285 VPWR VGND sg13g2_fill_2
XFILLER_32_907 VPWR VGND sg13g2_decap_8
XFILLER_25_970 VPWR VGND sg13g2_decap_8
XFILLER_43_288 VPWR VGND sg13g2_decap_8
XFILLER_12_620 VPWR VGND sg13g2_decap_8
XFILLER_7_112 VPWR VGND sg13g2_decap_8
XFILLER_12_697 VPWR VGND sg13g2_decap_8
XFILLER_40_995 VPWR VGND sg13g2_decap_8
XFILLER_8_657 VPWR VGND sg13g2_decap_8
XFILLER_7_189 VPWR VGND sg13g2_decap_8
XFILLER_4_885 VPWR VGND sg13g2_decap_8
XFILLER_3_395 VPWR VGND sg13g2_fill_2
XFILLER_39_539 VPWR VGND sg13g2_decap_8
XFILLER_19_263 VPWR VGND sg13g2_decap_8
XFILLER_16_970 VPWR VGND sg13g2_decap_8
XFILLER_34_266 VPWR VGND sg13g2_decap_8
XFILLER_35_767 VPWR VGND sg13g2_decap_8
XFILLER_15_480 VPWR VGND sg13g2_decap_8
XFILLER_31_951 VPWR VGND sg13g2_decap_8
XFILLER_30_472 VPWR VGND sg13g2_decap_8
XFILLER_33_1028 VPWR VGND sg13g2_fill_1
XFILLER_27_48 VPWR VGND sg13g2_decap_8
XFILLER_38_572 VPWR VGND sg13g2_decap_8
XFILLER_25_222 VPWR VGND sg13g2_decap_8
XFILLER_43_14 VPWR VGND sg13g2_decap_8
XFILLER_26_767 VPWR VGND sg13g2_decap_8
XFILLER_41_715 VPWR VGND sg13g2_decap_8
XFILLER_13_439 VPWR VGND sg13g2_decap_8
XFILLER_40_214 VPWR VGND sg13g2_decap_8
XFILLER_40_225 VPWR VGND sg13g2_fill_2
XFILLER_40_247 VPWR VGND sg13g2_decap_8
XFILLER_21_472 VPWR VGND sg13g2_decap_8
XFILLER_22_984 VPWR VGND sg13g2_decap_8
XFILLER_5_605 VPWR VGND sg13g2_decap_8
XFILLER_49_1024 VPWR VGND sg13g2_decap_4
XFILLER_4_137 VPWR VGND sg13g2_decap_8
XFILLER_0_343 VPWR VGND sg13g2_decap_8
XFILLER_1_866 VPWR VGND sg13g2_decap_8
XFILLER_48_358 VPWR VGND sg13g2_decap_8
XFILLER_17_712 VPWR VGND sg13g2_decap_8
XFILLER_29_561 VPWR VGND sg13g2_decap_8
XFILLER_44_542 VPWR VGND sg13g2_decap_8
XFILLER_16_222 VPWR VGND sg13g2_decap_8
XFILLER_17_81 VPWR VGND sg13g2_decap_8
XFILLER_17_789 VPWR VGND sg13g2_decap_8
X_585_ net67 VGND VPWR _125_ DP_4.matrix\[1\] clknet_5_2__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_704 VPWR VGND sg13g2_decap_8
XFILLER_31_203 VPWR VGND sg13g2_decap_8
XFILLER_8_421 VPWR VGND sg13g2_decap_8
XFILLER_13_984 VPWR VGND sg13g2_decap_8
XFILLER_9_955 VPWR VGND sg13g2_decap_8
XFILLER_40_792 VPWR VGND sg13g2_decap_8
XFILLER_4_682 VPWR VGND sg13g2_decap_8
XFILLER_48_881 VPWR VGND sg13g2_decap_8
XFILLER_35_564 VPWR VGND sg13g2_decap_8
Xclkbuf_5_1__f_clk clknet_4_0_0_clk clknet_5_1__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_23_737 VPWR VGND sg13g2_decap_8
XFILLER_13_39 VPWR VGND sg13g2_decap_8
XFILLER_38_14 VPWR VGND sg13g2_decap_8
XFILLER_38_69 VPWR VGND sg13g2_decap_8
XFILLER_45_306 VPWR VGND sg13g2_decap_8
XFILLER_26_564 VPWR VGND sg13g2_decap_8
XFILLER_13_203 VPWR VGND sg13g2_decap_8
X_370_ _218_ net143 net89 VPWR VGND sg13g2_nand2_1
XFILLER_41_512 VPWR VGND sg13g2_decap_8
XFILLER_10_921 VPWR VGND sg13g2_decap_8
XFILLER_16_1012 VPWR VGND sg13g2_decap_8
XFILLER_22_781 VPWR VGND sg13g2_decap_8
XFILLER_41_589 VPWR VGND sg13g2_decap_8
XFILLER_6_914 VPWR VGND sg13g2_decap_8
XFILLER_5_413 VPWR VGND sg13g2_decap_8
XFILLER_10_998 VPWR VGND sg13g2_decap_8
XFILLER_5_457 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_1_663 VPWR VGND sg13g2_decap_8
XFILLER_49_667 VPWR VGND sg13g2_decap_8
XFILLER_37_807 VPWR VGND sg13g2_decap_8
XFILLER_48_155 VPWR VGND sg13g2_decap_8
XFILLER_48_188 VPWR VGND sg13g2_fill_1
XFILLER_28_91 VPWR VGND sg13g2_decap_8
XFILLER_29_391 VPWR VGND sg13g2_decap_4
XFILLER_17_564 VPWR VGND sg13g2_decap_8
XFILLER_45_884 VPWR VGND sg13g2_decap_8
X_568_ net67 VGND VPWR _108_ DP_3.matrix\[9\] clknet_5_3__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_501 VPWR VGND sg13g2_decap_8
X_499_ net80 VGND VPWR _060_ mac2.products_ff\[85\] clknet_5_15__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_578 VPWR VGND sg13g2_decap_8
XFILLER_9_752 VPWR VGND sg13g2_decap_8
XFILLER_12_280 VPWR VGND sg13g2_decap_8
XFILLER_13_781 VPWR VGND sg13g2_decap_8
XFILLER_8_273 VPWR VGND sg13g2_decap_8
XFILLER_8_262 VPWR VGND sg13g2_fill_2
XFILLER_5_95 VPWR VGND sg13g2_decap_8
Xclkbuf_4_7_0_clk clknet_0_clk clknet_4_7_0_clk VPWR VGND sg13g2_buf_8
XFILLER_39_133 VPWR VGND sg13g2_fill_1
XFILLER_42_309 VPWR VGND sg13g2_decap_8
XFILLER_39_1001 VPWR VGND sg13g2_decap_8
XFILLER_35_361 VPWR VGND sg13g2_decap_8
XFILLER_36_884 VPWR VGND sg13g2_decap_8
XFILLER_11_718 VPWR VGND sg13g2_decap_8
XFILLER_46_1005 VPWR VGND sg13g2_decap_8
XFILLER_49_35 VPWR VGND sg13g2_decap_8
XFILLER_18_306 VPWR VGND sg13g2_decap_8
XFILLER_19_818 VPWR VGND sg13g2_decap_8
XFILLER_46_648 VPWR VGND sg13g2_decap_8
XFILLER_45_125 VPWR VGND sg13g2_decap_8
XFILLER_27_862 VPWR VGND sg13g2_decap_8
X_422_ net125 _116_ VPWR VGND sg13g2_buf_1
XFILLER_26_394 VPWR VGND sg13g2_decap_4
XFILLER_41_320 VPWR VGND sg13g2_decap_8
XFILLER_42_876 VPWR VGND sg13g2_decap_8
XFILLER_14_567 VPWR VGND sg13g2_decap_8
X_353_ _207_ _206_ _051_ VPWR VGND sg13g2_xor2_1
X_284_ net99 mac1.products_ff\[102\] _008_ VPWR VGND sg13g2_xor2_1
XFILLER_6_711 VPWR VGND sg13g2_decap_8
XFILLER_10_795 VPWR VGND sg13g2_decap_8
XFILLER_5_210 VPWR VGND sg13g2_decap_8
XFILLER_6_788 VPWR VGND sg13g2_decap_8
XFILLER_30_70 VPWR VGND sg13g2_decap_8
XFILLER_2_950 VPWR VGND sg13g2_decap_8
XFILLER_1_460 VPWR VGND sg13g2_decap_8
XFILLER_39_7 VPWR VGND sg13g2_decap_8
XFILLER_49_464 VPWR VGND sg13g2_decap_8
XFILLER_37_604 VPWR VGND sg13g2_decap_8
XFILLER_36_114 VPWR VGND sg13g2_decap_4
XFILLER_18_851 VPWR VGND sg13g2_decap_8
XFILLER_45_681 VPWR VGND sg13g2_decap_8
XFILLER_33_832 VPWR VGND sg13g2_decap_8
XFILLER_17_394 VPWR VGND sg13g2_decap_4
XFILLER_32_375 VPWR VGND sg13g2_decap_8
XFILLER_27_125 VPWR VGND sg13g2_decap_8
XFILLER_28_637 VPWR VGND sg13g2_decap_8
XFILLER_43_629 VPWR VGND sg13g2_decap_8
XFILLER_36_681 VPWR VGND sg13g2_decap_8
XFILLER_23_331 VPWR VGND sg13g2_decap_8
XFILLER_24_832 VPWR VGND sg13g2_decap_8
XFILLER_11_515 VPWR VGND sg13g2_decap_8
XFILLER_11_526 VPWR VGND sg13g2_fill_2
XFILLER_13_1026 VPWR VGND sg13g2_fill_2
XFILLER_2_202 VPWR VGND sg13g2_decap_8
XFILLER_4_4 VPWR VGND sg13g2_decap_8
XFILLER_3_769 VPWR VGND sg13g2_decap_8
XFILLER_2_279 VPWR VGND sg13g2_decap_8
XFILLER_47_924 VPWR VGND sg13g2_decap_8
XFILLER_19_615 VPWR VGND sg13g2_decap_8
XFILLER_46_401 VPWR VGND sg13g2_decap_4
XFILLER_46_445 VPWR VGND sg13g2_decap_8
XFILLER_18_147 VPWR VGND sg13g2_decap_8
XFILLER_34_629 VPWR VGND sg13g2_decap_8
XFILLER_26_191 VPWR VGND sg13g2_decap_8
XFILLER_42_673 VPWR VGND sg13g2_decap_8
XFILLER_15_876 VPWR VGND sg13g2_decap_8
XFILLER_25_81 VPWR VGND sg13g2_fill_2
X_405_ net59 _099_ VPWR VGND sg13g2_buf_1
X_336_ _196_ net152 net57 VPWR VGND sg13g2_nand2_1
XFILLER_30_857 VPWR VGND sg13g2_decap_8
X_267_ net3 _156_ _159_ VPWR VGND sg13g2_xnor2_1
XFILLER_10_592 VPWR VGND sg13g2_decap_8
XFILLER_6_585 VPWR VGND sg13g2_decap_8
XFILLER_49_261 VPWR VGND sg13g2_decap_8
XFILLER_38_957 VPWR VGND sg13g2_decap_8
XFILLER_37_467 VPWR VGND sg13g2_decap_8
XFILLER_24_117 VPWR VGND sg13g2_decap_8
XFILLER_21_813 VPWR VGND sg13g2_decap_8
XFILLER_32_150 VPWR VGND sg13g2_decap_8
XFILLER_20_312 VPWR VGND sg13g2_decap_8
XFILLER_20_356 VPWR VGND sg13g2_fill_1
XFILLER_32_194 VPWR VGND sg13g2_fill_2
XFILLER_21_39 VPWR VGND sg13g2_decap_8
XFILLER_0_728 VPWR VGND sg13g2_decap_8
XFILLER_47_209 VPWR VGND sg13g2_decap_8
XFILLER_46_14 VPWR VGND sg13g2_decap_8
XFILLER_29_946 VPWR VGND sg13g2_decap_8
XFILLER_44_927 VPWR VGND sg13g2_decap_8
XFILLER_28_478 VPWR VGND sg13g2_decap_8
XFILLER_12_802 VPWR VGND sg13g2_decap_8
XFILLER_23_172 VPWR VGND sg13g2_fill_2
XFILLER_12_879 VPWR VGND sg13g2_decap_8
XFILLER_8_839 VPWR VGND sg13g2_decap_8
XFILLER_7_327 VPWR VGND sg13g2_decap_8
XFILLER_11_367 VPWR VGND sg13g2_decap_8
XFILLER_3_555 VPWR VGND sg13g2_decap_4
XFILLER_3_533 VPWR VGND sg13g2_fill_1
XFILLER_38_209 VPWR VGND sg13g2_decap_8
XFILLER_47_721 VPWR VGND sg13g2_decap_8
XFILLER_46_231 VPWR VGND sg13g2_decap_8
XFILLER_47_798 VPWR VGND sg13g2_decap_8
XFILLER_35_949 VPWR VGND sg13g2_decap_8
XFILLER_34_437 VPWR VGND sg13g2_decap_8
XFILLER_15_673 VPWR VGND sg13g2_decap_8
XFILLER_43_993 VPWR VGND sg13g2_decap_8
XFILLER_42_470 VPWR VGND sg13g2_decap_8
XFILLER_14_183 VPWR VGND sg13g2_decap_4
XFILLER_30_654 VPWR VGND sg13g2_decap_8
X_319_ net168 VPWR _016_ VGND _142_ _144_ sg13g2_o21ai_1
XFILLER_7_883 VPWR VGND sg13g2_decap_8
XFILLER_38_754 VPWR VGND sg13g2_decap_8
XFILLER_25_437 VPWR VGND sg13g2_decap_8
XFILLER_26_949 VPWR VGND sg13g2_decap_8
XFILLER_37_286 VPWR VGND sg13g2_decap_4
XFILLER_21_610 VPWR VGND sg13g2_decap_8
XFILLER_34_993 VPWR VGND sg13g2_decap_8
XFILLER_21_687 VPWR VGND sg13g2_decap_8
XFILLER_20_186 VPWR VGND sg13g2_decap_8
XFILLER_0_525 VPWR VGND sg13g2_decap_8
XFILLER_29_743 VPWR VGND sg13g2_decap_8
XFILLER_44_724 VPWR VGND sg13g2_decap_8
XFILLER_28_253 VPWR VGND sg13g2_decap_8
XFILLER_43_245 VPWR VGND sg13g2_decap_8
XFILLER_16_459 VPWR VGND sg13g2_decap_8
XFILLER_19_1021 VPWR VGND sg13g2_decap_8
XFILLER_8_636 VPWR VGND sg13g2_decap_8
XFILLER_12_676 VPWR VGND sg13g2_decap_8
XFILLER_40_974 VPWR VGND sg13g2_decap_8
XFILLER_11_186 VPWR VGND sg13g2_fill_2
XFILLER_7_168 VPWR VGND sg13g2_decap_8
XFILLER_22_82 VPWR VGND sg13g2_fill_2
XFILLER_4_864 VPWR VGND sg13g2_decap_8
XFILLER_19_242 VPWR VGND sg13g2_decap_8
XFILLER_47_595 VPWR VGND sg13g2_decap_8
XFILLER_35_746 VPWR VGND sg13g2_decap_8
XFILLER_23_919 VPWR VGND sg13g2_decap_8
XFILLER_34_245 VPWR VGND sg13g2_decap_8
XFILLER_43_790 VPWR VGND sg13g2_decap_8
XFILLER_31_930 VPWR VGND sg13g2_decap_8
XFILLER_33_1007 VPWR VGND sg13g2_decap_8
XFILLER_8_95 VPWR VGND sg13g2_decap_8
XFILLER_7_680 VPWR VGND sg13g2_decap_8
XFILLER_38_551 VPWR VGND sg13g2_decap_8
XFILLER_26_746 VPWR VGND sg13g2_decap_8
XFILLER_13_407 VPWR VGND sg13g2_fill_2
XFILLER_13_418 VPWR VGND sg13g2_decap_8
XFILLER_22_963 VPWR VGND sg13g2_decap_8
XFILLER_34_790 VPWR VGND sg13g2_decap_8
XFILLER_21_451 VPWR VGND sg13g2_decap_8
XFILLER_49_1003 VPWR VGND sg13g2_decap_8
XFILLER_1_845 VPWR VGND sg13g2_decap_8
XFILLER_0_322 VPWR VGND sg13g2_decap_8
XFILLER_49_849 VPWR VGND sg13g2_decap_8
XFILLER_48_337 VPWR VGND sg13g2_decap_8
XFILLER_0_399 VPWR VGND sg13g2_decap_8
XFILLER_29_540 VPWR VGND sg13g2_decap_8
XFILLER_44_521 VPWR VGND sg13g2_decap_8
XFILLER_1_1027 VPWR VGND sg13g2_fill_2
XFILLER_17_60 VPWR VGND sg13g2_decap_8
XFILLER_17_768 VPWR VGND sg13g2_decap_8
X_584_ net67 VGND VPWR _124_ DP_4.matrix\[0\] clknet_5_8__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_598 VPWR VGND sg13g2_decap_8
XFILLER_13_963 VPWR VGND sg13g2_decap_8
XFILLER_31_259 VPWR VGND sg13g2_decap_8
XFILLER_9_934 VPWR VGND sg13g2_decap_8
XFILLER_40_771 VPWR VGND sg13g2_decap_8
XFILLER_33_81 VPWR VGND sg13g2_decap_8
XFILLER_8_477 VPWR VGND sg13g2_decap_8
XFILLER_4_661 VPWR VGND sg13g2_decap_8
XFILLER_39_348 VPWR VGND sg13g2_fill_1
XFILLER_48_860 VPWR VGND sg13g2_decap_8
XFILLER_35_543 VPWR VGND sg13g2_decap_8
XFILLER_23_716 VPWR VGND sg13g2_decap_8
XFILLER_22_259 VPWR VGND sg13g2_decap_4
XFILLER_13_18 VPWR VGND sg13g2_decap_8
XFILLER_30_281 VPWR VGND sg13g2_decap_8
XFILLER_39_882 VPWR VGND sg13g2_decap_8
XFILLER_26_543 VPWR VGND sg13g2_decap_8
XFILLER_38_392 VPWR VGND sg13g2_decap_8
XFILLER_14_749 VPWR VGND sg13g2_decap_8
XFILLER_10_900 VPWR VGND sg13g2_decap_8
XFILLER_22_760 VPWR VGND sg13g2_decap_8
XFILLER_41_568 VPWR VGND sg13g2_decap_8
XFILLER_10_977 VPWR VGND sg13g2_decap_8
XFILLER_21_292 VPWR VGND sg13g2_decap_8
XFILLER_1_642 VPWR VGND sg13g2_decap_8
XFILLER_49_646 VPWR VGND sg13g2_decap_8
XFILLER_48_134 VPWR VGND sg13g2_decap_8
XFILLER_0_196 VPWR VGND sg13g2_decap_8
XFILLER_23_1017 VPWR VGND sg13g2_decap_8
XFILLER_23_1028 VPWR VGND sg13g2_fill_1
XFILLER_28_70 VPWR VGND sg13g2_decap_8
XFILLER_29_370 VPWR VGND sg13g2_decap_8
XFILLER_45_863 VPWR VGND sg13g2_decap_8
X_567_ net68 VGND VPWR _107_ DP_3.matrix\[1\] clknet_5_8__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_395 VPWR VGND sg13g2_decap_8
XFILLER_32_557 VPWR VGND sg13g2_decap_8
X_498_ net80 VGND VPWR _037_ mac2.products_ff\[69\] clknet_5_14__leaf_clk sg13g2_dfrbpq_1
XFILLER_13_760 VPWR VGND sg13g2_decap_8
XFILLER_9_731 VPWR VGND sg13g2_decap_8
XFILLER_8_241 VPWR VGND sg13g2_decap_8
XFILLER_5_74 VPWR VGND sg13g2_decap_8
XFILLER_27_307 VPWR VGND sg13g2_fill_2
XFILLER_28_819 VPWR VGND sg13g2_decap_8
XFILLER_35_340 VPWR VGND sg13g2_decap_8
XFILLER_36_863 VPWR VGND sg13g2_decap_8
XFILLER_49_14 VPWR VGND sg13g2_decap_8
XFILLER_46_1028 VPWR VGND sg13g2_fill_1
XFILLER_46_627 VPWR VGND sg13g2_decap_8
XFILLER_45_104 VPWR VGND sg13g2_decap_8
XFILLER_27_841 VPWR VGND sg13g2_decap_8
X_421_ net58 _115_ VPWR VGND sg13g2_buf_1
XFILLER_26_373 VPWR VGND sg13g2_decap_8
XFILLER_42_855 VPWR VGND sg13g2_decap_8
X_352_ _207_ net139 net44 VPWR VGND sg13g2_nand2_1
XFILLER_14_546 VPWR VGND sg13g2_decap_8
X_283_ _009_ _166_ _167_ VPWR VGND sg13g2_xnor2_1
XFILLER_41_398 VPWR VGND sg13g2_decap_8
XFILLER_14_83 VPWR VGND sg13g2_decap_8
XFILLER_10_774 VPWR VGND sg13g2_decap_8
XFILLER_6_767 VPWR VGND sg13g2_decap_8
XFILLER_49_443 VPWR VGND sg13g2_decap_8
XFILLER_18_830 VPWR VGND sg13g2_decap_8
XFILLER_45_660 VPWR VGND sg13g2_decap_8
XFILLER_33_811 VPWR VGND sg13g2_decap_8
XFILLER_44_181 VPWR VGND sg13g2_decap_8
XFILLER_32_343 VPWR VGND sg13g2_decap_4
XFILLER_33_888 VPWR VGND sg13g2_decap_8
XFILLER_20_549 VPWR VGND sg13g2_decap_8
XFILLER_19_39 VPWR VGND sg13g2_decap_8
XFILLER_28_616 VPWR VGND sg13g2_decap_8
XFILLER_27_104 VPWR VGND sg13g2_decap_8
XFILLER_43_608 VPWR VGND sg13g2_decap_8
XFILLER_24_811 VPWR VGND sg13g2_decap_8
XFILLER_36_660 VPWR VGND sg13g2_decap_8
XFILLER_42_129 VPWR VGND sg13g2_decap_8
XFILLER_23_310 VPWR VGND sg13g2_decap_8
XFILLER_24_888 VPWR VGND sg13g2_decap_8
XFILLER_11_549 VPWR VGND sg13g2_decap_8
XFILLER_23_387 VPWR VGND sg13g2_decap_8
XFILLER_7_509 VPWR VGND sg13g2_decap_8
XFILLER_13_1005 VPWR VGND sg13g2_decap_8
XFILLER_3_748 VPWR VGND sg13g2_decap_8
XFILLER_2_258 VPWR VGND sg13g2_decap_8
XFILLER_47_903 VPWR VGND sg13g2_decap_8
XFILLER_46_424 VPWR VGND sg13g2_decap_8
XFILLER_18_126 VPWR VGND sg13g2_decap_8
XFILLER_34_608 VPWR VGND sg13g2_decap_8
XFILLER_15_855 VPWR VGND sg13g2_decap_8
XFILLER_26_170 VPWR VGND sg13g2_decap_8
XFILLER_42_652 VPWR VGND sg13g2_decap_8
X_404_ net150 _098_ VPWR VGND sg13g2_buf_1
XFILLER_25_60 VPWR VGND sg13g2_decap_8
X_335_ _195_ _194_ _039_ VPWR VGND sg13g2_xor2_1
XFILLER_14_398 VPWR VGND sg13g2_decap_8
XFILLER_30_836 VPWR VGND sg13g2_decap_8
X_266_ _159_ _158_ _157_ VPWR VGND sg13g2_nand2b_1
Xclkbuf_4_6_0_clk clknet_0_clk clknet_4_6_0_clk VPWR VGND sg13g2_buf_8
XFILLER_10_571 VPWR VGND sg13g2_decap_8
XFILLER_6_531 VPWR VGND sg13g2_decap_4
XFILLER_6_575 VPWR VGND sg13g2_fill_1
XFILLER_29_1023 VPWR VGND sg13g2_decap_4
XFILLER_49_240 VPWR VGND sg13g2_decap_8
XFILLER_2_53 VPWR VGND sg13g2_decap_8
XFILLER_38_936 VPWR VGND sg13g2_decap_8
XFILLER_37_446 VPWR VGND sg13g2_decap_8
XFILLER_46_991 VPWR VGND sg13g2_decap_8
XFILLER_33_685 VPWR VGND sg13g2_decap_8
XFILLER_21_869 VPWR VGND sg13g2_decap_8
XFILLER_21_18 VPWR VGND sg13g2_decap_8
XFILLER_0_707 VPWR VGND sg13g2_decap_8
XFILLER_29_925 VPWR VGND sg13g2_decap_8
XFILLER_44_906 VPWR VGND sg13g2_decap_8
XFILLER_23_151 VPWR VGND sg13g2_decap_8
XFILLER_24_685 VPWR VGND sg13g2_decap_8
XFILLER_8_818 VPWR VGND sg13g2_decap_8
XFILLER_7_306 VPWR VGND sg13g2_decap_8
XFILLER_11_346 VPWR VGND sg13g2_decap_8
XFILLER_12_858 VPWR VGND sg13g2_decap_8
XFILLER_47_700 VPWR VGND sg13g2_decap_8
XFILLER_4_1025 VPWR VGND sg13g2_decap_4
XFILLER_19_413 VPWR VGND sg13g2_decap_4
XFILLER_47_777 VPWR VGND sg13g2_decap_8
XFILLER_28_980 VPWR VGND sg13g2_decap_8
XFILLER_34_416 VPWR VGND sg13g2_decap_8
XFILLER_35_928 VPWR VGND sg13g2_decap_8
XFILLER_43_972 VPWR VGND sg13g2_decap_8
XFILLER_15_652 VPWR VGND sg13g2_decap_8
XFILLER_30_633 VPWR VGND sg13g2_decap_8
X_318_ net95 mac2.products_ff\[0\] _022_ VPWR VGND sg13g2_xor2_1
X_249_ _015_ _146_ _147_ VPWR VGND sg13g2_xnor2_1
XFILLER_7_862 VPWR VGND sg13g2_decap_8
XFILLER_38_733 VPWR VGND sg13g2_decap_8
XFILLER_26_928 VPWR VGND sg13g2_decap_8
XFILLER_37_265 VPWR VGND sg13g2_decap_8
XFILLER_34_972 VPWR VGND sg13g2_decap_8
XFILLER_33_482 VPWR VGND sg13g2_decap_8
XFILLER_40_419 VPWR VGND sg13g2_decap_4
XFILLER_20_110 VPWR VGND sg13g2_decap_4
XFILLER_20_165 VPWR VGND sg13g2_decap_8
XFILLER_21_666 VPWR VGND sg13g2_decap_8
XFILLER_10_1019 VPWR VGND sg13g2_decap_8
XFILLER_0_504 VPWR VGND sg13g2_decap_8
XFILLER_29_722 VPWR VGND sg13g2_decap_8
XFILLER_44_703 VPWR VGND sg13g2_decap_8
XFILLER_29_799 VPWR VGND sg13g2_decap_8
XFILLER_43_224 VPWR VGND sg13g2_decap_8
XFILLER_16_416 VPWR VGND sg13g2_decap_8
XFILLER_19_1000 VPWR VGND sg13g2_decap_8
XFILLER_24_460 VPWR VGND sg13g2_decap_8
XFILLER_31_419 VPWR VGND sg13g2_decap_8
XFILLER_12_655 VPWR VGND sg13g2_decap_8
XFILLER_40_953 VPWR VGND sg13g2_decap_8
XFILLER_8_615 VPWR VGND sg13g2_decap_8
XFILLER_7_147 VPWR VGND sg13g2_decap_8
XFILLER_22_72 VPWR VGND sg13g2_fill_1
XFILLER_4_843 VPWR VGND sg13g2_decap_8
XFILLER_3_320 VPWR VGND sg13g2_decap_8
XFILLER_3_397 VPWR VGND sg13g2_fill_1
XFILLER_3_375 VPWR VGND sg13g2_decap_8
XFILLER_26_1026 VPWR VGND sg13g2_fill_2
XFILLER_19_221 VPWR VGND sg13g2_decap_8
XFILLER_47_574 VPWR VGND sg13g2_decap_8
XFILLER_19_298 VPWR VGND sg13g2_decap_8
XFILLER_34_224 VPWR VGND sg13g2_decap_8
XFILLER_35_725 VPWR VGND sg13g2_decap_8
XFILLER_31_986 VPWR VGND sg13g2_decap_8
XFILLER_8_74 VPWR VGND sg13g2_decap_8
XFILLER_40_0 VPWR VGND sg13g2_decap_8
XFILLER_38_530 VPWR VGND sg13g2_decap_8
XFILLER_26_725 VPWR VGND sg13g2_decap_8
XFILLER_43_49 VPWR VGND sg13g2_decap_8
XFILLER_22_942 VPWR VGND sg13g2_decap_8
XFILLER_0_301 VPWR VGND sg13g2_decap_8
XFILLER_1_824 VPWR VGND sg13g2_decap_8
XFILLER_49_828 VPWR VGND sg13g2_decap_8
XFILLER_48_316 VPWR VGND sg13g2_decap_8
XFILLER_0_378 VPWR VGND sg13g2_decap_8
Xclkbuf_5_26__f_clk clknet_4_13_0_clk clknet_5_26__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_1_1006 VPWR VGND sg13g2_decap_8
XFILLER_44_500 VPWR VGND sg13g2_decap_8
XFILLER_17_747 VPWR VGND sg13g2_decap_8
XFILLER_29_596 VPWR VGND sg13g2_decap_8
X_583_ net62 VGND VPWR _123_ DP_3.matrix\[73\] clknet_5_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_577 VPWR VGND sg13g2_decap_8
XFILLER_32_739 VPWR VGND sg13g2_decap_8
XFILLER_13_942 VPWR VGND sg13g2_decap_8
XFILLER_24_290 VPWR VGND sg13g2_decap_8
XFILLER_31_238 VPWR VGND sg13g2_decap_8
XFILLER_9_913 VPWR VGND sg13g2_decap_8
XFILLER_12_441 VPWR VGND sg13g2_decap_8
XFILLER_12_452 VPWR VGND sg13g2_fill_1
XFILLER_33_60 VPWR VGND sg13g2_decap_8
XFILLER_40_750 VPWR VGND sg13g2_decap_8
XFILLER_8_456 VPWR VGND sg13g2_decap_8
XFILLER_4_640 VPWR VGND sg13g2_decap_8
Xhold1 mac2.products_ff\[136\] VPWR VGND net25 sg13g2_dlygate4sd3_1
XFILLER_12_4 VPWR VGND sg13g2_decap_8
XFILLER_39_327 VPWR VGND sg13g2_decap_8
XFILLER_35_522 VPWR VGND sg13g2_decap_8
XFILLER_35_599 VPWR VGND sg13g2_decap_8
XFILLER_22_249 VPWR VGND sg13g2_fill_1
XFILLER_30_260 VPWR VGND sg13g2_decap_8
XFILLER_31_783 VPWR VGND sg13g2_decap_8
XFILLER_1_109 VPWR VGND sg13g2_decap_8
XFILLER_46_809 VPWR VGND sg13g2_decap_8
XFILLER_39_861 VPWR VGND sg13g2_decap_8
XFILLER_26_522 VPWR VGND sg13g2_decap_8
XFILLER_14_728 VPWR VGND sg13g2_decap_8
XFILLER_26_599 VPWR VGND sg13g2_decap_8
XFILLER_41_547 VPWR VGND sg13g2_decap_8
XFILLER_9_209 VPWR VGND sg13g2_decap_8
XFILLER_21_271 VPWR VGND sg13g2_decap_8
XFILLER_10_956 VPWR VGND sg13g2_decap_8
XFILLER_6_949 VPWR VGND sg13g2_decap_8
XFILLER_1_621 VPWR VGND sg13g2_decap_8
XFILLER_49_625 VPWR VGND sg13g2_decap_8
XFILLER_0_175 VPWR VGND sg13g2_decap_8
XFILLER_1_698 VPWR VGND sg13g2_decap_8
XFILLER_36_319 VPWR VGND sg13g2_decap_8
XFILLER_45_842 VPWR VGND sg13g2_decap_8
XFILLER_17_533 VPWR VGND sg13g2_fill_2
XFILLER_44_374 VPWR VGND sg13g2_decap_8
X_566_ net67 VGND VPWR _106_ DP_3.matrix\[0\] clknet_5_2__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_536 VPWR VGND sg13g2_decap_8
XFILLER_9_710 VPWR VGND sg13g2_decap_8
X_497_ net80 VGND VPWR _036_ mac2.products_ff\[68\] clknet_5_13__leaf_clk sg13g2_dfrbpq_1
XFILLER_9_787 VPWR VGND sg13g2_decap_8
XFILLER_5_53 VPWR VGND sg13g2_decap_8
XFILLER_4_492 VPWR VGND sg13g2_decap_8
XFILLER_39_124 VPWR VGND sg13g2_decap_8
XFILLER_39_157 VPWR VGND sg13g2_decap_8
XFILLER_36_842 VPWR VGND sg13g2_decap_8
XFILLER_23_514 VPWR VGND sg13g2_decap_8
XFILLER_24_18 VPWR VGND sg13g2_fill_2
XFILLER_24_29 VPWR VGND sg13g2_fill_2
XFILLER_35_396 VPWR VGND sg13g2_decap_8
XFILLER_23_569 VPWR VGND sg13g2_decap_8
XFILLER_31_580 VPWR VGND sg13g2_decap_8
XFILLER_46_606 VPWR VGND sg13g2_decap_8
XFILLER_27_820 VPWR VGND sg13g2_decap_8
XFILLER_26_352 VPWR VGND sg13g2_decap_8
XFILLER_27_897 VPWR VGND sg13g2_decap_8
X_420_ net156 _114_ VPWR VGND sg13g2_buf_1
XFILLER_42_834 VPWR VGND sg13g2_decap_8
XFILLER_14_525 VPWR VGND sg13g2_decap_8
X_351_ _206_ net122 net87 VPWR VGND sg13g2_nand2_1
XFILLER_41_355 VPWR VGND sg13g2_decap_8
X_282_ mac1.products_ff\[120\] mac1.products_ff\[103\] _167_ VPWR VGND sg13g2_xor2_1
XFILLER_14_62 VPWR VGND sg13g2_decap_8
XFILLER_10_753 VPWR VGND sg13g2_decap_8
XFILLER_6_746 VPWR VGND sg13g2_decap_8
XFILLER_5_245 VPWR VGND sg13g2_decap_8
XFILLER_2_985 VPWR VGND sg13g2_decap_8
XFILLER_49_422 VPWR VGND sg13g2_decap_8
XFILLER_7_1023 VPWR VGND sg13g2_decap_4
XFILLER_1_495 VPWR VGND sg13g2_decap_8
XFILLER_49_499 VPWR VGND sg13g2_decap_8
XFILLER_37_639 VPWR VGND sg13g2_decap_8
XFILLER_18_886 VPWR VGND sg13g2_decap_8
XFILLER_44_160 VPWR VGND sg13g2_decap_8
X_549_ net83 VGND VPWR _089_ DP_2.matrix\[1\] clknet_5_28__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_867 VPWR VGND sg13g2_decap_8
XFILLER_20_528 VPWR VGND sg13g2_decap_8
XFILLER_9_584 VPWR VGND sg13g2_decap_8
XFILLER_19_18 VPWR VGND sg13g2_decap_8
XFILLER_42_108 VPWR VGND sg13g2_decap_8
XFILLER_35_182 VPWR VGND sg13g2_decap_8
XFILLER_23_366 VPWR VGND sg13g2_decap_8
XFILLER_24_867 VPWR VGND sg13g2_decap_8
XFILLER_13_1028 VPWR VGND sg13g2_fill_1
XFILLER_3_727 VPWR VGND sg13g2_decap_8
XFILLER_2_237 VPWR VGND sg13g2_decap_8
XFILLER_18_105 VPWR VGND sg13g2_decap_8
XFILLER_47_959 VPWR VGND sg13g2_decap_8
XFILLER_42_631 VPWR VGND sg13g2_decap_8
X_403_ net44 _097_ VPWR VGND sg13g2_buf_1
XFILLER_14_300 VPWR VGND sg13g2_decap_8
XFILLER_15_834 VPWR VGND sg13g2_decap_8
XFILLER_27_694 VPWR VGND sg13g2_decap_8
X_334_ _195_ net127 net43 VPWR VGND sg13g2_nand2_1
XFILLER_14_377 VPWR VGND sg13g2_decap_8
XFILLER_25_83 VPWR VGND sg13g2_fill_1
XFILLER_30_815 VPWR VGND sg13g2_decap_8
XFILLER_41_163 VPWR VGND sg13g2_decap_8
X_265_ VGND VPWR _158_ mac2.total_sum\[2\] mac1.total_sum\[2\] sg13g2_or2_1
XFILLER_41_185 VPWR VGND sg13g2_decap_8
XFILLER_10_550 VPWR VGND sg13g2_decap_8
XFILLER_6_510 VPWR VGND sg13g2_decap_8
XFILLER_41_82 VPWR VGND sg13g2_decap_8
XFILLER_44_7 VPWR VGND sg13g2_decap_8
XFILLER_29_1002 VPWR VGND sg13g2_decap_8
XFILLER_2_782 VPWR VGND sg13g2_decap_8
XFILLER_1_292 VPWR VGND sg13g2_decap_8
XFILLER_2_32 VPWR VGND sg13g2_decap_8
XFILLER_38_915 VPWR VGND sg13g2_decap_8
XFILLER_49_296 VPWR VGND sg13g2_decap_8
XFILLER_37_425 VPWR VGND sg13g2_decap_8
XFILLER_46_970 VPWR VGND sg13g2_decap_8
XFILLER_18_683 VPWR VGND sg13g2_decap_8
XFILLER_33_664 VPWR VGND sg13g2_decap_8
XFILLER_36_1017 VPWR VGND sg13g2_decap_8
XFILLER_36_1028 VPWR VGND sg13g2_fill_1
XFILLER_20_347 VPWR VGND sg13g2_decap_8
XFILLER_21_848 VPWR VGND sg13g2_decap_8
XFILLER_9_370 VPWR VGND sg13g2_fill_1
Xclkbuf_5_7__f_clk clknet_4_3_0_clk clknet_5_7__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_29_904 VPWR VGND sg13g2_decap_8
XFILLER_46_49 VPWR VGND sg13g2_decap_4
XFILLER_28_425 VPWR VGND sg13g2_decap_8
XFILLER_15_119 VPWR VGND sg13g2_decap_8
XFILLER_23_130 VPWR VGND sg13g2_decap_8
XFILLER_24_664 VPWR VGND sg13g2_decap_8
XFILLER_12_837 VPWR VGND sg13g2_decap_8
XFILLER_11_325 VPWR VGND sg13g2_decap_8
XFILLER_20_892 VPWR VGND sg13g2_decap_8
XFILLER_3_524 VPWR VGND sg13g2_fill_2
XFILLER_4_1004 VPWR VGND sg13g2_decap_8
XFILLER_47_756 VPWR VGND sg13g2_decap_8
XFILLER_19_469 VPWR VGND sg13g2_decap_8
XFILLER_35_907 VPWR VGND sg13g2_decap_8
XFILLER_46_277 VPWR VGND sg13g2_fill_2
XFILLER_27_480 VPWR VGND sg13g2_decap_8
XFILLER_43_951 VPWR VGND sg13g2_decap_8
XFILLER_15_631 VPWR VGND sg13g2_decap_8
XFILLER_36_93 VPWR VGND sg13g2_decap_8
XFILLER_30_612 VPWR VGND sg13g2_decap_8
X_317_ _023_ _184_ _185_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_689 VPWR VGND sg13g2_decap_8
XFILLER_10_380 VPWR VGND sg13g2_decap_8
XFILLER_7_841 VPWR VGND sg13g2_decap_8
X_248_ mac1.sum_lvl2_ff\[5\] mac1.sum_lvl2_ff\[1\] _147_ VPWR VGND sg13g2_xor2_1
XFILLER_10_391 VPWR VGND sg13g2_fill_2
XFILLER_6_384 VPWR VGND sg13g2_fill_2
XFILLER_38_712 VPWR VGND sg13g2_decap_8
XFILLER_26_907 VPWR VGND sg13g2_decap_8
XFILLER_37_244 VPWR VGND sg13g2_decap_8
XFILLER_38_789 VPWR VGND sg13g2_decap_8
XFILLER_18_491 VPWR VGND sg13g2_decap_8
XFILLER_34_951 VPWR VGND sg13g2_decap_8
XFILLER_21_645 VPWR VGND sg13g2_decap_8
XFILLER_20_144 VPWR VGND sg13g2_decap_8
XFILLER_29_701 VPWR VGND sg13g2_decap_8
Xclkbuf_4_5_0_clk clknet_0_clk clknet_4_5_0_clk VPWR VGND sg13g2_buf_8
XFILLER_17_929 VPWR VGND sg13g2_decap_8
XFILLER_29_778 VPWR VGND sg13g2_decap_8
XFILLER_43_203 VPWR VGND sg13g2_decap_8
XFILLER_44_759 VPWR VGND sg13g2_decap_8
XFILLER_25_984 VPWR VGND sg13g2_decap_8
XFILLER_12_634 VPWR VGND sg13g2_decap_8
XFILLER_40_932 VPWR VGND sg13g2_decap_8
XFILLER_11_144 VPWR VGND sg13g2_decap_8
XFILLER_7_126 VPWR VGND sg13g2_decap_8
XFILLER_11_188 VPWR VGND sg13g2_fill_1
XFILLER_22_84 VPWR VGND sg13g2_fill_1
XFILLER_4_822 VPWR VGND sg13g2_decap_8
XFILLER_4_899 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_26_1005 VPWR VGND sg13g2_decap_8
XFILLER_19_200 VPWR VGND sg13g2_decap_8
XFILLER_47_553 VPWR VGND sg13g2_decap_8
XFILLER_47_92 VPWR VGND sg13g2_decap_8
XFILLER_35_704 VPWR VGND sg13g2_decap_8
XFILLER_19_277 VPWR VGND sg13g2_decap_8
XFILLER_16_984 VPWR VGND sg13g2_decap_8
XFILLER_22_409 VPWR VGND sg13g2_decap_8
XFILLER_15_494 VPWR VGND sg13g2_decap_8
XFILLER_31_965 VPWR VGND sg13g2_decap_8
XFILLER_8_53 VPWR VGND sg13g2_decap_8
XFILLER_30_486 VPWR VGND sg13g2_decap_8
XFILLER_6_170 VPWR VGND sg13g2_fill_2
XFILLER_6_192 VPWR VGND sg13g2_decap_8
XFILLER_33_0 VPWR VGND sg13g2_decap_8
XFILLER_26_704 VPWR VGND sg13g2_decap_8
XFILLER_38_586 VPWR VGND sg13g2_decap_8
XFILLER_25_236 VPWR VGND sg13g2_decap_8
XFILLER_43_28 VPWR VGND sg13g2_decap_8
XFILLER_22_921 VPWR VGND sg13g2_decap_8
XFILLER_41_729 VPWR VGND sg13g2_decap_8
XFILLER_21_486 VPWR VGND sg13g2_decap_8
XFILLER_22_998 VPWR VGND sg13g2_decap_8
XFILLER_5_619 VPWR VGND sg13g2_decap_8
XFILLER_1_803 VPWR VGND sg13g2_decap_8
XFILLER_49_807 VPWR VGND sg13g2_decap_8
XFILLER_0_357 VPWR VGND sg13g2_decap_8
X_582_ net62 VGND VPWR _122_ DP_3.matrix\[72\] clknet_5_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_726 VPWR VGND sg13g2_decap_8
XFILLER_29_575 VPWR VGND sg13g2_decap_8
XFILLER_44_556 VPWR VGND sg13g2_decap_8
XFILLER_16_269 VPWR VGND sg13g2_decap_8
XFILLER_17_95 VPWR VGND sg13g2_decap_8
XFILLER_31_217 VPWR VGND sg13g2_decap_8
XFILLER_32_718 VPWR VGND sg13g2_decap_8
XFILLER_12_420 VPWR VGND sg13g2_decap_8
XFILLER_13_921 VPWR VGND sg13g2_decap_8
XFILLER_25_781 VPWR VGND sg13g2_decap_8
XFILLER_8_435 VPWR VGND sg13g2_decap_8
XFILLER_9_969 VPWR VGND sg13g2_decap_8
XFILLER_13_998 VPWR VGND sg13g2_decap_8
XFILLER_4_696 VPWR VGND sg13g2_decap_8
XFILLER_3_173 VPWR VGND sg13g2_decap_4
Xhold2 mac2.sum_lvl1_ff\[32\] VPWR VGND net26 sg13g2_dlygate4sd3_1
XFILLER_48_895 VPWR VGND sg13g2_decap_8
XFILLER_35_501 VPWR VGND sg13g2_decap_8
XFILLER_35_578 VPWR VGND sg13g2_decap_8
XFILLER_15_280 VPWR VGND sg13g2_fill_1
XFILLER_16_781 VPWR VGND sg13g2_decap_8
XFILLER_22_239 VPWR VGND sg13g2_fill_2
XFILLER_31_762 VPWR VGND sg13g2_decap_8
XFILLER_38_28 VPWR VGND sg13g2_decap_8
XFILLER_39_840 VPWR VGND sg13g2_decap_8
XFILLER_26_501 VPWR VGND sg13g2_decap_8
XFILLER_38_361 VPWR VGND sg13g2_decap_8
XFILLER_14_707 VPWR VGND sg13g2_decap_8
XFILLER_26_578 VPWR VGND sg13g2_decap_8
XFILLER_13_217 VPWR VGND sg13g2_decap_8
XFILLER_41_526 VPWR VGND sg13g2_decap_8
XFILLER_16_1026 VPWR VGND sg13g2_fill_2
XFILLER_10_935 VPWR VGND sg13g2_decap_8
XFILLER_22_795 VPWR VGND sg13g2_decap_8
XFILLER_6_928 VPWR VGND sg13g2_decap_8
XFILLER_1_600 VPWR VGND sg13g2_decap_8
XFILLER_49_604 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_1_677 VPWR VGND sg13g2_decap_8
XFILLER_48_169 VPWR VGND sg13g2_decap_8
XFILLER_45_821 VPWR VGND sg13g2_decap_8
XFILLER_45_898 VPWR VGND sg13g2_decap_8
XFILLER_44_353 VPWR VGND sg13g2_decap_8
X_565_ net61 VGND VPWR _105_ DP_2.matrix\[73\] clknet_5_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_515 VPWR VGND sg13g2_decap_8
X_496_ net68 VGND VPWR _059_ mac2.products_ff\[52\] clknet_5_8__leaf_clk sg13g2_dfrbpq_1
XFILLER_13_795 VPWR VGND sg13g2_decap_8
XFILLER_9_766 VPWR VGND sg13g2_decap_8
XFILLER_12_294 VPWR VGND sg13g2_decap_8
XFILLER_8_287 VPWR VGND sg13g2_fill_1
XFILLER_5_983 VPWR VGND sg13g2_decap_8
XFILLER_5_32 VPWR VGND sg13g2_decap_8
XFILLER_4_471 VPWR VGND sg13g2_decap_8
XFILLER_39_103 VPWR VGND sg13g2_decap_8
XFILLER_36_821 VPWR VGND sg13g2_decap_8
XFILLER_48_692 VPWR VGND sg13g2_decap_8
XFILLER_36_898 VPWR VGND sg13g2_decap_8
XFILLER_39_1015 VPWR VGND sg13g2_decap_8
XFILLER_35_375 VPWR VGND sg13g2_decap_8
XFILLER_3_909 VPWR VGND sg13g2_decap_8
XFILLER_46_1019 VPWR VGND sg13g2_decap_8
XFILLER_49_49 VPWR VGND sg13g2_decap_8
XFILLER_45_139 VPWR VGND sg13g2_decap_8
XFILLER_26_331 VPWR VGND sg13g2_decap_8
XFILLER_38_191 VPWR VGND sg13g2_fill_2
XFILLER_42_813 VPWR VGND sg13g2_decap_8
XFILLER_14_504 VPWR VGND sg13g2_decap_8
XFILLER_27_876 VPWR VGND sg13g2_decap_8
X_350_ _205_ _204_ _049_ VPWR VGND sg13g2_xor2_1
XFILLER_41_334 VPWR VGND sg13g2_decap_8
X_281_ _166_ net193 net99 VPWR VGND sg13g2_nand2_1
XFILLER_10_732 VPWR VGND sg13g2_decap_8
XFILLER_22_592 VPWR VGND sg13g2_decap_8
XFILLER_6_725 VPWR VGND sg13g2_decap_8
XFILLER_5_224 VPWR VGND sg13g2_decap_8
XFILLER_30_84 VPWR VGND sg13g2_decap_4
XFILLER_2_964 VPWR VGND sg13g2_decap_8
XFILLER_49_401 VPWR VGND sg13g2_decap_8
XFILLER_7_1002 VPWR VGND sg13g2_decap_8
XFILLER_1_474 VPWR VGND sg13g2_decap_8
XFILLER_49_478 VPWR VGND sg13g2_decap_8
XFILLER_37_618 VPWR VGND sg13g2_decap_8
XFILLER_36_139 VPWR VGND sg13g2_decap_8
XFILLER_17_342 VPWR VGND sg13g2_fill_2
XFILLER_18_865 VPWR VGND sg13g2_decap_8
XFILLER_45_695 VPWR VGND sg13g2_decap_8
X_548_ net79 VGND VPWR _088_ DP_2.matrix\[0\] clknet_5_28__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_323 VPWR VGND sg13g2_fill_2
XFILLER_33_846 VPWR VGND sg13g2_decap_8
X_479_ net75 VGND VPWR net174 mac1.sum_lvl2_ff\[5\] clknet_5_22__leaf_clk sg13g2_dfrbpq_1
XFILLER_20_507 VPWR VGND sg13g2_decap_8
XFILLER_32_389 VPWR VGND sg13g2_decap_8
XFILLER_13_592 VPWR VGND sg13g2_decap_8
XFILLER_41_890 VPWR VGND sg13g2_decap_8
XFILLER_9_563 VPWR VGND sg13g2_decap_8
XFILLER_5_780 VPWR VGND sg13g2_decap_8
XFILLER_27_139 VPWR VGND sg13g2_decap_8
XFILLER_24_846 VPWR VGND sg13g2_decap_8
XFILLER_35_161 VPWR VGND sg13g2_decap_8
XFILLER_36_695 VPWR VGND sg13g2_decap_8
XFILLER_23_345 VPWR VGND sg13g2_decap_8
XFILLER_3_706 VPWR VGND sg13g2_decap_8
XFILLER_2_216 VPWR VGND sg13g2_decap_8
XFILLER_47_938 VPWR VGND sg13g2_decap_8
XFILLER_19_629 VPWR VGND sg13g2_decap_8
XFILLER_46_459 VPWR VGND sg13g2_decap_8
XFILLER_33_109 VPWR VGND sg13g2_fill_1
XFILLER_42_610 VPWR VGND sg13g2_decap_8
X_402_ net122 _096_ VPWR VGND sg13g2_buf_1
XFILLER_15_813 VPWR VGND sg13g2_decap_8
XFILLER_27_673 VPWR VGND sg13g2_decap_8
XFILLER_14_356 VPWR VGND sg13g2_decap_8
XFILLER_42_687 VPWR VGND sg13g2_decap_8
X_333_ _194_ net140 net41 VPWR VGND sg13g2_nand2_1
XFILLER_41_142 VPWR VGND sg13g2_decap_8
X_264_ mac1.total_sum\[2\] mac2.total_sum\[2\] _157_ VPWR VGND sg13g2_and2_1
XFILLER_41_61 VPWR VGND sg13g2_decap_8
XFILLER_6_599 VPWR VGND sg13g2_decap_8
XFILLER_2_761 VPWR VGND sg13g2_decap_8
XFILLER_37_7 VPWR VGND sg13g2_decap_8
XFILLER_1_271 VPWR VGND sg13g2_decap_8
XFILLER_2_11 VPWR VGND sg13g2_decap_8
XFILLER_49_275 VPWR VGND sg13g2_decap_8
XFILLER_37_404 VPWR VGND sg13g2_decap_8
XFILLER_18_662 VPWR VGND sg13g2_decap_8
XFILLER_17_150 VPWR VGND sg13g2_fill_1
XFILLER_45_492 VPWR VGND sg13g2_decap_8
XFILLER_33_643 VPWR VGND sg13g2_decap_8
XFILLER_21_827 VPWR VGND sg13g2_decap_8
XFILLER_32_164 VPWR VGND sg13g2_decap_4
XFILLER_20_326 VPWR VGND sg13g2_decap_8
XFILLER_28_404 VPWR VGND sg13g2_decap_8
XFILLER_46_28 VPWR VGND sg13g2_decap_8
XFILLER_43_407 VPWR VGND sg13g2_decap_4
XFILLER_37_982 VPWR VGND sg13g2_decap_8
XFILLER_24_643 VPWR VGND sg13g2_decap_8
XFILLER_36_492 VPWR VGND sg13g2_decap_8
XFILLER_11_304 VPWR VGND sg13g2_decap_8
XFILLER_12_816 VPWR VGND sg13g2_decap_8
XFILLER_20_871 VPWR VGND sg13g2_decap_8
XFILLER_3_503 VPWR VGND sg13g2_decap_8
XFILLER_11_53 VPWR VGND sg13g2_decap_8
XFILLER_2_4 VPWR VGND sg13g2_decap_8
XFILLER_11_86 VPWR VGND sg13g2_decap_8
XFILLER_47_735 VPWR VGND sg13g2_decap_8
XFILLER_46_201 VPWR VGND sg13g2_decap_8
XFILLER_19_448 VPWR VGND sg13g2_decap_8
XFILLER_46_245 VPWR VGND sg13g2_decap_8
XFILLER_43_930 VPWR VGND sg13g2_decap_8
XFILLER_15_610 VPWR VGND sg13g2_decap_8
XFILLER_36_72 VPWR VGND sg13g2_decap_8
XFILLER_14_153 VPWR VGND sg13g2_decap_8
XFILLER_15_687 VPWR VGND sg13g2_decap_8
XFILLER_42_484 VPWR VGND sg13g2_decap_8
X_316_ mac2.products_ff\[18\] mac2.products_ff\[1\] _185_ VPWR VGND sg13g2_xor2_1
XFILLER_30_668 VPWR VGND sg13g2_decap_8
X_247_ net153 mac1.sum_lvl2_ff\[0\] _014_ VPWR VGND sg13g2_xor2_1
XFILLER_7_820 VPWR VGND sg13g2_decap_8
XFILLER_11_893 VPWR VGND sg13g2_decap_8
XFILLER_7_897 VPWR VGND sg13g2_decap_8
XFILLER_6_363 VPWR VGND sg13g2_decap_8
XFILLER_37_212 VPWR VGND sg13g2_decap_8
XFILLER_37_223 VPWR VGND sg13g2_fill_1
XFILLER_38_768 VPWR VGND sg13g2_decap_8
XFILLER_19_993 VPWR VGND sg13g2_decap_8
XFILLER_34_930 VPWR VGND sg13g2_decap_8
XFILLER_33_451 VPWR VGND sg13g2_decap_8
XFILLER_21_624 VPWR VGND sg13g2_decap_8
XFILLER_0_539 VPWR VGND sg13g2_decap_8
XFILLER_17_908 VPWR VGND sg13g2_decap_8
XFILLER_29_757 VPWR VGND sg13g2_decap_8
XFILLER_44_738 VPWR VGND sg13g2_decap_8
XFILLER_28_267 VPWR VGND sg13g2_decap_8
XFILLER_43_259 VPWR VGND sg13g2_fill_2
XFILLER_12_613 VPWR VGND sg13g2_decap_8
XFILLER_25_963 VPWR VGND sg13g2_decap_8
XFILLER_40_911 VPWR VGND sg13g2_decap_8
XFILLER_7_105 VPWR VGND sg13g2_decap_8
XFILLER_40_988 VPWR VGND sg13g2_decap_8
XFILLER_4_801 VPWR VGND sg13g2_decap_8
XFILLER_22_96 VPWR VGND sg13g2_decap_8
XFILLER_4_878 VPWR VGND sg13g2_decap_8
XFILLER_26_1028 VPWR VGND sg13g2_fill_1
XFILLER_47_532 VPWR VGND sg13g2_decap_8
XFILLER_19_256 VPWR VGND sg13g2_decap_8
XFILLER_16_963 VPWR VGND sg13g2_decap_8
XFILLER_34_259 VPWR VGND sg13g2_decap_8
XFILLER_15_473 VPWR VGND sg13g2_decap_8
XFILLER_31_944 VPWR VGND sg13g2_decap_8
XFILLER_8_32 VPWR VGND sg13g2_decap_8
XFILLER_30_432 VPWR VGND sg13g2_decap_8
XFILLER_30_465 VPWR VGND sg13g2_decap_8
XFILLER_11_690 VPWR VGND sg13g2_decap_8
XFILLER_7_694 VPWR VGND sg13g2_decap_8
XFILLER_38_565 VPWR VGND sg13g2_decap_8
XFILLER_25_215 VPWR VGND sg13g2_decap_8
XFILLER_19_790 VPWR VGND sg13g2_decap_8
XFILLER_22_900 VPWR VGND sg13g2_decap_8
XFILLER_40_207 VPWR VGND sg13g2_decap_8
XFILLER_41_708 VPWR VGND sg13g2_decap_8
XFILLER_22_977 VPWR VGND sg13g2_decap_8
XFILLER_33_292 VPWR VGND sg13g2_decap_8
XFILLER_21_465 VPWR VGND sg13g2_decap_8
XFILLER_49_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_1017 VPWR VGND sg13g2_decap_8
XFILLER_0_336 VPWR VGND sg13g2_decap_8
XFILLER_1_859 VPWR VGND sg13g2_decap_8
XFILLER_17_705 VPWR VGND sg13g2_decap_8
XFILLER_29_554 VPWR VGND sg13g2_decap_8
X_581_ net82 VGND VPWR _121_ DP_3.matrix\[64\] clknet_5_27__leaf_clk sg13g2_dfrbpq_1
XFILLER_16_215 VPWR VGND sg13g2_decap_8
XFILLER_44_535 VPWR VGND sg13g2_decap_8
XFILLER_17_74 VPWR VGND sg13g2_decap_8
XFILLER_13_900 VPWR VGND sg13g2_decap_8
XFILLER_25_760 VPWR VGND sg13g2_decap_8
XFILLER_13_977 VPWR VGND sg13g2_decap_8
XFILLER_8_414 VPWR VGND sg13g2_decap_8
XFILLER_9_948 VPWR VGND sg13g2_decap_8
XFILLER_33_95 VPWR VGND sg13g2_decap_8
XFILLER_40_785 VPWR VGND sg13g2_decap_8
XFILLER_4_675 VPWR VGND sg13g2_decap_8
XFILLER_3_152 VPWR VGND sg13g2_decap_8
Xhold3 mac1.products_ff\[136\] VPWR VGND net27 sg13g2_dlygate4sd3_1
XFILLER_48_874 VPWR VGND sg13g2_decap_8
XFILLER_35_557 VPWR VGND sg13g2_decap_8
XFILLER_16_760 VPWR VGND sg13g2_decap_8
XFILLER_31_741 VPWR VGND sg13g2_decap_8
XFILLER_30_295 VPWR VGND sg13g2_decap_8
Xclkbuf_4_4_0_clk clknet_0_clk clknet_4_4_0_clk VPWR VGND sg13g2_buf_8
XFILLER_7_491 VPWR VGND sg13g2_fill_2
XFILLER_38_340 VPWR VGND sg13g2_decap_8
XFILLER_39_896 VPWR VGND sg13g2_decap_8
XFILLER_26_557 VPWR VGND sg13g2_decap_8
XFILLER_41_505 VPWR VGND sg13g2_decap_8
XFILLER_16_1005 VPWR VGND sg13g2_decap_8
XFILLER_10_914 VPWR VGND sg13g2_decap_8
XFILLER_22_774 VPWR VGND sg13g2_decap_8
XFILLER_6_907 VPWR VGND sg13g2_decap_8
XFILLER_5_406 VPWR VGND sg13g2_decap_8
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_1_656 VPWR VGND sg13g2_decap_8
XFILLER_48_148 VPWR VGND sg13g2_decap_8
XFILLER_45_800 VPWR VGND sg13g2_decap_8
XFILLER_28_84 VPWR VGND sg13g2_decap_8
XFILLER_44_332 VPWR VGND sg13g2_decap_8
XFILLER_29_384 VPWR VGND sg13g2_decap_8
XFILLER_29_395 VPWR VGND sg13g2_fill_2
XFILLER_45_877 VPWR VGND sg13g2_decap_8
X_564_ net60 VGND VPWR _104_ DP_2.matrix\[72\] clknet_5_4__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_579 VPWR VGND sg13g2_fill_1
X_495_ net68 VGND VPWR _058_ mac2.products_ff\[51\] clknet_5_9__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_72 VPWR VGND sg13g2_decap_4
XFILLER_9_745 VPWR VGND sg13g2_decap_8
XFILLER_13_774 VPWR VGND sg13g2_decap_8
XFILLER_8_255 VPWR VGND sg13g2_decap_8
XFILLER_12_273 VPWR VGND sg13g2_decap_8
XFILLER_40_582 VPWR VGND sg13g2_decap_8
XFILLER_5_11 VPWR VGND sg13g2_decap_8
XFILLER_5_962 VPWR VGND sg13g2_decap_8
XFILLER_4_450 VPWR VGND sg13g2_decap_8
XFILLER_5_88 VPWR VGND sg13g2_decap_8
XFILLER_48_671 VPWR VGND sg13g2_decap_8
XFILLER_36_800 VPWR VGND sg13g2_decap_8
XFILLER_35_354 VPWR VGND sg13g2_decap_8
XFILLER_36_877 VPWR VGND sg13g2_decap_8
XFILLER_49_28 VPWR VGND sg13g2_decap_8
XFILLER_45_118 VPWR VGND sg13g2_decap_8
XFILLER_26_310 VPWR VGND sg13g2_decap_8
XFILLER_27_855 VPWR VGND sg13g2_decap_8
XFILLER_38_170 VPWR VGND sg13g2_decap_8
XFILLER_39_693 VPWR VGND sg13g2_decap_8
XFILLER_26_387 VPWR VGND sg13g2_decap_8
XFILLER_26_398 VPWR VGND sg13g2_fill_1
XFILLER_41_313 VPWR VGND sg13g2_decap_8
XFILLER_42_869 VPWR VGND sg13g2_decap_8
X_280_ net113 mac1.products_ff\[85\] _006_ VPWR VGND sg13g2_xor2_1
XFILLER_10_711 VPWR VGND sg13g2_decap_8
XFILLER_14_31 VPWR VGND sg13g2_fill_2
XFILLER_22_571 VPWR VGND sg13g2_decap_8
XFILLER_10_788 VPWR VGND sg13g2_decap_8
XFILLER_6_704 VPWR VGND sg13g2_decap_8
XFILLER_5_203 VPWR VGND sg13g2_decap_8
XFILLER_14_97 VPWR VGND sg13g2_decap_8
XFILLER_30_63 VPWR VGND sg13g2_decap_8
XFILLER_2_943 VPWR VGND sg13g2_decap_8
XFILLER_1_453 VPWR VGND sg13g2_decap_8
XFILLER_49_457 VPWR VGND sg13g2_decap_8
XFILLER_36_107 VPWR VGND sg13g2_decap_8
XFILLER_17_321 VPWR VGND sg13g2_decap_8
XFILLER_18_844 VPWR VGND sg13g2_decap_8
XFILLER_36_118 VPWR VGND sg13g2_fill_1
XFILLER_45_674 VPWR VGND sg13g2_decap_8
X_547_ net61 VGND VPWR _087_ DP_1.matrix\[73\] clknet_5_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_387 VPWR VGND sg13g2_decap_8
XFILLER_32_302 VPWR VGND sg13g2_decap_8
XFILLER_33_825 VPWR VGND sg13g2_decap_8
XFILLER_44_195 VPWR VGND sg13g2_decap_8
X_478_ net73 VGND VPWR net162 mac1.sum_lvl2_ff\[4\] clknet_5_17__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_368 VPWR VGND sg13g2_decap_8
XFILLER_9_542 VPWR VGND sg13g2_decap_8
XFILLER_27_118 VPWR VGND sg13g2_decap_8
XFILLER_24_825 VPWR VGND sg13g2_decap_8
XFILLER_36_674 VPWR VGND sg13g2_decap_8
XFILLER_23_324 VPWR VGND sg13g2_decap_8
XFILLER_11_508 VPWR VGND sg13g2_decap_8
XFILLER_13_1019 VPWR VGND sg13g2_decap_8
XFILLER_31_390 VPWR VGND sg13g2_decap_4
XFILLER_47_917 VPWR VGND sg13g2_decap_8
XFILLER_46_405 VPWR VGND sg13g2_fill_1
XFILLER_19_608 VPWR VGND sg13g2_decap_8
XFILLER_46_438 VPWR VGND sg13g2_decap_8
XFILLER_27_652 VPWR VGND sg13g2_decap_8
X_401_ net53 _095_ VPWR VGND sg13g2_buf_1
XFILLER_15_869 VPWR VGND sg13g2_decap_8
XFILLER_26_184 VPWR VGND sg13g2_decap_8
XFILLER_42_666 VPWR VGND sg13g2_decap_8
X_332_ _158_ _156_ _157_ net4 VPWR VGND sg13g2_a21o_2
XFILLER_25_74 VPWR VGND sg13g2_decap_8
X_263_ _153_ VPWR _156_ VGND _152_ _154_ sg13g2_o21ai_1
XFILLER_23_891 VPWR VGND sg13g2_decap_8
XFILLER_41_40 VPWR VGND sg13g2_decap_8
XFILLER_10_585 VPWR VGND sg13g2_decap_8
XFILLER_2_740 VPWR VGND sg13g2_decap_8
XFILLER_1_250 VPWR VGND sg13g2_decap_8
XFILLER_49_254 VPWR VGND sg13g2_decap_8
XFILLER_2_67 VPWR VGND sg13g2_fill_2
XFILLER_18_641 VPWR VGND sg13g2_decap_8
XFILLER_45_471 VPWR VGND sg13g2_decap_8
XFILLER_33_622 VPWR VGND sg13g2_decap_8
XFILLER_20_305 VPWR VGND sg13g2_decap_8
XFILLER_21_806 VPWR VGND sg13g2_decap_8
XFILLER_32_143 VPWR VGND sg13g2_decap_8
XFILLER_32_176 VPWR VGND sg13g2_fill_1
XFILLER_33_699 VPWR VGND sg13g2_decap_8
XFILLER_29_939 VPWR VGND sg13g2_decap_8
XFILLER_37_961 VPWR VGND sg13g2_decap_8
XFILLER_24_622 VPWR VGND sg13g2_decap_8
XFILLER_23_165 VPWR VGND sg13g2_decap_8
XFILLER_24_699 VPWR VGND sg13g2_decap_8
XFILLER_20_850 VPWR VGND sg13g2_decap_8
XFILLER_3_526 VPWR VGND sg13g2_fill_1
XFILLER_3_559 VPWR VGND sg13g2_fill_1
XFILLER_47_714 VPWR VGND sg13g2_decap_8
XFILLER_46_224 VPWR VGND sg13g2_decap_8
XFILLER_28_994 VPWR VGND sg13g2_decap_8
XFILLER_43_986 VPWR VGND sg13g2_decap_8
XFILLER_42_463 VPWR VGND sg13g2_decap_8
XFILLER_14_132 VPWR VGND sg13g2_decap_8
XFILLER_15_666 VPWR VGND sg13g2_decap_8
XFILLER_14_176 VPWR VGND sg13g2_decap_8
XFILLER_14_187 VPWR VGND sg13g2_fill_2
X_315_ _184_ net191 net95 VPWR VGND sg13g2_nand2_1
XFILLER_30_647 VPWR VGND sg13g2_decap_8
X_246_ _146_ net197 net153 VPWR VGND sg13g2_nand2_1
XFILLER_11_872 VPWR VGND sg13g2_decap_8
XFILLER_7_876 VPWR VGND sg13g2_decap_8
XFILLER_42_1023 VPWR VGND sg13g2_decap_4
XFILLER_28_4 VPWR VGND sg13g2_decap_8
XFILLER_38_747 VPWR VGND sg13g2_decap_8
XFILLER_19_972 VPWR VGND sg13g2_decap_8
XFILLER_37_279 VPWR VGND sg13g2_decap_8
XFILLER_21_603 VPWR VGND sg13g2_decap_8
XFILLER_34_986 VPWR VGND sg13g2_decap_8
XFILLER_20_102 VPWR VGND sg13g2_decap_4
XFILLER_33_496 VPWR VGND sg13g2_decap_8
XFILLER_20_179 VPWR VGND sg13g2_decap_8
Xclkbuf_5_15__f_clk clknet_4_7_0_clk clknet_5_15__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_0_518 VPWR VGND sg13g2_decap_8
XFILLER_29_736 VPWR VGND sg13g2_decap_8
XFILLER_28_246 VPWR VGND sg13g2_decap_8
XFILLER_44_717 VPWR VGND sg13g2_decap_8
XFILLER_43_238 VPWR VGND sg13g2_decap_8
XFILLER_25_942 VPWR VGND sg13g2_decap_8
XFILLER_19_1014 VPWR VGND sg13g2_decap_8
XFILLER_11_113 VPWR VGND sg13g2_decap_4
XFILLER_24_474 VPWR VGND sg13g2_fill_2
XFILLER_8_629 VPWR VGND sg13g2_decap_8
XFILLER_12_669 VPWR VGND sg13g2_decap_8
XFILLER_40_967 VPWR VGND sg13g2_decap_8
XFILLER_4_857 VPWR VGND sg13g2_decap_8
XFILLER_3_334 VPWR VGND sg13g2_decap_8
XFILLER_3_389 VPWR VGND sg13g2_fill_2
XFILLER_47_511 VPWR VGND sg13g2_decap_8
XFILLER_19_235 VPWR VGND sg13g2_decap_8
XFILLER_47_588 VPWR VGND sg13g2_decap_8
XFILLER_35_739 VPWR VGND sg13g2_decap_8
XFILLER_16_942 VPWR VGND sg13g2_decap_8
XFILLER_28_791 VPWR VGND sg13g2_decap_8
XFILLER_34_238 VPWR VGND sg13g2_decap_8
XFILLER_15_452 VPWR VGND sg13g2_decap_8
XFILLER_43_783 VPWR VGND sg13g2_decap_8
XFILLER_30_411 VPWR VGND sg13g2_decap_8
XFILLER_31_923 VPWR VGND sg13g2_decap_8
XFILLER_8_11 VPWR VGND sg13g2_decap_8
X_229_ _143_ net167 mac1.sum_lvl3_ff\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_8_88 VPWR VGND sg13g2_decap_8
XFILLER_7_673 VPWR VGND sg13g2_decap_8
XFILLER_38_544 VPWR VGND sg13g2_decap_8
XFILLER_25_205 VPWR VGND sg13g2_fill_1
XFILLER_26_739 VPWR VGND sg13g2_decap_8
XFILLER_33_271 VPWR VGND sg13g2_decap_8
XFILLER_34_783 VPWR VGND sg13g2_decap_8
XFILLER_21_444 VPWR VGND sg13g2_decap_8
XFILLER_22_956 VPWR VGND sg13g2_decap_8
XFILLER_0_315 VPWR VGND sg13g2_decap_8
XFILLER_1_838 VPWR VGND sg13g2_decap_8
XFILLER_29_533 VPWR VGND sg13g2_decap_8
X_580_ net82 VGND VPWR _120_ DP_3.matrix\[63\] clknet_5_30__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_514 VPWR VGND sg13g2_decap_8
XFILLER_17_53 VPWR VGND sg13g2_decap_8
XFILLER_9_927 VPWR VGND sg13g2_decap_8
XFILLER_13_956 VPWR VGND sg13g2_decap_8
XFILLER_40_764 VPWR VGND sg13g2_decap_8
XFILLER_33_74 VPWR VGND sg13g2_decap_8
XFILLER_3_120 VPWR VGND sg13g2_decap_4
XFILLER_4_654 VPWR VGND sg13g2_decap_8
XFILLER_0_882 VPWR VGND sg13g2_decap_8
Xhold4 mac2.sum_lvl1_ff\[33\] VPWR VGND net28 sg13g2_dlygate4sd3_1
XFILLER_48_853 VPWR VGND sg13g2_decap_8
XFILLER_35_536 VPWR VGND sg13g2_decap_8
XFILLER_23_709 VPWR VGND sg13g2_decap_8
XFILLER_43_580 VPWR VGND sg13g2_decap_8
XFILLER_22_208 VPWR VGND sg13g2_decap_4
XFILLER_31_720 VPWR VGND sg13g2_decap_8
XFILLER_31_797 VPWR VGND sg13g2_decap_8
XFILLER_30_274 VPWR VGND sg13g2_decap_8
XFILLER_8_993 VPWR VGND sg13g2_decap_8
XFILLER_39_875 VPWR VGND sg13g2_decap_8
XFILLER_26_536 VPWR VGND sg13g2_decap_8
XFILLER_34_580 VPWR VGND sg13g2_decap_8
XFILLER_22_753 VPWR VGND sg13g2_decap_8
XFILLER_16_1028 VPWR VGND sg13g2_fill_1
XFILLER_21_285 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_1_635 VPWR VGND sg13g2_decap_8
XFILLER_49_639 VPWR VGND sg13g2_decap_8
XFILLER_48_105 VPWR VGND sg13g2_fill_2
XFILLER_0_189 VPWR VGND sg13g2_decap_8
XFILLER_28_63 VPWR VGND sg13g2_decap_8
XFILLER_29_363 VPWR VGND sg13g2_decap_8
XFILLER_45_856 VPWR VGND sg13g2_decap_8
XFILLER_44_311 VPWR VGND sg13g2_decap_8
X_563_ net76 VGND VPWR _103_ DP_2.matrix\[64\] clknet_5_21__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_388 VPWR VGND sg13g2_decap_8
X_494_ net68 VGND VPWR _067_ mac2.products_ff\[35\] clknet_5_10__leaf_clk sg13g2_dfrbpq_1
XFILLER_13_753 VPWR VGND sg13g2_decap_8
XFILLER_9_724 VPWR VGND sg13g2_decap_8
XFILLER_40_561 VPWR VGND sg13g2_decap_8
XFILLER_5_941 VPWR VGND sg13g2_decap_8
XFILLER_5_67 VPWR VGND sg13g2_decap_8
XFILLER_48_650 VPWR VGND sg13g2_decap_8
XFILLER_10_4 VPWR VGND sg13g2_decap_8
XFILLER_35_333 VPWR VGND sg13g2_decap_8
XFILLER_36_856 VPWR VGND sg13g2_decap_8
XFILLER_23_528 VPWR VGND sg13g2_decap_8
XFILLER_31_594 VPWR VGND sg13g2_decap_8
XFILLER_8_790 VPWR VGND sg13g2_decap_8
XFILLER_39_672 VPWR VGND sg13g2_decap_8
XFILLER_27_834 VPWR VGND sg13g2_decap_8
XFILLER_42_848 VPWR VGND sg13g2_decap_8
XFILLER_14_539 VPWR VGND sg13g2_decap_8
XFILLER_26_366 VPWR VGND sg13g2_decap_8
XFILLER_22_550 VPWR VGND sg13g2_decap_8
XFILLER_14_76 VPWR VGND sg13g2_decap_8
XFILLER_10_767 VPWR VGND sg13g2_decap_8
XFILLER_5_259 VPWR VGND sg13g2_fill_1
XFILLER_2_922 VPWR VGND sg13g2_decap_8
XFILLER_1_432 VPWR VGND sg13g2_decap_8
XFILLER_2_999 VPWR VGND sg13g2_decap_8
XFILLER_49_436 VPWR VGND sg13g2_decap_8
XFILLER_39_62 VPWR VGND sg13g2_decap_8
Xclkbuf_4_3_0_clk clknet_0_clk clknet_4_3_0_clk VPWR VGND sg13g2_buf_8
XFILLER_17_300 VPWR VGND sg13g2_decap_8
XFILLER_18_823 VPWR VGND sg13g2_decap_8
XFILLER_45_653 VPWR VGND sg13g2_decap_8
XFILLER_33_804 VPWR VGND sg13g2_decap_8
XFILLER_44_174 VPWR VGND sg13g2_decap_8
X_546_ net60 VGND VPWR _086_ DP_1.matrix\[72\] clknet_5_4__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_336 VPWR VGND sg13g2_decap_8
XFILLER_32_347 VPWR VGND sg13g2_fill_1
X_477_ net74 VGND VPWR net176 mac1.sum_lvl2_ff\[1\] clknet_5_19__leaf_clk sg13g2_dfrbpq_1
XFILLER_9_521 VPWR VGND sg13g2_fill_1
XFILLER_13_572 VPWR VGND sg13g2_fill_2
XFILLER_9_598 VPWR VGND sg13g2_decap_8
XFILLER_45_1010 VPWR VGND sg13g2_decap_8
XFILLER_4_270 VPWR VGND sg13g2_decap_4
XFILLER_28_609 VPWR VGND sg13g2_decap_8
XFILLER_24_804 VPWR VGND sg13g2_decap_8
XFILLER_36_653 VPWR VGND sg13g2_decap_8
XFILLER_23_303 VPWR VGND sg13g2_decap_8
XFILLER_35_196 VPWR VGND sg13g2_decap_8
XFILLER_46_417 VPWR VGND sg13g2_decap_8
XFILLER_18_119 VPWR VGND sg13g2_decap_8
XFILLER_27_631 VPWR VGND sg13g2_decap_8
XFILLER_39_491 VPWR VGND sg13g2_decap_4
X_400_ net160 _094_ VPWR VGND sg13g2_buf_1
XFILLER_26_163 VPWR VGND sg13g2_decap_8
X_331_ _193_ _192_ _037_ VPWR VGND sg13g2_xor2_1
XFILLER_42_645 VPWR VGND sg13g2_decap_8
XFILLER_14_314 VPWR VGND sg13g2_decap_4
XFILLER_15_848 VPWR VGND sg13g2_decap_8
XFILLER_25_53 VPWR VGND sg13g2_decap_8
XFILLER_23_870 VPWR VGND sg13g2_decap_8
XFILLER_30_829 VPWR VGND sg13g2_decap_8
X_262_ net2 _152_ _155_ VPWR VGND sg13g2_xnor2_1
XFILLER_41_177 VPWR VGND sg13g2_decap_4
XFILLER_10_564 VPWR VGND sg13g2_decap_8
XFILLER_6_535 VPWR VGND sg13g2_fill_2
XFILLER_6_524 VPWR VGND sg13g2_decap_8
XFILLER_6_568 VPWR VGND sg13g2_decap_8
XFILLER_29_1016 VPWR VGND sg13g2_decap_8
XFILLER_29_1027 VPWR VGND sg13g2_fill_2
XFILLER_49_233 VPWR VGND sg13g2_decap_8
XFILLER_2_796 VPWR VGND sg13g2_decap_8
XFILLER_2_46 VPWR VGND sg13g2_decap_8
XFILLER_38_929 VPWR VGND sg13g2_decap_8
XFILLER_18_620 VPWR VGND sg13g2_decap_8
XFILLER_37_439 VPWR VGND sg13g2_decap_8
XFILLER_46_984 VPWR VGND sg13g2_decap_8
XFILLER_45_450 VPWR VGND sg13g2_decap_8
XFILLER_33_601 VPWR VGND sg13g2_decap_8
XFILLER_18_697 VPWR VGND sg13g2_decap_8
XFILLER_32_122 VPWR VGND sg13g2_decap_8
X_529_ net60 VGND VPWR net172 mac2.total_sum\[2\] clknet_5_6__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_678 VPWR VGND sg13g2_decap_8
XFILLER_9_384 VPWR VGND sg13g2_fill_2
XFILLER_49_0 VPWR VGND sg13g2_decap_8
XFILLER_29_918 VPWR VGND sg13g2_decap_8
XFILLER_37_940 VPWR VGND sg13g2_decap_8
XFILLER_24_601 VPWR VGND sg13g2_decap_8
XFILLER_23_144 VPWR VGND sg13g2_decap_8
XFILLER_24_678 VPWR VGND sg13g2_decap_8
XFILLER_11_339 VPWR VGND sg13g2_decap_8
XFILLER_11_11 VPWR VGND sg13g2_decap_8
XFILLER_4_1018 VPWR VGND sg13g2_decap_8
XFILLER_19_406 VPWR VGND sg13g2_decap_8
XFILLER_19_417 VPWR VGND sg13g2_fill_2
XFILLER_28_973 VPWR VGND sg13g2_decap_8
XFILLER_14_111 VPWR VGND sg13g2_decap_8
XFILLER_15_645 VPWR VGND sg13g2_decap_8
XFILLER_43_965 VPWR VGND sg13g2_decap_8
XFILLER_42_442 VPWR VGND sg13g2_decap_8
XFILLER_30_626 VPWR VGND sg13g2_decap_8
X_314_ net136 mac2.sum_lvl1_ff\[16\] _032_ VPWR VGND sg13g2_xor2_1
XFILLER_11_851 VPWR VGND sg13g2_decap_8
X_245_ net132 net119 _064_ VPWR VGND sg13g2_and2_1
XFILLER_7_855 VPWR VGND sg13g2_decap_8
XFILLER_6_332 VPWR VGND sg13g2_decap_4
XFILLER_2_560 VPWR VGND sg13g2_fill_1
XFILLER_42_7 VPWR VGND sg13g2_decap_8
XFILLER_2_593 VPWR VGND sg13g2_decap_8
XFILLER_42_1002 VPWR VGND sg13g2_decap_8
XFILLER_38_726 VPWR VGND sg13g2_decap_8
XFILLER_19_951 VPWR VGND sg13g2_decap_8
XFILLER_18_461 VPWR VGND sg13g2_fill_1
XFILLER_37_258 VPWR VGND sg13g2_decap_8
XFILLER_46_781 VPWR VGND sg13g2_decap_8
XFILLER_34_965 VPWR VGND sg13g2_decap_8
XFILLER_20_114 VPWR VGND sg13g2_fill_1
XFILLER_21_659 VPWR VGND sg13g2_decap_8
XFILLER_20_158 VPWR VGND sg13g2_decap_8
XFILLER_29_715 VPWR VGND sg13g2_decap_8
XFILLER_43_217 VPWR VGND sg13g2_decap_8
XFILLER_25_921 VPWR VGND sg13g2_decap_8
XFILLER_36_280 VPWR VGND sg13g2_fill_2
XFILLER_24_453 VPWR VGND sg13g2_decap_8
XFILLER_25_998 VPWR VGND sg13g2_decap_8
XFILLER_40_946 VPWR VGND sg13g2_decap_8
XFILLER_8_608 VPWR VGND sg13g2_decap_8
XFILLER_12_648 VPWR VGND sg13g2_decap_8
XFILLER_11_158 VPWR VGND sg13g2_fill_1
XFILLER_22_32 VPWR VGND sg13g2_decap_4
XFILLER_4_836 VPWR VGND sg13g2_decap_8
XFILLER_3_313 VPWR VGND sg13g2_decap_8
XFILLER_3_368 VPWR VGND sg13g2_decap_8
XFILLER_26_1019 VPWR VGND sg13g2_decap_8
XFILLER_19_214 VPWR VGND sg13g2_decap_8
XFILLER_47_567 VPWR VGND sg13g2_decap_8
XFILLER_28_770 VPWR VGND sg13g2_decap_8
XFILLER_35_718 VPWR VGND sg13g2_decap_8
XFILLER_16_921 VPWR VGND sg13g2_decap_8
XFILLER_34_217 VPWR VGND sg13g2_decap_8
XFILLER_43_762 VPWR VGND sg13g2_decap_8
Xclkbuf_5_21__f_clk clknet_4_10_0_clk clknet_5_21__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_15_431 VPWR VGND sg13g2_decap_8
XFILLER_31_902 VPWR VGND sg13g2_decap_8
XFILLER_16_998 VPWR VGND sg13g2_decap_8
XFILLER_31_979 VPWR VGND sg13g2_decap_8
XFILLER_8_67 VPWR VGND sg13g2_decap_8
XFILLER_7_652 VPWR VGND sg13g2_decap_8
X_228_ net127 net140 _038_ VPWR VGND sg13g2_and2_1
XFILLER_10_180 VPWR VGND sg13g2_decap_4
XFILLER_38_523 VPWR VGND sg13g2_decap_8
XFILLER_26_718 VPWR VGND sg13g2_decap_8
XFILLER_34_762 VPWR VGND sg13g2_decap_8
XFILLER_22_935 VPWR VGND sg13g2_decap_8
XFILLER_33_250 VPWR VGND sg13g2_decap_8
XFILLER_30_990 VPWR VGND sg13g2_decap_8
XFILLER_1_817 VPWR VGND sg13g2_decap_8
XFILLER_48_309 VPWR VGND sg13g2_decap_8
XFILLER_17_21 VPWR VGND sg13g2_decap_8
XFILLER_29_589 VPWR VGND sg13g2_decap_8
XFILLER_13_935 VPWR VGND sg13g2_decap_8
XFILLER_24_250 VPWR VGND sg13g2_decap_8
XFILLER_25_795 VPWR VGND sg13g2_decap_8
XFILLER_9_906 VPWR VGND sg13g2_decap_8
XFILLER_12_434 VPWR VGND sg13g2_decap_8
XFILLER_24_283 VPWR VGND sg13g2_decap_8
XFILLER_33_31 VPWR VGND sg13g2_decap_4
XFILLER_40_743 VPWR VGND sg13g2_decap_8
XFILLER_32_1012 VPWR VGND sg13g2_decap_8
XFILLER_33_53 VPWR VGND sg13g2_decap_8
XFILLER_8_449 VPWR VGND sg13g2_decap_8
XFILLER_4_633 VPWR VGND sg13g2_decap_8
XFILLER_0_861 VPWR VGND sg13g2_decap_8
XFILLER_39_309 VPWR VGND sg13g2_fill_2
XFILLER_48_832 VPWR VGND sg13g2_decap_8
Xhold5 mac2.products_ff\[137\] VPWR VGND net29 sg13g2_dlygate4sd3_1
XFILLER_47_353 VPWR VGND sg13g2_decap_4
XFILLER_47_375 VPWR VGND sg13g2_decap_4
XFILLER_35_515 VPWR VGND sg13g2_decap_8
XFILLER_16_795 VPWR VGND sg13g2_decap_8
XFILLER_30_253 VPWR VGND sg13g2_decap_8
XFILLER_31_776 VPWR VGND sg13g2_decap_8
XFILLER_8_972 VPWR VGND sg13g2_decap_8
XFILLER_31_0 VPWR VGND sg13g2_decap_8
XFILLER_39_854 VPWR VGND sg13g2_decap_8
XFILLER_26_515 VPWR VGND sg13g2_decap_8
XFILLER_38_375 VPWR VGND sg13g2_decap_4
XFILLER_22_732 VPWR VGND sg13g2_decap_8
XFILLER_21_264 VPWR VGND sg13g2_decap_8
XFILLER_10_949 VPWR VGND sg13g2_decap_8
XFILLER_1_614 VPWR VGND sg13g2_decap_8
XFILLER_49_618 VPWR VGND sg13g2_decap_8
XFILLER_0_168 VPWR VGND sg13g2_decap_8
XFILLER_29_320 VPWR VGND sg13g2_fill_2
XFILLER_45_835 VPWR VGND sg13g2_decap_8
X_562_ net75 VGND VPWR _102_ DP_2.matrix\[63\] clknet_5_21__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_559 VPWR VGND sg13g2_fill_2
XFILLER_44_367 VPWR VGND sg13g2_decap_8
XFILLER_32_529 VPWR VGND sg13g2_decap_8
X_493_ net70 VGND VPWR _066_ mac2.products_ff\[34\] clknet_5_11__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_63 VPWR VGND sg13g2_decap_4
XFILLER_13_732 VPWR VGND sg13g2_decap_8
XFILLER_25_592 VPWR VGND sg13g2_decap_8
XFILLER_9_703 VPWR VGND sg13g2_decap_8
XFILLER_12_253 VPWR VGND sg13g2_decap_4
XFILLER_40_540 VPWR VGND sg13g2_decap_8
XFILLER_5_920 VPWR VGND sg13g2_decap_8
XFILLER_5_46 VPWR VGND sg13g2_decap_8
XFILLER_5_997 VPWR VGND sg13g2_decap_8
XFILLER_4_485 VPWR VGND sg13g2_decap_8
XFILLER_39_117 VPWR VGND sg13g2_decap_8
XFILLER_35_301 VPWR VGND sg13g2_fill_2
XFILLER_35_312 VPWR VGND sg13g2_decap_8
XFILLER_36_835 VPWR VGND sg13g2_decap_8
XFILLER_23_507 VPWR VGND sg13g2_decap_8
XFILLER_35_389 VPWR VGND sg13g2_decap_8
XFILLER_31_573 VPWR VGND sg13g2_decap_8
XFILLER_39_651 VPWR VGND sg13g2_decap_8
XFILLER_27_813 VPWR VGND sg13g2_decap_8
XFILLER_26_345 VPWR VGND sg13g2_decap_8
XFILLER_42_827 VPWR VGND sg13g2_decap_8
XFILLER_14_518 VPWR VGND sg13g2_decap_8
XFILLER_14_11 VPWR VGND sg13g2_decap_8
XFILLER_41_348 VPWR VGND sg13g2_decap_8
XFILLER_14_33 VPWR VGND sg13g2_fill_1
XFILLER_14_55 VPWR VGND sg13g2_decap_8
XFILLER_10_746 VPWR VGND sg13g2_decap_8
XFILLER_6_739 VPWR VGND sg13g2_decap_8
XFILLER_30_21 VPWR VGND sg13g2_decap_8
XFILLER_5_238 VPWR VGND sg13g2_decap_8
XFILLER_2_901 VPWR VGND sg13g2_decap_8
XFILLER_1_411 VPWR VGND sg13g2_decap_8
XFILLER_49_415 VPWR VGND sg13g2_decap_8
XFILLER_7_1016 VPWR VGND sg13g2_decap_8
XFILLER_2_978 VPWR VGND sg13g2_decap_8
XFILLER_7_1027 VPWR VGND sg13g2_fill_2
XFILLER_1_488 VPWR VGND sg13g2_decap_8
XFILLER_18_802 VPWR VGND sg13g2_decap_8
XFILLER_39_96 VPWR VGND sg13g2_decap_8
XFILLER_29_172 VPWR VGND sg13g2_decap_8
XFILLER_45_632 VPWR VGND sg13g2_decap_8
XFILLER_18_879 VPWR VGND sg13g2_decap_8
XFILLER_44_153 VPWR VGND sg13g2_decap_8
X_545_ net76 VGND VPWR _085_ DP_1.matrix\[64\] clknet_5_21__leaf_clk sg13g2_dfrbpq_1
X_476_ net73 VGND VPWR net146 mac1.sum_lvl2_ff\[0\] clknet_5_19__leaf_clk sg13g2_dfrbpq_1
XFILLER_13_562 VPWR VGND sg13g2_fill_1
XFILLER_9_577 VPWR VGND sg13g2_decap_8
XFILLER_5_794 VPWR VGND sg13g2_decap_8
XFILLER_49_982 VPWR VGND sg13g2_decap_8
XFILLER_36_632 VPWR VGND sg13g2_decap_8
XFILLER_35_175 VPWR VGND sg13g2_decap_8
XFILLER_23_359 VPWR VGND sg13g2_decap_8
XFILLER_32_893 VPWR VGND sg13g2_decap_8
XFILLER_27_610 VPWR VGND sg13g2_decap_8
XFILLER_15_827 VPWR VGND sg13g2_decap_8
Xclkbuf_5_2__f_clk clknet_4_1_0_clk clknet_5_2__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_27_687 VPWR VGND sg13g2_decap_8
XFILLER_42_624 VPWR VGND sg13g2_decap_8
X_330_ _193_ net156 net52 VPWR VGND sg13g2_nand2_1
XFILLER_25_32 VPWR VGND sg13g2_decap_8
XFILLER_30_808 VPWR VGND sg13g2_decap_8
XFILLER_41_156 VPWR VGND sg13g2_decap_8
X_261_ mac2.total_sum\[1\] mac1.total_sum\[1\] _155_ VPWR VGND sg13g2_xor2_1
XFILLER_10_543 VPWR VGND sg13g2_decap_8
XFILLER_22_381 VPWR VGND sg13g2_decap_8
XFILLER_6_503 VPWR VGND sg13g2_decap_8
XFILLER_41_75 VPWR VGND sg13g2_decap_8
XFILLER_2_775 VPWR VGND sg13g2_decap_8
XFILLER_49_212 VPWR VGND sg13g2_decap_8
XFILLER_1_285 VPWR VGND sg13g2_decap_8
XFILLER_2_25 VPWR VGND sg13g2_decap_8
XFILLER_38_908 VPWR VGND sg13g2_decap_8
XFILLER_49_289 VPWR VGND sg13g2_decap_8
XFILLER_37_418 VPWR VGND sg13g2_decap_8
XFILLER_46_963 VPWR VGND sg13g2_decap_8
XFILLER_18_676 VPWR VGND sg13g2_decap_8
XFILLER_32_101 VPWR VGND sg13g2_decap_8
X_528_ net60 VGND VPWR net202 mac2.total_sum\[1\] clknet_5_6__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_657 VPWR VGND sg13g2_decap_8
XFILLER_14_882 VPWR VGND sg13g2_decap_8
X_459_ net77 VGND VPWR _053_ mac1.products_ff\[86\] clknet_5_29__leaf_clk sg13g2_dfrbpq_1
XFILLER_5_591 VPWR VGND sg13g2_decap_8
XFILLER_28_418 VPWR VGND sg13g2_decap_8
XFILLER_37_996 VPWR VGND sg13g2_decap_8
XFILLER_23_101 VPWR VGND sg13g2_decap_8
XFILLER_24_657 VPWR VGND sg13g2_decap_8
XFILLER_11_318 VPWR VGND sg13g2_decap_8
XFILLER_32_690 VPWR VGND sg13g2_decap_8
XFILLER_20_885 VPWR VGND sg13g2_decap_8
Xclkbuf_4_2_0_clk clknet_0_clk clknet_4_2_0_clk VPWR VGND sg13g2_buf_8
XFILLER_3_517 VPWR VGND sg13g2_decap_8
XFILLER_11_67 VPWR VGND sg13g2_fill_2
XFILLER_46_215 VPWR VGND sg13g2_decap_4
XFILLER_47_749 VPWR VGND sg13g2_decap_8
XFILLER_28_952 VPWR VGND sg13g2_decap_8
XFILLER_46_259 VPWR VGND sg13g2_decap_8
XFILLER_43_944 VPWR VGND sg13g2_decap_8
XFILLER_42_421 VPWR VGND sg13g2_decap_8
XFILLER_15_624 VPWR VGND sg13g2_decap_8
XFILLER_27_473 VPWR VGND sg13g2_decap_8
XFILLER_36_86 VPWR VGND sg13g2_decap_8
XFILLER_30_605 VPWR VGND sg13g2_decap_8
XFILLER_42_498 VPWR VGND sg13g2_decap_8
X_313_ _033_ _182_ _183_ VPWR VGND sg13g2_xnor2_1
XFILLER_11_830 VPWR VGND sg13g2_decap_8
X_244_ net144 net143 _062_ VPWR VGND sg13g2_and2_1
XFILLER_7_834 VPWR VGND sg13g2_decap_8
XFILLER_6_311 VPWR VGND sg13g2_decap_8
XFILLER_10_373 VPWR VGND sg13g2_decap_8
XFILLER_6_377 VPWR VGND sg13g2_decap_8
XFILLER_2_572 VPWR VGND sg13g2_decap_8
XFILLER_35_7 VPWR VGND sg13g2_decap_8
XFILLER_38_705 VPWR VGND sg13g2_decap_8
XFILLER_19_930 VPWR VGND sg13g2_decap_8
XFILLER_37_237 VPWR VGND sg13g2_decap_8
XFILLER_46_760 VPWR VGND sg13g2_decap_8
XFILLER_34_944 VPWR VGND sg13g2_decap_8
XFILLER_45_292 VPWR VGND sg13g2_decap_8
XFILLER_21_638 VPWR VGND sg13g2_decap_8
XFILLER_33_465 VPWR VGND sg13g2_decap_4
XFILLER_20_137 VPWR VGND sg13g2_decap_8
XFILLER_25_900 VPWR VGND sg13g2_decap_8
XFILLER_37_793 VPWR VGND sg13g2_decap_8
XFILLER_24_432 VPWR VGND sg13g2_decap_8
XFILLER_25_977 VPWR VGND sg13g2_decap_8
XFILLER_12_627 VPWR VGND sg13g2_decap_8
XFILLER_40_925 VPWR VGND sg13g2_decap_8
XFILLER_7_119 VPWR VGND sg13g2_decap_8
XFILLER_22_11 VPWR VGND sg13g2_decap_8
XFILLER_20_682 VPWR VGND sg13g2_decap_8
XFILLER_4_815 VPWR VGND sg13g2_decap_8
XFILLER_47_546 VPWR VGND sg13g2_decap_8
XFILLER_47_63 VPWR VGND sg13g2_decap_4
XFILLER_47_85 VPWR VGND sg13g2_decap_8
XFILLER_16_900 VPWR VGND sg13g2_decap_8
XFILLER_15_410 VPWR VGND sg13g2_decap_8
XFILLER_43_741 VPWR VGND sg13g2_decap_8
XFILLER_16_977 VPWR VGND sg13g2_decap_8
XFILLER_42_262 VPWR VGND sg13g2_decap_8
XFILLER_15_487 VPWR VGND sg13g2_decap_8
XFILLER_42_295 VPWR VGND sg13g2_decap_8
XFILLER_31_958 VPWR VGND sg13g2_decap_8
XFILLER_8_46 VPWR VGND sg13g2_decap_8
XFILLER_30_479 VPWR VGND sg13g2_decap_8
XFILLER_7_631 VPWR VGND sg13g2_decap_8
X_227_ net156 net131 _036_ VPWR VGND sg13g2_and2_1
XFILLER_6_185 VPWR VGND sg13g2_decap_8
XFILLER_6_163 VPWR VGND sg13g2_decap_8
XFILLER_3_881 VPWR VGND sg13g2_decap_8
XFILLER_38_502 VPWR VGND sg13g2_decap_8
XFILLER_38_579 VPWR VGND sg13g2_decap_8
XFILLER_25_229 VPWR VGND sg13g2_decap_8
XFILLER_18_292 VPWR VGND sg13g2_decap_8
XFILLER_34_741 VPWR VGND sg13g2_decap_8
XFILLER_22_914 VPWR VGND sg13g2_decap_8
XFILLER_21_479 VPWR VGND sg13g2_decap_8
XFILLER_17_719 VPWR VGND sg13g2_decap_8
XFILLER_29_568 VPWR VGND sg13g2_decap_8
XFILLER_44_549 VPWR VGND sg13g2_decap_8
XFILLER_17_88 VPWR VGND sg13g2_decap_8
XFILLER_37_590 VPWR VGND sg13g2_decap_8
XFILLER_13_914 VPWR VGND sg13g2_decap_8
XFILLER_25_774 VPWR VGND sg13g2_decap_8
XFILLER_33_21 VPWR VGND sg13g2_decap_4
XFILLER_40_722 VPWR VGND sg13g2_decap_8
XFILLER_8_428 VPWR VGND sg13g2_decap_8
XFILLER_40_799 VPWR VGND sg13g2_decap_8
XFILLER_4_612 VPWR VGND sg13g2_decap_8
XFILLER_4_689 VPWR VGND sg13g2_decap_8
XFILLER_3_166 VPWR VGND sg13g2_decap_8
XFILLER_0_840 VPWR VGND sg13g2_decap_8
XFILLER_48_811 VPWR VGND sg13g2_decap_8
Xhold6 mac1.sum_lvl2_ff\[9\] VPWR VGND net30 sg13g2_dlygate4sd3_1
XFILLER_48_888 VPWR VGND sg13g2_decap_8
XFILLER_47_332 VPWR VGND sg13g2_decap_8
XFILLER_16_774 VPWR VGND sg13g2_decap_8
XFILLER_15_273 VPWR VGND sg13g2_decap_8
XFILLER_30_232 VPWR VGND sg13g2_decap_8
XFILLER_31_755 VPWR VGND sg13g2_decap_8
XFILLER_12_991 VPWR VGND sg13g2_decap_8
XFILLER_8_951 VPWR VGND sg13g2_decap_8
XFILLER_7_450 VPWR VGND sg13g2_decap_8
XFILLER_39_833 VPWR VGND sg13g2_decap_8
XFILLER_38_354 VPWR VGND sg13g2_decap_8
XFILLER_0_1022 VPWR VGND sg13g2_decap_8
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_22_711 VPWR VGND sg13g2_decap_8
XFILLER_41_519 VPWR VGND sg13g2_decap_8
XFILLER_10_928 VPWR VGND sg13g2_decap_8
XFILLER_16_1019 VPWR VGND sg13g2_decap_8
XFILLER_22_788 VPWR VGND sg13g2_decap_8
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_45_814 VPWR VGND sg13g2_decap_8
X_561_ net74 VGND VPWR _101_ DP_2.matrix\[55\] clknet_5_17__leaf_clk sg13g2_dfrbpq_1
XFILLER_28_98 VPWR VGND sg13g2_decap_8
XFILLER_44_346 VPWR VGND sg13g2_fill_2
XFILLER_44_42 VPWR VGND sg13g2_decap_8
XFILLER_13_711 VPWR VGND sg13g2_decap_8
X_492_ net69 VGND VPWR _041_ mac2.products_ff\[18\] clknet_5_2__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_508 VPWR VGND sg13g2_decap_8
XFILLER_25_571 VPWR VGND sg13g2_decap_8
XFILLER_8_203 VPWR VGND sg13g2_fill_2
XFILLER_12_232 VPWR VGND sg13g2_decap_8
XFILLER_9_759 VPWR VGND sg13g2_decap_8
XFILLER_12_287 VPWR VGND sg13g2_decap_8
XFILLER_13_788 VPWR VGND sg13g2_decap_8
XFILLER_40_596 VPWR VGND sg13g2_decap_8
XFILLER_5_976 VPWR VGND sg13g2_decap_8
XFILLER_5_25 VPWR VGND sg13g2_decap_8
XFILLER_4_464 VPWR VGND sg13g2_decap_8
XFILLER_48_685 VPWR VGND sg13g2_decap_8
XFILLER_47_162 VPWR VGND sg13g2_decap_4
XFILLER_36_814 VPWR VGND sg13g2_decap_8
XFILLER_47_195 VPWR VGND sg13g2_decap_8
XFILLER_39_1008 VPWR VGND sg13g2_decap_8
XFILLER_16_560 VPWR VGND sg13g2_fill_1
XFILLER_35_368 VPWR VGND sg13g2_decap_8
XFILLER_31_552 VPWR VGND sg13g2_decap_8
XFILLER_22_1012 VPWR VGND sg13g2_decap_8
XFILLER_39_630 VPWR VGND sg13g2_decap_8
XFILLER_26_324 VPWR VGND sg13g2_decap_8
XFILLER_27_869 VPWR VGND sg13g2_decap_8
XFILLER_38_184 VPWR VGND sg13g2_decap_8
XFILLER_42_806 VPWR VGND sg13g2_decap_8
XFILLER_41_327 VPWR VGND sg13g2_decap_8
XFILLER_10_725 VPWR VGND sg13g2_decap_8
XFILLER_22_585 VPWR VGND sg13g2_decap_8
XFILLER_6_718 VPWR VGND sg13g2_decap_8
XFILLER_5_217 VPWR VGND sg13g2_decap_8
XFILLER_30_33 VPWR VGND sg13g2_fill_2
XFILLER_30_77 VPWR VGND sg13g2_decap_8
XFILLER_2_957 VPWR VGND sg13g2_decap_8
XFILLER_1_467 VPWR VGND sg13g2_decap_8
XFILLER_45_611 VPWR VGND sg13g2_decap_8
XFILLER_29_151 VPWR VGND sg13g2_decap_8
XFILLER_17_335 VPWR VGND sg13g2_decap_8
XFILLER_18_858 VPWR VGND sg13g2_decap_8
XFILLER_29_195 VPWR VGND sg13g2_fill_2
XFILLER_45_688 VPWR VGND sg13g2_decap_8
XFILLER_44_132 VPWR VGND sg13g2_decap_8
X_544_ net76 VGND VPWR _084_ DP_1.matrix\[63\] clknet_5_21__leaf_clk sg13g2_dfrbpq_1
X_475_ net64 VGND VPWR net33 mac1.sum_lvl1_ff\[33\] clknet_5_5__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_316 VPWR VGND sg13g2_decap_8
XFILLER_33_839 VPWR VGND sg13g2_decap_8
XFILLER_13_541 VPWR VGND sg13g2_decap_8
XFILLER_13_552 VPWR VGND sg13g2_fill_2
XFILLER_9_512 VPWR VGND sg13g2_decap_8
XFILLER_13_585 VPWR VGND sg13g2_decap_8
XFILLER_41_883 VPWR VGND sg13g2_decap_8
XFILLER_9_556 VPWR VGND sg13g2_decap_8
XFILLER_5_773 VPWR VGND sg13g2_decap_8
XFILLER_49_961 VPWR VGND sg13g2_decap_8
XFILLER_36_611 VPWR VGND sg13g2_decap_8
XFILLER_48_482 VPWR VGND sg13g2_decap_8
XFILLER_35_110 VPWR VGND sg13g2_decap_8
XFILLER_35_154 VPWR VGND sg13g2_decap_8
XFILLER_36_688 VPWR VGND sg13g2_decap_8
XFILLER_17_880 VPWR VGND sg13g2_decap_8
XFILLER_23_338 VPWR VGND sg13g2_decap_8
XFILLER_24_839 VPWR VGND sg13g2_decap_8
XFILLER_31_371 VPWR VGND sg13g2_decap_8
XFILLER_32_872 VPWR VGND sg13g2_decap_8
XFILLER_2_209 VPWR VGND sg13g2_decap_8
XFILLER_42_603 VPWR VGND sg13g2_decap_8
XFILLER_15_806 VPWR VGND sg13g2_decap_8
XFILLER_25_11 VPWR VGND sg13g2_decap_8
XFILLER_27_666 VPWR VGND sg13g2_decap_8
XFILLER_26_198 VPWR VGND sg13g2_decap_8
XFILLER_14_349 VPWR VGND sg13g2_decap_8
XFILLER_41_135 VPWR VGND sg13g2_decap_8
X_260_ mac1.total_sum\[1\] mac2.total_sum\[1\] _154_ VPWR VGND sg13g2_nor2_1
XFILLER_22_360 VPWR VGND sg13g2_decap_8
XFILLER_10_522 VPWR VGND sg13g2_decap_8
XFILLER_41_54 VPWR VGND sg13g2_decap_8
XFILLER_10_599 VPWR VGND sg13g2_decap_8
XFILLER_2_754 VPWR VGND sg13g2_decap_8
XFILLER_1_264 VPWR VGND sg13g2_decap_8
XFILLER_49_268 VPWR VGND sg13g2_decap_8
XFILLER_46_942 VPWR VGND sg13g2_decap_8
XFILLER_17_143 VPWR VGND sg13g2_decap_8
XFILLER_18_655 VPWR VGND sg13g2_decap_8
XFILLER_45_485 VPWR VGND sg13g2_decap_8
X_527_ net60 VGND VPWR net116 mac2.total_sum\[0\] clknet_5_6__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_636 VPWR VGND sg13g2_decap_8
XFILLER_14_861 VPWR VGND sg13g2_decap_8
X_458_ net78 VGND VPWR _052_ mac1.products_ff\[85\] clknet_5_22__leaf_clk sg13g2_dfrbpq_1
XFILLER_20_319 VPWR VGND sg13g2_decap_8
XFILLER_32_157 VPWR VGND sg13g2_decap_8
X_389_ net54 _083_ VPWR VGND sg13g2_buf_1
XFILLER_13_382 VPWR VGND sg13g2_decap_8
XFILLER_41_680 VPWR VGND sg13g2_decap_8
XFILLER_36_441 VPWR VGND sg13g2_decap_8
XFILLER_36_463 VPWR VGND sg13g2_decap_4
XFILLER_37_975 VPWR VGND sg13g2_decap_8
XFILLER_24_636 VPWR VGND sg13g2_decap_8
XFILLER_36_485 VPWR VGND sg13g2_decap_8
XFILLER_12_809 VPWR VGND sg13g2_decap_8
XFILLER_20_864 VPWR VGND sg13g2_decap_8
XFILLER_11_79 VPWR VGND sg13g2_decap_8
XFILLER_47_728 VPWR VGND sg13g2_decap_8
XFILLER_46_238 VPWR VGND sg13g2_decap_8
XFILLER_28_931 VPWR VGND sg13g2_decap_8
XFILLER_15_603 VPWR VGND sg13g2_decap_8
XFILLER_27_452 VPWR VGND sg13g2_decap_8
XFILLER_43_923 VPWR VGND sg13g2_decap_8
XFILLER_42_400 VPWR VGND sg13g2_decap_8
XFILLER_36_65 VPWR VGND sg13g2_decap_8
XFILLER_14_146 VPWR VGND sg13g2_decap_8
XFILLER_42_477 VPWR VGND sg13g2_decap_8
X_312_ mac2.sum_lvl1_ff\[25\] mac2.sum_lvl1_ff\[17\] _183_ VPWR VGND sg13g2_xor2_1
X_243_ net125 net158 _060_ VPWR VGND sg13g2_and2_1
XFILLER_10_352 VPWR VGND sg13g2_decap_8
XFILLER_7_813 VPWR VGND sg13g2_decap_8
XFILLER_11_886 VPWR VGND sg13g2_decap_8
XFILLER_22_190 VPWR VGND sg13g2_fill_1
XFILLER_6_356 VPWR VGND sg13g2_decap_8
XFILLER_37_205 VPWR VGND sg13g2_decap_8
XFILLER_18_452 VPWR VGND sg13g2_decap_8
XFILLER_19_986 VPWR VGND sg13g2_decap_8
XFILLER_45_271 VPWR VGND sg13g2_decap_8
XFILLER_34_923 VPWR VGND sg13g2_decap_8
XFILLER_21_617 VPWR VGND sg13g2_decap_8
XFILLER_9_172 VPWR VGND sg13g2_decap_8
XFILLER_24_411 VPWR VGND sg13g2_decap_8
XFILLER_37_772 VPWR VGND sg13g2_decap_8
XFILLER_25_956 VPWR VGND sg13g2_decap_8
XFILLER_40_904 VPWR VGND sg13g2_decap_8
XFILLER_12_606 VPWR VGND sg13g2_decap_8
XFILLER_19_1028 VPWR VGND sg13g2_fill_1
XFILLER_20_661 VPWR VGND sg13g2_decap_8
XFILLER_22_89 VPWR VGND sg13g2_decap_8
XFILLER_47_525 VPWR VGND sg13g2_decap_8
XFILLER_47_42 VPWR VGND sg13g2_decap_8
XFILLER_19_249 VPWR VGND sg13g2_decap_8
XFILLER_43_720 VPWR VGND sg13g2_decap_8
XFILLER_16_956 VPWR VGND sg13g2_decap_8
XFILLER_27_282 VPWR VGND sg13g2_decap_8
XFILLER_42_241 VPWR VGND sg13g2_decap_8
XFILLER_15_466 VPWR VGND sg13g2_decap_8
XFILLER_31_937 VPWR VGND sg13g2_decap_8
XFILLER_43_797 VPWR VGND sg13g2_decap_8
XFILLER_30_425 VPWR VGND sg13g2_decap_8
XFILLER_30_447 VPWR VGND sg13g2_fill_2
XFILLER_8_25 VPWR VGND sg13g2_decap_8
XFILLER_30_458 VPWR VGND sg13g2_decap_8
X_226_ net141 net121 _034_ VPWR VGND sg13g2_and2_1
XFILLER_7_610 VPWR VGND sg13g2_decap_8
XFILLER_11_683 VPWR VGND sg13g2_decap_8
XFILLER_6_131 VPWR VGND sg13g2_decap_8
XFILLER_6_120 VPWR VGND sg13g2_fill_2
XFILLER_7_687 VPWR VGND sg13g2_decap_8
XFILLER_3_860 VPWR VGND sg13g2_decap_8
XFILLER_2_370 VPWR VGND sg13g2_decap_4
XFILLER_26_4 VPWR VGND sg13g2_decap_8
Xclkbuf_4_1_0_clk clknet_0_clk clknet_4_1_0_clk VPWR VGND sg13g2_buf_8
XFILLER_38_558 VPWR VGND sg13g2_decap_8
XFILLER_19_783 VPWR VGND sg13g2_decap_8
XFILLER_34_720 VPWR VGND sg13g2_decap_8
XFILLER_18_271 VPWR VGND sg13g2_decap_8
XFILLER_33_285 VPWR VGND sg13g2_decap_8
XFILLER_34_797 VPWR VGND sg13g2_decap_8
XFILLER_21_458 VPWR VGND sg13g2_decap_8
XFILLER_0_329 VPWR VGND sg13g2_decap_8
XFILLER_29_547 VPWR VGND sg13g2_decap_8
XFILLER_44_528 VPWR VGND sg13g2_decap_8
XFILLER_16_208 VPWR VGND sg13g2_decap_8
XFILLER_17_67 VPWR VGND sg13g2_decap_8
XFILLER_25_753 VPWR VGND sg13g2_decap_8
XFILLER_40_701 VPWR VGND sg13g2_decap_8
XFILLER_40_778 VPWR VGND sg13g2_decap_8
XFILLER_21_981 VPWR VGND sg13g2_decap_8
XFILLER_33_88 VPWR VGND sg13g2_decap_8
XFILLER_3_101 VPWR VGND sg13g2_decap_4
XFILLER_4_668 VPWR VGND sg13g2_decap_8
XFILLER_3_145 VPWR VGND sg13g2_decap_8
XFILLER_47_311 VPWR VGND sg13g2_decap_8
Xhold7 mac1.sum_lvl1_ff\[33\] VPWR VGND net31 sg13g2_dlygate4sd3_1
XFILLER_0_896 VPWR VGND sg13g2_decap_8
XFILLER_48_867 VPWR VGND sg13g2_decap_8
XFILLER_15_252 VPWR VGND sg13g2_decap_8
XFILLER_16_753 VPWR VGND sg13g2_decap_8
XFILLER_43_594 VPWR VGND sg13g2_decap_8
XFILLER_30_211 VPWR VGND sg13g2_decap_8
XFILLER_31_734 VPWR VGND sg13g2_decap_8
XFILLER_8_930 VPWR VGND sg13g2_decap_8
XFILLER_12_970 VPWR VGND sg13g2_decap_8
XFILLER_30_288 VPWR VGND sg13g2_decap_8
XFILLER_7_484 VPWR VGND sg13g2_decap_8
XFILLER_48_1021 VPWR VGND sg13g2_decap_8
XFILLER_39_812 VPWR VGND sg13g2_decap_8
XFILLER_17_0 VPWR VGND sg13g2_decap_8
XFILLER_38_333 VPWR VGND sg13g2_decap_8
XFILLER_0_1001 VPWR VGND sg13g2_decap_8
XFILLER_39_889 VPWR VGND sg13g2_decap_8
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_19_580 VPWR VGND sg13g2_decap_8
XFILLER_38_399 VPWR VGND sg13g2_decap_8
XFILLER_34_594 VPWR VGND sg13g2_decap_8
XFILLER_10_907 VPWR VGND sg13g2_decap_8
XFILLER_22_767 VPWR VGND sg13g2_decap_8
XFILLER_21_299 VPWR VGND sg13g2_decap_8
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_1_649 VPWR VGND sg13g2_decap_8
XFILLER_28_11 VPWR VGND sg13g2_decap_8
XFILLER_28_33 VPWR VGND sg13g2_fill_2
XFILLER_29_322 VPWR VGND sg13g2_fill_1
X_560_ net73 VGND VPWR _100_ DP_2.matrix\[54\] clknet_5_17__leaf_clk sg13g2_dfrbpq_1
XFILLER_28_77 VPWR VGND sg13g2_decap_8
XFILLER_29_377 VPWR VGND sg13g2_decap_8
XFILLER_44_325 VPWR VGND sg13g2_decap_8
XFILLER_44_21 VPWR VGND sg13g2_decap_8
X_491_ net69 VGND VPWR _040_ mac2.products_ff\[17\] clknet_5_3__leaf_clk sg13g2_dfrbpq_1
XFILLER_25_550 VPWR VGND sg13g2_decap_8
XFILLER_44_87 VPWR VGND sg13g2_fill_2
XFILLER_44_76 VPWR VGND sg13g2_fill_2
XFILLER_44_98 VPWR VGND sg13g2_decap_4
XFILLER_13_767 VPWR VGND sg13g2_decap_8
XFILLER_9_738 VPWR VGND sg13g2_decap_8
XFILLER_12_266 VPWR VGND sg13g2_decap_8
XFILLER_40_575 VPWR VGND sg13g2_decap_8
XFILLER_8_248 VPWR VGND sg13g2_decap_8
XFILLER_5_955 VPWR VGND sg13g2_decap_8
XFILLER_4_443 VPWR VGND sg13g2_decap_8
XFILLER_0_693 VPWR VGND sg13g2_decap_8
XFILLER_48_664 VPWR VGND sg13g2_decap_8
XFILLER_47_141 VPWR VGND sg13g2_decap_8
XFILLER_35_347 VPWR VGND sg13g2_decap_8
XFILLER_44_892 VPWR VGND sg13g2_decap_8
XFILLER_31_531 VPWR VGND sg13g2_decap_8
XFILLER_26_303 VPWR VGND sg13g2_decap_8
XFILLER_38_152 VPWR VGND sg13g2_decap_4
XFILLER_39_686 VPWR VGND sg13g2_decap_8
XFILLER_27_848 VPWR VGND sg13g2_decap_8
XFILLER_10_704 VPWR VGND sg13g2_decap_8
XFILLER_22_564 VPWR VGND sg13g2_decap_8
XFILLER_30_56 VPWR VGND sg13g2_decap_8
XFILLER_2_936 VPWR VGND sg13g2_decap_8
XFILLER_1_446 VPWR VGND sg13g2_decap_8
XFILLER_39_21 VPWR VGND sg13g2_decap_8
XFILLER_39_32 VPWR VGND sg13g2_fill_2
XFILLER_17_314 VPWR VGND sg13g2_decap_8
XFILLER_18_837 VPWR VGND sg13g2_decap_8
XFILLER_45_667 VPWR VGND sg13g2_decap_8
X_543_ net73 VGND VPWR _083_ DP_1.matrix\[55\] clknet_5_17__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_818 VPWR VGND sg13g2_decap_8
XFILLER_44_188 VPWR VGND sg13g2_decap_8
X_474_ net61 VGND VPWR net27 mac1.sum_lvl1_ff\[32\] clknet_5_4__leaf_clk sg13g2_dfrbpq_1
XFILLER_38_1020 VPWR VGND sg13g2_decap_8
XFILLER_13_520 VPWR VGND sg13g2_decap_8
XFILLER_41_862 VPWR VGND sg13g2_decap_8
XFILLER_9_535 VPWR VGND sg13g2_decap_8
XFILLER_5_752 VPWR VGND sg13g2_decap_8
XFILLER_45_1024 VPWR VGND sg13g2_decap_4
Xclkbuf_5_27__f_clk clknet_4_13_0_clk clknet_5_27__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_49_940 VPWR VGND sg13g2_decap_8
XFILLER_0_490 VPWR VGND sg13g2_decap_8
XFILLER_48_461 VPWR VGND sg13g2_decap_8
XFILLER_24_818 VPWR VGND sg13g2_decap_8
XFILLER_35_144 VPWR VGND sg13g2_fill_1
XFILLER_36_667 VPWR VGND sg13g2_decap_8
XFILLER_23_317 VPWR VGND sg13g2_decap_8
XFILLER_16_380 VPWR VGND sg13g2_fill_1
XFILLER_32_851 VPWR VGND sg13g2_decap_8
XFILLER_31_350 VPWR VGND sg13g2_decap_8
XFILLER_31_394 VPWR VGND sg13g2_fill_2
XFILLER_39_461 VPWR VGND sg13g2_decap_8
XFILLER_27_645 VPWR VGND sg13g2_decap_8
XFILLER_39_472 VPWR VGND sg13g2_fill_2
XFILLER_26_122 VPWR VGND sg13g2_decap_8
XFILLER_26_177 VPWR VGND sg13g2_decap_8
XFILLER_42_659 VPWR VGND sg13g2_decap_8
XFILLER_25_67 VPWR VGND sg13g2_decap_8
XFILLER_10_501 VPWR VGND sg13g2_decap_8
XFILLER_23_884 VPWR VGND sg13g2_decap_8
XFILLER_41_11 VPWR VGND sg13g2_fill_2
XFILLER_10_578 VPWR VGND sg13g2_decap_8
XFILLER_2_733 VPWR VGND sg13g2_decap_8
XFILLER_1_243 VPWR VGND sg13g2_decap_8
XFILLER_49_247 VPWR VGND sg13g2_decap_8
XFILLER_46_921 VPWR VGND sg13g2_decap_8
XFILLER_18_634 VPWR VGND sg13g2_decap_8
XFILLER_45_464 VPWR VGND sg13g2_decap_8
XFILLER_46_998 VPWR VGND sg13g2_decap_8
X_526_ net65 VGND VPWR net34 mac2.sum_lvl3_ff\[3\] clknet_5_7__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_615 VPWR VGND sg13g2_decap_8
XFILLER_14_840 VPWR VGND sg13g2_decap_8
XFILLER_32_136 VPWR VGND sg13g2_decap_8
X_457_ net77 VGND VPWR _051_ mac1.products_ff\[69\] clknet_5_23__leaf_clk sg13g2_dfrbpq_1
X_388_ net151 _082_ VPWR VGND sg13g2_buf_1
XFILLER_12_1012 VPWR VGND sg13g2_decap_8
XFILLER_37_954 VPWR VGND sg13g2_decap_8
XFILLER_24_615 VPWR VGND sg13g2_decap_8
XFILLER_23_158 VPWR VGND sg13g2_decap_8
XFILLER_20_843 VPWR VGND sg13g2_decap_8
XFILLER_11_69 VPWR VGND sg13g2_fill_1
XFILLER_47_707 VPWR VGND sg13g2_decap_8
Xclkbuf_5_10__f_clk clknet_4_5_0_clk clknet_5_10__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_28_910 VPWR VGND sg13g2_decap_8
XFILLER_43_902 VPWR VGND sg13g2_decap_8
XFILLER_27_431 VPWR VGND sg13g2_decap_8
XFILLER_36_44 VPWR VGND sg13g2_fill_2
XFILLER_28_987 VPWR VGND sg13g2_decap_8
XFILLER_43_979 VPWR VGND sg13g2_decap_8
XFILLER_14_125 VPWR VGND sg13g2_decap_8
XFILLER_15_659 VPWR VGND sg13g2_decap_8
XFILLER_42_456 VPWR VGND sg13g2_decap_8
XFILLER_14_169 VPWR VGND sg13g2_fill_2
XFILLER_35_1012 VPWR VGND sg13g2_decap_8
X_311_ _182_ net189 net136 VPWR VGND sg13g2_nand2_1
XFILLER_23_681 VPWR VGND sg13g2_decap_8
X_242_ net149 net155 _058_ VPWR VGND sg13g2_and2_1
XFILLER_10_331 VPWR VGND sg13g2_decap_8
XFILLER_11_865 VPWR VGND sg13g2_decap_8
XFILLER_7_869 VPWR VGND sg13g2_decap_8
XFILLER_42_1016 VPWR VGND sg13g2_decap_8
XFILLER_42_1027 VPWR VGND sg13g2_fill_2
XFILLER_18_431 VPWR VGND sg13g2_decap_8
XFILLER_19_965 VPWR VGND sg13g2_decap_8
XFILLER_34_902 VPWR VGND sg13g2_decap_8
XFILLER_46_795 VPWR VGND sg13g2_decap_8
XFILLER_18_475 VPWR VGND sg13g2_fill_2
XFILLER_33_423 VPWR VGND sg13g2_fill_1
XFILLER_34_979 VPWR VGND sg13g2_decap_8
X_509_ net70 VGND VPWR net110 mac2.sum_lvl1_ff\[8\] clknet_5_12__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_489 VPWR VGND sg13g2_decap_8
XFILLER_9_151 VPWR VGND sg13g2_decap_8
XFILLER_9_195 VPWR VGND sg13g2_decap_8
XFILLER_47_0 VPWR VGND sg13g2_decap_8
XFILLER_29_729 VPWR VGND sg13g2_decap_8
XFILLER_3_1021 VPWR VGND sg13g2_decap_8
XFILLER_28_239 VPWR VGND sg13g2_decap_8
XFILLER_37_751 VPWR VGND sg13g2_decap_8
XFILLER_24_401 VPWR VGND sg13g2_fill_2
XFILLER_25_935 VPWR VGND sg13g2_decap_8
XFILLER_19_1007 VPWR VGND sg13g2_decap_8
XFILLER_24_467 VPWR VGND sg13g2_decap_8
XFILLER_11_106 VPWR VGND sg13g2_decap_8
XFILLER_20_640 VPWR VGND sg13g2_decap_8
XFILLER_3_327 VPWR VGND sg13g2_decap_8
XFILLER_47_504 VPWR VGND sg13g2_decap_8
XFILLER_47_21 VPWR VGND sg13g2_decap_8
XFILLER_19_228 VPWR VGND sg13g2_decap_8
XFILLER_16_935 VPWR VGND sg13g2_decap_8
XFILLER_27_261 VPWR VGND sg13g2_decap_8
XFILLER_28_784 VPWR VGND sg13g2_decap_8
XFILLER_42_220 VPWR VGND sg13g2_decap_8
XFILLER_15_445 VPWR VGND sg13g2_decap_8
XFILLER_43_776 VPWR VGND sg13g2_decap_8
XFILLER_30_404 VPWR VGND sg13g2_decap_8
XFILLER_31_916 VPWR VGND sg13g2_decap_8
X_225_ net165 mac1.sum_lvl3_ff\[0\] _017_ VPWR VGND sg13g2_xor2_1
XFILLER_11_662 VPWR VGND sg13g2_decap_8
XFILLER_7_666 VPWR VGND sg13g2_decap_8
XFILLER_12_90 VPWR VGND sg13g2_decap_8
XFILLER_40_7 VPWR VGND sg13g2_decap_8
XFILLER_19_4 VPWR VGND sg13g2_decap_8
XFILLER_38_537 VPWR VGND sg13g2_decap_8
XFILLER_18_250 VPWR VGND sg13g2_decap_8
XFILLER_19_762 VPWR VGND sg13g2_decap_8
XFILLER_46_592 VPWR VGND sg13g2_decap_8
XFILLER_34_776 VPWR VGND sg13g2_decap_8
XFILLER_21_437 VPWR VGND sg13g2_decap_8
XFILLER_22_949 VPWR VGND sg13g2_decap_8
XFILLER_33_264 VPWR VGND sg13g2_decap_8
XFILLER_0_308 VPWR VGND sg13g2_decap_8
XFILLER_29_526 VPWR VGND sg13g2_decap_8
XFILLER_44_507 VPWR VGND sg13g2_decap_8
XFILLER_17_46 VPWR VGND sg13g2_decap_8
XFILLER_25_732 VPWR VGND sg13g2_decap_8
XFILLER_13_949 VPWR VGND sg13g2_decap_8
XFILLER_24_264 VPWR VGND sg13g2_decap_4
XFILLER_12_448 VPWR VGND sg13g2_decap_4
XFILLER_24_297 VPWR VGND sg13g2_decap_8
XFILLER_33_67 VPWR VGND sg13g2_decap_8
XFILLER_40_757 VPWR VGND sg13g2_decap_8
XFILLER_21_960 VPWR VGND sg13g2_decap_8
XFILLER_32_1026 VPWR VGND sg13g2_fill_2
XFILLER_4_647 VPWR VGND sg13g2_decap_8
Xclkbuf_5_8__f_clk clknet_4_4_0_clk clknet_5_8__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_0_875 VPWR VGND sg13g2_decap_8
XFILLER_48_846 VPWR VGND sg13g2_decap_8
Xhold8 mac2.sum_lvl2_ff\[8\] VPWR VGND net32 sg13g2_dlygate4sd3_1
XFILLER_35_529 VPWR VGND sg13g2_decap_8
XFILLER_16_732 VPWR VGND sg13g2_decap_8
XFILLER_28_581 VPWR VGND sg13g2_decap_8
XFILLER_15_231 VPWR VGND sg13g2_decap_8
XFILLER_43_573 VPWR VGND sg13g2_decap_8
XFILLER_31_713 VPWR VGND sg13g2_decap_8
XFILLER_30_267 VPWR VGND sg13g2_decap_8
XFILLER_11_470 VPWR VGND sg13g2_decap_8
XFILLER_8_986 VPWR VGND sg13g2_decap_8
XFILLER_48_1000 VPWR VGND sg13g2_decap_8
XFILLER_38_312 VPWR VGND sg13g2_decap_8
XFILLER_39_868 VPWR VGND sg13g2_decap_8
XFILLER_26_529 VPWR VGND sg13g2_decap_8
XFILLER_21_212 VPWR VGND sg13g2_decap_8
XFILLER_34_573 VPWR VGND sg13g2_decap_8
XFILLER_22_746 VPWR VGND sg13g2_decap_8
XFILLER_9_80 VPWR VGND sg13g2_fill_2
XFILLER_21_278 VPWR VGND sg13g2_decap_8
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_1_628 VPWR VGND sg13g2_decap_8
XFILLER_28_56 VPWR VGND sg13g2_decap_8
XFILLER_44_304 VPWR VGND sg13g2_decap_8
XFILLER_17_529 VPWR VGND sg13g2_decap_4
XFILLER_29_356 VPWR VGND sg13g2_decap_8
XFILLER_45_849 VPWR VGND sg13g2_decap_8
XFILLER_44_348 VPWR VGND sg13g2_fill_1
X_490_ net67 VGND VPWR _065_ mac2.products_ff\[1\] clknet_5_9__leaf_clk sg13g2_dfrbpq_1
XFILLER_9_717 VPWR VGND sg13g2_decap_8
XFILLER_13_746 VPWR VGND sg13g2_decap_8
XFILLER_40_554 VPWR VGND sg13g2_decap_8
XFILLER_5_934 VPWR VGND sg13g2_decap_8
Xclkbuf_4_0_0_clk clknet_0_clk clknet_4_0_0_clk VPWR VGND sg13g2_buf_8
XFILLER_4_499 VPWR VGND sg13g2_decap_8
XFILLER_0_672 VPWR VGND sg13g2_decap_8
XFILLER_48_643 VPWR VGND sg13g2_decap_8
XFILLER_29_890 VPWR VGND sg13g2_decap_8
XFILLER_35_326 VPWR VGND sg13g2_decap_8
XFILLER_36_849 VPWR VGND sg13g2_decap_8
XFILLER_44_871 VPWR VGND sg13g2_decap_8
XFILLER_31_510 VPWR VGND sg13g2_decap_8
XFILLER_31_587 VPWR VGND sg13g2_decap_8
XFILLER_8_783 VPWR VGND sg13g2_decap_8
XFILLER_27_827 VPWR VGND sg13g2_decap_8
XFILLER_38_131 VPWR VGND sg13g2_decap_8
XFILLER_39_665 VPWR VGND sg13g2_decap_8
XFILLER_26_359 VPWR VGND sg13g2_decap_8
XFILLER_35_893 VPWR VGND sg13g2_decap_8
XFILLER_14_25 VPWR VGND sg13g2_fill_2
XFILLER_22_543 VPWR VGND sg13g2_decap_8
XFILLER_14_69 VPWR VGND sg13g2_decap_8
XFILLER_30_35 VPWR VGND sg13g2_fill_1
XFILLER_2_915 VPWR VGND sg13g2_decap_8
XFILLER_1_425 VPWR VGND sg13g2_decap_8
XFILLER_49_429 VPWR VGND sg13g2_decap_8
XFILLER_39_55 VPWR VGND sg13g2_decap_8
XFILLER_29_120 VPWR VGND sg13g2_decap_8
XFILLER_18_816 VPWR VGND sg13g2_decap_8
XFILLER_45_646 VPWR VGND sg13g2_decap_8
XFILLER_29_186 VPWR VGND sg13g2_fill_1
X_542_ net73 VGND VPWR _082_ DP_1.matrix\[54\] clknet_5_16__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_167 VPWR VGND sg13g2_decap_8
X_473_ net75 VGND VPWR net194 mac1.sum_lvl1_ff\[25\] clknet_5_20__leaf_clk sg13g2_dfrbpq_1
XFILLER_26_893 VPWR VGND sg13g2_decap_8
XFILLER_32_329 VPWR VGND sg13g2_decap_8
XFILLER_41_841 VPWR VGND sg13g2_decap_8
XFILLER_5_731 VPWR VGND sg13g2_decap_8
XFILLER_4_274 VPWR VGND sg13g2_fill_1
XFILLER_4_263 VPWR VGND sg13g2_decap_8
XFILLER_45_1003 VPWR VGND sg13g2_decap_8
XFILLER_1_992 VPWR VGND sg13g2_decap_8
XFILLER_48_440 VPWR VGND sg13g2_decap_8
XFILLER_49_996 VPWR VGND sg13g2_decap_8
XFILLER_36_646 VPWR VGND sg13g2_decap_8
XFILLER_35_189 VPWR VGND sg13g2_decap_8
XFILLER_32_830 VPWR VGND sg13g2_decap_8
XFILLER_8_580 VPWR VGND sg13g2_decap_8
XFILLER_6_81 VPWR VGND sg13g2_decap_8
XFILLER_27_624 VPWR VGND sg13g2_decap_8
XFILLER_39_484 VPWR VGND sg13g2_decap_8
XFILLER_39_495 VPWR VGND sg13g2_fill_2
XFILLER_42_638 VPWR VGND sg13g2_decap_8
XFILLER_14_307 VPWR VGND sg13g2_decap_8
XFILLER_26_156 VPWR VGND sg13g2_decap_8
XFILLER_25_46 VPWR VGND sg13g2_decap_8
XFILLER_35_690 VPWR VGND sg13g2_decap_8
XFILLER_23_863 VPWR VGND sg13g2_decap_8
XFILLER_22_395 VPWR VGND sg13g2_decap_8
XFILLER_10_557 VPWR VGND sg13g2_decap_8
XFILLER_6_517 VPWR VGND sg13g2_decap_8
XFILLER_41_89 VPWR VGND sg13g2_decap_4
XFILLER_2_712 VPWR VGND sg13g2_decap_8
XFILLER_29_1009 VPWR VGND sg13g2_decap_8
XFILLER_1_222 VPWR VGND sg13g2_decap_8
XFILLER_2_789 VPWR VGND sg13g2_decap_8
XFILLER_49_226 VPWR VGND sg13g2_decap_8
XFILLER_1_299 VPWR VGND sg13g2_decap_8
XFILLER_2_39 VPWR VGND sg13g2_decap_8
XFILLER_46_900 VPWR VGND sg13g2_decap_8
XFILLER_18_613 VPWR VGND sg13g2_decap_8
XFILLER_46_977 VPWR VGND sg13g2_decap_8
XFILLER_45_443 VPWR VGND sg13g2_decap_8
X_525_ net62 VGND VPWR net32 mac2.sum_lvl3_ff\[2\] clknet_5_6__leaf_clk sg13g2_dfrbpq_1
XFILLER_26_690 VPWR VGND sg13g2_decap_8
XFILLER_32_115 VPWR VGND sg13g2_decap_8
XFILLER_13_351 VPWR VGND sg13g2_decap_8
X_456_ net78 VGND VPWR _050_ mac1.products_ff\[68\] clknet_5_22__leaf_clk sg13g2_dfrbpq_1
XFILLER_14_896 VPWR VGND sg13g2_decap_8
X_387_ net105 _081_ VPWR VGND sg13g2_buf_1
XFILLER_9_399 VPWR VGND sg13g2_decap_8
XFILLER_49_793 VPWR VGND sg13g2_decap_8
XFILLER_48_270 VPWR VGND sg13g2_fill_2
XFILLER_36_410 VPWR VGND sg13g2_decap_8
XFILLER_37_933 VPWR VGND sg13g2_decap_8
XFILLER_48_281 VPWR VGND sg13g2_decap_8
XFILLER_23_115 VPWR VGND sg13g2_fill_1
XFILLER_23_137 VPWR VGND sg13g2_decap_8
XFILLER_20_822 VPWR VGND sg13g2_decap_8
XFILLER_20_899 VPWR VGND sg13g2_decap_8
XFILLER_27_410 VPWR VGND sg13g2_decap_8
XFILLER_28_966 VPWR VGND sg13g2_decap_8
XFILLER_39_281 VPWR VGND sg13g2_decap_8
XFILLER_14_104 VPWR VGND sg13g2_decap_8
XFILLER_27_487 VPWR VGND sg13g2_decap_8
XFILLER_43_958 VPWR VGND sg13g2_decap_8
XFILLER_42_435 VPWR VGND sg13g2_decap_8
XFILLER_15_638 VPWR VGND sg13g2_decap_8
XFILLER_27_498 VPWR VGND sg13g2_decap_4
X_310_ net123 mac2.products_ff\[119\] _028_ VPWR VGND sg13g2_xor2_1
XFILLER_23_660 VPWR VGND sg13g2_decap_8
XFILLER_30_619 VPWR VGND sg13g2_decap_8
XFILLER_10_310 VPWR VGND sg13g2_decap_8
X_241_ net135 net126 _056_ VPWR VGND sg13g2_and2_1
XFILLER_11_844 VPWR VGND sg13g2_decap_8
XFILLER_7_848 VPWR VGND sg13g2_decap_8
XFILLER_6_325 VPWR VGND sg13g2_decap_8
XFILLER_10_387 VPWR VGND sg13g2_decap_4
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_2_553 VPWR VGND sg13g2_decap_8
XFILLER_2_586 VPWR VGND sg13g2_decap_8
XFILLER_38_719 VPWR VGND sg13g2_decap_8
XFILLER_19_944 VPWR VGND sg13g2_decap_8
XFILLER_46_774 VPWR VGND sg13g2_decap_8
XFILLER_33_402 VPWR VGND sg13g2_decap_8
XFILLER_18_498 VPWR VGND sg13g2_decap_8
XFILLER_34_958 VPWR VGND sg13g2_decap_8
X_508_ net71 VGND VPWR net192 mac2.sum_lvl1_ff\[1\] clknet_5_9__leaf_clk sg13g2_dfrbpq_1
X_439_ net52 _133_ VPWR VGND sg13g2_buf_1
XFILLER_14_693 VPWR VGND sg13g2_decap_8
XFILLER_9_130 VPWR VGND sg13g2_decap_8
XFILLER_5_380 VPWR VGND sg13g2_decap_8
XFILLER_3_60 VPWR VGND sg13g2_decap_8
XFILLER_29_708 VPWR VGND sg13g2_decap_8
XFILLER_3_1000 VPWR VGND sg13g2_decap_8
XFILLER_49_590 VPWR VGND sg13g2_decap_8
XFILLER_37_730 VPWR VGND sg13g2_decap_8
XFILLER_25_914 VPWR VGND sg13g2_decap_8
XFILLER_36_251 VPWR VGND sg13g2_fill_2
XFILLER_24_446 VPWR VGND sg13g2_decap_8
XFILLER_40_939 VPWR VGND sg13g2_decap_8
XFILLER_22_25 VPWR VGND sg13g2_decap_8
XFILLER_20_696 VPWR VGND sg13g2_decap_8
XFILLER_4_829 VPWR VGND sg13g2_decap_8
XFILLER_3_306 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_19_207 VPWR VGND sg13g2_decap_8
XFILLER_47_99 VPWR VGND sg13g2_decap_4
XFILLER_16_914 VPWR VGND sg13g2_decap_8
XFILLER_27_240 VPWR VGND sg13g2_decap_8
XFILLER_28_763 VPWR VGND sg13g2_decap_8
XFILLER_15_424 VPWR VGND sg13g2_decap_8
XFILLER_43_755 VPWR VGND sg13g2_decap_8
X_224_ _142_ net203 net165 VPWR VGND sg13g2_nand2_1
XFILLER_11_641 VPWR VGND sg13g2_decap_8
XFILLER_10_184 VPWR VGND sg13g2_fill_2
XFILLER_10_173 VPWR VGND sg13g2_decap_8
XFILLER_7_645 VPWR VGND sg13g2_decap_8
XFILLER_6_199 VPWR VGND sg13g2_decap_8
XFILLER_3_895 VPWR VGND sg13g2_decap_8
XFILLER_33_7 VPWR VGND sg13g2_decap_8
XFILLER_38_516 VPWR VGND sg13g2_decap_8
XFILLER_19_741 VPWR VGND sg13g2_decap_8
XFILLER_46_571 VPWR VGND sg13g2_decap_8
XFILLER_33_243 VPWR VGND sg13g2_decap_8
XFILLER_34_755 VPWR VGND sg13g2_decap_8
XFILLER_22_928 VPWR VGND sg13g2_decap_8
XFILLER_14_490 VPWR VGND sg13g2_decap_8
XFILLER_30_983 VPWR VGND sg13g2_decap_8
XFILLER_25_1012 VPWR VGND sg13g2_decap_8
XFILLER_17_14 VPWR VGND sg13g2_decap_8
XFILLER_25_711 VPWR VGND sg13g2_decap_8
XFILLER_24_243 VPWR VGND sg13g2_decap_8
XFILLER_12_427 VPWR VGND sg13g2_decap_8
XFILLER_13_928 VPWR VGND sg13g2_decap_8
XFILLER_25_788 VPWR VGND sg13g2_decap_8
XFILLER_40_736 VPWR VGND sg13g2_decap_8
XFILLER_33_35 VPWR VGND sg13g2_fill_2
XFILLER_33_46 VPWR VGND sg13g2_decap_8
XFILLER_32_1005 VPWR VGND sg13g2_decap_8
XFILLER_20_493 VPWR VGND sg13g2_decap_8
XFILLER_4_626 VPWR VGND sg13g2_decap_8
XFILLER_0_854 VPWR VGND sg13g2_decap_8
XFILLER_48_825 VPWR VGND sg13g2_decap_8
Xhold9 mac1.products_ff\[137\] VPWR VGND net33 sg13g2_dlygate4sd3_1
XFILLER_47_346 VPWR VGND sg13g2_fill_2
XFILLER_47_379 VPWR VGND sg13g2_fill_1
XFILLER_47_368 VPWR VGND sg13g2_decap_8
XFILLER_47_357 VPWR VGND sg13g2_fill_2
XFILLER_28_560 VPWR VGND sg13g2_decap_8
XFILLER_35_508 VPWR VGND sg13g2_decap_8
XFILLER_16_711 VPWR VGND sg13g2_decap_8
XFILLER_43_552 VPWR VGND sg13g2_decap_8
XFILLER_16_788 VPWR VGND sg13g2_decap_8
XFILLER_30_246 VPWR VGND sg13g2_decap_8
XFILLER_31_769 VPWR VGND sg13g2_decap_8
XFILLER_8_965 VPWR VGND sg13g2_decap_8
XFILLER_3_692 VPWR VGND sg13g2_decap_8
XFILLER_39_847 VPWR VGND sg13g2_decap_8
XFILLER_26_508 VPWR VGND sg13g2_decap_8
XFILLER_38_368 VPWR VGND sg13g2_decap_8
XFILLER_38_379 VPWR VGND sg13g2_fill_1
XFILLER_34_552 VPWR VGND sg13g2_decap_8
XFILLER_22_725 VPWR VGND sg13g2_decap_8
XFILLER_21_224 VPWR VGND sg13g2_decap_4
XFILLER_21_257 VPWR VGND sg13g2_decap_8
XFILLER_30_780 VPWR VGND sg13g2_decap_8
XFILLER_1_607 VPWR VGND sg13g2_decap_8
XFILLER_28_35 VPWR VGND sg13g2_fill_1
XFILLER_29_313 VPWR VGND sg13g2_decap_8
XFILLER_45_828 VPWR VGND sg13g2_decap_8
XFILLER_38_880 VPWR VGND sg13g2_decap_8
XFILLER_37_390 VPWR VGND sg13g2_decap_8
XFILLER_44_67 VPWR VGND sg13g2_fill_1
XFILLER_44_56 VPWR VGND sg13g2_decap_8
XFILLER_13_725 VPWR VGND sg13g2_decap_8
XFILLER_25_585 VPWR VGND sg13g2_decap_8
XFILLER_40_511 VPWR VGND sg13g2_decap_4
XFILLER_44_89 VPWR VGND sg13g2_fill_1
XFILLER_40_533 VPWR VGND sg13g2_decap_8
XFILLER_12_246 VPWR VGND sg13g2_decap_8
XFILLER_12_257 VPWR VGND sg13g2_fill_1
XFILLER_5_913 VPWR VGND sg13g2_decap_8
XFILLER_4_401 VPWR VGND sg13g2_decap_8
XFILLER_5_39 VPWR VGND sg13g2_decap_8
XFILLER_4_478 VPWR VGND sg13g2_decap_8
XFILLER_0_651 VPWR VGND sg13g2_decap_8
XFILLER_48_622 VPWR VGND sg13g2_decap_8
XFILLER_36_828 VPWR VGND sg13g2_decap_8
XFILLER_48_699 VPWR VGND sg13g2_decap_8
XFILLER_44_850 VPWR VGND sg13g2_decap_8
XFILLER_28_390 VPWR VGND sg13g2_decap_8
XFILLER_16_574 VPWR VGND sg13g2_decap_4
XFILLER_43_393 VPWR VGND sg13g2_decap_8
XFILLER_31_566 VPWR VGND sg13g2_decap_8
XFILLER_8_762 VPWR VGND sg13g2_decap_8
XFILLER_11_290 VPWR VGND sg13g2_decap_8
XFILLER_7_272 VPWR VGND sg13g2_decap_8
XFILLER_4_990 VPWR VGND sg13g2_decap_8
XFILLER_39_644 VPWR VGND sg13g2_decap_8
XFILLER_22_1026 VPWR VGND sg13g2_fill_2
XFILLER_27_806 VPWR VGND sg13g2_decap_8
XFILLER_26_338 VPWR VGND sg13g2_decap_8
XFILLER_35_872 VPWR VGND sg13g2_decap_8
XFILLER_22_522 VPWR VGND sg13g2_decap_8
XFILLER_10_739 VPWR VGND sg13g2_decap_8
XFILLER_22_599 VPWR VGND sg13g2_decap_8
XFILLER_30_14 VPWR VGND sg13g2_decap_8
XFILLER_1_404 VPWR VGND sg13g2_decap_8
XFILLER_49_408 VPWR VGND sg13g2_decap_8
XFILLER_7_1009 VPWR VGND sg13g2_decap_8
XFILLER_39_34 VPWR VGND sg13g2_fill_1
XFILLER_45_625 VPWR VGND sg13g2_decap_8
XFILLER_29_165 VPWR VGND sg13g2_decap_8
X_541_ net83 VGND VPWR _081_ DP_1.matrix\[46\] clknet_5_28__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_146 VPWR VGND sg13g2_decap_8
X_472_ net75 VGND VPWR net100 mac1.sum_lvl1_ff\[24\] clknet_5_20__leaf_clk sg13g2_dfrbpq_1
XFILLER_26_872 VPWR VGND sg13g2_decap_8
XFILLER_41_820 VPWR VGND sg13g2_decap_8
XFILLER_13_599 VPWR VGND sg13g2_decap_8
XFILLER_41_897 VPWR VGND sg13g2_decap_8
XFILLER_5_710 VPWR VGND sg13g2_decap_8
XFILLER_5_787 VPWR VGND sg13g2_decap_8
XFILLER_1_971 VPWR VGND sg13g2_decap_8
XFILLER_49_975 VPWR VGND sg13g2_decap_8
XFILLER_48_496 VPWR VGND sg13g2_decap_8
XFILLER_36_625 VPWR VGND sg13g2_decap_8
XFILLER_35_124 VPWR VGND sg13g2_fill_2
XFILLER_35_168 VPWR VGND sg13g2_decap_8
XFILLER_17_894 VPWR VGND sg13g2_decap_8
XFILLER_32_886 VPWR VGND sg13g2_decap_8
XFILLER_31_385 VPWR VGND sg13g2_fill_1
XFILLER_6_60 VPWR VGND sg13g2_decap_8
XFILLER_27_603 VPWR VGND sg13g2_decap_8
XFILLER_42_617 VPWR VGND sg13g2_decap_8
XFILLER_25_25 VPWR VGND sg13g2_decap_8
XFILLER_23_842 VPWR VGND sg13g2_decap_8
XFILLER_41_149 VPWR VGND sg13g2_decap_8
XFILLER_22_374 VPWR VGND sg13g2_decap_8
XFILLER_10_536 VPWR VGND sg13g2_decap_8
XFILLER_41_68 VPWR VGND sg13g2_decap_8
XFILLER_1_201 VPWR VGND sg13g2_decap_8
XFILLER_9_4 VPWR VGND sg13g2_decap_8
XFILLER_49_205 VPWR VGND sg13g2_decap_8
XFILLER_2_768 VPWR VGND sg13g2_decap_8
XFILLER_1_278 VPWR VGND sg13g2_decap_8
XFILLER_2_18 VPWR VGND sg13g2_decap_8
XFILLER_17_102 VPWR VGND sg13g2_decap_8
XFILLER_46_956 VPWR VGND sg13g2_decap_8
XFILLER_45_422 VPWR VGND sg13g2_decap_8
XFILLER_18_669 VPWR VGND sg13g2_decap_8
X_524_ net65 VGND VPWR net200 mac2.sum_lvl3_ff\[1\] clknet_5_7__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_499 VPWR VGND sg13g2_decap_8
X_455_ net65 VGND VPWR _049_ mac1.products_ff\[52\] clknet_5_24__leaf_clk sg13g2_dfrbpq_1
XFILLER_14_875 VPWR VGND sg13g2_decap_8
X_386_ net138 _080_ VPWR VGND sg13g2_buf_1
XFILLER_41_694 VPWR VGND sg13g2_decap_8
XFILLER_13_396 VPWR VGND sg13g2_decap_8
XFILLER_49_772 VPWR VGND sg13g2_decap_8
XFILLER_37_912 VPWR VGND sg13g2_decap_8
XFILLER_36_455 VPWR VGND sg13g2_decap_4
XFILLER_37_989 VPWR VGND sg13g2_decap_8
XFILLER_17_691 VPWR VGND sg13g2_decap_8
XFILLER_36_499 VPWR VGND sg13g2_decap_8
XFILLER_20_801 VPWR VGND sg13g2_decap_8
XFILLER_32_683 VPWR VGND sg13g2_decap_8
XFILLER_31_182 VPWR VGND sg13g2_fill_2
XFILLER_20_878 VPWR VGND sg13g2_decap_8
XFILLER_46_219 VPWR VGND sg13g2_fill_1
XFILLER_46_208 VPWR VGND sg13g2_decap_8
XFILLER_28_945 VPWR VGND sg13g2_decap_8
XFILLER_36_46 VPWR VGND sg13g2_fill_1
XFILLER_15_617 VPWR VGND sg13g2_decap_8
XFILLER_27_466 VPWR VGND sg13g2_decap_8
XFILLER_36_79 VPWR VGND sg13g2_decap_8
XFILLER_43_937 VPWR VGND sg13g2_decap_8
XFILLER_42_414 VPWR VGND sg13g2_decap_8
X_240_ net120 net151 _054_ VPWR VGND sg13g2_and2_1
XFILLER_11_823 VPWR VGND sg13g2_decap_8
XFILLER_10_366 VPWR VGND sg13g2_decap_8
XFILLER_7_827 VPWR VGND sg13g2_decap_8
XFILLER_6_304 VPWR VGND sg13g2_decap_8
XFILLER_2_565 VPWR VGND sg13g2_decap_8
XFILLER_19_923 VPWR VGND sg13g2_decap_8
XFILLER_37_219 VPWR VGND sg13g2_decap_4
XFILLER_46_753 VPWR VGND sg13g2_decap_8
XFILLER_18_411 VPWR VGND sg13g2_decap_8
XFILLER_18_422 VPWR VGND sg13g2_fill_1
XFILLER_45_241 VPWR VGND sg13g2_decap_8
XFILLER_18_477 VPWR VGND sg13g2_fill_1
XFILLER_45_285 VPWR VGND sg13g2_decap_8
XFILLER_34_937 VPWR VGND sg13g2_decap_8
X_507_ net71 VGND VPWR net96 mac2.sum_lvl1_ff\[0\] clknet_5_12__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_458 VPWR VGND sg13g2_decap_8
XFILLER_42_981 VPWR VGND sg13g2_decap_8
XFILLER_14_672 VPWR VGND sg13g2_decap_8
X_438_ net131 _132_ VPWR VGND sg13g2_buf_1
X_369_ _217_ _216_ _061_ VPWR VGND sg13g2_xor2_1
XFILLER_13_182 VPWR VGND sg13g2_decap_8
XFILLER_9_186 VPWR VGND sg13g2_fill_1
XFILLER_6_893 VPWR VGND sg13g2_decap_8
XFILLER_3_94 VPWR VGND sg13g2_decap_8
XFILLER_36_230 VPWR VGND sg13g2_decap_8
XFILLER_37_786 VPWR VGND sg13g2_decap_8
XFILLER_24_425 VPWR VGND sg13g2_decap_8
XFILLER_40_918 VPWR VGND sg13g2_decap_8
XFILLER_32_480 VPWR VGND sg13g2_decap_8
XFILLER_20_675 VPWR VGND sg13g2_decap_8
XFILLER_4_808 VPWR VGND sg13g2_decap_8
XFILLER_47_539 VPWR VGND sg13g2_decap_8
XFILLER_47_78 VPWR VGND sg13g2_decap_8
XFILLER_47_67 VPWR VGND sg13g2_fill_2
XFILLER_47_56 VPWR VGND sg13g2_decap_8
XFILLER_28_742 VPWR VGND sg13g2_decap_8
XFILLER_43_734 VPWR VGND sg13g2_decap_8
XFILLER_15_403 VPWR VGND sg13g2_decap_8
XFILLER_27_296 VPWR VGND sg13g2_decap_8
XFILLER_42_255 VPWR VGND sg13g2_decap_8
XFILLER_42_288 VPWR VGND sg13g2_decap_8
XFILLER_8_39 VPWR VGND sg13g2_decap_8
X_223_ net118 net133 _068_ VPWR VGND sg13g2_and2_1
XFILLER_11_620 VPWR VGND sg13g2_decap_8
XFILLER_10_152 VPWR VGND sg13g2_decap_8
XFILLER_7_624 VPWR VGND sg13g2_decap_8
XFILLER_11_697 VPWR VGND sg13g2_decap_8
XFILLER_6_145 VPWR VGND sg13g2_decap_4
XFILLER_3_874 VPWR VGND sg13g2_decap_8
XFILLER_19_720 VPWR VGND sg13g2_decap_8
XFILLER_46_550 VPWR VGND sg13g2_decap_8
XFILLER_18_285 VPWR VGND sg13g2_decap_8
XFILLER_19_797 VPWR VGND sg13g2_decap_8
XFILLER_34_734 VPWR VGND sg13g2_decap_8
XFILLER_22_907 VPWR VGND sg13g2_decap_8
XFILLER_15_981 VPWR VGND sg13g2_decap_8
XFILLER_33_299 VPWR VGND sg13g2_fill_2
XFILLER_30_962 VPWR VGND sg13g2_decap_8
XFILLER_6_690 VPWR VGND sg13g2_decap_8
XFILLER_37_583 VPWR VGND sg13g2_decap_8
XFILLER_13_907 VPWR VGND sg13g2_decap_8
XFILLER_24_222 VPWR VGND sg13g2_decap_8
XFILLER_25_767 VPWR VGND sg13g2_decap_8
XFILLER_33_14 VPWR VGND sg13g2_decap_8
XFILLER_33_25 VPWR VGND sg13g2_fill_2
XFILLER_40_715 VPWR VGND sg13g2_decap_8
XFILLER_32_1028 VPWR VGND sg13g2_fill_1
XFILLER_20_472 VPWR VGND sg13g2_decap_8
XFILLER_21_995 VPWR VGND sg13g2_decap_8
XFILLER_4_605 VPWR VGND sg13g2_decap_8
XFILLER_3_115 VPWR VGND sg13g2_fill_1
XFILLER_3_159 VPWR VGND sg13g2_decap_8
XFILLER_0_833 VPWR VGND sg13g2_decap_8
XFILLER_48_804 VPWR VGND sg13g2_decap_8
XFILLER_47_325 VPWR VGND sg13g2_decap_8
XFILLER_43_531 VPWR VGND sg13g2_decap_8
XFILLER_16_767 VPWR VGND sg13g2_decap_8
XFILLER_15_266 VPWR VGND sg13g2_decap_8
XFILLER_30_225 VPWR VGND sg13g2_decap_8
XFILLER_31_748 VPWR VGND sg13g2_decap_8
XFILLER_8_944 VPWR VGND sg13g2_decap_8
XFILLER_12_984 VPWR VGND sg13g2_decap_8
XFILLER_7_443 VPWR VGND sg13g2_decap_8
XFILLER_3_671 VPWR VGND sg13g2_decap_8
XFILLER_24_4 VPWR VGND sg13g2_decap_8
XFILLER_39_826 VPWR VGND sg13g2_decap_8
XFILLER_38_347 VPWR VGND sg13g2_decap_8
XFILLER_0_1015 VPWR VGND sg13g2_decap_8
XFILLER_46_380 VPWR VGND sg13g2_fill_2
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_19_594 VPWR VGND sg13g2_decap_8
XFILLER_34_531 VPWR VGND sg13g2_decap_8
XFILLER_22_704 VPWR VGND sg13g2_decap_8
XFILLER_28_25 VPWR VGND sg13g2_decap_4
XFILLER_45_807 VPWR VGND sg13g2_decap_8
XFILLER_44_339 VPWR VGND sg13g2_decap_8
XFILLER_44_35 VPWR VGND sg13g2_decap_8
XFILLER_13_704 VPWR VGND sg13g2_decap_8
XFILLER_25_564 VPWR VGND sg13g2_decap_8
XFILLER_12_225 VPWR VGND sg13g2_decap_8
XFILLER_21_792 VPWR VGND sg13g2_decap_8
XFILLER_40_589 VPWR VGND sg13g2_decap_8
Xclkbuf_5_16__f_clk clknet_4_8_0_clk clknet_5_16__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_20_291 VPWR VGND sg13g2_decap_8
XFILLER_5_18 VPWR VGND sg13g2_decap_8
XFILLER_5_969 VPWR VGND sg13g2_decap_8
XFILLER_4_457 VPWR VGND sg13g2_decap_8
XFILLER_0_630 VPWR VGND sg13g2_decap_8
XFILLER_48_601 VPWR VGND sg13g2_decap_8
XFILLER_48_678 VPWR VGND sg13g2_decap_8
XFILLER_47_155 VPWR VGND sg13g2_decap_8
XFILLER_36_807 VPWR VGND sg13g2_decap_8
XFILLER_47_166 VPWR VGND sg13g2_fill_2
XFILLER_16_520 VPWR VGND sg13g2_decap_8
XFILLER_16_531 VPWR VGND sg13g2_fill_2
XFILLER_43_372 VPWR VGND sg13g2_decap_8
XFILLER_31_545 VPWR VGND sg13g2_decap_8
XFILLER_8_741 VPWR VGND sg13g2_decap_8
XFILLER_12_781 VPWR VGND sg13g2_decap_8
XFILLER_15_1023 VPWR VGND sg13g2_decap_4
XFILLER_7_251 VPWR VGND sg13g2_decap_8
XFILLER_22_1005 VPWR VGND sg13g2_decap_8
XFILLER_39_623 VPWR VGND sg13g2_decap_8
XFILLER_26_317 VPWR VGND sg13g2_decap_8
XFILLER_38_177 VPWR VGND sg13g2_fill_2
XFILLER_35_851 VPWR VGND sg13g2_decap_8
XFILLER_34_372 VPWR VGND sg13g2_decap_8
XFILLER_10_718 VPWR VGND sg13g2_decap_8
XFILLER_22_578 VPWR VGND sg13g2_decap_8
XFILLER_45_604 VPWR VGND sg13g2_decap_8
XFILLER_29_144 VPWR VGND sg13g2_decap_8
XFILLER_17_328 VPWR VGND sg13g2_decap_8
X_540_ net77 VGND VPWR _080_ DP_1.matrix\[45\] clknet_5_29__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_114 VPWR VGND sg13g2_fill_2
XFILLER_26_851 VPWR VGND sg13g2_decap_8
X_471_ net77 VGND VPWR net188 mac1.sum_lvl1_ff\[17\] clknet_5_22__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_309 VPWR VGND sg13g2_decap_8
XFILLER_13_534 VPWR VGND sg13g2_decap_8
XFILLER_9_505 VPWR VGND sg13g2_decap_8
XFILLER_41_876 VPWR VGND sg13g2_decap_8
XFILLER_9_549 VPWR VGND sg13g2_decap_8
XFILLER_13_578 VPWR VGND sg13g2_decap_8
XFILLER_40_364 VPWR VGND sg13g2_decap_8
XFILLER_5_766 VPWR VGND sg13g2_decap_8
XFILLER_4_243 VPWR VGND sg13g2_decap_4
XFILLER_20_81 VPWR VGND sg13g2_decap_8
XFILLER_1_950 VPWR VGND sg13g2_decap_8
XFILLER_49_954 VPWR VGND sg13g2_decap_8
XFILLER_48_475 VPWR VGND sg13g2_decap_8
Xhold90 DP_4.matrix\[72\] VPWR VGND net140 sg13g2_dlygate4sd3_1
XFILLER_36_604 VPWR VGND sg13g2_decap_8
XFILLER_17_873 VPWR VGND sg13g2_decap_8
XFILLER_43_180 VPWR VGND sg13g2_decap_4
XFILLER_32_865 VPWR VGND sg13g2_decap_8
XFILLER_31_364 VPWR VGND sg13g2_decap_8
XFILLER_39_420 VPWR VGND sg13g2_fill_1
XFILLER_27_659 VPWR VGND sg13g2_decap_8
XFILLER_23_821 VPWR VGND sg13g2_decap_8
XFILLER_41_106 VPWR VGND sg13g2_fill_2
XFILLER_34_180 VPWR VGND sg13g2_decap_8
XFILLER_10_515 VPWR VGND sg13g2_decap_8
XFILLER_22_353 VPWR VGND sg13g2_decap_8
XFILLER_23_898 VPWR VGND sg13g2_decap_8
XFILLER_41_47 VPWR VGND sg13g2_decap_8
XFILLER_2_747 VPWR VGND sg13g2_decap_8
XFILLER_1_257 VPWR VGND sg13g2_decap_8
XFILLER_46_935 VPWR VGND sg13g2_decap_8
XFILLER_18_648 VPWR VGND sg13g2_decap_8
XFILLER_45_478 VPWR VGND sg13g2_decap_8
X_523_ net65 VGND VPWR net164 mac2.sum_lvl3_ff\[0\] clknet_5_7__leaf_clk sg13g2_dfrbpq_1
X_454_ net65 VGND VPWR _048_ mac1.products_ff\[51\] clknet_5_25__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_629 VPWR VGND sg13g2_decap_8
XFILLER_14_854 VPWR VGND sg13g2_decap_8
XFILLER_25_191 VPWR VGND sg13g2_decap_8
X_385_ net87 _079_ VPWR VGND sg13g2_buf_1
XFILLER_41_673 VPWR VGND sg13g2_decap_8
XFILLER_12_1026 VPWR VGND sg13g2_fill_2
XFILLER_31_91 VPWR VGND sg13g2_decap_8
Xoutput1 net1 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_49_751 VPWR VGND sg13g2_decap_8
XFILLER_37_968 VPWR VGND sg13g2_decap_8
XFILLER_36_467 VPWR VGND sg13g2_fill_2
XFILLER_36_478 VPWR VGND sg13g2_decap_8
XFILLER_17_670 VPWR VGND sg13g2_decap_8
XFILLER_24_629 VPWR VGND sg13g2_decap_8
XFILLER_31_161 VPWR VGND sg13g2_decap_8
XFILLER_32_662 VPWR VGND sg13g2_decap_8
XFILLER_20_857 VPWR VGND sg13g2_decap_8
XFILLER_28_1022 VPWR VGND sg13g2_decap_8
XFILLER_28_924 VPWR VGND sg13g2_decap_8
XFILLER_36_14 VPWR VGND sg13g2_fill_2
XFILLER_43_916 VPWR VGND sg13g2_decap_8
XFILLER_27_445 VPWR VGND sg13g2_decap_8
XFILLER_14_139 VPWR VGND sg13g2_decap_8
XFILLER_10_301 VPWR VGND sg13g2_decap_4
XFILLER_11_802 VPWR VGND sg13g2_decap_8
XFILLER_35_1026 VPWR VGND sg13g2_fill_2
XFILLER_7_806 VPWR VGND sg13g2_decap_8
XFILLER_22_183 VPWR VGND sg13g2_decap_8
XFILLER_22_194 VPWR VGND sg13g2_decap_8
XFILLER_23_695 VPWR VGND sg13g2_decap_8
XFILLER_10_345 VPWR VGND sg13g2_decap_8
XFILLER_11_879 VPWR VGND sg13g2_decap_8
XFILLER_6_349 VPWR VGND sg13g2_decap_8
XFILLER_2_511 VPWR VGND sg13g2_decap_8
XFILLER_19_902 VPWR VGND sg13g2_decap_8
XFILLER_46_732 VPWR VGND sg13g2_decap_8
XFILLER_45_220 VPWR VGND sg13g2_decap_8
XFILLER_18_445 VPWR VGND sg13g2_decap_8
XFILLER_19_979 VPWR VGND sg13g2_decap_8
XFILLER_34_916 VPWR VGND sg13g2_decap_8
XFILLER_45_264 VPWR VGND sg13g2_decap_8
X_506_ net62 VGND VPWR _039_ mac2.products_ff\[137\] clknet_5_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_42_960 VPWR VGND sg13g2_decap_8
XFILLER_14_651 VPWR VGND sg13g2_decap_8
X_437_ net49 _131_ VPWR VGND sg13g2_buf_1
X_368_ _217_ net125 net39 VPWR VGND sg13g2_nand2_1
XFILLER_9_165 VPWR VGND sg13g2_decap_8
X_299_ _176_ net179 net109 VPWR VGND sg13g2_nand2_1
XFILLER_6_872 VPWR VGND sg13g2_decap_8
XFILLER_36_253 VPWR VGND sg13g2_fill_1
XFILLER_37_765 VPWR VGND sg13g2_decap_8
XFILLER_25_949 VPWR VGND sg13g2_decap_8
XFILLER_33_993 VPWR VGND sg13g2_decap_8
XFILLER_20_654 VPWR VGND sg13g2_decap_8
XFILLER_47_518 VPWR VGND sg13g2_decap_8
XFILLER_47_35 VPWR VGND sg13g2_decap_8
XFILLER_28_721 VPWR VGND sg13g2_decap_8
XFILLER_43_713 VPWR VGND sg13g2_decap_8
XFILLER_16_949 VPWR VGND sg13g2_decap_8
XFILLER_27_275 VPWR VGND sg13g2_decap_8
XFILLER_28_798 VPWR VGND sg13g2_decap_8
XFILLER_42_234 VPWR VGND sg13g2_decap_8
XFILLER_15_459 VPWR VGND sg13g2_decap_8
XFILLER_30_418 VPWR VGND sg13g2_decap_8
X_222_ net148 net130 _066_ VPWR VGND sg13g2_and2_1
XFILLER_8_18 VPWR VGND sg13g2_decap_8
XFILLER_24_993 VPWR VGND sg13g2_decap_8
XFILLER_10_131 VPWR VGND sg13g2_decap_8
XFILLER_7_603 VPWR VGND sg13g2_decap_8
XFILLER_11_676 VPWR VGND sg13g2_decap_8
XFILLER_6_102 VPWR VGND sg13g2_decap_8
XFILLER_3_853 VPWR VGND sg13g2_decap_8
XFILLER_2_363 VPWR VGND sg13g2_decap_8
XFILLER_2_374 VPWR VGND sg13g2_fill_2
XFILLER_19_776 VPWR VGND sg13g2_decap_8
XFILLER_18_264 VPWR VGND sg13g2_decap_8
XFILLER_34_713 VPWR VGND sg13g2_decap_8
XFILLER_33_234 VPWR VGND sg13g2_decap_4
XFILLER_15_960 VPWR VGND sg13g2_decap_8
XFILLER_33_278 VPWR VGND sg13g2_decap_8
XFILLER_30_941 VPWR VGND sg13g2_decap_8
XFILLER_45_0 VPWR VGND sg13g2_decap_8
XFILLER_24_201 VPWR VGND sg13g2_decap_8
XFILLER_37_562 VPWR VGND sg13g2_decap_8
XFILLER_25_746 VPWR VGND sg13g2_decap_8
XFILLER_33_790 VPWR VGND sg13g2_decap_8
XFILLER_20_451 VPWR VGND sg13g2_decap_8
XFILLER_21_974 VPWR VGND sg13g2_decap_8
XFILLER_3_105 VPWR VGND sg13g2_fill_2
XFILLER_3_138 VPWR VGND sg13g2_decap_8
XFILLER_0_812 VPWR VGND sg13g2_decap_8
XFILLER_47_304 VPWR VGND sg13g2_decap_8
XFILLER_0_889 VPWR VGND sg13g2_decap_8
XFILLER_47_348 VPWR VGND sg13g2_fill_1
XFILLER_43_510 VPWR VGND sg13g2_decap_8
XFILLER_15_212 VPWR VGND sg13g2_fill_2
XFILLER_16_746 VPWR VGND sg13g2_decap_8
XFILLER_28_595 VPWR VGND sg13g2_decap_8
XFILLER_43_587 VPWR VGND sg13g2_decap_8
XFILLER_15_245 VPWR VGND sg13g2_decap_8
XFILLER_30_204 VPWR VGND sg13g2_decap_8
XFILLER_31_727 VPWR VGND sg13g2_decap_8
XFILLER_24_790 VPWR VGND sg13g2_decap_8
XFILLER_8_923 VPWR VGND sg13g2_decap_8
XFILLER_12_963 VPWR VGND sg13g2_decap_8
XFILLER_7_422 VPWR VGND sg13g2_decap_8
XFILLER_7_477 VPWR VGND sg13g2_decap_8
XFILLER_48_1014 VPWR VGND sg13g2_decap_8
XFILLER_3_650 VPWR VGND sg13g2_decap_8
XFILLER_39_805 VPWR VGND sg13g2_decap_8
XFILLER_38_326 VPWR VGND sg13g2_decap_8
XFILLER_47_882 VPWR VGND sg13g2_decap_8
XFILLER_19_573 VPWR VGND sg13g2_decap_8
XFILLER_34_510 VPWR VGND sg13g2_decap_8
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_34_587 VPWR VGND sg13g2_decap_8
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_44_318 VPWR VGND sg13g2_decap_8
XFILLER_44_14 VPWR VGND sg13g2_decap_8
XFILLER_25_543 VPWR VGND sg13g2_decap_8
XFILLER_40_568 VPWR VGND sg13g2_decap_8
XFILLER_21_771 VPWR VGND sg13g2_decap_8
XFILLER_20_270 VPWR VGND sg13g2_decap_8
XFILLER_5_948 VPWR VGND sg13g2_decap_8
XFILLER_4_436 VPWR VGND sg13g2_decap_8
XFILLER_0_686 VPWR VGND sg13g2_decap_8
XFILLER_48_657 VPWR VGND sg13g2_decap_8
XFILLER_47_134 VPWR VGND sg13g2_decap_8
XFILLER_18_81 VPWR VGND sg13g2_decap_4
XFILLER_44_885 VPWR VGND sg13g2_decap_8
XFILLER_43_351 VPWR VGND sg13g2_decap_8
XFILLER_31_524 VPWR VGND sg13g2_decap_8
XFILLER_15_1002 VPWR VGND sg13g2_decap_8
XFILLER_8_720 VPWR VGND sg13g2_decap_8
XFILLER_12_760 VPWR VGND sg13g2_decap_8
XFILLER_7_230 VPWR VGND sg13g2_decap_8
XFILLER_8_797 VPWR VGND sg13g2_decap_8
XFILLER_39_602 VPWR VGND sg13g2_decap_8
XFILLER_22_1028 VPWR VGND sg13g2_fill_1
XFILLER_38_145 VPWR VGND sg13g2_decap_8
XFILLER_38_156 VPWR VGND sg13g2_fill_1
XFILLER_39_679 VPWR VGND sg13g2_decap_8
XFILLER_19_392 VPWR VGND sg13g2_decap_8
XFILLER_35_830 VPWR VGND sg13g2_decap_8
Xclkbuf_5_22__f_clk clknet_4_11_0_clk clknet_5_22__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_34_351 VPWR VGND sg13g2_decap_8
XFILLER_22_557 VPWR VGND sg13g2_decap_8
XFILLER_30_49 VPWR VGND sg13g2_decap_8
XFILLER_2_929 VPWR VGND sg13g2_decap_8
XFILLER_1_439 VPWR VGND sg13g2_decap_8
XFILLER_39_14 VPWR VGND sg13g2_decap_8
XFILLER_17_307 VPWR VGND sg13g2_decap_8
XFILLER_26_830 VPWR VGND sg13g2_decap_8
X_470_ net77 VGND VPWR net114 mac1.sum_lvl1_ff\[16\] clknet_5_22__leaf_clk sg13g2_dfrbpq_1
XFILLER_25_351 VPWR VGND sg13g2_decap_8
XFILLER_38_1013 VPWR VGND sg13g2_decap_8
XFILLER_13_513 VPWR VGND sg13g2_decap_8
XFILLER_41_855 VPWR VGND sg13g2_decap_8
XFILLER_40_398 VPWR VGND sg13g2_decap_8
XFILLER_4_200 VPWR VGND sg13g2_decap_8
XFILLER_5_745 VPWR VGND sg13g2_decap_8
XFILLER_20_60 VPWR VGND sg13g2_decap_8
XFILLER_45_1017 VPWR VGND sg13g2_decap_8
XFILLER_45_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_933 VPWR VGND sg13g2_decap_8
XFILLER_48_454 VPWR VGND sg13g2_decap_8
XFILLER_0_483 VPWR VGND sg13g2_decap_8
Xhold91 DP_3.matrix\[63\] VPWR VGND net141 sg13g2_dlygate4sd3_1
Xhold80 DP_4.matrix\[18\] VPWR VGND net130 sg13g2_dlygate4sd3_1
XFILLER_35_126 VPWR VGND sg13g2_fill_1
XFILLER_17_852 VPWR VGND sg13g2_decap_8
X_599_ net82 VGND VPWR _139_ DP_4.matrix\[64\] clknet_5_30__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_90 VPWR VGND sg13g2_decap_8
XFILLER_44_682 VPWR VGND sg13g2_decap_8
XFILLER_16_362 VPWR VGND sg13g2_decap_8
XFILLER_32_844 VPWR VGND sg13g2_decap_8
XFILLER_8_594 VPWR VGND sg13g2_decap_8
XFILLER_6_95 VPWR VGND sg13g2_decap_8
XFILLER_26_115 VPWR VGND sg13g2_decap_8
XFILLER_27_638 VPWR VGND sg13g2_decap_8
XFILLER_23_800 VPWR VGND sg13g2_decap_8
XFILLER_22_332 VPWR VGND sg13g2_decap_8
XFILLER_23_877 VPWR VGND sg13g2_decap_8
XFILLER_2_726 VPWR VGND sg13g2_decap_8
XFILLER_1_236 VPWR VGND sg13g2_decap_8
XFILLER_46_914 VPWR VGND sg13g2_decap_8
XFILLER_18_627 VPWR VGND sg13g2_decap_8
XFILLER_45_457 VPWR VGND sg13g2_decap_8
X_522_ net63 VGND VPWR net28 mac2.sum_lvl2_ff\[9\] clknet_5_3__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_608 VPWR VGND sg13g2_decap_8
XFILLER_14_833 VPWR VGND sg13g2_decap_8
X_453_ net65 VGND VPWR _047_ mac1.products_ff\[35\] clknet_5_25__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_129 VPWR VGND sg13g2_decap_8
XFILLER_25_170 VPWR VGND sg13g2_decap_8
XFILLER_41_652 VPWR VGND sg13g2_decap_8
XFILLER_9_325 VPWR VGND sg13g2_decap_4
XFILLER_13_365 VPWR VGND sg13g2_decap_4
X_384_ net139 _078_ VPWR VGND sg13g2_buf_1
XFILLER_40_173 VPWR VGND sg13g2_fill_2
XFILLER_12_1005 VPWR VGND sg13g2_decap_8
XFILLER_5_520 VPWR VGND sg13g2_decap_8
XFILLER_31_70 VPWR VGND sg13g2_decap_8
XFILLER_5_553 VPWR VGND sg13g2_decap_8
XFILLER_49_7 VPWR VGND sg13g2_decap_8
Xoutput2 net2 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_49_730 VPWR VGND sg13g2_decap_8
XFILLER_0_280 VPWR VGND sg13g2_decap_8
XFILLER_48_295 VPWR VGND sg13g2_decap_8
XFILLER_36_424 VPWR VGND sg13g2_decap_4
XFILLER_37_947 VPWR VGND sg13g2_decap_8
XFILLER_24_608 VPWR VGND sg13g2_decap_8
XFILLER_32_641 VPWR VGND sg13g2_decap_8
XFILLER_31_140 VPWR VGND sg13g2_decap_8
XFILLER_20_836 VPWR VGND sg13g2_decap_8
XFILLER_31_184 VPWR VGND sg13g2_fill_1
XFILLER_9_892 VPWR VGND sg13g2_decap_8
XFILLER_11_18 VPWR VGND sg13g2_decap_4
XFILLER_28_1001 VPWR VGND sg13g2_decap_8
XFILLER_28_903 VPWR VGND sg13g2_decap_8
XFILLER_27_424 VPWR VGND sg13g2_decap_8
XFILLER_39_295 VPWR VGND sg13g2_decap_8
XFILLER_14_118 VPWR VGND sg13g2_decap_8
XFILLER_42_449 VPWR VGND sg13g2_decap_8
XFILLER_23_674 VPWR VGND sg13g2_decap_8
XFILLER_35_1005 VPWR VGND sg13g2_decap_8
XFILLER_10_324 VPWR VGND sg13g2_decap_8
XFILLER_11_858 VPWR VGND sg13g2_decap_8
XFILLER_22_162 VPWR VGND sg13g2_decap_8
XFILLER_42_1009 VPWR VGND sg13g2_decap_8
XFILLER_46_711 VPWR VGND sg13g2_decap_8
XFILLER_19_958 VPWR VGND sg13g2_decap_8
XFILLER_46_788 VPWR VGND sg13g2_decap_8
X_505_ net62 VGND VPWR _038_ mac2.products_ff\[136\] clknet_5_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_416 VPWR VGND sg13g2_decap_8
XFILLER_14_630 VPWR VGND sg13g2_decap_8
XFILLER_26_81 VPWR VGND sg13g2_decap_8
XFILLER_13_151 VPWR VGND sg13g2_decap_8
X_436_ net155 _130_ VPWR VGND sg13g2_buf_1
X_367_ _216_ net158 net102 VPWR VGND sg13g2_nand2_1
XFILLER_41_482 VPWR VGND sg13g2_decap_8
XFILLER_42_80 VPWR VGND sg13g2_decap_8
XFILLER_9_144 VPWR VGND sg13g2_decap_8
X_298_ net115 mac2.sum_lvl3_ff\[2\] _020_ VPWR VGND sg13g2_xor2_1
XFILLER_6_851 VPWR VGND sg13g2_decap_8
XFILLER_5_394 VPWR VGND sg13g2_decap_8
XFILLER_3_1014 VPWR VGND sg13g2_decap_8
XFILLER_37_744 VPWR VGND sg13g2_decap_8
XFILLER_18_991 VPWR VGND sg13g2_decap_8
XFILLER_25_928 VPWR VGND sg13g2_decap_8
XFILLER_36_276 VPWR VGND sg13g2_decap_4
XFILLER_17_490 VPWR VGND sg13g2_fill_2
XFILLER_36_298 VPWR VGND sg13g2_decap_8
XFILLER_33_972 VPWR VGND sg13g2_decap_8
XFILLER_20_633 VPWR VGND sg13g2_decap_8
XFILLER_47_14 VPWR VGND sg13g2_decap_8
XFILLER_28_700 VPWR VGND sg13g2_decap_8
XFILLER_27_210 VPWR VGND sg13g2_fill_2
XFILLER_28_777 VPWR VGND sg13g2_decap_8
XFILLER_16_928 VPWR VGND sg13g2_decap_8
XFILLER_27_254 VPWR VGND sg13g2_decap_8
XFILLER_43_769 VPWR VGND sg13g2_decap_8
XFILLER_42_213 VPWR VGND sg13g2_decap_8
XFILLER_15_438 VPWR VGND sg13g2_decap_8
XFILLER_31_909 VPWR VGND sg13g2_decap_8
XFILLER_24_972 VPWR VGND sg13g2_decap_8
XFILLER_11_655 VPWR VGND sg13g2_decap_8
XFILLER_7_659 VPWR VGND sg13g2_decap_8
XFILLER_12_83 VPWR VGND sg13g2_decap_8
XFILLER_3_832 VPWR VGND sg13g2_decap_8
XFILLER_2_342 VPWR VGND sg13g2_decap_8
XFILLER_18_243 VPWR VGND sg13g2_decap_8
XFILLER_19_755 VPWR VGND sg13g2_decap_8
Xclkbuf_5_3__f_clk clknet_4_1_0_clk clknet_5_3__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_46_585 VPWR VGND sg13g2_decap_8
XFILLER_34_769 VPWR VGND sg13g2_decap_8
XFILLER_21_408 VPWR VGND sg13g2_fill_2
XFILLER_33_257 VPWR VGND sg13g2_decap_8
XFILLER_30_920 VPWR VGND sg13g2_decap_8
X_419_ net50 _113_ VPWR VGND sg13g2_buf_1
XFILLER_30_997 VPWR VGND sg13g2_decap_8
XFILLER_38_0 VPWR VGND sg13g2_decap_8
XFILLER_25_1026 VPWR VGND sg13g2_fill_2
XFILLER_29_519 VPWR VGND sg13g2_decap_8
XFILLER_17_28 VPWR VGND sg13g2_fill_2
XFILLER_37_541 VPWR VGND sg13g2_decap_8
XFILLER_17_39 VPWR VGND sg13g2_decap_8
XFILLER_25_725 VPWR VGND sg13g2_decap_8
XFILLER_24_257 VPWR VGND sg13g2_decap_8
XFILLER_24_268 VPWR VGND sg13g2_fill_2
XFILLER_20_430 VPWR VGND sg13g2_decap_8
XFILLER_21_953 VPWR VGND sg13g2_decap_8
XFILLER_32_1019 VPWR VGND sg13g2_decap_8
XFILLER_0_868 VPWR VGND sg13g2_decap_8
XFILLER_48_839 VPWR VGND sg13g2_decap_8
XFILLER_16_725 VPWR VGND sg13g2_decap_8
XFILLER_28_574 VPWR VGND sg13g2_decap_8
XFILLER_15_224 VPWR VGND sg13g2_decap_8
XFILLER_43_566 VPWR VGND sg13g2_decap_8
XFILLER_31_706 VPWR VGND sg13g2_decap_8
XFILLER_8_902 VPWR VGND sg13g2_decap_8
XFILLER_12_942 VPWR VGND sg13g2_decap_8
XFILLER_7_401 VPWR VGND sg13g2_fill_1
XFILLER_11_463 VPWR VGND sg13g2_decap_8
XFILLER_8_979 VPWR VGND sg13g2_decap_8
XFILLER_31_7 VPWR VGND sg13g2_decap_8
XFILLER_38_305 VPWR VGND sg13g2_decap_8
XFILLER_47_861 VPWR VGND sg13g2_decap_8
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_19_552 VPWR VGND sg13g2_decap_8
XFILLER_46_382 VPWR VGND sg13g2_fill_1
XFILLER_34_566 VPWR VGND sg13g2_decap_8
XFILLER_21_205 VPWR VGND sg13g2_decap_8
XFILLER_22_739 VPWR VGND sg13g2_decap_8
XFILLER_9_62 VPWR VGND sg13g2_decap_8
XFILLER_9_95 VPWR VGND sg13g2_decap_8
XFILLER_30_794 VPWR VGND sg13g2_decap_8
Xclkbuf_4_15_0_clk clknet_0_clk clknet_4_15_0_clk VPWR VGND sg13g2_buf_8
XFILLER_29_327 VPWR VGND sg13g2_fill_2
XFILLER_28_49 VPWR VGND sg13g2_decap_8
XFILLER_25_522 VPWR VGND sg13g2_decap_8
XFILLER_38_894 VPWR VGND sg13g2_decap_8
XFILLER_13_739 VPWR VGND sg13g2_decap_8
XFILLER_25_599 VPWR VGND sg13g2_decap_8
XFILLER_21_750 VPWR VGND sg13g2_decap_8
XFILLER_40_547 VPWR VGND sg13g2_decap_8
XFILLER_5_927 VPWR VGND sg13g2_decap_8
XFILLER_0_665 VPWR VGND sg13g2_decap_8
XFILLER_48_636 VPWR VGND sg13g2_decap_8
XFILLER_18_60 VPWR VGND sg13g2_decap_8
XFILLER_29_883 VPWR VGND sg13g2_decap_8
XFILLER_35_319 VPWR VGND sg13g2_decap_8
XFILLER_44_864 VPWR VGND sg13g2_decap_8
XFILLER_43_330 VPWR VGND sg13g2_decap_8
XFILLER_31_503 VPWR VGND sg13g2_decap_8
XFILLER_8_776 VPWR VGND sg13g2_decap_8
XFILLER_7_286 VPWR VGND sg13g2_decap_8
XFILLER_38_124 VPWR VGND sg13g2_decap_8
XFILLER_39_658 VPWR VGND sg13g2_decap_8
XFILLER_38_179 VPWR VGND sg13g2_fill_1
XFILLER_19_360 VPWR VGND sg13g2_decap_4
XFILLER_34_330 VPWR VGND sg13g2_decap_8
XFILLER_14_18 VPWR VGND sg13g2_decap_8
XFILLER_35_886 VPWR VGND sg13g2_decap_8
XFILLER_22_536 VPWR VGND sg13g2_decap_8
XFILLER_30_591 VPWR VGND sg13g2_decap_8
XFILLER_30_28 VPWR VGND sg13g2_fill_1
XFILLER_2_908 VPWR VGND sg13g2_decap_8
XFILLER_1_418 VPWR VGND sg13g2_decap_8
XFILLER_39_48 VPWR VGND sg13g2_decap_8
XFILLER_18_809 VPWR VGND sg13g2_decap_8
XFILLER_29_113 VPWR VGND sg13g2_decap_8
XFILLER_29_179 VPWR VGND sg13g2_decap_8
XFILLER_45_639 VPWR VGND sg13g2_decap_8
XFILLER_38_691 VPWR VGND sg13g2_decap_8
XFILLER_25_330 VPWR VGND sg13g2_decap_8
XFILLER_26_886 VPWR VGND sg13g2_decap_8
XFILLER_41_834 VPWR VGND sg13g2_decap_8
XFILLER_13_558 VPWR VGND sg13g2_decap_4
XFILLER_25_396 VPWR VGND sg13g2_decap_8
XFILLER_5_724 VPWR VGND sg13g2_decap_8
XFILLER_4_256 VPWR VGND sg13g2_decap_8
XFILLER_49_912 VPWR VGND sg13g2_decap_8
XFILLER_0_462 VPWR VGND sg13g2_decap_8
XFILLER_1_985 VPWR VGND sg13g2_decap_8
XFILLER_48_433 VPWR VGND sg13g2_decap_8
XFILLER_49_989 VPWR VGND sg13g2_decap_8
Xhold70 DP_2.matrix\[54\] VPWR VGND net120 sg13g2_dlygate4sd3_1
Xhold92 DP_2.matrix\[0\] VPWR VGND net142 sg13g2_dlygate4sd3_1
Xhold81 DP_4.matrix\[36\] VPWR VGND net131 sg13g2_dlygate4sd3_1
XFILLER_17_831 VPWR VGND sg13g2_decap_8
XFILLER_29_680 VPWR VGND sg13g2_decap_8
XFILLER_36_639 VPWR VGND sg13g2_decap_8
XFILLER_16_341 VPWR VGND sg13g2_decap_8
X_598_ net82 VGND VPWR _138_ DP_4.matrix\[63\] clknet_5_27__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_661 VPWR VGND sg13g2_decap_8
XFILLER_32_823 VPWR VGND sg13g2_decap_8
XFILLER_31_322 VPWR VGND sg13g2_fill_2
XFILLER_8_573 VPWR VGND sg13g2_decap_8
XFILLER_6_74 VPWR VGND sg13g2_decap_8
XFILLER_6_1012 VPWR VGND sg13g2_decap_8
XFILLER_27_617 VPWR VGND sg13g2_decap_8
XFILLER_39_477 VPWR VGND sg13g2_decap_8
XFILLER_26_149 VPWR VGND sg13g2_decap_8
XFILLER_25_39 VPWR VGND sg13g2_decap_8
XFILLER_35_683 VPWR VGND sg13g2_decap_8
XFILLER_23_856 VPWR VGND sg13g2_decap_8
XFILLER_22_388 VPWR VGND sg13g2_decap_8
XFILLER_2_705 VPWR VGND sg13g2_decap_8
XFILLER_1_215 VPWR VGND sg13g2_decap_8
XFILLER_49_219 VPWR VGND sg13g2_decap_8
XFILLER_18_606 VPWR VGND sg13g2_decap_8
XFILLER_45_436 VPWR VGND sg13g2_decap_8
XFILLER_17_116 VPWR VGND sg13g2_decap_4
X_521_ net63 VGND VPWR net26 mac2.sum_lvl2_ff\[8\] clknet_5_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_14_812 VPWR VGND sg13g2_decap_8
X_452_ net85 VGND VPWR _046_ mac1.products_ff\[34\] clknet_5_18__leaf_clk sg13g2_dfrbpq_1
XFILLER_26_683 VPWR VGND sg13g2_decap_8
XFILLER_32_108 VPWR VGND sg13g2_decap_8
X_383_ net47 _077_ VPWR VGND sg13g2_buf_1
XFILLER_41_631 VPWR VGND sg13g2_decap_8
XFILLER_13_344 VPWR VGND sg13g2_decap_8
XFILLER_14_889 VPWR VGND sg13g2_decap_8
XFILLER_40_152 VPWR VGND sg13g2_decap_8
XFILLER_12_1028 VPWR VGND sg13g2_fill_1
XFILLER_5_598 VPWR VGND sg13g2_decap_8
Xoutput3 net3 uo_out[2] VPWR VGND sg13g2_buf_1
XFILLER_1_782 VPWR VGND sg13g2_decap_8
XFILLER_49_786 VPWR VGND sg13g2_decap_8
XFILLER_37_926 VPWR VGND sg13g2_decap_8
XFILLER_48_263 VPWR VGND sg13g2_decap_8
XFILLER_36_403 VPWR VGND sg13g2_decap_8
XFILLER_23_108 VPWR VGND sg13g2_decap_8
XFILLER_32_620 VPWR VGND sg13g2_decap_8
XFILLER_20_815 VPWR VGND sg13g2_decap_8
XFILLER_32_697 VPWR VGND sg13g2_decap_8
XFILLER_9_871 VPWR VGND sg13g2_decap_8
XFILLER_31_196 VPWR VGND sg13g2_decap_8
XFILLER_28_959 VPWR VGND sg13g2_decap_8
XFILLER_36_16 VPWR VGND sg13g2_fill_1
XFILLER_42_428 VPWR VGND sg13g2_decap_8
XFILLER_35_480 VPWR VGND sg13g2_fill_1
XFILLER_22_141 VPWR VGND sg13g2_decap_8
XFILLER_23_653 VPWR VGND sg13g2_decap_8
XFILLER_35_1028 VPWR VGND sg13g2_fill_1
XFILLER_11_837 VPWR VGND sg13g2_decap_8
XFILLER_6_318 VPWR VGND sg13g2_decap_8
XFILLER_2_546 VPWR VGND sg13g2_decap_8
XFILLER_2_579 VPWR VGND sg13g2_decap_8
XFILLER_19_937 VPWR VGND sg13g2_decap_8
XFILLER_46_767 VPWR VGND sg13g2_decap_8
XFILLER_45_255 VPWR VGND sg13g2_decap_4
X_504_ net82 VGND VPWR _035_ mac2.products_ff\[120\] clknet_5_30__leaf_clk sg13g2_dfrbpq_1
XFILLER_26_60 VPWR VGND sg13g2_decap_8
XFILLER_27_981 VPWR VGND sg13g2_decap_8
XFILLER_45_299 VPWR VGND sg13g2_decap_8
XFILLER_26_480 VPWR VGND sg13g2_decap_8
X_435_ net45 _129_ VPWR VGND sg13g2_buf_1
XFILLER_13_130 VPWR VGND sg13g2_decap_8
XFILLER_42_995 VPWR VGND sg13g2_decap_8
XFILLER_9_123 VPWR VGND sg13g2_decap_8
XFILLER_14_686 VPWR VGND sg13g2_decap_8
X_366_ _215_ _214_ _059_ VPWR VGND sg13g2_xor2_1
XFILLER_41_461 VPWR VGND sg13g2_decap_8
XFILLER_13_196 VPWR VGND sg13g2_decap_8
X_297_ _021_ _172_ _175_ VPWR VGND sg13g2_xnor2_1
XFILLER_6_830 VPWR VGND sg13g2_decap_8
XFILLER_5_373 VPWR VGND sg13g2_decap_8
XFILLER_3_53 VPWR VGND sg13g2_decap_8
XFILLER_49_583 VPWR VGND sg13g2_decap_8
XFILLER_37_723 VPWR VGND sg13g2_decap_8
XFILLER_25_907 VPWR VGND sg13g2_decap_8
XFILLER_36_244 VPWR VGND sg13g2_decap_8
XFILLER_18_970 VPWR VGND sg13g2_decap_8
XFILLER_24_439 VPWR VGND sg13g2_decap_8
XFILLER_33_951 VPWR VGND sg13g2_decap_8
XFILLER_20_612 VPWR VGND sg13g2_decap_8
XFILLER_22_18 VPWR VGND sg13g2_decap_8
XFILLER_32_494 VPWR VGND sg13g2_decap_8
XFILLER_20_689 VPWR VGND sg13g2_decap_8
XFILLER_16_907 VPWR VGND sg13g2_decap_8
XFILLER_27_233 VPWR VGND sg13g2_decap_8
XFILLER_28_756 VPWR VGND sg13g2_decap_8
XFILLER_15_417 VPWR VGND sg13g2_decap_8
XFILLER_43_748 VPWR VGND sg13g2_decap_8
XFILLER_42_269 VPWR VGND sg13g2_fill_1
XFILLER_24_951 VPWR VGND sg13g2_decap_8
XFILLER_11_634 VPWR VGND sg13g2_decap_8
XFILLER_10_166 VPWR VGND sg13g2_decap_8
XFILLER_7_638 VPWR VGND sg13g2_decap_8
XFILLER_12_62 VPWR VGND sg13g2_decap_8
XFILLER_3_811 VPWR VGND sg13g2_decap_8
XFILLER_2_321 VPWR VGND sg13g2_decap_8
XFILLER_3_888 VPWR VGND sg13g2_decap_8
XFILLER_38_509 VPWR VGND sg13g2_decap_8
XFILLER_19_734 VPWR VGND sg13g2_decap_8
XFILLER_46_564 VPWR VGND sg13g2_decap_8
XFILLER_18_299 VPWR VGND sg13g2_decap_8
XFILLER_34_748 VPWR VGND sg13g2_decap_8
XFILLER_18_1012 VPWR VGND sg13g2_decap_8
XFILLER_42_792 VPWR VGND sg13g2_decap_8
XFILLER_14_461 VPWR VGND sg13g2_decap_8
XFILLER_15_995 VPWR VGND sg13g2_decap_8
X_418_ net149 _112_ VPWR VGND sg13g2_buf_1
X_349_ _205_ net117 net53 VPWR VGND sg13g2_nand2_1
XFILLER_30_976 VPWR VGND sg13g2_decap_8
XFILLER_25_1005 VPWR VGND sg13g2_decap_8
XFILLER_49_380 VPWR VGND sg13g2_decap_8
XFILLER_37_520 VPWR VGND sg13g2_decap_8
XFILLER_25_704 VPWR VGND sg13g2_decap_8
XFILLER_24_236 VPWR VGND sg13g2_decap_8
XFILLER_37_597 VPWR VGND sg13g2_decap_8
XFILLER_21_932 VPWR VGND sg13g2_decap_8
XFILLER_40_729 VPWR VGND sg13g2_decap_8
XFILLER_20_486 VPWR VGND sg13g2_decap_8
XFILLER_4_619 VPWR VGND sg13g2_decap_8
XFILLER_0_847 VPWR VGND sg13g2_decap_8
XFILLER_48_818 VPWR VGND sg13g2_decap_8
XFILLER_47_339 VPWR VGND sg13g2_decap_8
XFILLER_16_704 VPWR VGND sg13g2_decap_8
XFILLER_28_553 VPWR VGND sg13g2_decap_8
XFILLER_15_214 VPWR VGND sg13g2_fill_1
XFILLER_43_545 VPWR VGND sg13g2_decap_8
XFILLER_12_921 VPWR VGND sg13g2_decap_8
XFILLER_11_442 VPWR VGND sg13g2_decap_8
XFILLER_30_239 VPWR VGND sg13g2_decap_8
XFILLER_12_998 VPWR VGND sg13g2_decap_8
XFILLER_23_61 VPWR VGND sg13g2_fill_1
XFILLER_8_958 VPWR VGND sg13g2_decap_8
XFILLER_7_457 VPWR VGND sg13g2_fill_2
XFILLER_23_94 VPWR VGND sg13g2_decap_8
XFILLER_3_685 VPWR VGND sg13g2_decap_8
XFILLER_47_840 VPWR VGND sg13g2_decap_8
XFILLER_48_91 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_46_394 VPWR VGND sg13g2_decap_8
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_22_718 VPWR VGND sg13g2_decap_8
XFILLER_34_545 VPWR VGND sg13g2_decap_8
XFILLER_21_228 VPWR VGND sg13g2_fill_2
XFILLER_15_792 VPWR VGND sg13g2_decap_8
XFILLER_30_773 VPWR VGND sg13g2_decap_8
XFILLER_29_306 VPWR VGND sg13g2_decap_8
XFILLER_38_873 VPWR VGND sg13g2_decap_8
XFILLER_37_383 VPWR VGND sg13g2_decap_8
XFILLER_44_49 VPWR VGND sg13g2_decap_8
XFILLER_13_718 VPWR VGND sg13g2_decap_8
XFILLER_25_578 VPWR VGND sg13g2_decap_8
XFILLER_40_515 VPWR VGND sg13g2_fill_2
XFILLER_40_526 VPWR VGND sg13g2_decap_8
XFILLER_12_239 VPWR VGND sg13g2_decap_8
XFILLER_5_906 VPWR VGND sg13g2_decap_8
XFILLER_0_644 VPWR VGND sg13g2_decap_8
XFILLER_48_615 VPWR VGND sg13g2_decap_8
XFILLER_29_862 VPWR VGND sg13g2_decap_8
XFILLER_44_843 VPWR VGND sg13g2_decap_8
XFILLER_28_383 VPWR VGND sg13g2_decap_8
XFILLER_43_386 VPWR VGND sg13g2_decap_8
XFILLER_16_578 VPWR VGND sg13g2_fill_1
XFILLER_31_559 VPWR VGND sg13g2_decap_8
XFILLER_34_82 VPWR VGND sg13g2_decap_8
XFILLER_8_755 VPWR VGND sg13g2_decap_8
XFILLER_7_210 VPWR VGND sg13g2_decap_8
XFILLER_11_283 VPWR VGND sg13g2_decap_8
XFILLER_12_795 VPWR VGND sg13g2_decap_8
XFILLER_7_265 VPWR VGND sg13g2_decap_8
XFILLER_4_983 VPWR VGND sg13g2_decap_8
XFILLER_3_471 VPWR VGND sg13g2_decap_8
XFILLER_22_4 VPWR VGND sg13g2_decap_8
XFILLER_22_1019 VPWR VGND sg13g2_decap_8
XFILLER_39_637 VPWR VGND sg13g2_decap_8
XFILLER_35_865 VPWR VGND sg13g2_decap_8
XFILLER_22_515 VPWR VGND sg13g2_decap_8
XFILLER_30_570 VPWR VGND sg13g2_decap_8
XFILLER_45_618 VPWR VGND sg13g2_decap_8
XFILLER_29_158 VPWR VGND sg13g2_decap_8
XFILLER_38_670 VPWR VGND sg13g2_decap_8
XFILLER_44_139 VPWR VGND sg13g2_decap_8
XFILLER_26_865 VPWR VGND sg13g2_decap_8
XFILLER_37_191 VPWR VGND sg13g2_decap_8
XFILLER_41_813 VPWR VGND sg13g2_decap_8
XFILLER_13_548 VPWR VGND sg13g2_decap_4
XFILLER_40_312 VPWR VGND sg13g2_decap_8
XFILLER_9_519 VPWR VGND sg13g2_fill_2
XFILLER_5_703 VPWR VGND sg13g2_decap_8
XFILLER_20_95 VPWR VGND sg13g2_decap_8
XFILLER_0_441 VPWR VGND sg13g2_decap_8
XFILLER_1_964 VPWR VGND sg13g2_decap_8
XFILLER_49_968 VPWR VGND sg13g2_decap_8
Xhold71 DP_4.matrix\[63\] VPWR VGND net121 sg13g2_dlygate4sd3_1
Xhold82 DP_3.matrix\[0\] VPWR VGND net132 sg13g2_dlygate4sd3_1
Xhold60 _024_ VPWR VGND net110 sg13g2_dlygate4sd3_1
XFILLER_36_618 VPWR VGND sg13g2_decap_8
XFILLER_48_489 VPWR VGND sg13g2_decap_8
XFILLER_17_810 VPWR VGND sg13g2_decap_8
XFILLER_35_117 VPWR VGND sg13g2_decap_8
Xhold93 DP_4.matrix\[54\] VPWR VGND net143 sg13g2_dlygate4sd3_1
XFILLER_44_640 VPWR VGND sg13g2_decap_8
XFILLER_17_887 VPWR VGND sg13g2_decap_8
XFILLER_31_301 VPWR VGND sg13g2_decap_8
XFILLER_32_802 VPWR VGND sg13g2_decap_8
X_597_ net83 VGND VPWR _137_ DP_4.matrix\[55\] clknet_5_31__leaf_clk sg13g2_dfrbpq_1
XFILLER_31_378 VPWR VGND sg13g2_decap_8
XFILLER_32_879 VPWR VGND sg13g2_decap_8
XFILLER_12_570 VPWR VGND sg13g2_fill_2
Xclkbuf_4_14_0_clk clknet_0_clk clknet_4_14_0_clk VPWR VGND sg13g2_buf_8
XFILLER_40_890 VPWR VGND sg13g2_decap_8
XFILLER_8_552 VPWR VGND sg13g2_decap_8
XFILLER_12_592 VPWR VGND sg13g2_decap_8
XFILLER_6_53 VPWR VGND sg13g2_decap_8
XFILLER_4_780 VPWR VGND sg13g2_decap_8
XFILLER_25_18 VPWR VGND sg13g2_decap_8
XFILLER_35_662 VPWR VGND sg13g2_decap_8
XFILLER_23_835 VPWR VGND sg13g2_decap_8
XFILLER_34_194 VPWR VGND sg13g2_fill_2
XFILLER_22_367 VPWR VGND sg13g2_decap_8
XFILLER_10_529 VPWR VGND sg13g2_decap_8
XFILLER_46_949 VPWR VGND sg13g2_decap_8
XFILLER_45_415 VPWR VGND sg13g2_decap_8
X_520_ net79 VGND VPWR net190 mac2.sum_lvl2_ff\[5\] clknet_5_13__leaf_clk sg13g2_dfrbpq_1
XFILLER_26_662 VPWR VGND sg13g2_decap_8
X_451_ net81 VGND VPWR _045_ mac1.products_ff\[18\] clknet_5_26__leaf_clk sg13g2_dfrbpq_1
XFILLER_13_334 VPWR VGND sg13g2_fill_1
X_382_ net117 _076_ VPWR VGND sg13g2_buf_1
XFILLER_41_610 VPWR VGND sg13g2_decap_8
XFILLER_14_868 VPWR VGND sg13g2_decap_8
XFILLER_40_131 VPWR VGND sg13g2_decap_8
XFILLER_9_338 VPWR VGND sg13g2_decap_4
XFILLER_13_389 VPWR VGND sg13g2_decap_8
XFILLER_41_687 VPWR VGND sg13g2_decap_8
Xoutput4 net4 uo_out[3] VPWR VGND sg13g2_buf_1
XFILLER_1_761 VPWR VGND sg13g2_decap_8
XFILLER_49_765 VPWR VGND sg13g2_decap_8
XFILLER_48_253 VPWR VGND sg13g2_decap_4
XFILLER_37_905 VPWR VGND sg13g2_decap_8
XFILLER_36_448 VPWR VGND sg13g2_decap_8
XFILLER_45_982 VPWR VGND sg13g2_decap_8
XFILLER_16_183 VPWR VGND sg13g2_fill_2
XFILLER_17_684 VPWR VGND sg13g2_decap_8
XFILLER_16_194 VPWR VGND sg13g2_fill_1
XFILLER_32_676 VPWR VGND sg13g2_decap_8
XFILLER_31_175 VPWR VGND sg13g2_decap_8
XFILLER_9_850 VPWR VGND sg13g2_decap_8
XFILLER_39_253 VPWR VGND sg13g2_fill_2
XFILLER_28_938 VPWR VGND sg13g2_decap_8
XFILLER_27_459 VPWR VGND sg13g2_decap_8
XFILLER_42_407 VPWR VGND sg13g2_decap_8
XFILLER_36_982 VPWR VGND sg13g2_decap_8
XFILLER_23_632 VPWR VGND sg13g2_decap_8
XFILLER_11_816 VPWR VGND sg13g2_decap_8
XFILLER_10_359 VPWR VGND sg13g2_decap_8
XFILLER_19_916 VPWR VGND sg13g2_decap_8
XFILLER_45_201 VPWR VGND sg13g2_decap_4
XFILLER_18_404 VPWR VGND sg13g2_decap_8
XFILLER_46_746 VPWR VGND sg13g2_decap_8
XFILLER_45_234 VPWR VGND sg13g2_decap_8
XFILLER_18_459 VPWR VGND sg13g2_fill_2
XFILLER_45_278 VPWR VGND sg13g2_decap_8
XFILLER_27_960 VPWR VGND sg13g2_decap_8
X_503_ net82 VGND VPWR _034_ mac2.products_ff\[119\] clknet_5_27__leaf_clk sg13g2_dfrbpq_1
X_434_ net130 _128_ VPWR VGND sg13g2_buf_1
XFILLER_42_974 VPWR VGND sg13g2_decap_8
XFILLER_14_665 VPWR VGND sg13g2_decap_8
XFILLER_9_102 VPWR VGND sg13g2_decap_8
XFILLER_13_175 VPWR VGND sg13g2_decap_8
X_365_ _215_ net149 net49 VPWR VGND sg13g2_nand2_1
X_296_ mac2.sum_lvl3_ff\[1\] net170 _175_ VPWR VGND sg13g2_xor2_1
XFILLER_9_179 VPWR VGND sg13g2_decap_8
XFILLER_10_893 VPWR VGND sg13g2_decap_8
XFILLER_6_886 VPWR VGND sg13g2_decap_8
XFILLER_5_352 VPWR VGND sg13g2_decap_8
XFILLER_3_32 VPWR VGND sg13g2_decap_8
XFILLER_49_562 VPWR VGND sg13g2_decap_8
XFILLER_37_702 VPWR VGND sg13g2_decap_8
XFILLER_36_223 VPWR VGND sg13g2_decap_8
XFILLER_24_418 VPWR VGND sg13g2_decap_8
XFILLER_37_779 VPWR VGND sg13g2_decap_8
XFILLER_17_492 VPWR VGND sg13g2_fill_1
XFILLER_33_930 VPWR VGND sg13g2_decap_8
XFILLER_32_473 VPWR VGND sg13g2_decap_8
XFILLER_20_668 VPWR VGND sg13g2_decap_8
Xclkbuf_5_28__f_clk clknet_4_14_0_clk clknet_5_28__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_47_49 VPWR VGND sg13g2_decap_8
XFILLER_28_735 VPWR VGND sg13g2_decap_8
XFILLER_43_727 VPWR VGND sg13g2_decap_8
XFILLER_24_930 VPWR VGND sg13g2_decap_8
XFILLER_27_289 VPWR VGND sg13g2_decap_8
XFILLER_42_248 VPWR VGND sg13g2_decap_8
XFILLER_11_613 VPWR VGND sg13g2_decap_8
XFILLER_23_462 VPWR VGND sg13g2_decap_8
XFILLER_10_145 VPWR VGND sg13g2_decap_8
XFILLER_7_617 VPWR VGND sg13g2_decap_8
XFILLER_6_116 VPWR VGND sg13g2_decap_4
XFILLER_6_149 VPWR VGND sg13g2_fill_1
XFILLER_6_138 VPWR VGND sg13g2_decap_8
XFILLER_12_41 VPWR VGND sg13g2_decap_8
XFILLER_2_300 VPWR VGND sg13g2_decap_8
XFILLER_3_867 VPWR VGND sg13g2_decap_8
XFILLER_19_713 VPWR VGND sg13g2_decap_8
XFILLER_46_543 VPWR VGND sg13g2_decap_8
XFILLER_37_71 VPWR VGND sg13g2_decap_8
XFILLER_18_278 VPWR VGND sg13g2_decap_8
XFILLER_34_727 VPWR VGND sg13g2_decap_8
XFILLER_14_440 VPWR VGND sg13g2_decap_8
X_417_ net56 _111_ VPWR VGND sg13g2_buf_1
XFILLER_42_771 VPWR VGND sg13g2_decap_8
XFILLER_15_974 VPWR VGND sg13g2_decap_8
X_348_ _204_ net160 net47 VPWR VGND sg13g2_nand2_1
XFILLER_30_955 VPWR VGND sg13g2_decap_8
XFILLER_10_690 VPWR VGND sg13g2_decap_8
X_279_ _007_ _164_ _165_ VPWR VGND sg13g2_xnor2_1
XFILLER_6_683 VPWR VGND sg13g2_decap_8
XFILLER_5_182 VPWR VGND sg13g2_decap_8
XFILLER_25_1028 VPWR VGND sg13g2_fill_1
XFILLER_37_576 VPWR VGND sg13g2_decap_8
XFILLER_24_215 VPWR VGND sg13g2_decap_8
XFILLER_40_708 VPWR VGND sg13g2_decap_8
XFILLER_21_911 VPWR VGND sg13g2_decap_8
XFILLER_32_281 VPWR VGND sg13g2_decap_8
XFILLER_20_465 VPWR VGND sg13g2_decap_8
XFILLER_21_988 VPWR VGND sg13g2_decap_8
XFILLER_0_826 VPWR VGND sg13g2_decap_8
XFILLER_47_318 VPWR VGND sg13g2_decap_8
XFILLER_28_532 VPWR VGND sg13g2_decap_8
XFILLER_43_524 VPWR VGND sg13g2_decap_8
XFILLER_15_259 VPWR VGND sg13g2_decap_8
XFILLER_12_900 VPWR VGND sg13g2_decap_8
XFILLER_30_218 VPWR VGND sg13g2_decap_8
XFILLER_8_937 VPWR VGND sg13g2_decap_8
XFILLER_12_977 VPWR VGND sg13g2_decap_8
XFILLER_7_436 VPWR VGND sg13g2_decap_8
XFILLER_48_1028 VPWR VGND sg13g2_fill_1
XFILLER_3_664 VPWR VGND sg13g2_decap_8
XFILLER_2_130 VPWR VGND sg13g2_decap_8
XFILLER_2_174 VPWR VGND sg13g2_fill_1
Xclkbuf_5_11__f_clk clknet_4_5_0_clk clknet_5_11__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_48_70 VPWR VGND sg13g2_decap_8
XFILLER_39_819 VPWR VGND sg13g2_decap_8
XFILLER_17_7 VPWR VGND sg13g2_decap_8
XFILLER_0_1008 VPWR VGND sg13g2_decap_8
XFILLER_47_896 VPWR VGND sg13g2_decap_8
XFILLER_46_373 VPWR VGND sg13g2_decap_8
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_19_587 VPWR VGND sg13g2_decap_8
XFILLER_34_524 VPWR VGND sg13g2_decap_8
XFILLER_15_771 VPWR VGND sg13g2_decap_8
XFILLER_30_752 VPWR VGND sg13g2_decap_8
XFILLER_31_1021 VPWR VGND sg13g2_decap_8
XFILLER_7_981 VPWR VGND sg13g2_decap_8
XFILLER_43_0 VPWR VGND sg13g2_decap_8
XFILLER_9_1011 VPWR VGND sg13g2_decap_8
XFILLER_28_18 VPWR VGND sg13g2_decap_8
XFILLER_29_329 VPWR VGND sg13g2_fill_1
XFILLER_38_852 VPWR VGND sg13g2_decap_8
XFILLER_37_362 VPWR VGND sg13g2_decap_8
XFILLER_44_28 VPWR VGND sg13g2_decap_8
XFILLER_25_557 VPWR VGND sg13g2_decap_8
XFILLER_12_218 VPWR VGND sg13g2_decap_8
XFILLER_20_284 VPWR VGND sg13g2_decap_8
XFILLER_21_785 VPWR VGND sg13g2_decap_8
XFILLER_0_623 VPWR VGND sg13g2_decap_8
XFILLER_29_841 VPWR VGND sg13g2_decap_8
XFILLER_47_148 VPWR VGND sg13g2_decap_8
XFILLER_44_822 VPWR VGND sg13g2_decap_8
XFILLER_28_362 VPWR VGND sg13g2_decap_8
XFILLER_44_899 VPWR VGND sg13g2_decap_8
XFILLER_43_365 VPWR VGND sg13g2_decap_8
XFILLER_31_538 VPWR VGND sg13g2_decap_8
XFILLER_34_61 VPWR VGND sg13g2_decap_8
XFILLER_12_774 VPWR VGND sg13g2_decap_8
XFILLER_15_1016 VPWR VGND sg13g2_decap_8
XFILLER_15_1027 VPWR VGND sg13g2_fill_2
XFILLER_8_734 VPWR VGND sg13g2_decap_8
XFILLER_11_251 VPWR VGND sg13g2_decap_8
XFILLER_7_244 VPWR VGND sg13g2_decap_8
XFILLER_4_962 VPWR VGND sg13g2_decap_8
XFILLER_3_450 VPWR VGND sg13g2_decap_8
XFILLER_39_616 VPWR VGND sg13g2_decap_8
XFILLER_15_4 VPWR VGND sg13g2_decap_8
XFILLER_38_104 VPWR VGND sg13g2_decap_4
XFILLER_47_693 VPWR VGND sg13g2_decap_8
XFILLER_34_310 VPWR VGND sg13g2_decap_8
XFILLER_35_844 VPWR VGND sg13g2_decap_8
XFILLER_34_365 VPWR VGND sg13g2_decap_8
XFILLER_44_107 VPWR VGND sg13g2_decap_8
XFILLER_26_844 VPWR VGND sg13g2_decap_8
XFILLER_37_170 VPWR VGND sg13g2_decap_8
XFILLER_25_365 VPWR VGND sg13g2_decap_4
XFILLER_38_1027 VPWR VGND sg13g2_fill_2
XFILLER_13_527 VPWR VGND sg13g2_decap_8
XFILLER_40_357 VPWR VGND sg13g2_decap_8
XFILLER_41_869 VPWR VGND sg13g2_decap_8
XFILLER_21_560 VPWR VGND sg13g2_fill_1
XFILLER_5_759 VPWR VGND sg13g2_decap_8
XFILLER_20_74 VPWR VGND sg13g2_decap_8
XFILLER_0_420 VPWR VGND sg13g2_decap_8
XFILLER_1_943 VPWR VGND sg13g2_decap_8
XFILLER_49_947 VPWR VGND sg13g2_decap_8
Xhold50 _008_ VPWR VGND net100 sg13g2_dlygate4sd3_1
XFILLER_0_497 VPWR VGND sg13g2_decap_8
XFILLER_29_61 VPWR VGND sg13g2_decap_8
XFILLER_48_468 VPWR VGND sg13g2_decap_8
Xhold83 DP_1.matrix\[72\] VPWR VGND net133 sg13g2_dlygate4sd3_1
Xhold72 DP_2.matrix\[36\] VPWR VGND net122 sg13g2_dlygate4sd3_1
Xhold61 mac1.products_ff\[51\] VPWR VGND net111 sg13g2_dlygate4sd3_1
Xhold94 DP_3.matrix\[54\] VPWR VGND net144 sg13g2_dlygate4sd3_1
XFILLER_17_866 VPWR VGND sg13g2_decap_8
XFILLER_16_376 VPWR VGND sg13g2_decap_4
X_596_ net84 VGND VPWR _136_ DP_4.matrix\[54\] clknet_5_28__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_696 VPWR VGND sg13g2_decap_8
XFILLER_43_173 VPWR VGND sg13g2_decap_8
XFILLER_31_324 VPWR VGND sg13g2_fill_1
XFILLER_32_858 VPWR VGND sg13g2_decap_8
XFILLER_31_357 VPWR VGND sg13g2_decap_8
XFILLER_8_531 VPWR VGND sg13g2_decap_8
XFILLER_6_32 VPWR VGND sg13g2_decap_8
Xclkbuf_5_9__f_clk clknet_4_4_0_clk clknet_5_9__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_39_413 VPWR VGND sg13g2_decap_8
XFILLER_39_468 VPWR VGND sg13g2_decap_4
XFILLER_47_490 VPWR VGND sg13g2_decap_8
XFILLER_26_129 VPWR VGND sg13g2_decap_8
XFILLER_35_641 VPWR VGND sg13g2_decap_8
XFILLER_23_814 VPWR VGND sg13g2_decap_8
XFILLER_22_302 VPWR VGND sg13g2_fill_2
XFILLER_10_508 VPWR VGND sg13g2_decap_8
XFILLER_22_346 VPWR VGND sg13g2_decap_8
XFILLER_46_928 VPWR VGND sg13g2_decap_8
XFILLER_39_980 VPWR VGND sg13g2_decap_8
XFILLER_17_129 VPWR VGND sg13g2_fill_1
XFILLER_26_641 VPWR VGND sg13g2_decap_8
X_450_ net74 VGND VPWR _044_ mac1.products_ff\[17\] clknet_5_25__leaf_clk sg13g2_dfrbpq_1
XFILLER_13_302 VPWR VGND sg13g2_decap_8
X_381_ net55 _075_ VPWR VGND sg13g2_buf_1
XFILLER_14_847 VPWR VGND sg13g2_decap_8
XFILLER_25_184 VPWR VGND sg13g2_decap_8
XFILLER_9_306 VPWR VGND sg13g2_fill_2
XFILLER_41_666 VPWR VGND sg13g2_decap_8
XFILLER_15_85 VPWR VGND sg13g2_decap_8
XFILLER_12_1019 VPWR VGND sg13g2_decap_8
XFILLER_31_84 VPWR VGND sg13g2_decap_8
XFILLER_1_740 VPWR VGND sg13g2_decap_8
XFILLER_49_744 VPWR VGND sg13g2_decap_8
XFILLER_48_232 VPWR VGND sg13g2_decap_8
XFILLER_0_294 VPWR VGND sg13g2_decap_8
XFILLER_45_961 VPWR VGND sg13g2_decap_8
XFILLER_17_663 VPWR VGND sg13g2_decap_8
XFILLER_44_493 VPWR VGND sg13g2_decap_8
XFILLER_16_162 VPWR VGND sg13g2_decap_8
XFILLER_32_655 VPWR VGND sg13g2_decap_8
X_579_ net83 VGND VPWR _119_ DP_3.matrix\[55\] clknet_5_29__leaf_clk sg13g2_dfrbpq_1
XFILLER_31_154 VPWR VGND sg13g2_decap_8
XFILLER_8_383 VPWR VGND sg13g2_decap_4
XFILLER_28_1015 VPWR VGND sg13g2_decap_8
XFILLER_39_210 VPWR VGND sg13g2_decap_8
XFILLER_39_221 VPWR VGND sg13g2_fill_1
XFILLER_28_917 VPWR VGND sg13g2_decap_8
XFILLER_43_909 VPWR VGND sg13g2_decap_8
XFILLER_27_438 VPWR VGND sg13g2_decap_8
XFILLER_36_961 VPWR VGND sg13g2_decap_8
XFILLER_23_611 VPWR VGND sg13g2_decap_8
XFILLER_35_1019 VPWR VGND sg13g2_decap_8
XFILLER_10_305 VPWR VGND sg13g2_fill_1
XFILLER_22_176 VPWR VGND sg13g2_decap_8
XFILLER_23_688 VPWR VGND sg13g2_decap_8
XFILLER_10_338 VPWR VGND sg13g2_decap_8
Xclkbuf_4_13_0_clk clknet_0_clk clknet_4_13_0_clk VPWR VGND sg13g2_buf_8
XFILLER_46_725 VPWR VGND sg13g2_decap_8
XFILLER_18_438 VPWR VGND sg13g2_decap_8
XFILLER_34_909 VPWR VGND sg13g2_decap_8
X_502_ net84 VGND VPWR _063_ mac2.products_ff\[103\] clknet_5_31__leaf_clk sg13g2_dfrbpq_1
X_433_ net42 _127_ VPWR VGND sg13g2_buf_1
XFILLER_42_953 VPWR VGND sg13g2_decap_8
XFILLER_14_644 VPWR VGND sg13g2_decap_8
X_364_ _214_ net155 net50 VPWR VGND sg13g2_nand2_1
XFILLER_9_158 VPWR VGND sg13g2_decap_8
X_295_ net170 mac2.sum_lvl3_ff\[1\] _174_ VPWR VGND sg13g2_nor2_1
XFILLER_42_94 VPWR VGND sg13g2_decap_8
XFILLER_10_872 VPWR VGND sg13g2_decap_8
XFILLER_5_331 VPWR VGND sg13g2_decap_8
XFILLER_6_865 VPWR VGND sg13g2_decap_8
XFILLER_47_7 VPWR VGND sg13g2_decap_8
XFILLER_3_11 VPWR VGND sg13g2_decap_8
XFILLER_49_541 VPWR VGND sg13g2_decap_8
XFILLER_36_202 VPWR VGND sg13g2_decap_8
XFILLER_3_1028 VPWR VGND sg13g2_fill_1
XFILLER_37_758 VPWR VGND sg13g2_decap_8
XFILLER_44_290 VPWR VGND sg13g2_decap_8
XFILLER_32_452 VPWR VGND sg13g2_decap_8
XFILLER_33_986 VPWR VGND sg13g2_decap_8
XFILLER_20_647 VPWR VGND sg13g2_decap_8
XFILLER_47_28 VPWR VGND sg13g2_decap_8
XFILLER_28_714 VPWR VGND sg13g2_decap_8
XFILLER_41_1023 VPWR VGND sg13g2_decap_4
XFILLER_43_706 VPWR VGND sg13g2_decap_8
XFILLER_27_268 VPWR VGND sg13g2_decap_8
XFILLER_42_227 VPWR VGND sg13g2_decap_8
XFILLER_24_986 VPWR VGND sg13g2_decap_8
XFILLER_10_124 VPWR VGND sg13g2_decap_8
XFILLER_11_669 VPWR VGND sg13g2_decap_8
XFILLER_12_97 VPWR VGND sg13g2_decap_8
XFILLER_3_846 VPWR VGND sg13g2_decap_8
XFILLER_2_356 VPWR VGND sg13g2_decap_8
XFILLER_46_522 VPWR VGND sg13g2_decap_8
XFILLER_18_202 VPWR VGND sg13g2_decap_8
XFILLER_37_50 VPWR VGND sg13g2_decap_8
XFILLER_18_257 VPWR VGND sg13g2_decap_8
XFILLER_19_769 VPWR VGND sg13g2_decap_8
XFILLER_34_706 VPWR VGND sg13g2_decap_8
XFILLER_46_599 VPWR VGND sg13g2_decap_8
XFILLER_33_227 VPWR VGND sg13g2_decap_8
XFILLER_42_750 VPWR VGND sg13g2_decap_8
XFILLER_15_953 VPWR VGND sg13g2_decap_8
XFILLER_33_238 VPWR VGND sg13g2_fill_1
X_416_ net148 _110_ VPWR VGND sg13g2_buf_1
X_347_ _203_ _202_ _047_ VPWR VGND sg13g2_xor2_1
XFILLER_30_934 VPWR VGND sg13g2_decap_8
X_278_ mac1.products_ff\[69\] mac1.products_ff\[86\] _165_ VPWR VGND sg13g2_xor2_1
XFILLER_6_662 VPWR VGND sg13g2_decap_8
XFILLER_5_161 VPWR VGND sg13g2_decap_8
XFILLER_37_555 VPWR VGND sg13g2_decap_8
XFILLER_25_739 VPWR VGND sg13g2_decap_8
XFILLER_33_783 VPWR VGND sg13g2_decap_8
XFILLER_20_444 VPWR VGND sg13g2_decap_8
XFILLER_21_967 VPWR VGND sg13g2_decap_8
XFILLER_0_805 VPWR VGND sg13g2_decap_8
XFILLER_43_503 VPWR VGND sg13g2_decap_8
XFILLER_15_205 VPWR VGND sg13g2_decap_8
XFILLER_16_739 VPWR VGND sg13g2_decap_8
XFILLER_28_588 VPWR VGND sg13g2_decap_8
XFILLER_15_238 VPWR VGND sg13g2_decap_8
XFILLER_12_956 VPWR VGND sg13g2_decap_8
XFILLER_23_282 VPWR VGND sg13g2_decap_8
XFILLER_24_783 VPWR VGND sg13g2_decap_8
XFILLER_8_916 VPWR VGND sg13g2_decap_8
XFILLER_7_415 VPWR VGND sg13g2_decap_8
XFILLER_23_52 VPWR VGND sg13g2_decap_8
XFILLER_11_477 VPWR VGND sg13g2_decap_8
XFILLER_7_459 VPWR VGND sg13g2_fill_1
XFILLER_48_1007 VPWR VGND sg13g2_decap_8
XFILLER_3_643 VPWR VGND sg13g2_decap_8
XFILLER_38_319 VPWR VGND sg13g2_decap_8
XFILLER_19_533 VPWR VGND sg13g2_fill_2
XFILLER_47_875 VPWR VGND sg13g2_decap_8
XFILLER_19_566 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_15_750 VPWR VGND sg13g2_decap_8
XFILLER_21_219 VPWR VGND sg13g2_fill_1
XFILLER_30_731 VPWR VGND sg13g2_decap_8
XFILLER_9_76 VPWR VGND sg13g2_decap_4
XFILLER_14_293 VPWR VGND sg13g2_decap_8
XFILLER_31_1000 VPWR VGND sg13g2_decap_8
XFILLER_7_960 VPWR VGND sg13g2_decap_8
XFILLER_6_481 VPWR VGND sg13g2_fill_1
XFILLER_36_0 VPWR VGND sg13g2_decap_8
XFILLER_38_831 VPWR VGND sg13g2_decap_8
XFILLER_25_536 VPWR VGND sg13g2_decap_8
XFILLER_33_580 VPWR VGND sg13g2_decap_8
XFILLER_21_764 VPWR VGND sg13g2_decap_8
XFILLER_20_263 VPWR VGND sg13g2_decap_8
XFILLER_4_429 VPWR VGND sg13g2_decap_8
XFILLER_0_602 VPWR VGND sg13g2_decap_8
XFILLER_0_679 VPWR VGND sg13g2_decap_8
XFILLER_29_820 VPWR VGND sg13g2_decap_8
XFILLER_44_801 VPWR VGND sg13g2_decap_8
XFILLER_18_74 VPWR VGND sg13g2_decap_8
XFILLER_29_897 VPWR VGND sg13g2_decap_8
XFILLER_43_344 VPWR VGND sg13g2_decap_8
XFILLER_44_878 VPWR VGND sg13g2_decap_8
XFILLER_31_517 VPWR VGND sg13g2_decap_8
XFILLER_24_580 VPWR VGND sg13g2_decap_8
XFILLER_34_51 VPWR VGND sg13g2_fill_1
XFILLER_8_713 VPWR VGND sg13g2_decap_8
XFILLER_11_230 VPWR VGND sg13g2_decap_8
XFILLER_12_753 VPWR VGND sg13g2_decap_8
XFILLER_4_941 VPWR VGND sg13g2_decap_8
XFILLER_38_138 VPWR VGND sg13g2_decap_8
XFILLER_47_672 VPWR VGND sg13g2_decap_8
XFILLER_35_823 VPWR VGND sg13g2_decap_8
XFILLER_19_385 VPWR VGND sg13g2_decap_8
XFILLER_34_344 VPWR VGND sg13g2_decap_8
XFILLER_26_823 VPWR VGND sg13g2_decap_8
XFILLER_13_506 VPWR VGND sg13g2_decap_8
XFILLER_25_344 VPWR VGND sg13g2_decap_8
XFILLER_38_1006 VPWR VGND sg13g2_decap_8
XFILLER_41_848 VPWR VGND sg13g2_decap_8
XFILLER_5_738 VPWR VGND sg13g2_decap_8
XFILLER_20_53 VPWR VGND sg13g2_decap_8
XFILLER_1_922 VPWR VGND sg13g2_decap_8
XFILLER_49_926 VPWR VGND sg13g2_decap_8
Xhold40 DP_2.matrix\[55\] VPWR VGND net90 sg13g2_dlygate4sd3_1
XFILLER_0_476 VPWR VGND sg13g2_decap_8
XFILLER_1_999 VPWR VGND sg13g2_decap_8
XFILLER_48_447 VPWR VGND sg13g2_decap_8
Xhold62 _004_ VPWR VGND net112 sg13g2_dlygate4sd3_1
Xhold51 DP_4.matrix\[1\] VPWR VGND net101 sg13g2_dlygate4sd3_1
Xhold73 mac2.products_ff\[102\] VPWR VGND net123 sg13g2_dlygate4sd3_1
Xhold84 DP_1.matrix\[18\] VPWR VGND net134 sg13g2_dlygate4sd3_1
Xhold95 mac1.sum_lvl1_ff\[0\] VPWR VGND net145 sg13g2_dlygate4sd3_1
XFILLER_17_845 VPWR VGND sg13g2_decap_8
XFILLER_29_694 VPWR VGND sg13g2_decap_8
X_595_ net80 VGND VPWR _135_ DP_4.matrix\[46\] clknet_5_15__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_675 VPWR VGND sg13g2_decap_8
XFILLER_43_141 VPWR VGND sg13g2_decap_8
XFILLER_16_355 VPWR VGND sg13g2_decap_8
XFILLER_43_163 VPWR VGND sg13g2_fill_1
XFILLER_32_837 VPWR VGND sg13g2_decap_8
XFILLER_43_196 VPWR VGND sg13g2_decap_8
XFILLER_8_587 VPWR VGND sg13g2_decap_8
XFILLER_6_11 VPWR VGND sg13g2_decap_8
XFILLER_6_88 VPWR VGND sg13g2_decap_8
XFILLER_3_292 VPWR VGND sg13g2_decap_8
XFILLER_6_1026 VPWR VGND sg13g2_fill_2
XFILLER_26_108 VPWR VGND sg13g2_decap_8
XFILLER_35_620 VPWR VGND sg13g2_decap_8
XFILLER_19_193 VPWR VGND sg13g2_decap_8
XFILLER_35_697 VPWR VGND sg13g2_decap_8
XFILLER_34_196 VPWR VGND sg13g2_fill_1
XFILLER_31_881 VPWR VGND sg13g2_decap_8
XFILLER_2_719 VPWR VGND sg13g2_decap_8
XFILLER_1_229 VPWR VGND sg13g2_decap_8
XFILLER_46_907 VPWR VGND sg13g2_decap_8
Xheichips25_template_20 VPWR VGND uio_oe[3] sg13g2_tiehi
XFILLER_26_620 VPWR VGND sg13g2_decap_8
XFILLER_14_826 VPWR VGND sg13g2_decap_8
X_380_ net134 _074_ VPWR VGND sg13g2_buf_1
XFILLER_25_163 VPWR VGND sg13g2_decap_8
XFILLER_26_697 VPWR VGND sg13g2_decap_8
XFILLER_13_358 VPWR VGND sg13g2_decap_8
XFILLER_41_645 VPWR VGND sg13g2_decap_8
XFILLER_9_318 VPWR VGND sg13g2_decap_8
XFILLER_40_166 VPWR VGND sg13g2_decap_8
XFILLER_5_513 VPWR VGND sg13g2_decap_8
XFILLER_5_546 VPWR VGND sg13g2_decap_8
XFILLER_31_63 VPWR VGND sg13g2_decap_8
XFILLER_49_723 VPWR VGND sg13g2_decap_8
XFILLER_0_273 VPWR VGND sg13g2_decap_8
XFILLER_1_796 VPWR VGND sg13g2_decap_8
XFILLER_36_417 VPWR VGND sg13g2_decap_8
XFILLER_48_288 VPWR VGND sg13g2_decap_8
XFILLER_45_940 VPWR VGND sg13g2_decap_8
XFILLER_17_642 VPWR VGND sg13g2_decap_8
XFILLER_44_472 VPWR VGND sg13g2_decap_8
X_578_ net83 VGND VPWR _118_ DP_3.matrix\[54\] clknet_5_31__leaf_clk sg13g2_dfrbpq_1
XFILLER_16_185 VPWR VGND sg13g2_fill_1
XFILLER_31_133 VPWR VGND sg13g2_decap_8
XFILLER_32_634 VPWR VGND sg13g2_decap_8
XFILLER_20_829 VPWR VGND sg13g2_decap_8
XFILLER_9_885 VPWR VGND sg13g2_decap_8
.ends

