magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755170679
<< metal1 >>
rect 576 38576 99360 38600
rect 576 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 95072 38576
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95440 38536 99360 38576
rect 576 38512 99360 38536
rect 37315 38240 37373 38241
rect 37315 38200 37324 38240
rect 37364 38200 37373 38240
rect 37315 38199 37373 38200
rect 36643 37988 36701 37989
rect 36643 37948 36652 37988
rect 36692 37948 36701 37988
rect 36643 37947 36701 37948
rect 576 37820 99360 37844
rect 576 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 93832 37820
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 94200 37780 99360 37820
rect 576 37756 99360 37780
rect 37603 37652 37661 37653
rect 37603 37612 37612 37652
rect 37652 37612 37661 37652
rect 37603 37611 37661 37612
rect 9475 37484 9533 37485
rect 9475 37444 9484 37484
rect 9524 37444 9533 37484
rect 9475 37443 9533 37444
rect 20715 37484 20757 37493
rect 20715 37444 20716 37484
rect 20756 37444 20757 37484
rect 20715 37435 20757 37444
rect 10339 37400 10397 37401
rect 10339 37360 10348 37400
rect 10388 37360 10397 37400
rect 10339 37359 10397 37360
rect 18691 37400 18749 37401
rect 18691 37360 18700 37400
rect 18740 37360 18749 37400
rect 18691 37359 18749 37360
rect 19555 37400 19613 37401
rect 19555 37360 19564 37400
rect 19604 37360 19613 37400
rect 19555 37359 19613 37360
rect 20899 37400 20957 37401
rect 20899 37360 20908 37400
rect 20948 37360 20957 37400
rect 20899 37359 20957 37360
rect 25411 37400 25469 37401
rect 25411 37360 25420 37400
rect 25460 37360 25469 37400
rect 25411 37359 25469 37360
rect 35587 37400 35645 37401
rect 35587 37360 35596 37400
rect 35636 37360 35645 37400
rect 35587 37359 35645 37360
rect 36451 37400 36509 37401
rect 36451 37360 36460 37400
rect 36500 37360 36509 37400
rect 36451 37359 36509 37360
rect 18315 37316 18357 37325
rect 18315 37276 18316 37316
rect 18356 37276 18357 37316
rect 18315 37267 18357 37276
rect 35211 37316 35253 37325
rect 35211 37276 35212 37316
rect 35252 37276 35253 37316
rect 35211 37267 35253 37276
rect 9291 37232 9333 37241
rect 9291 37192 9292 37232
rect 9332 37192 9333 37232
rect 9291 37183 9333 37192
rect 9667 37232 9725 37233
rect 9667 37192 9676 37232
rect 9716 37192 9725 37232
rect 9667 37191 9725 37192
rect 21571 37232 21629 37233
rect 21571 37192 21580 37232
rect 21620 37192 21629 37232
rect 21571 37191 21629 37192
rect 24739 37232 24797 37233
rect 24739 37192 24748 37232
rect 24788 37192 24797 37232
rect 24739 37191 24797 37192
rect 576 37064 99360 37088
rect 576 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 95072 37064
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95440 37024 99360 37064
rect 576 37000 99360 37024
rect 11779 36896 11837 36897
rect 11779 36856 11788 36896
rect 11828 36856 11837 36896
rect 11779 36855 11837 36856
rect 9387 36812 9429 36821
rect 9387 36772 9388 36812
rect 9428 36772 9429 36812
rect 9387 36763 9429 36772
rect 7267 36728 7325 36729
rect 7267 36688 7276 36728
rect 7316 36688 7325 36728
rect 7267 36687 7325 36688
rect 9763 36728 9821 36729
rect 9763 36688 9772 36728
rect 9812 36688 9821 36728
rect 9763 36687 9821 36688
rect 10627 36728 10685 36729
rect 10627 36688 10636 36728
rect 10676 36688 10685 36728
rect 10627 36687 10685 36688
rect 18795 36728 18837 36737
rect 18795 36688 18796 36728
rect 18836 36688 18837 36728
rect 18795 36679 18837 36688
rect 19171 36728 19229 36729
rect 19171 36688 19180 36728
rect 19220 36688 19229 36728
rect 19171 36687 19229 36688
rect 20035 36728 20093 36729
rect 20035 36688 20044 36728
rect 20084 36688 20093 36728
rect 20035 36687 20093 36688
rect 21379 36728 21437 36729
rect 21379 36688 21388 36728
rect 21428 36688 21437 36728
rect 21379 36687 21437 36688
rect 24555 36728 24597 36737
rect 24555 36688 24556 36728
rect 24596 36688 24597 36728
rect 24555 36679 24597 36688
rect 24931 36728 24989 36729
rect 24931 36688 24940 36728
rect 24980 36688 24989 36728
rect 24931 36687 24989 36688
rect 25795 36728 25853 36729
rect 25795 36688 25804 36728
rect 25844 36688 25853 36728
rect 25795 36687 25853 36688
rect 32803 36728 32861 36729
rect 32803 36688 32812 36728
rect 32852 36688 32861 36728
rect 32803 36687 32861 36688
rect 36555 36728 36597 36737
rect 36555 36688 36556 36728
rect 36596 36688 36597 36728
rect 36555 36679 36597 36688
rect 36931 36728 36989 36729
rect 36931 36688 36940 36728
rect 36980 36688 36989 36728
rect 36931 36687 36989 36688
rect 37795 36728 37853 36729
rect 37795 36688 37804 36728
rect 37844 36688 37853 36728
rect 37795 36687 37853 36688
rect 5827 36644 5885 36645
rect 5827 36604 5836 36644
rect 5876 36604 5885 36644
rect 5827 36603 5885 36604
rect 21195 36644 21237 36653
rect 21195 36604 21196 36644
rect 21236 36604 21237 36644
rect 21195 36595 21237 36604
rect 31363 36644 31421 36645
rect 31363 36604 31372 36644
rect 31412 36604 31421 36644
rect 31363 36603 31421 36604
rect 5643 36560 5685 36569
rect 5643 36520 5644 36560
rect 5684 36520 5685 36560
rect 5643 36511 5685 36520
rect 6595 36560 6653 36561
rect 6595 36520 6604 36560
rect 6644 36520 6653 36560
rect 6595 36519 6653 36520
rect 31179 36560 31221 36569
rect 31179 36520 31180 36560
rect 31220 36520 31221 36560
rect 31179 36511 31221 36520
rect 32131 36560 32189 36561
rect 32131 36520 32140 36560
rect 32180 36520 32189 36560
rect 32131 36519 32189 36520
rect 38947 36560 39005 36561
rect 38947 36520 38956 36560
rect 38996 36520 39005 36560
rect 38947 36519 39005 36520
rect 22051 36476 22109 36477
rect 22051 36436 22060 36476
rect 22100 36436 22109 36476
rect 22051 36435 22109 36436
rect 26947 36476 27005 36477
rect 26947 36436 26956 36476
rect 26996 36436 27005 36476
rect 26947 36435 27005 36436
rect 576 36308 99360 36332
rect 576 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 93832 36308
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 94200 36268 99360 36308
rect 576 36244 99360 36268
rect 7075 36140 7133 36141
rect 7075 36100 7084 36140
rect 7124 36100 7133 36140
rect 7075 36099 7133 36100
rect 19275 36140 19317 36149
rect 19275 36100 19276 36140
rect 19316 36100 19317 36140
rect 19275 36091 19317 36100
rect 19851 36140 19893 36149
rect 19851 36100 19852 36140
rect 19892 36100 19893 36140
rect 19851 36091 19893 36100
rect 25987 36140 26045 36141
rect 25987 36100 25996 36140
rect 26036 36100 26045 36140
rect 25987 36099 26045 36100
rect 32611 36140 32669 36141
rect 32611 36100 32620 36140
rect 32660 36100 32669 36140
rect 32611 36099 32669 36100
rect 35211 36140 35253 36149
rect 35211 36100 35212 36140
rect 35252 36100 35253 36140
rect 35211 36091 35253 36100
rect 36459 36140 36501 36149
rect 36459 36100 36460 36140
rect 36500 36100 36501 36140
rect 36459 36091 36501 36100
rect 19459 35972 19517 35973
rect 19459 35932 19468 35972
rect 19508 35932 19517 35972
rect 19459 35931 19517 35932
rect 20035 35972 20093 35973
rect 20035 35932 20044 35972
rect 20084 35932 20093 35972
rect 20035 35931 20093 35932
rect 23203 35972 23261 35973
rect 23203 35932 23212 35972
rect 23252 35932 23261 35972
rect 23203 35931 23261 35932
rect 35395 35972 35453 35973
rect 35395 35932 35404 35972
rect 35444 35932 35453 35972
rect 35395 35931 35453 35932
rect 36642 35972 36700 35973
rect 36642 35932 36651 35972
rect 36691 35932 36700 35972
rect 36642 35931 36700 35932
rect 36843 35972 36885 35981
rect 36843 35932 36844 35972
rect 36884 35932 36885 35972
rect 36843 35923 36885 35932
rect 4683 35888 4725 35897
rect 4683 35848 4684 35888
rect 4724 35848 4725 35888
rect 4683 35839 4725 35848
rect 5059 35888 5117 35889
rect 5059 35848 5068 35888
rect 5108 35848 5117 35888
rect 5059 35847 5117 35848
rect 5923 35888 5981 35889
rect 5923 35848 5932 35888
rect 5972 35848 5981 35888
rect 5923 35847 5981 35848
rect 9187 35888 9245 35889
rect 9187 35848 9196 35888
rect 9236 35848 9245 35888
rect 9187 35847 9245 35848
rect 9387 35888 9429 35897
rect 9387 35848 9388 35888
rect 9428 35848 9429 35888
rect 9387 35839 9429 35848
rect 9955 35888 10013 35889
rect 9955 35848 9964 35888
rect 10004 35848 10013 35888
rect 9955 35847 10013 35848
rect 10819 35888 10877 35889
rect 10819 35848 10828 35888
rect 10868 35848 10877 35888
rect 10819 35847 10877 35848
rect 22155 35888 22197 35897
rect 22155 35848 22156 35888
rect 22196 35848 22197 35888
rect 22155 35839 22197 35848
rect 22339 35888 22397 35889
rect 22339 35848 22348 35888
rect 22388 35848 22397 35888
rect 22339 35847 22397 35848
rect 23971 35888 24029 35889
rect 23971 35848 23980 35888
rect 24020 35848 24029 35888
rect 23971 35847 24029 35848
rect 24835 35888 24893 35889
rect 24835 35848 24844 35888
rect 24884 35848 24893 35888
rect 24835 35847 24893 35848
rect 26851 35888 26909 35889
rect 26851 35848 26860 35888
rect 26900 35848 26909 35888
rect 26851 35847 26909 35848
rect 30219 35888 30261 35897
rect 30219 35848 30220 35888
rect 30260 35848 30261 35888
rect 30219 35839 30261 35848
rect 30595 35888 30653 35889
rect 30595 35848 30604 35888
rect 30644 35848 30653 35888
rect 30595 35847 30653 35848
rect 31459 35888 31517 35889
rect 31459 35848 31468 35888
rect 31508 35848 31517 35888
rect 31459 35847 31517 35848
rect 36067 35888 36125 35889
rect 36067 35848 36076 35888
rect 36116 35848 36125 35888
rect 36067 35847 36125 35848
rect 36267 35888 36309 35897
rect 36267 35848 36268 35888
rect 36308 35848 36309 35888
rect 36267 35839 36309 35848
rect 37507 35888 37565 35889
rect 37507 35848 37516 35888
rect 37556 35848 37565 35888
rect 37507 35847 37565 35848
rect 9291 35804 9333 35813
rect 9291 35764 9292 35804
rect 9332 35764 9333 35804
rect 9291 35755 9333 35764
rect 9579 35804 9621 35813
rect 9579 35764 9580 35804
rect 9620 35764 9621 35804
rect 9579 35755 9621 35764
rect 22251 35804 22293 35813
rect 22251 35764 22252 35804
rect 22292 35764 22293 35804
rect 22251 35755 22293 35764
rect 23595 35804 23637 35813
rect 23595 35764 23596 35804
rect 23636 35764 23637 35804
rect 23595 35755 23637 35764
rect 36171 35804 36213 35813
rect 36171 35764 36172 35804
rect 36212 35764 36213 35804
rect 36171 35755 36213 35764
rect 11971 35720 12029 35721
rect 11971 35680 11980 35720
rect 12020 35680 12029 35720
rect 11971 35679 12029 35680
rect 23403 35720 23445 35729
rect 23403 35680 23404 35720
rect 23444 35680 23445 35720
rect 23403 35671 23445 35680
rect 26179 35720 26237 35721
rect 26179 35680 26188 35720
rect 26228 35680 26237 35720
rect 26179 35679 26237 35680
rect 576 35552 99360 35576
rect 576 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 95072 35552
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95440 35512 99360 35552
rect 576 35488 99360 35512
rect 9483 35384 9525 35393
rect 9483 35344 9484 35384
rect 9524 35344 9525 35384
rect 9483 35335 9525 35344
rect 25219 35384 25277 35385
rect 25219 35344 25228 35384
rect 25268 35344 25277 35384
rect 25219 35343 25277 35344
rect 7371 35300 7413 35309
rect 7371 35260 7372 35300
rect 7412 35260 7413 35300
rect 7371 35251 7413 35260
rect 22147 35300 22205 35301
rect 22147 35260 22156 35300
rect 22196 35260 22205 35300
rect 22147 35259 22205 35260
rect 36259 35300 36317 35301
rect 36259 35260 36268 35300
rect 36308 35260 36317 35300
rect 36259 35259 36317 35260
rect 5835 35216 5877 35225
rect 5835 35176 5836 35216
rect 5876 35176 5877 35216
rect 5835 35167 5877 35176
rect 6499 35216 6557 35217
rect 6499 35176 6508 35216
rect 6548 35176 6557 35216
rect 6499 35175 6557 35176
rect 7275 35216 7317 35225
rect 7275 35176 7276 35216
rect 7316 35176 7317 35216
rect 7275 35167 7317 35176
rect 7459 35216 7517 35217
rect 7459 35176 7468 35216
rect 7508 35176 7517 35216
rect 7459 35175 7517 35176
rect 10339 35216 10397 35217
rect 10339 35176 10348 35216
rect 10388 35176 10397 35216
rect 10339 35175 10397 35176
rect 21291 35216 21333 35225
rect 21291 35176 21292 35216
rect 21332 35176 21333 35216
rect 21291 35167 21333 35176
rect 21475 35216 21533 35217
rect 21475 35176 21484 35216
rect 21524 35176 21533 35216
rect 21475 35175 21533 35176
rect 21667 35216 21725 35217
rect 21667 35176 21676 35216
rect 21716 35176 21725 35216
rect 21667 35175 21725 35176
rect 22051 35216 22109 35217
rect 22051 35176 22060 35216
rect 22100 35176 22109 35216
rect 22051 35175 22109 35176
rect 25315 35216 25373 35217
rect 25315 35176 25324 35216
rect 25364 35176 25373 35216
rect 25315 35175 25373 35176
rect 32899 35216 32957 35217
rect 32899 35176 32908 35216
rect 32948 35176 32957 35216
rect 32899 35175 32957 35176
rect 33099 35216 33141 35225
rect 33099 35176 33100 35216
rect 33140 35176 33141 35216
rect 33099 35167 33141 35176
rect 33195 35216 33237 35225
rect 33195 35176 33196 35216
rect 33236 35176 33237 35216
rect 33195 35167 33237 35176
rect 33283 35216 33341 35217
rect 33283 35176 33292 35216
rect 33332 35176 33341 35216
rect 33283 35175 33341 35176
rect 35779 35216 35837 35217
rect 35779 35176 35788 35216
rect 35828 35176 35837 35216
rect 35779 35175 35837 35176
rect 36163 35216 36221 35217
rect 36163 35176 36172 35216
rect 36212 35176 36221 35216
rect 36163 35175 36221 35176
rect 5059 35132 5117 35133
rect 5059 35092 5068 35132
rect 5108 35092 5117 35132
rect 5059 35091 5117 35092
rect 9283 35132 9341 35133
rect 9283 35092 9292 35132
rect 9332 35092 9341 35132
rect 9283 35091 9341 35092
rect 9675 35132 9717 35141
rect 9675 35092 9676 35132
rect 9716 35092 9717 35132
rect 9675 35083 9717 35092
rect 24835 35132 24893 35133
rect 24835 35092 24844 35132
rect 24884 35092 24893 35132
rect 24835 35091 24893 35092
rect 31459 35132 31517 35133
rect 31459 35092 31468 35132
rect 31508 35092 31517 35132
rect 31459 35091 31517 35092
rect 32235 35132 32277 35141
rect 32235 35092 32236 35132
rect 32276 35092 32277 35132
rect 32235 35083 32277 35092
rect 21387 35048 21429 35057
rect 21387 35008 21388 35048
rect 21428 35008 21429 35048
rect 21387 34999 21429 35008
rect 24651 35048 24693 35057
rect 24651 35008 24652 35048
rect 24692 35008 24693 35048
rect 24651 34999 24693 35008
rect 4875 34964 4917 34973
rect 4875 34924 4876 34964
rect 4916 34924 4917 34964
rect 4875 34915 4917 34924
rect 25507 34964 25565 34965
rect 25507 34924 25516 34964
rect 25556 34924 25565 34964
rect 25507 34923 25565 34924
rect 31275 34964 31317 34973
rect 31275 34924 31276 34964
rect 31316 34924 31317 34964
rect 31275 34915 31317 34924
rect 576 34796 99360 34820
rect 576 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 93832 34796
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 94200 34756 99360 34796
rect 576 34732 99360 34756
rect 6307 34628 6365 34629
rect 6307 34588 6316 34628
rect 6356 34588 6365 34628
rect 6307 34587 6365 34588
rect 20331 34628 20373 34637
rect 20331 34588 20332 34628
rect 20372 34588 20373 34628
rect 20331 34579 20373 34588
rect 32707 34628 32765 34629
rect 32707 34588 32716 34628
rect 32756 34588 32765 34628
rect 32707 34587 32765 34588
rect 16875 34460 16917 34469
rect 16875 34420 16876 34460
rect 16916 34420 16917 34460
rect 16875 34411 16917 34420
rect 3915 34376 3957 34385
rect 3915 34336 3916 34376
rect 3956 34336 3957 34376
rect 3915 34327 3957 34336
rect 4291 34376 4349 34377
rect 4291 34336 4300 34376
rect 4340 34336 4349 34376
rect 4291 34335 4349 34336
rect 5155 34376 5213 34377
rect 5155 34336 5164 34376
rect 5204 34336 5213 34376
rect 5155 34335 5213 34336
rect 8035 34376 8093 34377
rect 8035 34336 8044 34376
rect 8084 34336 8093 34376
rect 8035 34335 8093 34336
rect 8419 34376 8477 34377
rect 8419 34336 8428 34376
rect 8468 34336 8477 34376
rect 8419 34335 8477 34336
rect 8707 34376 8765 34377
rect 8707 34336 8716 34376
rect 8756 34336 8765 34376
rect 8707 34335 8765 34336
rect 14851 34376 14909 34377
rect 14851 34336 14860 34376
rect 14900 34336 14909 34376
rect 14851 34335 14909 34336
rect 15715 34376 15773 34377
rect 15715 34336 15724 34376
rect 15764 34336 15773 34376
rect 15715 34335 15773 34336
rect 17731 34376 17789 34377
rect 17731 34336 17740 34376
rect 17780 34336 17789 34376
rect 17731 34335 17789 34336
rect 20803 34376 20861 34377
rect 20803 34336 20812 34376
rect 20852 34336 20861 34376
rect 20803 34335 20861 34336
rect 30315 34376 30357 34385
rect 30315 34336 30316 34376
rect 30356 34336 30357 34376
rect 30315 34327 30357 34336
rect 30691 34376 30749 34377
rect 30691 34336 30700 34376
rect 30740 34336 30749 34376
rect 30691 34335 30749 34336
rect 31555 34376 31613 34377
rect 31555 34336 31564 34376
rect 31604 34336 31613 34376
rect 31555 34335 31613 34336
rect 33859 34376 33917 34377
rect 33859 34336 33868 34376
rect 33908 34336 33917 34376
rect 33859 34335 33917 34336
rect 37323 34376 37365 34385
rect 37323 34336 37324 34376
rect 37364 34336 37365 34376
rect 37323 34327 37365 34336
rect 37699 34376 37757 34377
rect 37699 34336 37708 34376
rect 37748 34336 37757 34376
rect 37699 34335 37757 34336
rect 38563 34376 38621 34377
rect 38563 34336 38572 34376
rect 38612 34336 38621 34376
rect 38563 34335 38621 34336
rect 14475 34292 14517 34301
rect 14475 34252 14476 34292
rect 14516 34252 14517 34292
rect 14475 34243 14517 34252
rect 7939 34208 7997 34209
rect 7939 34168 7948 34208
rect 7988 34168 7997 34208
rect 7939 34167 7997 34168
rect 8227 34208 8285 34209
rect 8227 34168 8236 34208
rect 8276 34168 8285 34208
rect 8227 34167 8285 34168
rect 8907 34208 8949 34217
rect 8907 34168 8908 34208
rect 8948 34168 8949 34208
rect 8907 34159 8949 34168
rect 17059 34208 17117 34209
rect 17059 34168 17068 34208
rect 17108 34168 17117 34208
rect 17059 34167 17117 34168
rect 20331 34208 20373 34217
rect 20331 34168 20332 34208
rect 20372 34168 20373 34208
rect 20331 34159 20373 34168
rect 33763 34208 33821 34209
rect 33763 34168 33772 34208
rect 33812 34168 33821 34208
rect 33763 34167 33821 34168
rect 34051 34208 34109 34209
rect 34051 34168 34060 34208
rect 34100 34168 34109 34208
rect 34051 34167 34109 34168
rect 39715 34208 39773 34209
rect 39715 34168 39724 34208
rect 39764 34168 39773 34208
rect 39715 34167 39773 34168
rect 576 34040 99360 34064
rect 576 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 95072 34040
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95440 34000 99360 34040
rect 576 33976 99360 34000
rect 10723 33704 10781 33705
rect 10723 33664 10732 33704
rect 10772 33664 10781 33704
rect 10723 33663 10781 33664
rect 11107 33704 11165 33705
rect 11107 33664 11116 33704
rect 11156 33664 11165 33704
rect 11107 33663 11165 33664
rect 12067 33704 12125 33705
rect 12067 33664 12076 33704
rect 12116 33664 12125 33704
rect 12067 33663 12125 33664
rect 14955 33704 14997 33713
rect 14955 33664 14956 33704
rect 14996 33664 14997 33704
rect 14955 33655 14997 33664
rect 15331 33704 15389 33705
rect 15331 33664 15340 33704
rect 15380 33664 15389 33704
rect 15331 33663 15389 33664
rect 16195 33704 16253 33705
rect 16195 33664 16204 33704
rect 16244 33664 16253 33704
rect 16195 33663 16253 33664
rect 17539 33704 17597 33705
rect 17539 33664 17548 33704
rect 17588 33664 17597 33704
rect 17539 33663 17597 33664
rect 24259 33704 24317 33705
rect 24259 33664 24268 33704
rect 24308 33664 24317 33704
rect 24259 33663 24317 33664
rect 24547 33704 24605 33705
rect 24547 33664 24556 33704
rect 24596 33664 24605 33704
rect 24547 33663 24605 33664
rect 47491 33704 47549 33705
rect 47491 33664 47500 33704
rect 47540 33664 47549 33704
rect 47491 33663 47549 33664
rect 17355 33620 17397 33629
rect 17355 33580 17356 33620
rect 17396 33580 17397 33620
rect 17355 33571 17397 33580
rect 11403 33536 11445 33545
rect 11403 33496 11404 33536
rect 11444 33496 11445 33536
rect 11403 33487 11445 33496
rect 18211 33452 18269 33453
rect 18211 33412 18220 33452
rect 18260 33412 18269 33452
rect 18211 33411 18269 33412
rect 25035 33452 25077 33461
rect 25035 33412 25036 33452
rect 25076 33412 25077 33452
rect 25035 33403 25077 33412
rect 46819 33452 46877 33453
rect 46819 33412 46828 33452
rect 46868 33412 46877 33452
rect 46819 33411 46877 33412
rect 576 33284 99360 33308
rect 576 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 18232 33284
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18600 33244 33352 33284
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33720 33244 48472 33284
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48840 33244 63592 33284
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63960 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 93832 33284
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 94200 33244 99360 33284
rect 576 33220 99360 33244
rect 15435 33116 15477 33125
rect 15435 33076 15436 33116
rect 15476 33076 15477 33116
rect 15435 33067 15477 33076
rect 15915 33116 15957 33125
rect 15915 33076 15916 33116
rect 15956 33076 15957 33116
rect 15915 33067 15957 33076
rect 47779 33116 47837 33117
rect 47779 33076 47788 33116
rect 47828 33076 47837 33116
rect 47779 33075 47837 33076
rect 43371 33032 43413 33041
rect 43371 32992 43372 33032
rect 43412 32992 43413 33032
rect 43371 32983 43413 32992
rect 15619 32948 15677 32949
rect 15619 32908 15628 32948
rect 15668 32908 15677 32948
rect 15619 32907 15677 32908
rect 16099 32948 16157 32949
rect 16099 32908 16108 32948
rect 16148 32908 16157 32948
rect 16099 32907 16157 32908
rect 43555 32948 43613 32949
rect 43555 32908 43564 32948
rect 43604 32908 43613 32948
rect 43555 32907 43613 32908
rect 44331 32948 44373 32957
rect 44331 32908 44332 32948
rect 44372 32908 44373 32948
rect 44331 32899 44373 32908
rect 6499 32864 6557 32865
rect 6499 32824 6508 32864
rect 6548 32824 6557 32864
rect 6499 32823 6557 32824
rect 7459 32864 7517 32865
rect 7459 32824 7468 32864
rect 7508 32824 7517 32864
rect 7459 32823 7517 32824
rect 8811 32864 8853 32873
rect 8811 32824 8812 32864
rect 8852 32824 8853 32864
rect 8811 32815 8853 32824
rect 9187 32864 9245 32865
rect 9187 32824 9196 32864
rect 9236 32824 9245 32864
rect 9187 32823 9245 32824
rect 10051 32864 10109 32865
rect 10051 32824 10060 32864
rect 10100 32824 10109 32864
rect 10051 32823 10109 32824
rect 21771 32864 21813 32873
rect 21771 32824 21772 32864
rect 21812 32824 21813 32864
rect 21771 32815 21813 32824
rect 22147 32864 22205 32865
rect 22147 32824 22156 32864
rect 22196 32824 22205 32864
rect 22147 32823 22205 32824
rect 23011 32864 23069 32865
rect 23011 32824 23020 32864
rect 23060 32824 23069 32864
rect 23011 32823 23069 32824
rect 25611 32864 25653 32873
rect 25611 32824 25612 32864
rect 25652 32824 25653 32864
rect 25611 32815 25653 32824
rect 25987 32864 26045 32865
rect 25987 32824 25996 32864
rect 26036 32824 26045 32864
rect 25987 32823 26045 32824
rect 26851 32864 26909 32865
rect 26851 32824 26860 32864
rect 26900 32824 26909 32864
rect 26851 32823 26909 32824
rect 36931 32864 36989 32865
rect 36931 32824 36940 32864
rect 36980 32824 36989 32864
rect 36931 32823 36989 32824
rect 44995 32864 45053 32865
rect 44995 32824 45004 32864
rect 45044 32824 45053 32864
rect 44995 32823 45053 32824
rect 45763 32864 45821 32865
rect 45763 32824 45772 32864
rect 45812 32824 45821 32864
rect 45763 32823 45821 32824
rect 46627 32864 46685 32865
rect 46627 32824 46636 32864
rect 46676 32824 46685 32864
rect 46627 32823 46685 32824
rect 45387 32780 45429 32789
rect 45387 32740 45388 32780
rect 45428 32740 45429 32780
rect 45387 32731 45429 32740
rect 6987 32696 7029 32705
rect 6987 32656 6988 32696
rect 7028 32656 7029 32696
rect 6987 32647 7029 32656
rect 11203 32696 11261 32697
rect 11203 32656 11212 32696
rect 11252 32656 11261 32696
rect 11203 32655 11261 32656
rect 24163 32696 24221 32697
rect 24163 32656 24172 32696
rect 24212 32656 24221 32696
rect 24163 32655 24221 32656
rect 28003 32696 28061 32697
rect 28003 32656 28012 32696
rect 28052 32656 28061 32696
rect 28003 32655 28061 32656
rect 37603 32696 37661 32697
rect 37603 32656 37612 32696
rect 37652 32656 37661 32696
rect 37603 32655 37661 32656
rect 576 32528 99360 32552
rect 576 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 19472 32528
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19840 32488 34592 32528
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34960 32488 49712 32528
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 50080 32488 64832 32528
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 65200 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 95072 32528
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95440 32488 99360 32528
rect 576 32464 99360 32488
rect 44899 32360 44957 32361
rect 44899 32320 44908 32360
rect 44948 32320 44957 32360
rect 44899 32319 44957 32320
rect 45483 32360 45525 32369
rect 45483 32320 45484 32360
rect 45524 32320 45525 32360
rect 45483 32311 45525 32320
rect 8811 32276 8853 32285
rect 8811 32236 8812 32276
rect 8852 32236 8853 32276
rect 8811 32227 8853 32236
rect 33867 32276 33909 32285
rect 33867 32236 33868 32276
rect 33908 32236 33909 32276
rect 33867 32227 33909 32236
rect 38083 32276 38141 32277
rect 38083 32236 38092 32276
rect 38132 32236 38141 32276
rect 38083 32235 38141 32236
rect 39907 32276 39965 32277
rect 39907 32236 39916 32276
rect 39956 32236 39965 32276
rect 39907 32235 39965 32236
rect 42507 32276 42549 32285
rect 42507 32236 42508 32276
rect 42548 32236 42549 32276
rect 42507 32227 42549 32236
rect 9187 32192 9245 32193
rect 9187 32152 9196 32192
rect 9236 32152 9245 32192
rect 9187 32151 9245 32152
rect 10051 32192 10109 32193
rect 10051 32152 10060 32192
rect 10100 32152 10109 32192
rect 10051 32151 10109 32152
rect 16971 32192 17013 32201
rect 16971 32152 16972 32192
rect 17012 32152 17013 32192
rect 16971 32143 17013 32152
rect 17155 32192 17213 32193
rect 17155 32152 17164 32192
rect 17204 32152 17213 32192
rect 17155 32151 17213 32152
rect 34243 32192 34301 32193
rect 34243 32152 34252 32192
rect 34292 32152 34301 32192
rect 34243 32151 34301 32152
rect 35107 32192 35165 32193
rect 35107 32152 35116 32192
rect 35156 32152 35165 32192
rect 35107 32151 35165 32152
rect 37227 32192 37269 32201
rect 37227 32152 37228 32192
rect 37268 32152 37269 32192
rect 37227 32143 37269 32152
rect 37411 32192 37469 32193
rect 37411 32152 37420 32192
rect 37460 32152 37469 32192
rect 37411 32151 37469 32152
rect 37603 32192 37661 32193
rect 37603 32152 37612 32192
rect 37652 32152 37661 32192
rect 37603 32151 37661 32152
rect 37987 32192 38045 32193
rect 37987 32152 37996 32192
rect 38036 32152 38045 32192
rect 37987 32151 38045 32152
rect 40003 32192 40061 32193
rect 40003 32152 40012 32192
rect 40052 32152 40061 32192
rect 40003 32151 40061 32152
rect 40387 32192 40445 32193
rect 40387 32152 40396 32192
rect 40436 32152 40445 32192
rect 40387 32151 40445 32152
rect 42883 32192 42941 32193
rect 42883 32152 42892 32192
rect 42932 32152 42941 32192
rect 42883 32151 42941 32152
rect 43747 32192 43805 32193
rect 43747 32152 43756 32192
rect 43796 32152 43805 32192
rect 43747 32151 43805 32152
rect 36267 32108 36309 32117
rect 36267 32068 36268 32108
rect 36308 32068 36309 32108
rect 36267 32059 36309 32068
rect 45667 32108 45725 32109
rect 45667 32068 45676 32108
rect 45716 32068 45725 32108
rect 45667 32067 45725 32068
rect 11203 31940 11261 31941
rect 11203 31900 11212 31940
rect 11252 31900 11261 31940
rect 11203 31899 11261 31900
rect 17067 31940 17109 31949
rect 17067 31900 17068 31940
rect 17108 31900 17109 31940
rect 17067 31891 17109 31900
rect 37323 31940 37365 31949
rect 37323 31900 37324 31940
rect 37364 31900 37365 31940
rect 37323 31891 37365 31900
rect 576 31772 99360 31796
rect 576 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 18232 31772
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18600 31732 33352 31772
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33720 31732 48472 31772
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48840 31732 63592 31772
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63960 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 93832 31772
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 94200 31732 99360 31772
rect 576 31708 99360 31732
rect 38275 31604 38333 31605
rect 38275 31564 38284 31604
rect 38324 31564 38333 31604
rect 38275 31563 38333 31564
rect 22347 31520 22389 31529
rect 22347 31480 22348 31520
rect 22388 31480 22389 31520
rect 22347 31471 22389 31480
rect 33771 31520 33813 31529
rect 33771 31480 33772 31520
rect 33812 31480 33813 31520
rect 33771 31471 33813 31480
rect 37131 31520 37173 31529
rect 37131 31480 37132 31520
rect 37172 31480 37173 31520
rect 37131 31471 37173 31480
rect 38467 31436 38525 31437
rect 38467 31396 38476 31436
rect 38516 31396 38525 31436
rect 38467 31395 38525 31396
rect 3907 31352 3965 31353
rect 3907 31312 3916 31352
rect 3956 31312 3965 31352
rect 3907 31311 3965 31312
rect 4867 31352 4925 31353
rect 4867 31312 4876 31352
rect 4916 31312 4925 31352
rect 4867 31311 4925 31312
rect 11779 31352 11837 31353
rect 11779 31312 11788 31352
rect 11828 31312 11837 31352
rect 11779 31311 11837 31312
rect 22627 31352 22685 31353
rect 22627 31312 22636 31352
rect 22676 31312 22685 31352
rect 22627 31311 22685 31312
rect 23875 31352 23933 31353
rect 23875 31312 23884 31352
rect 23924 31312 23933 31352
rect 23875 31311 23933 31312
rect 24163 31352 24221 31353
rect 24163 31312 24172 31352
rect 24212 31312 24221 31352
rect 24163 31311 24221 31312
rect 27619 31352 27677 31353
rect 27619 31312 27628 31352
rect 27668 31312 27677 31352
rect 27619 31311 27677 31312
rect 31171 31352 31229 31353
rect 31171 31312 31180 31352
rect 31220 31312 31229 31352
rect 31171 31311 31229 31312
rect 33091 31352 33149 31353
rect 33091 31312 33100 31352
rect 33140 31312 33149 31352
rect 33091 31311 33149 31312
rect 34051 31352 34109 31353
rect 34051 31312 34060 31352
rect 34100 31312 34109 31352
rect 34051 31311 34109 31312
rect 36163 31352 36221 31353
rect 36163 31312 36172 31352
rect 36212 31312 36221 31352
rect 36163 31311 36221 31312
rect 36451 31352 36509 31353
rect 36451 31312 36460 31352
rect 36500 31312 36509 31352
rect 36451 31311 36509 31312
rect 37411 31352 37469 31353
rect 37411 31312 37420 31352
rect 37460 31312 37469 31352
rect 37411 31311 37469 31312
rect 37603 31352 37661 31353
rect 37603 31312 37612 31352
rect 37652 31312 37661 31352
rect 37603 31311 37661 31312
rect 38755 31352 38813 31353
rect 38755 31312 38764 31352
rect 38804 31312 38813 31352
rect 38755 31311 38813 31312
rect 38859 31352 38901 31361
rect 38859 31312 38860 31352
rect 38900 31312 38901 31352
rect 38859 31303 38901 31312
rect 44515 31352 44573 31353
rect 44515 31312 44524 31352
rect 44564 31312 44573 31352
rect 44515 31311 44573 31312
rect 11107 31184 11165 31185
rect 11107 31144 11116 31184
rect 11156 31144 11165 31184
rect 11107 31143 11165 31144
rect 24363 31184 24405 31193
rect 24363 31144 24364 31184
rect 24404 31144 24405 31184
rect 24363 31135 24405 31144
rect 26947 31184 27005 31185
rect 26947 31144 26956 31184
rect 26996 31144 27005 31184
rect 26947 31143 27005 31144
rect 30499 31184 30557 31185
rect 30499 31144 30508 31184
rect 30548 31144 30557 31184
rect 30499 31143 30557 31144
rect 35491 31184 35549 31185
rect 35491 31144 35500 31184
rect 35540 31144 35549 31184
rect 35491 31143 35549 31144
rect 44323 31184 44381 31185
rect 44323 31144 44332 31184
rect 44372 31144 44381 31184
rect 44323 31143 44381 31144
rect 44611 31184 44669 31185
rect 44611 31144 44620 31184
rect 44660 31144 44669 31184
rect 44611 31143 44669 31144
rect 576 31016 99360 31040
rect 576 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 19472 31016
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19840 30976 34592 31016
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34960 30976 49712 31016
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 50080 30976 64832 31016
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 65200 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 95072 31016
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95440 30976 99360 31016
rect 576 30952 99360 30976
rect 18211 30848 18269 30849
rect 18211 30808 18220 30848
rect 18260 30808 18269 30848
rect 18211 30807 18269 30808
rect 22531 30848 22589 30849
rect 22531 30808 22540 30848
rect 22580 30808 22589 30848
rect 22531 30807 22589 30808
rect 30403 30848 30461 30849
rect 30403 30808 30412 30848
rect 30452 30808 30461 30848
rect 30403 30807 30461 30808
rect 34635 30848 34677 30857
rect 34635 30808 34636 30848
rect 34676 30808 34677 30848
rect 34635 30799 34677 30808
rect 35971 30848 36029 30849
rect 35971 30808 35980 30848
rect 36020 30808 36029 30848
rect 35971 30807 36029 30808
rect 39427 30848 39485 30849
rect 39427 30808 39436 30848
rect 39476 30808 39485 30848
rect 39427 30807 39485 30808
rect 17923 30764 17981 30765
rect 17923 30724 17932 30764
rect 17972 30724 17981 30764
rect 17923 30723 17981 30724
rect 20139 30764 20181 30773
rect 20139 30724 20140 30764
rect 20180 30724 20181 30764
rect 20139 30715 20181 30724
rect 32811 30764 32853 30773
rect 32811 30724 32812 30764
rect 32852 30724 32853 30764
rect 32811 30715 32853 30724
rect 41835 30764 41877 30773
rect 41835 30724 41836 30764
rect 41876 30724 41877 30764
rect 41835 30715 41877 30724
rect 45475 30764 45533 30765
rect 45475 30724 45484 30764
rect 45524 30724 45533 30764
rect 45475 30723 45533 30724
rect 2859 30680 2901 30689
rect 2859 30640 2860 30680
rect 2900 30640 2901 30680
rect 2859 30631 2901 30640
rect 3235 30680 3293 30681
rect 3235 30640 3244 30680
rect 3284 30640 3293 30680
rect 3235 30639 3293 30640
rect 4099 30680 4157 30681
rect 4099 30640 4108 30680
rect 4148 30640 4157 30680
rect 4099 30639 4157 30640
rect 6115 30680 6173 30681
rect 6115 30640 6124 30680
rect 6164 30640 6173 30680
rect 6115 30639 6173 30640
rect 16203 30680 16245 30689
rect 16203 30640 16204 30680
rect 16244 30640 16245 30680
rect 16203 30631 16245 30640
rect 16867 30680 16925 30681
rect 16867 30640 16876 30680
rect 16916 30640 16925 30680
rect 16867 30639 16925 30640
rect 17067 30680 17109 30689
rect 17067 30640 17068 30680
rect 17108 30640 17109 30680
rect 17067 30631 17109 30640
rect 17251 30680 17309 30681
rect 17251 30640 17260 30680
rect 17300 30640 17309 30680
rect 17251 30639 17309 30640
rect 17443 30680 17501 30681
rect 17443 30640 17452 30680
rect 17492 30640 17501 30680
rect 17443 30639 17501 30640
rect 17731 30680 17789 30681
rect 17731 30640 17740 30680
rect 17780 30640 17789 30680
rect 17731 30639 17789 30640
rect 18307 30680 18365 30681
rect 18307 30640 18316 30680
rect 18356 30640 18365 30680
rect 18307 30639 18365 30640
rect 20515 30680 20573 30681
rect 20515 30640 20524 30680
rect 20564 30640 20573 30680
rect 20515 30639 20573 30640
rect 21379 30680 21437 30681
rect 21379 30640 21388 30680
rect 21428 30640 21437 30680
rect 21379 30639 21437 30640
rect 24259 30680 24317 30681
rect 24259 30640 24268 30680
rect 24308 30640 24317 30680
rect 24259 30639 24317 30640
rect 24939 30680 24981 30689
rect 24939 30640 24940 30680
rect 24980 30640 24981 30680
rect 24939 30631 24981 30640
rect 25123 30680 25181 30681
rect 25123 30640 25132 30680
rect 25172 30640 25181 30680
rect 25123 30639 25181 30640
rect 25227 30680 25269 30689
rect 25227 30640 25228 30680
rect 25268 30640 25269 30680
rect 25227 30631 25269 30640
rect 25323 30680 25365 30689
rect 25323 30640 25324 30680
rect 25364 30640 25365 30680
rect 25323 30631 25365 30640
rect 25707 30680 25749 30689
rect 25707 30640 25708 30680
rect 25748 30640 25749 30680
rect 25707 30631 25749 30640
rect 25795 30680 25853 30681
rect 25795 30640 25804 30680
rect 25844 30640 25853 30680
rect 25795 30639 25853 30640
rect 26755 30680 26813 30681
rect 26755 30640 26764 30680
rect 26804 30640 26813 30680
rect 26755 30639 26813 30640
rect 31555 30680 31613 30681
rect 31555 30640 31564 30680
rect 31604 30640 31613 30680
rect 31555 30639 31613 30640
rect 32419 30680 32477 30681
rect 32419 30640 32428 30680
rect 32468 30640 32477 30680
rect 32419 30639 32477 30640
rect 34147 30680 34205 30681
rect 34147 30640 34156 30680
rect 34196 30640 34205 30680
rect 34147 30639 34205 30640
rect 35107 30680 35165 30681
rect 35107 30640 35116 30680
rect 35156 30640 35165 30680
rect 35107 30639 35165 30640
rect 35779 30680 35837 30681
rect 35779 30640 35788 30680
rect 35828 30640 35837 30680
rect 35779 30639 35837 30640
rect 37123 30680 37181 30681
rect 37123 30640 37132 30680
rect 37172 30640 37181 30680
rect 37123 30639 37181 30640
rect 37987 30680 38045 30681
rect 37987 30640 37996 30680
rect 38036 30640 38045 30680
rect 37987 30639 38045 30640
rect 38379 30680 38421 30689
rect 38379 30640 38380 30680
rect 38420 30640 38421 30680
rect 38379 30631 38421 30640
rect 40579 30680 40637 30681
rect 40579 30640 40588 30680
rect 40628 30640 40637 30680
rect 40579 30639 40637 30640
rect 41443 30680 41501 30681
rect 41443 30640 41452 30680
rect 41492 30640 41501 30680
rect 41443 30639 41501 30640
rect 44995 30680 45053 30681
rect 44995 30640 45004 30680
rect 45044 30640 45053 30680
rect 44995 30639 45053 30640
rect 45379 30680 45437 30681
rect 45379 30640 45388 30680
rect 45428 30640 45437 30680
rect 45379 30639 45437 30640
rect 46435 30680 46493 30681
rect 46435 30640 46444 30680
rect 46484 30640 46493 30680
rect 46435 30639 46493 30640
rect 46539 30680 46581 30689
rect 46539 30640 46540 30680
rect 46580 30640 46581 30680
rect 46539 30631 46581 30640
rect 46635 30680 46677 30689
rect 46635 30640 46636 30680
rect 46676 30640 46677 30680
rect 46635 30631 46677 30640
rect 49219 30680 49277 30681
rect 49219 30640 49228 30680
rect 49268 30640 49277 30680
rect 49219 30639 49277 30640
rect 5259 30596 5301 30605
rect 5259 30556 5260 30596
rect 5300 30556 5301 30596
rect 5259 30547 5301 30556
rect 15427 30596 15485 30597
rect 15427 30556 15436 30596
rect 15476 30556 15485 30596
rect 15427 30555 15485 30556
rect 26083 30596 26141 30597
rect 26083 30556 26092 30596
rect 26132 30556 26141 30596
rect 26083 30555 26141 30556
rect 47491 30596 47549 30597
rect 47491 30556 47500 30596
rect 47540 30556 47549 30596
rect 47491 30555 47549 30556
rect 48555 30596 48597 30605
rect 48555 30556 48556 30596
rect 48596 30556 48597 30596
rect 48555 30547 48597 30556
rect 17163 30512 17205 30521
rect 17163 30472 17164 30512
rect 17204 30472 17205 30512
rect 17163 30463 17205 30472
rect 5443 30428 5501 30429
rect 5443 30388 5452 30428
rect 5492 30388 5501 30428
rect 5443 30387 5501 30388
rect 15243 30428 15285 30437
rect 15243 30388 15244 30428
rect 15284 30388 15285 30428
rect 15243 30379 15285 30388
rect 18499 30428 18557 30429
rect 18499 30388 18508 30428
rect 18548 30388 18557 30428
rect 18499 30387 18557 30388
rect 27427 30428 27485 30429
rect 27427 30388 27436 30428
rect 27476 30388 27485 30428
rect 27427 30387 27485 30388
rect 47307 30428 47349 30437
rect 47307 30388 47308 30428
rect 47348 30388 47349 30428
rect 47307 30379 47349 30388
rect 576 30260 99360 30284
rect 576 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 18232 30260
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18600 30220 33352 30260
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33720 30220 48472 30260
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48840 30220 63592 30260
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63960 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 93832 30260
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 94200 30220 99360 30260
rect 576 30196 99360 30220
rect 3915 30092 3957 30101
rect 3915 30052 3916 30092
rect 3956 30052 3957 30092
rect 3915 30043 3957 30052
rect 9675 30092 9717 30101
rect 9675 30052 9676 30092
rect 9716 30052 9717 30092
rect 9675 30043 9717 30052
rect 16771 30092 16829 30093
rect 16771 30052 16780 30092
rect 16820 30052 16829 30092
rect 16771 30051 16829 30052
rect 17251 30092 17309 30093
rect 17251 30052 17260 30092
rect 17300 30052 17309 30092
rect 17251 30051 17309 30052
rect 23203 30092 23261 30093
rect 23203 30052 23212 30092
rect 23252 30052 23261 30092
rect 23203 30051 23261 30052
rect 44907 30092 44949 30101
rect 44907 30052 44908 30092
rect 44948 30052 44949 30092
rect 44907 30043 44949 30052
rect 49315 30092 49373 30093
rect 49315 30052 49324 30092
rect 49364 30052 49373 30092
rect 49315 30051 49373 30052
rect 45579 30008 45621 30017
rect 45579 29968 45580 30008
rect 45620 29968 45621 30008
rect 45579 29959 45621 29968
rect 3715 29924 3773 29925
rect 3715 29884 3724 29924
rect 3764 29884 3773 29924
rect 3715 29883 3773 29884
rect 4099 29924 4157 29925
rect 4099 29884 4108 29924
rect 4148 29884 4157 29924
rect 4099 29883 4157 29884
rect 4587 29924 4629 29933
rect 4587 29884 4588 29924
rect 4628 29884 4629 29924
rect 4587 29875 4629 29884
rect 29739 29924 29781 29933
rect 29739 29884 29740 29924
rect 29780 29884 29781 29924
rect 29739 29875 29781 29884
rect 5251 29840 5309 29841
rect 5251 29800 5260 29840
rect 5300 29800 5309 29840
rect 5251 29799 5309 29800
rect 10147 29840 10205 29841
rect 10147 29800 10156 29840
rect 10196 29800 10205 29840
rect 10147 29799 10205 29800
rect 10531 29840 10589 29841
rect 10531 29800 10540 29840
rect 10580 29800 10589 29840
rect 10531 29799 10589 29800
rect 10915 29840 10973 29841
rect 10915 29800 10924 29840
rect 10964 29800 10973 29840
rect 10915 29799 10973 29800
rect 14379 29840 14421 29849
rect 14379 29800 14380 29840
rect 14420 29800 14421 29840
rect 14379 29791 14421 29800
rect 14755 29840 14813 29841
rect 14755 29800 14764 29840
rect 14804 29800 14813 29840
rect 14755 29799 14813 29800
rect 15619 29840 15677 29841
rect 15619 29800 15628 29840
rect 15668 29800 15677 29840
rect 15619 29799 15677 29800
rect 17923 29840 17981 29841
rect 17923 29800 17932 29840
rect 17972 29800 17981 29840
rect 17923 29799 17981 29800
rect 20811 29840 20853 29849
rect 20811 29800 20812 29840
rect 20852 29800 20853 29840
rect 20811 29791 20853 29800
rect 21187 29840 21245 29841
rect 21187 29800 21196 29840
rect 21236 29800 21245 29840
rect 21187 29799 21245 29800
rect 22051 29840 22109 29841
rect 22051 29800 22060 29840
rect 22100 29800 22109 29840
rect 22051 29799 22109 29800
rect 25315 29840 25373 29841
rect 25315 29800 25324 29840
rect 25364 29800 25373 29840
rect 25315 29799 25373 29800
rect 25603 29840 25661 29841
rect 25603 29800 25612 29840
rect 25652 29800 25661 29840
rect 25603 29799 25661 29800
rect 26083 29840 26141 29841
rect 26083 29800 26092 29840
rect 26132 29800 26141 29840
rect 26083 29799 26141 29800
rect 27043 29840 27101 29841
rect 27043 29800 27052 29840
rect 27092 29800 27101 29840
rect 27043 29799 27101 29800
rect 27339 29840 27381 29849
rect 27339 29800 27340 29840
rect 27380 29800 27381 29840
rect 27339 29791 27381 29800
rect 27715 29840 27773 29841
rect 27715 29800 27724 29840
rect 27764 29800 27773 29840
rect 27715 29799 27773 29800
rect 28579 29840 28637 29841
rect 28579 29800 28588 29840
rect 28628 29800 28637 29840
rect 28579 29799 28637 29800
rect 30019 29840 30077 29841
rect 30019 29800 30028 29840
rect 30068 29800 30077 29840
rect 30019 29799 30077 29800
rect 30403 29840 30461 29841
rect 30403 29800 30412 29840
rect 30452 29800 30461 29840
rect 30403 29799 30461 29800
rect 39619 29840 39677 29841
rect 39619 29800 39628 29840
rect 39668 29800 39677 29840
rect 39619 29799 39677 29800
rect 44515 29840 44573 29841
rect 44515 29800 44524 29840
rect 44564 29800 44573 29840
rect 44515 29799 44573 29800
rect 44811 29840 44853 29849
rect 44811 29800 44812 29840
rect 44852 29800 44853 29840
rect 44811 29791 44853 29800
rect 44995 29840 45053 29841
rect 44995 29800 45004 29840
rect 45044 29800 45053 29840
rect 44995 29799 45053 29800
rect 45283 29840 45341 29841
rect 45283 29800 45292 29840
rect 45332 29800 45341 29840
rect 45283 29799 45341 29800
rect 46923 29840 46965 29849
rect 46923 29800 46924 29840
rect 46964 29800 46965 29840
rect 46923 29791 46965 29800
rect 47299 29840 47357 29841
rect 47299 29800 47308 29840
rect 47348 29800 47357 29840
rect 47299 29799 47357 29800
rect 48163 29840 48221 29841
rect 48163 29800 48172 29840
rect 48212 29800 48221 29840
rect 48163 29799 48221 29800
rect 3531 29672 3573 29681
rect 3531 29632 3532 29672
rect 3572 29632 3573 29672
rect 3531 29623 3573 29632
rect 11019 29672 11061 29681
rect 11019 29632 11020 29672
rect 11060 29632 11061 29672
rect 11019 29623 11061 29632
rect 25803 29672 25845 29681
rect 25803 29632 25804 29672
rect 25844 29632 25845 29672
rect 25803 29623 25845 29632
rect 30507 29672 30549 29681
rect 30507 29632 30508 29672
rect 30548 29632 30549 29672
rect 30507 29623 30549 29632
rect 40291 29672 40349 29673
rect 40291 29632 40300 29672
rect 40340 29632 40349 29672
rect 40291 29631 40349 29632
rect 45771 29672 45813 29681
rect 45771 29632 45772 29672
rect 45812 29632 45813 29672
rect 45771 29623 45813 29632
rect 576 29504 99360 29528
rect 576 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 19472 29504
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19840 29464 34592 29504
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34960 29464 49712 29504
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 50080 29464 64832 29504
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 65200 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 95072 29504
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95440 29464 99360 29504
rect 576 29440 99360 29464
rect 5155 29336 5213 29337
rect 5155 29296 5164 29336
rect 5204 29296 5213 29336
rect 5155 29295 5213 29296
rect 10243 29336 10301 29337
rect 10243 29296 10252 29336
rect 10292 29296 10301 29336
rect 10243 29295 10301 29296
rect 15051 29336 15093 29345
rect 15051 29296 15052 29336
rect 15092 29296 15093 29336
rect 15051 29287 15093 29296
rect 17827 29336 17885 29337
rect 17827 29296 17836 29336
rect 17876 29296 17885 29336
rect 17827 29295 17885 29296
rect 44803 29336 44861 29337
rect 44803 29296 44812 29336
rect 44852 29296 44861 29336
rect 44803 29295 44861 29296
rect 2763 29252 2805 29261
rect 2763 29212 2764 29252
rect 2804 29212 2805 29252
rect 2763 29203 2805 29212
rect 3139 29168 3197 29169
rect 3139 29128 3148 29168
rect 3188 29128 3197 29168
rect 3139 29127 3197 29128
rect 4003 29168 4061 29169
rect 4003 29128 4012 29168
rect 4052 29128 4061 29168
rect 4003 29127 4061 29128
rect 7851 29168 7893 29177
rect 7851 29128 7852 29168
rect 7892 29128 7893 29168
rect 7851 29119 7893 29128
rect 8227 29168 8285 29169
rect 8227 29128 8236 29168
rect 8276 29128 8285 29168
rect 8227 29127 8285 29128
rect 9091 29168 9149 29169
rect 9091 29128 9100 29168
rect 9140 29128 9149 29168
rect 9091 29127 9149 29128
rect 11875 29168 11933 29169
rect 11875 29128 11884 29168
rect 11924 29128 11933 29168
rect 11875 29127 11933 29128
rect 15435 29168 15477 29177
rect 15435 29128 15436 29168
rect 15476 29128 15477 29168
rect 15435 29119 15477 29128
rect 15811 29168 15869 29169
rect 15811 29128 15820 29168
rect 15860 29128 15869 29168
rect 15811 29127 15869 29128
rect 16675 29168 16733 29169
rect 16675 29128 16684 29168
rect 16724 29128 16733 29168
rect 16675 29127 16733 29128
rect 22147 29168 22205 29169
rect 22147 29128 22156 29168
rect 22196 29128 22205 29168
rect 22147 29127 22205 29128
rect 23107 29168 23165 29169
rect 23107 29128 23116 29168
rect 23156 29128 23165 29168
rect 23107 29127 23165 29128
rect 26083 29168 26141 29169
rect 26083 29128 26092 29168
rect 26132 29128 26141 29168
rect 26083 29127 26141 29128
rect 30595 29168 30653 29169
rect 30595 29128 30604 29168
rect 30644 29128 30653 29168
rect 30595 29127 30653 29128
rect 39907 29168 39965 29169
rect 39907 29128 39916 29168
rect 39956 29128 39965 29168
rect 39907 29127 39965 29128
rect 40867 29168 40925 29169
rect 40867 29128 40876 29168
rect 40916 29128 40925 29168
rect 40867 29127 40925 29128
rect 45475 29168 45533 29169
rect 45475 29128 45484 29168
rect 45524 29128 45533 29168
rect 45475 29127 45533 29128
rect 15235 29084 15293 29085
rect 15235 29044 15244 29084
rect 15284 29044 15293 29084
rect 15235 29043 15293 29044
rect 44611 29084 44669 29085
rect 44611 29044 44620 29084
rect 44660 29044 44669 29084
rect 44611 29043 44669 29044
rect 22635 29000 22677 29009
rect 22635 28960 22636 29000
rect 22676 28960 22677 29000
rect 22635 28951 22677 28960
rect 40395 29000 40437 29009
rect 40395 28960 40396 29000
rect 40436 28960 40437 29000
rect 40395 28951 40437 28960
rect 11203 28916 11261 28917
rect 11203 28876 11212 28916
rect 11252 28876 11261 28916
rect 11203 28875 11261 28876
rect 26755 28916 26813 28917
rect 26755 28876 26764 28916
rect 26804 28876 26813 28916
rect 26755 28875 26813 28876
rect 29923 28916 29981 28917
rect 29923 28876 29932 28916
rect 29972 28876 29981 28916
rect 29923 28875 29981 28876
rect 44427 28916 44469 28925
rect 44427 28876 44428 28916
rect 44468 28876 44469 28916
rect 44427 28867 44469 28876
rect 576 28748 99360 28772
rect 576 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 18232 28748
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18600 28708 33352 28748
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33720 28708 48472 28748
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48840 28708 63592 28748
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63960 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 93832 28748
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 94200 28708 99360 28748
rect 576 28684 99360 28708
rect 16203 28580 16245 28589
rect 16203 28540 16204 28580
rect 16244 28540 16245 28580
rect 16203 28531 16245 28540
rect 40491 28580 40533 28589
rect 40491 28540 40492 28580
rect 40532 28540 40533 28580
rect 40491 28531 40533 28540
rect 46915 28580 46973 28581
rect 46915 28540 46924 28580
rect 46964 28540 46973 28580
rect 46915 28539 46973 28540
rect 19947 28496 19989 28505
rect 19947 28456 19948 28496
rect 19988 28456 19989 28496
rect 19947 28447 19989 28456
rect 40299 28496 40341 28505
rect 40299 28456 40300 28496
rect 40340 28456 40341 28496
rect 40299 28447 40341 28456
rect 16387 28412 16445 28413
rect 16387 28372 16396 28412
rect 16436 28372 16445 28412
rect 16387 28371 16445 28372
rect 19267 28412 19325 28413
rect 19267 28372 19276 28412
rect 19316 28372 19325 28412
rect 19267 28371 19325 28372
rect 28771 28412 28829 28413
rect 28771 28372 28780 28412
rect 28820 28372 28829 28412
rect 28771 28371 28829 28372
rect 19651 28328 19709 28329
rect 19651 28288 19660 28328
rect 19700 28288 19709 28328
rect 19651 28287 19709 28288
rect 20611 28328 20669 28329
rect 20611 28288 20620 28328
rect 20660 28288 20669 28328
rect 20611 28287 20669 28288
rect 27139 28328 27197 28329
rect 27139 28288 27148 28328
rect 27188 28288 27197 28328
rect 27139 28287 27197 28288
rect 29059 28328 29117 28329
rect 29059 28288 29068 28328
rect 29108 28288 29117 28328
rect 29059 28287 29117 28288
rect 29163 28328 29205 28337
rect 29163 28288 29164 28328
rect 29204 28288 29205 28328
rect 29163 28279 29205 28288
rect 32899 28328 32957 28329
rect 32899 28288 32908 28328
rect 32948 28288 32957 28328
rect 32899 28287 32957 28288
rect 33859 28328 33917 28329
rect 33859 28288 33868 28328
rect 33908 28288 33917 28328
rect 33859 28287 33917 28288
rect 40963 28328 41021 28329
rect 40963 28288 40972 28328
rect 41012 28288 41021 28328
rect 40963 28287 41021 28288
rect 44523 28328 44565 28337
rect 44523 28288 44524 28328
rect 44564 28288 44565 28328
rect 44523 28279 44565 28288
rect 44899 28328 44957 28329
rect 44899 28288 44908 28328
rect 44948 28288 44957 28328
rect 44899 28287 44957 28288
rect 45763 28328 45821 28329
rect 45763 28288 45772 28328
rect 45812 28288 45821 28328
rect 45763 28287 45821 28288
rect 26467 28160 26525 28161
rect 26467 28120 26476 28160
rect 26516 28120 26525 28160
rect 26467 28119 26525 28120
rect 576 27992 99360 28016
rect 576 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 19472 27992
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19840 27952 34592 27992
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34960 27952 49712 27992
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 50080 27952 64832 27992
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 65200 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 95072 27992
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95440 27952 99360 27992
rect 576 27928 99360 27952
rect 4963 27824 5021 27825
rect 4963 27784 4972 27824
rect 5012 27784 5021 27824
rect 4963 27783 5021 27784
rect 4299 27740 4341 27749
rect 4299 27700 4300 27740
rect 4340 27700 4341 27740
rect 4299 27691 4341 27700
rect 4683 27740 4725 27749
rect 4683 27700 4684 27740
rect 4724 27700 4725 27740
rect 4683 27691 4725 27700
rect 5923 27740 5981 27741
rect 5923 27700 5932 27740
rect 5972 27700 5981 27740
rect 5923 27699 5981 27700
rect 26187 27740 26229 27749
rect 26187 27700 26188 27740
rect 26228 27700 26229 27740
rect 26187 27691 26229 27700
rect 4203 27656 4245 27665
rect 4203 27616 4204 27656
rect 4244 27616 4245 27656
rect 4203 27607 4245 27616
rect 4387 27656 4445 27657
rect 4387 27616 4396 27656
rect 4436 27616 4445 27656
rect 4387 27615 4445 27616
rect 4587 27656 4629 27665
rect 4587 27616 4588 27656
rect 4628 27616 4629 27656
rect 4587 27607 4629 27616
rect 4771 27656 4829 27657
rect 4771 27616 4780 27656
rect 4820 27616 4829 27656
rect 4771 27615 4829 27616
rect 5059 27656 5117 27657
rect 5059 27616 5068 27656
rect 5108 27616 5117 27656
rect 5059 27615 5117 27616
rect 5443 27656 5501 27657
rect 5443 27616 5452 27656
rect 5492 27616 5501 27656
rect 5443 27615 5501 27616
rect 5731 27656 5789 27657
rect 5731 27616 5740 27656
rect 5780 27616 5789 27656
rect 5731 27615 5789 27616
rect 9763 27656 9821 27657
rect 9763 27616 9772 27656
rect 9812 27616 9821 27656
rect 9763 27615 9821 27616
rect 11107 27656 11165 27657
rect 11107 27616 11116 27656
rect 11156 27616 11165 27656
rect 11107 27615 11165 27616
rect 11203 27656 11261 27657
rect 11203 27616 11212 27656
rect 11252 27616 11261 27656
rect 11203 27615 11261 27616
rect 11587 27656 11645 27657
rect 11587 27616 11596 27656
rect 11636 27616 11645 27656
rect 11587 27615 11645 27616
rect 26563 27656 26621 27657
rect 26563 27616 26572 27656
rect 26612 27616 26621 27656
rect 26563 27615 26621 27616
rect 27427 27656 27485 27657
rect 27427 27616 27436 27656
rect 27476 27616 27485 27656
rect 27427 27615 27485 27616
rect 28771 27656 28829 27657
rect 28771 27616 28780 27656
rect 28820 27616 28829 27656
rect 28771 27615 28829 27616
rect 33667 27656 33725 27657
rect 33667 27616 33676 27656
rect 33716 27616 33725 27656
rect 33667 27615 33725 27616
rect 34531 27656 34589 27657
rect 34531 27616 34540 27656
rect 34580 27616 34589 27656
rect 34531 27615 34589 27616
rect 34923 27656 34965 27665
rect 34923 27616 34924 27656
rect 34964 27616 34965 27656
rect 34923 27607 34965 27616
rect 39619 27656 39677 27657
rect 39619 27616 39628 27656
rect 39668 27616 39677 27656
rect 39619 27615 39677 27616
rect 40483 27656 40541 27657
rect 40483 27616 40492 27656
rect 40532 27616 40541 27656
rect 40483 27615 40541 27616
rect 40875 27656 40917 27665
rect 40875 27616 40876 27656
rect 40916 27616 40917 27656
rect 40875 27607 40917 27616
rect 11395 27572 11453 27573
rect 11395 27532 11404 27572
rect 11444 27532 11453 27572
rect 11395 27531 11453 27532
rect 28587 27572 28629 27581
rect 28587 27532 28588 27572
rect 28628 27532 28629 27572
rect 28587 27523 28629 27532
rect 5251 27404 5309 27405
rect 5251 27364 5260 27404
rect 5300 27364 5309 27404
rect 5251 27363 5309 27364
rect 9483 27404 9525 27413
rect 9483 27364 9484 27404
rect 9524 27364 9525 27404
rect 9483 27355 9525 27364
rect 12259 27404 12317 27405
rect 12259 27364 12268 27404
rect 12308 27364 12317 27404
rect 12259 27363 12317 27364
rect 29443 27404 29501 27405
rect 29443 27364 29452 27404
rect 29492 27364 29501 27404
rect 29443 27363 29501 27364
rect 32515 27404 32573 27405
rect 32515 27364 32524 27404
rect 32564 27364 32573 27404
rect 32515 27363 32573 27364
rect 38475 27404 38517 27413
rect 38475 27364 38476 27404
rect 38516 27364 38517 27404
rect 38475 27355 38517 27364
rect 576 27236 99360 27260
rect 576 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 18232 27236
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18600 27196 33352 27236
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33720 27196 48472 27236
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48840 27196 63592 27236
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63960 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 93832 27236
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 94200 27196 99360 27236
rect 576 27172 99360 27196
rect 4195 27068 4253 27069
rect 4195 27028 4204 27068
rect 4244 27028 4253 27068
rect 4195 27027 4253 27028
rect 5059 27068 5117 27069
rect 5059 27028 5068 27068
rect 5108 27028 5117 27068
rect 5059 27027 5117 27028
rect 11115 27068 11157 27077
rect 11115 27028 11116 27068
rect 11156 27028 11157 27068
rect 11115 27019 11157 27028
rect 28779 27068 28821 27077
rect 28779 27028 28780 27068
rect 28820 27028 28821 27068
rect 28779 27019 28821 27028
rect 3427 26900 3485 26901
rect 3427 26860 3436 26900
rect 3476 26860 3485 26900
rect 3427 26859 3485 26860
rect 3811 26900 3869 26901
rect 3811 26860 3820 26900
rect 3860 26860 3869 26900
rect 3811 26859 3869 26860
rect 42699 26900 42741 26909
rect 42699 26860 42700 26900
rect 42740 26860 42741 26900
rect 42699 26851 42741 26860
rect 4867 26816 4925 26817
rect 4867 26776 4876 26816
rect 4916 26776 4925 26816
rect 4867 26775 4925 26776
rect 5731 26816 5789 26817
rect 5731 26776 5740 26816
rect 5780 26776 5789 26816
rect 5731 26775 5789 26776
rect 10147 26816 10205 26817
rect 10147 26776 10156 26816
rect 10196 26776 10205 26816
rect 10147 26775 10205 26776
rect 11011 26816 11069 26817
rect 11011 26776 11020 26816
rect 11060 26776 11069 26816
rect 11011 26775 11069 26776
rect 11211 26816 11253 26825
rect 11211 26776 11212 26816
rect 11252 26776 11253 26816
rect 11211 26767 11253 26776
rect 28683 26816 28725 26825
rect 28683 26776 28684 26816
rect 28724 26776 28725 26816
rect 28683 26767 28725 26776
rect 28867 26816 28925 26817
rect 28867 26776 28876 26816
rect 28916 26776 28925 26816
rect 28867 26775 28925 26776
rect 33187 26816 33245 26817
rect 33187 26776 33196 26816
rect 33236 26776 33245 26816
rect 33187 26775 33245 26776
rect 34435 26816 34493 26817
rect 34435 26776 34444 26816
rect 34484 26776 34493 26816
rect 34435 26775 34493 26776
rect 35299 26816 35357 26817
rect 35299 26776 35308 26816
rect 35348 26776 35357 26816
rect 35299 26775 35357 26776
rect 40675 26816 40733 26817
rect 40675 26776 40684 26816
rect 40724 26776 40733 26816
rect 40675 26775 40733 26776
rect 41539 26816 41597 26817
rect 41539 26776 41548 26816
rect 41588 26776 41597 26816
rect 41539 26775 41597 26776
rect 42883 26816 42941 26817
rect 42883 26776 42892 26816
rect 42932 26776 42941 26816
rect 42883 26775 42941 26776
rect 34059 26732 34101 26741
rect 34059 26692 34060 26732
rect 34100 26692 34101 26732
rect 34059 26683 34101 26692
rect 40299 26732 40341 26741
rect 40299 26692 40300 26732
rect 40340 26692 40341 26732
rect 40299 26683 40341 26692
rect 3243 26648 3285 26657
rect 3243 26608 3244 26648
rect 3284 26608 3285 26648
rect 3243 26599 3285 26608
rect 3627 26648 3669 26657
rect 3627 26608 3628 26648
rect 3668 26608 3669 26648
rect 3627 26599 3669 26608
rect 10819 26648 10877 26649
rect 10819 26608 10828 26648
rect 10868 26608 10877 26648
rect 10819 26607 10877 26608
rect 33859 26648 33917 26649
rect 33859 26608 33868 26648
rect 33908 26608 33917 26648
rect 33859 26607 33917 26608
rect 36451 26648 36509 26649
rect 36451 26608 36460 26648
rect 36500 26608 36509 26648
rect 36451 26607 36509 26608
rect 43555 26648 43613 26649
rect 43555 26608 43564 26648
rect 43604 26608 43613 26648
rect 43555 26607 43613 26608
rect 576 26480 99360 26504
rect 576 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 19472 26480
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19840 26440 34592 26480
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34960 26440 49712 26480
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 50080 26440 64832 26480
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 65200 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 95072 26480
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95440 26440 99360 26480
rect 576 26416 99360 26440
rect 4867 26312 4925 26313
rect 4867 26272 4876 26312
rect 4916 26272 4925 26312
rect 4867 26271 4925 26272
rect 9475 26312 9533 26313
rect 9475 26272 9484 26312
rect 9524 26272 9533 26312
rect 9475 26271 9533 26272
rect 33579 26312 33621 26321
rect 33579 26272 33580 26312
rect 33620 26272 33621 26312
rect 33579 26263 33621 26272
rect 34059 26312 34101 26321
rect 34059 26272 34060 26312
rect 34100 26272 34101 26312
rect 34059 26263 34101 26272
rect 41451 26312 41493 26321
rect 41451 26272 41452 26312
rect 41492 26272 41493 26312
rect 41451 26263 41493 26272
rect 43947 26312 43989 26321
rect 43947 26272 43948 26312
rect 43988 26272 43989 26312
rect 43947 26263 43989 26272
rect 2475 26228 2517 26237
rect 2475 26188 2476 26228
rect 2516 26188 2517 26228
rect 2475 26179 2517 26188
rect 7083 26228 7125 26237
rect 7083 26188 7084 26228
rect 7124 26188 7125 26228
rect 7083 26179 7125 26188
rect 10531 26228 10589 26229
rect 10531 26188 10540 26228
rect 10580 26188 10589 26228
rect 10531 26187 10589 26188
rect 11691 26228 11733 26237
rect 11691 26188 11692 26228
rect 11732 26188 11733 26228
rect 11691 26179 11733 26188
rect 23979 26228 24021 26237
rect 23979 26188 23980 26228
rect 24020 26188 24021 26228
rect 23979 26179 24021 26188
rect 28675 26228 28733 26229
rect 28675 26188 28684 26228
rect 28724 26188 28733 26228
rect 28675 26187 28733 26188
rect 2851 26144 2909 26145
rect 2851 26104 2860 26144
rect 2900 26104 2909 26144
rect 2851 26103 2909 26104
rect 3715 26144 3773 26145
rect 3715 26104 3724 26144
rect 3764 26104 3773 26144
rect 3715 26103 3773 26104
rect 7459 26144 7517 26145
rect 7459 26104 7468 26144
rect 7508 26104 7517 26144
rect 7459 26103 7517 26104
rect 8323 26144 8381 26145
rect 8323 26104 8332 26144
rect 8372 26104 8381 26144
rect 8323 26103 8381 26104
rect 10051 26144 10109 26145
rect 10051 26104 10060 26144
rect 10100 26104 10109 26144
rect 10051 26103 10109 26104
rect 10435 26144 10493 26145
rect 10435 26104 10444 26144
rect 10484 26104 10493 26144
rect 10435 26103 10493 26104
rect 10819 26144 10877 26145
rect 10819 26104 10828 26144
rect 10868 26104 10877 26144
rect 10819 26103 10877 26104
rect 12067 26144 12125 26145
rect 12067 26104 12076 26144
rect 12116 26104 12125 26144
rect 12067 26103 12125 26104
rect 12931 26144 12989 26145
rect 12931 26104 12940 26144
rect 12980 26104 12989 26144
rect 12931 26103 12989 26104
rect 17827 26144 17885 26145
rect 17827 26104 17836 26144
rect 17876 26104 17885 26144
rect 17827 26103 17885 26104
rect 18507 26144 18549 26153
rect 18507 26104 18508 26144
rect 18548 26104 18549 26144
rect 18507 26095 18549 26104
rect 18699 26144 18741 26153
rect 18699 26104 18700 26144
rect 18740 26104 18741 26144
rect 18699 26095 18741 26104
rect 19075 26144 19133 26145
rect 19075 26104 19084 26144
rect 19124 26104 19133 26144
rect 19075 26103 19133 26104
rect 19939 26144 19997 26145
rect 19939 26104 19948 26144
rect 19988 26104 19997 26144
rect 19939 26103 19997 26104
rect 22723 26144 22781 26145
rect 22723 26104 22732 26144
rect 22772 26104 22781 26144
rect 22723 26103 22781 26104
rect 23587 26144 23645 26145
rect 23587 26104 23596 26144
rect 23636 26104 23645 26144
rect 23587 26103 23645 26104
rect 28387 26144 28445 26145
rect 28387 26104 28396 26144
rect 28436 26104 28445 26144
rect 28387 26103 28445 26104
rect 28771 26144 28829 26145
rect 28771 26104 28780 26144
rect 28820 26104 28829 26144
rect 28771 26103 28829 26104
rect 29155 26144 29213 26145
rect 29155 26104 29164 26144
rect 29204 26104 29213 26144
rect 29155 26103 29213 26104
rect 35107 26144 35165 26145
rect 35107 26104 35116 26144
rect 35156 26104 35165 26144
rect 35107 26103 35165 26104
rect 35587 26144 35645 26145
rect 35587 26104 35596 26144
rect 35636 26104 35645 26144
rect 35587 26103 35645 26104
rect 36547 26144 36605 26145
rect 36547 26104 36556 26144
rect 36596 26104 36605 26144
rect 36547 26103 36605 26104
rect 44419 26144 44477 26145
rect 44419 26104 44428 26144
rect 44468 26104 44477 26144
rect 44419 26103 44477 26104
rect 47011 26144 47069 26145
rect 47011 26104 47020 26144
rect 47060 26104 47069 26144
rect 47011 26103 47069 26104
rect 33379 26060 33437 26061
rect 33379 26020 33388 26060
rect 33428 26020 33437 26060
rect 33379 26019 33437 26020
rect 34243 26060 34301 26061
rect 34243 26020 34252 26060
rect 34292 26020 34301 26060
rect 34243 26019 34301 26020
rect 41635 26060 41693 26061
rect 41635 26020 41644 26060
rect 41684 26020 41693 26060
rect 41635 26019 41693 26020
rect 11491 25892 11549 25893
rect 11491 25852 11500 25892
rect 11540 25852 11549 25892
rect 11491 25851 11549 25852
rect 14083 25892 14141 25893
rect 14083 25852 14092 25892
rect 14132 25852 14141 25892
rect 14083 25851 14141 25852
rect 21091 25892 21149 25893
rect 21091 25852 21100 25892
rect 21140 25852 21149 25892
rect 21091 25851 21149 25852
rect 21571 25892 21629 25893
rect 21571 25852 21580 25892
rect 21620 25852 21629 25892
rect 21571 25851 21629 25852
rect 27715 25892 27773 25893
rect 27715 25852 27724 25892
rect 27764 25852 27773 25892
rect 27715 25851 27773 25852
rect 34435 25892 34493 25893
rect 34435 25852 34444 25892
rect 34484 25852 34493 25892
rect 34435 25851 34493 25852
rect 46339 25892 46397 25893
rect 46339 25852 46348 25892
rect 46388 25852 46397 25892
rect 46339 25851 46397 25852
rect 576 25724 99360 25748
rect 576 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 18232 25724
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18600 25684 33352 25724
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33720 25684 48472 25724
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48840 25684 63592 25724
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63960 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 93832 25724
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 94200 25684 99360 25724
rect 576 25660 99360 25684
rect 4771 25556 4829 25557
rect 4771 25516 4780 25556
rect 4820 25516 4829 25556
rect 4771 25515 4829 25516
rect 6123 25556 6165 25565
rect 6123 25516 6124 25556
rect 6164 25516 6165 25556
rect 6123 25507 6165 25516
rect 16875 25556 16917 25565
rect 16875 25516 16876 25556
rect 16916 25516 16917 25556
rect 16875 25507 16917 25516
rect 28971 25556 29013 25565
rect 28971 25516 28972 25556
rect 29012 25516 29013 25556
rect 28971 25507 29013 25516
rect 47587 25556 47645 25557
rect 47587 25516 47596 25556
rect 47636 25516 47645 25556
rect 47587 25515 47645 25516
rect 24555 25472 24597 25481
rect 24555 25432 24556 25472
rect 24596 25432 24597 25472
rect 24555 25423 24597 25432
rect 2379 25304 2421 25313
rect 2379 25264 2380 25304
rect 2420 25264 2421 25304
rect 2379 25255 2421 25264
rect 2755 25304 2813 25305
rect 2755 25264 2764 25304
rect 2804 25264 2813 25304
rect 2755 25263 2813 25264
rect 3619 25304 3677 25305
rect 3619 25264 3628 25304
rect 3668 25264 3677 25304
rect 3619 25263 3677 25264
rect 5827 25304 5885 25305
rect 5827 25264 5836 25304
rect 5876 25264 5885 25304
rect 5827 25263 5885 25264
rect 6787 25304 6845 25305
rect 6787 25264 6796 25304
rect 6836 25264 6845 25304
rect 6787 25263 6845 25264
rect 11403 25304 11445 25313
rect 11403 25264 11404 25304
rect 11444 25264 11445 25304
rect 11403 25255 11445 25264
rect 11779 25304 11837 25305
rect 11779 25264 11788 25304
rect 11828 25264 11837 25304
rect 11779 25263 11837 25264
rect 12643 25304 12701 25305
rect 12643 25264 12652 25304
rect 12692 25264 12701 25304
rect 12643 25263 12701 25264
rect 16587 25304 16629 25313
rect 16587 25264 16588 25304
rect 16628 25264 16629 25304
rect 16587 25255 16629 25264
rect 16675 25304 16733 25305
rect 16675 25264 16684 25304
rect 16724 25264 16733 25304
rect 16675 25263 16733 25264
rect 21763 25304 21821 25305
rect 21763 25264 21772 25304
rect 21812 25264 21821 25304
rect 21763 25263 21821 25264
rect 22051 25304 22109 25305
rect 22051 25264 22060 25304
rect 22100 25264 22109 25304
rect 22051 25263 22109 25264
rect 24259 25304 24317 25305
rect 24259 25264 24268 25304
rect 24308 25264 24317 25304
rect 24259 25263 24317 25264
rect 28779 25304 28821 25313
rect 28779 25264 28780 25304
rect 28820 25264 28821 25304
rect 28779 25255 28821 25264
rect 29635 25304 29693 25305
rect 29635 25264 29644 25304
rect 29684 25264 29693 25304
rect 29635 25263 29693 25264
rect 45571 25304 45629 25305
rect 45571 25264 45580 25304
rect 45620 25264 45629 25304
rect 45571 25263 45629 25264
rect 46435 25304 46493 25305
rect 46435 25264 46444 25304
rect 46484 25264 46493 25304
rect 46435 25263 46493 25264
rect 25123 25220 25181 25221
rect 25123 25180 25132 25220
rect 25172 25180 25181 25220
rect 25123 25179 25181 25180
rect 45195 25220 45237 25229
rect 45195 25180 45196 25220
rect 45236 25180 45237 25220
rect 45195 25171 45237 25180
rect 13795 25136 13853 25137
rect 13795 25096 13804 25136
rect 13844 25096 13853 25136
rect 13795 25095 13853 25096
rect 22251 25136 22293 25145
rect 22251 25096 22252 25136
rect 22292 25096 22293 25136
rect 22251 25087 22293 25096
rect 576 24968 99360 24992
rect 576 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 19472 24968
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19840 24928 34592 24968
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34960 24928 49712 24968
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 50080 24928 64832 24968
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 65200 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 95072 24968
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95440 24928 99360 24968
rect 576 24904 99360 24928
rect 16587 24800 16629 24809
rect 16587 24760 16588 24800
rect 16628 24760 16629 24800
rect 16587 24751 16629 24760
rect 45099 24800 45141 24809
rect 45099 24760 45100 24800
rect 45140 24760 45141 24800
rect 45099 24751 45141 24760
rect 12739 24716 12797 24717
rect 12739 24676 12748 24716
rect 12788 24676 12797 24716
rect 12739 24675 12797 24676
rect 16971 24716 17013 24725
rect 16971 24676 16972 24716
rect 17012 24676 17013 24716
rect 16971 24667 17013 24676
rect 22923 24716 22965 24725
rect 22923 24676 22924 24716
rect 22964 24676 22965 24716
rect 22923 24667 22965 24676
rect 27147 24716 27189 24725
rect 27147 24676 27148 24716
rect 27188 24676 27189 24716
rect 27147 24667 27189 24676
rect 11875 24632 11933 24633
rect 11875 24592 11884 24632
rect 11924 24592 11933 24632
rect 11875 24591 11933 24592
rect 15235 24632 15293 24633
rect 15235 24592 15244 24632
rect 15284 24592 15293 24632
rect 15235 24591 15293 24592
rect 16099 24632 16157 24633
rect 16099 24592 16108 24632
rect 16148 24592 16157 24632
rect 16099 24591 16157 24592
rect 16387 24632 16445 24633
rect 16387 24592 16396 24632
rect 16436 24592 16445 24632
rect 16387 24591 16445 24592
rect 16867 24632 16925 24633
rect 16867 24592 16876 24632
rect 16916 24592 16925 24632
rect 16867 24591 16925 24592
rect 17067 24632 17109 24641
rect 17067 24592 17068 24632
rect 17108 24592 17109 24632
rect 17067 24583 17109 24592
rect 20907 24632 20949 24641
rect 20907 24592 20908 24632
rect 20948 24592 20949 24632
rect 20907 24583 20949 24592
rect 21091 24632 21149 24633
rect 21091 24592 21100 24632
rect 21140 24592 21149 24632
rect 21091 24591 21149 24592
rect 23587 24632 23645 24633
rect 23587 24592 23596 24632
rect 23636 24592 23645 24632
rect 23587 24591 23645 24592
rect 25891 24632 25949 24633
rect 25891 24592 25900 24632
rect 25940 24592 25949 24632
rect 25891 24591 25949 24592
rect 26755 24632 26813 24633
rect 26755 24592 26764 24632
rect 26804 24592 26813 24632
rect 26755 24591 26813 24592
rect 33859 24632 33917 24633
rect 33859 24592 33868 24632
rect 33908 24592 33917 24632
rect 33859 24591 33917 24592
rect 34059 24632 34101 24641
rect 34059 24592 34060 24632
rect 34100 24592 34101 24632
rect 34059 24583 34101 24592
rect 35115 24632 35157 24641
rect 35115 24592 35116 24632
rect 35156 24592 35157 24632
rect 35115 24583 35157 24592
rect 43363 24632 43421 24633
rect 43363 24592 43372 24632
rect 43412 24592 43421 24632
rect 43363 24591 43421 24592
rect 43563 24632 43605 24641
rect 43563 24592 43564 24632
rect 43604 24592 43605 24632
rect 43563 24583 43605 24592
rect 46155 24632 46197 24641
rect 46155 24592 46156 24632
rect 46196 24592 46197 24632
rect 46155 24583 46197 24592
rect 46539 24632 46581 24641
rect 46539 24592 46540 24632
rect 46580 24592 46581 24632
rect 46539 24583 46581 24592
rect 46915 24632 46973 24633
rect 46915 24592 46924 24632
rect 46964 24592 46973 24632
rect 46915 24591 46973 24592
rect 47779 24632 47837 24633
rect 47779 24592 47788 24632
rect 47828 24592 47837 24632
rect 47779 24591 47837 24592
rect 24747 24548 24789 24557
rect 24747 24508 24748 24548
rect 24788 24508 24789 24548
rect 24747 24499 24789 24508
rect 31459 24548 31517 24549
rect 31459 24508 31468 24548
rect 31508 24508 31517 24548
rect 31459 24507 31517 24508
rect 44899 24548 44957 24549
rect 44899 24508 44908 24548
rect 44948 24508 44957 24548
rect 44899 24507 44957 24508
rect 12171 24464 12213 24473
rect 12171 24424 12172 24464
rect 12212 24424 12213 24464
rect 12171 24415 12213 24424
rect 15907 24464 15965 24465
rect 15907 24424 15916 24464
rect 15956 24424 15965 24464
rect 15907 24423 15965 24424
rect 21003 24380 21045 24389
rect 21003 24340 21004 24380
rect 21044 24340 21045 24380
rect 21003 24331 21045 24340
rect 31275 24380 31317 24389
rect 31275 24340 31276 24380
rect 31316 24340 31317 24380
rect 31275 24331 31317 24340
rect 33963 24380 34005 24389
rect 33963 24340 33964 24380
rect 34004 24340 34005 24380
rect 33963 24331 34005 24340
rect 34923 24380 34965 24389
rect 34923 24340 34924 24380
rect 34964 24340 34965 24380
rect 34923 24331 34965 24340
rect 43467 24380 43509 24389
rect 43467 24340 43468 24380
rect 43508 24340 43509 24380
rect 43467 24331 43509 24340
rect 45963 24380 46005 24389
rect 45963 24340 45964 24380
rect 46004 24340 46005 24380
rect 45963 24331 46005 24340
rect 48931 24380 48989 24381
rect 48931 24340 48940 24380
rect 48980 24340 48989 24380
rect 48931 24339 48989 24340
rect 576 24212 99360 24236
rect 576 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 18232 24212
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18600 24172 33352 24212
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33720 24172 48472 24212
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48840 24172 63592 24212
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63960 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 93832 24212
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 94200 24172 99360 24212
rect 576 24148 99360 24172
rect 16867 24044 16925 24045
rect 16867 24004 16876 24044
rect 16916 24004 16925 24044
rect 16867 24003 16925 24004
rect 46347 24044 46389 24053
rect 46347 24004 46348 24044
rect 46388 24004 46389 24044
rect 46347 23995 46389 24004
rect 21475 23960 21533 23961
rect 21475 23920 21484 23960
rect 21524 23920 21533 23960
rect 21475 23919 21533 23920
rect 20331 23876 20373 23885
rect 20331 23836 20332 23876
rect 20372 23836 20373 23876
rect 20331 23827 20373 23836
rect 46147 23876 46205 23877
rect 46147 23836 46156 23876
rect 46196 23836 46205 23876
rect 46147 23835 46205 23836
rect 47691 23876 47733 23885
rect 47691 23836 47692 23876
rect 47732 23836 47733 23876
rect 47691 23827 47733 23836
rect 15427 23792 15485 23793
rect 15427 23752 15436 23792
rect 15476 23752 15485 23792
rect 15427 23751 15485 23752
rect 15811 23792 15869 23793
rect 15811 23752 15820 23792
rect 15860 23752 15869 23792
rect 15811 23751 15869 23752
rect 16195 23792 16253 23793
rect 16195 23752 16204 23792
rect 16244 23752 16253 23792
rect 16195 23751 16253 23752
rect 17059 23792 17117 23793
rect 17059 23752 17068 23792
rect 17108 23752 17117 23792
rect 17059 23751 17117 23752
rect 18307 23792 18365 23793
rect 18307 23752 18316 23792
rect 18356 23752 18365 23792
rect 18307 23751 18365 23752
rect 19171 23792 19229 23793
rect 19171 23752 19180 23792
rect 19220 23752 19229 23792
rect 19171 23751 19229 23752
rect 20803 23792 20861 23793
rect 20803 23752 20812 23792
rect 20852 23752 20861 23792
rect 20803 23751 20861 23752
rect 21955 23792 22013 23793
rect 21955 23752 21964 23792
rect 22004 23752 22013 23792
rect 21955 23751 22013 23752
rect 22059 23792 22101 23801
rect 22059 23752 22060 23792
rect 22100 23752 22101 23792
rect 22059 23743 22101 23752
rect 30219 23792 30261 23801
rect 30219 23752 30220 23792
rect 30260 23752 30261 23792
rect 30219 23743 30261 23752
rect 30595 23792 30653 23793
rect 30595 23752 30604 23792
rect 30644 23752 30653 23792
rect 30595 23751 30653 23752
rect 31459 23792 31517 23793
rect 31459 23752 31468 23792
rect 31508 23752 31517 23792
rect 31459 23751 31517 23752
rect 34827 23792 34869 23801
rect 34827 23752 34828 23792
rect 34868 23752 34869 23792
rect 34827 23743 34869 23752
rect 34923 23792 34965 23801
rect 34923 23752 34924 23792
rect 34964 23752 34965 23792
rect 34923 23743 34965 23752
rect 35011 23792 35069 23793
rect 35011 23752 35020 23792
rect 35060 23752 35069 23792
rect 35011 23751 35069 23752
rect 35203 23792 35261 23793
rect 35203 23752 35212 23792
rect 35252 23752 35261 23792
rect 35203 23751 35261 23752
rect 35491 23792 35549 23793
rect 35491 23752 35500 23792
rect 35540 23752 35549 23792
rect 35491 23751 35549 23752
rect 39907 23792 39965 23793
rect 39907 23752 39916 23792
rect 39956 23752 39965 23792
rect 39907 23751 39965 23752
rect 42019 23792 42077 23793
rect 42019 23752 42028 23792
rect 42068 23752 42077 23792
rect 42019 23751 42077 23752
rect 42883 23792 42941 23793
rect 42883 23752 42892 23792
rect 42932 23752 42941 23792
rect 42883 23751 42941 23752
rect 43459 23792 43517 23793
rect 43459 23752 43468 23792
rect 43508 23752 43517 23792
rect 43459 23751 43517 23752
rect 43843 23792 43901 23793
rect 43843 23752 43852 23792
rect 43892 23752 43901 23792
rect 43843 23751 43901 23752
rect 45475 23792 45533 23793
rect 45475 23752 45484 23792
rect 45524 23752 45533 23792
rect 45475 23751 45533 23752
rect 45579 23792 45621 23801
rect 45579 23752 45580 23792
rect 45620 23752 45621 23792
rect 45579 23743 45621 23752
rect 45675 23792 45717 23801
rect 45675 23752 45676 23792
rect 45716 23752 45717 23792
rect 45675 23743 45717 23752
rect 48355 23792 48413 23793
rect 48355 23752 48364 23792
rect 48404 23752 48413 23792
rect 48355 23751 48413 23752
rect 15907 23708 15965 23709
rect 15907 23668 15916 23708
rect 15956 23668 15965 23708
rect 15907 23667 15965 23668
rect 17739 23708 17781 23717
rect 17739 23668 17740 23708
rect 17780 23668 17781 23708
rect 17739 23659 17781 23668
rect 17931 23708 17973 23717
rect 17931 23668 17932 23708
rect 17972 23668 17973 23708
rect 17931 23659 17973 23668
rect 43275 23708 43317 23717
rect 43275 23668 43276 23708
rect 43316 23668 43317 23708
rect 43275 23659 43317 23668
rect 21675 23624 21717 23633
rect 21675 23584 21676 23624
rect 21716 23584 21717 23624
rect 21675 23575 21717 23584
rect 32611 23624 32669 23625
rect 32611 23584 32620 23624
rect 32660 23584 32669 23624
rect 32611 23583 32669 23584
rect 35691 23624 35733 23633
rect 35691 23584 35692 23624
rect 35732 23584 35733 23624
rect 35691 23575 35733 23584
rect 40579 23624 40637 23625
rect 40579 23584 40588 23624
rect 40628 23584 40637 23624
rect 40579 23583 40637 23584
rect 40867 23624 40925 23625
rect 40867 23584 40876 23624
rect 40916 23584 40925 23624
rect 40867 23583 40925 23584
rect 43947 23624 43989 23633
rect 43947 23584 43948 23624
rect 43988 23584 43989 23624
rect 43947 23575 43989 23584
rect 576 23456 99360 23480
rect 576 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 19472 23456
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19840 23416 34592 23456
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34960 23416 49712 23456
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 50080 23416 64832 23456
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 65200 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 95072 23456
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95440 23416 99360 23456
rect 576 23392 99360 23416
rect 34435 23288 34493 23289
rect 34435 23248 34444 23288
rect 34484 23248 34493 23288
rect 34435 23247 34493 23248
rect 39235 23288 39293 23289
rect 39235 23248 39244 23288
rect 39284 23248 39293 23288
rect 39235 23247 39293 23248
rect 20707 23204 20765 23205
rect 20707 23164 20716 23204
rect 20756 23164 20765 23204
rect 20707 23163 20765 23164
rect 36843 23204 36885 23213
rect 36843 23164 36844 23204
rect 36884 23164 36885 23204
rect 36843 23155 36885 23164
rect 40291 23204 40349 23205
rect 40291 23164 40300 23204
rect 40340 23164 40349 23204
rect 40291 23163 40349 23164
rect 2083 23120 2141 23121
rect 2083 23080 2092 23120
rect 2132 23080 2141 23120
rect 2083 23079 2141 23080
rect 6115 23120 6173 23121
rect 6115 23080 6124 23120
rect 6164 23080 6173 23120
rect 6115 23079 6173 23080
rect 20899 23120 20957 23121
rect 20899 23080 20908 23120
rect 20948 23080 20957 23120
rect 20899 23079 20957 23080
rect 21187 23120 21245 23121
rect 21187 23080 21196 23120
rect 21236 23080 21245 23120
rect 21187 23079 21245 23080
rect 28195 23120 28253 23121
rect 28195 23080 28204 23120
rect 28244 23080 28253 23120
rect 28195 23079 28253 23080
rect 33763 23120 33821 23121
rect 33763 23080 33772 23120
rect 33812 23080 33821 23120
rect 33763 23079 33821 23080
rect 37219 23120 37277 23121
rect 37219 23080 37228 23120
rect 37268 23080 37277 23120
rect 37219 23079 37277 23080
rect 38083 23120 38141 23121
rect 38083 23080 38092 23120
rect 38132 23080 38141 23120
rect 38083 23079 38141 23080
rect 40483 23120 40541 23121
rect 40483 23080 40492 23120
rect 40532 23080 40541 23120
rect 40483 23079 40541 23080
rect 40771 23120 40829 23121
rect 40771 23080 40780 23120
rect 40820 23080 40829 23120
rect 40771 23079 40829 23080
rect 2947 23036 3005 23037
rect 2947 22996 2956 23036
rect 2996 22996 3005 23036
rect 2947 22995 3005 22996
rect 4483 23036 4541 23037
rect 4483 22996 4492 23036
rect 4532 22996 4541 23036
rect 4483 22995 4541 22996
rect 2755 22868 2813 22869
rect 2755 22828 2764 22868
rect 2804 22828 2813 22868
rect 2755 22827 2813 22828
rect 3147 22868 3189 22877
rect 3147 22828 3148 22868
rect 3188 22828 3189 22868
rect 3147 22819 3189 22828
rect 4299 22868 4341 22877
rect 4299 22828 4300 22868
rect 4340 22828 4341 22868
rect 4299 22819 4341 22828
rect 5443 22868 5501 22869
rect 5443 22828 5452 22868
rect 5492 22828 5501 22868
rect 5443 22827 5501 22828
rect 27523 22868 27581 22869
rect 27523 22828 27532 22868
rect 27572 22828 27581 22868
rect 27523 22827 27581 22828
rect 34435 22868 34493 22869
rect 34435 22828 34444 22868
rect 34484 22828 34493 22868
rect 34435 22827 34493 22828
rect 576 22700 99360 22724
rect 576 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 18232 22700
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18600 22660 33352 22700
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33720 22660 48472 22700
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48840 22660 63592 22700
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63960 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 93832 22700
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 94200 22660 99360 22700
rect 576 22636 99360 22660
rect 1219 22532 1277 22533
rect 1219 22492 1228 22532
rect 1268 22492 1277 22532
rect 1219 22491 1277 22492
rect 6211 22532 6269 22533
rect 6211 22492 6220 22532
rect 6260 22492 6269 22532
rect 6211 22491 6269 22492
rect 16003 22532 16061 22533
rect 16003 22492 16012 22532
rect 16052 22492 16061 22532
rect 16003 22491 16061 22492
rect 28099 22532 28157 22533
rect 28099 22492 28108 22532
rect 28148 22492 28157 22532
rect 28099 22491 28157 22492
rect 49611 22532 49653 22541
rect 49611 22492 49612 22532
rect 49652 22492 49653 22532
rect 49611 22483 49653 22492
rect 651 22448 693 22457
rect 651 22408 652 22448
rect 692 22408 693 22448
rect 651 22399 693 22408
rect 34243 22448 34301 22449
rect 34243 22408 34252 22448
rect 34292 22408 34301 22448
rect 34243 22407 34301 22408
rect 33475 22364 33533 22365
rect 33475 22324 33484 22364
rect 33524 22324 33533 22364
rect 33475 22323 33533 22324
rect 2371 22280 2429 22281
rect 2371 22240 2380 22280
rect 2420 22240 2429 22280
rect 2371 22239 2429 22240
rect 3235 22280 3293 22281
rect 3235 22240 3244 22280
rect 3284 22240 3293 22280
rect 3235 22239 3293 22240
rect 3627 22280 3669 22289
rect 3627 22240 3628 22280
rect 3668 22240 3669 22280
rect 3627 22231 3669 22240
rect 3819 22280 3861 22289
rect 3819 22240 3820 22280
rect 3860 22240 3861 22280
rect 3819 22231 3861 22240
rect 4195 22280 4253 22281
rect 4195 22240 4204 22280
rect 4244 22240 4253 22280
rect 4195 22239 4253 22240
rect 5059 22280 5117 22281
rect 5059 22240 5068 22280
rect 5108 22240 5117 22280
rect 5059 22239 5117 22240
rect 9955 22280 10013 22281
rect 9955 22240 9964 22280
rect 10004 22240 10013 22280
rect 9955 22239 10013 22240
rect 13987 22280 14045 22281
rect 13987 22240 13996 22280
rect 14036 22240 14045 22280
rect 13987 22239 14045 22240
rect 14851 22280 14909 22281
rect 14851 22240 14860 22280
rect 14900 22240 14909 22280
rect 14851 22239 14909 22240
rect 21955 22280 22013 22281
rect 21955 22240 21964 22280
rect 22004 22240 22013 22280
rect 21955 22239 22013 22240
rect 26083 22280 26141 22281
rect 26083 22240 26092 22280
rect 26132 22240 26141 22280
rect 26083 22239 26141 22240
rect 26947 22280 27005 22281
rect 26947 22240 26956 22280
rect 26996 22240 27005 22280
rect 26947 22239 27005 22240
rect 34915 22280 34973 22281
rect 34915 22240 34924 22280
rect 34964 22240 34973 22280
rect 34915 22239 34973 22240
rect 35203 22280 35261 22281
rect 35203 22240 35212 22280
rect 35252 22240 35261 22280
rect 35203 22239 35261 22240
rect 41059 22280 41117 22281
rect 41059 22240 41068 22280
rect 41108 22240 41117 22280
rect 41059 22239 41117 22240
rect 44995 22280 45053 22281
rect 44995 22240 45004 22280
rect 45044 22240 45053 22280
rect 44995 22239 45053 22240
rect 49315 22280 49373 22281
rect 49315 22240 49324 22280
rect 49364 22240 49373 22280
rect 49315 22239 49373 22240
rect 50275 22280 50333 22281
rect 50275 22240 50284 22280
rect 50324 22240 50333 22280
rect 50275 22239 50333 22240
rect 13611 22196 13653 22205
rect 13611 22156 13612 22196
rect 13652 22156 13653 22196
rect 13611 22147 13653 22156
rect 25707 22196 25749 22205
rect 25707 22156 25708 22196
rect 25748 22156 25749 22196
rect 25707 22147 25749 22156
rect 9483 22112 9525 22121
rect 9483 22072 9484 22112
rect 9524 22072 9525 22112
rect 9483 22063 9525 22072
rect 21283 22112 21341 22113
rect 21283 22072 21292 22112
rect 21332 22072 21341 22112
rect 21283 22071 21341 22072
rect 33291 22112 33333 22121
rect 33291 22072 33292 22112
rect 33332 22072 33333 22112
rect 33291 22063 33333 22072
rect 35107 22112 35165 22113
rect 35107 22072 35116 22112
rect 35156 22072 35165 22112
rect 35107 22071 35165 22072
rect 35395 22112 35453 22113
rect 35395 22072 35404 22112
rect 35444 22072 35453 22112
rect 35395 22071 35453 22072
rect 40387 22112 40445 22113
rect 40387 22072 40396 22112
rect 40436 22072 40445 22112
rect 40387 22071 40445 22072
rect 44899 22112 44957 22113
rect 44899 22072 44908 22112
rect 44948 22072 44957 22112
rect 44899 22071 44957 22072
rect 45187 22112 45245 22113
rect 45187 22072 45196 22112
rect 45236 22072 45245 22112
rect 45187 22071 45245 22072
rect 576 21944 99360 21968
rect 576 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 19472 21944
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19840 21904 34592 21944
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34960 21904 49712 21944
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 50080 21904 64832 21944
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 65200 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 95072 21944
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95440 21904 99360 21944
rect 576 21880 99360 21904
rect 13699 21776 13757 21777
rect 13699 21736 13708 21776
rect 13748 21736 13757 21776
rect 13699 21735 13757 21736
rect 34819 21776 34877 21777
rect 34819 21736 34828 21776
rect 34868 21736 34877 21776
rect 34819 21735 34877 21736
rect 32427 21692 32469 21701
rect 32427 21652 32428 21692
rect 32468 21652 32469 21692
rect 32427 21643 32469 21652
rect 36267 21692 36309 21701
rect 36267 21652 36268 21692
rect 36308 21652 36309 21692
rect 36267 21643 36309 21652
rect 4491 21608 4533 21617
rect 4491 21568 4492 21608
rect 4532 21568 4533 21608
rect 4491 21559 4533 21568
rect 4675 21608 4733 21609
rect 4675 21568 4684 21608
rect 4724 21568 4733 21608
rect 4675 21567 4733 21568
rect 8043 21608 8085 21617
rect 8043 21568 8044 21608
rect 8084 21568 8085 21608
rect 8043 21559 8085 21568
rect 8419 21608 8477 21609
rect 8419 21568 8428 21608
rect 8468 21568 8477 21608
rect 8419 21567 8477 21568
rect 9283 21608 9341 21609
rect 9283 21568 9292 21608
rect 9332 21568 9341 21608
rect 9283 21567 9341 21568
rect 11011 21608 11069 21609
rect 11011 21568 11020 21608
rect 11060 21568 11069 21608
rect 11011 21567 11069 21568
rect 13027 21608 13085 21609
rect 13027 21568 13036 21608
rect 13076 21568 13085 21608
rect 13027 21567 13085 21568
rect 14755 21608 14813 21609
rect 14755 21568 14764 21608
rect 14804 21568 14813 21608
rect 14755 21567 14813 21568
rect 15715 21608 15773 21609
rect 15715 21568 15724 21608
rect 15764 21568 15773 21608
rect 15715 21567 15773 21568
rect 20995 21608 21053 21609
rect 20995 21568 21004 21608
rect 21044 21568 21053 21608
rect 20995 21567 21053 21568
rect 25803 21608 25845 21617
rect 25803 21568 25804 21608
rect 25844 21568 25845 21608
rect 25803 21559 25845 21568
rect 26179 21608 26237 21609
rect 26179 21568 26188 21608
rect 26228 21568 26237 21608
rect 26179 21567 26237 21568
rect 27043 21608 27101 21609
rect 27043 21568 27052 21608
rect 27092 21568 27101 21608
rect 27043 21567 27101 21568
rect 29059 21608 29117 21609
rect 29059 21568 29068 21608
rect 29108 21568 29117 21608
rect 29059 21567 29117 21568
rect 31171 21608 31229 21609
rect 31171 21568 31180 21608
rect 31220 21568 31229 21608
rect 31171 21567 31229 21568
rect 32131 21608 32189 21609
rect 32131 21568 32140 21608
rect 32180 21568 32189 21608
rect 32131 21567 32189 21568
rect 32803 21608 32861 21609
rect 32803 21568 32812 21608
rect 32852 21568 32861 21608
rect 32803 21567 32861 21568
rect 33667 21608 33725 21609
rect 33667 21568 33676 21608
rect 33716 21568 33725 21608
rect 33667 21567 33725 21568
rect 36643 21608 36701 21609
rect 36643 21568 36652 21608
rect 36692 21568 36701 21608
rect 36643 21567 36701 21568
rect 37507 21608 37565 21609
rect 37507 21568 37516 21608
rect 37556 21568 37565 21608
rect 37507 21567 37565 21568
rect 38947 21608 39005 21609
rect 38947 21568 38956 21608
rect 38996 21568 39005 21608
rect 38947 21567 39005 21568
rect 43075 21608 43133 21609
rect 43075 21568 43084 21608
rect 43124 21568 43133 21608
rect 43075 21567 43133 21568
rect 44035 21608 44093 21609
rect 44035 21568 44044 21608
rect 44084 21568 44093 21608
rect 44035 21567 44093 21568
rect 44427 21608 44469 21617
rect 44427 21568 44428 21608
rect 44468 21568 44469 21608
rect 44427 21559 44469 21568
rect 44803 21608 44861 21609
rect 44803 21568 44812 21608
rect 44852 21568 44861 21608
rect 44803 21567 44861 21568
rect 45667 21608 45725 21609
rect 45667 21568 45676 21608
rect 45716 21568 45725 21608
rect 45667 21567 45725 21568
rect 10443 21524 10485 21533
rect 10443 21484 10444 21524
rect 10484 21484 10485 21524
rect 10443 21475 10485 21484
rect 28203 21524 28245 21533
rect 28203 21484 28204 21524
rect 28244 21484 28245 21524
rect 28203 21475 28245 21484
rect 38667 21524 38709 21533
rect 38667 21484 38668 21524
rect 38708 21484 38709 21524
rect 38667 21475 38709 21484
rect 15243 21440 15285 21449
rect 15243 21400 15244 21440
rect 15284 21400 15285 21440
rect 15243 21391 15285 21400
rect 31467 21440 31509 21449
rect 31467 21400 31468 21440
rect 31508 21400 31509 21440
rect 31467 21391 31509 21400
rect 43755 21440 43797 21449
rect 43755 21400 43756 21440
rect 43796 21400 43797 21440
rect 43755 21391 43797 21400
rect 4587 21356 4629 21365
rect 4587 21316 4588 21356
rect 4628 21316 4629 21356
rect 4587 21307 4629 21316
rect 11683 21356 11741 21357
rect 11683 21316 11692 21356
rect 11732 21316 11741 21356
rect 11683 21315 11741 21316
rect 20323 21356 20381 21357
rect 20323 21316 20332 21356
rect 20372 21316 20381 21356
rect 20323 21315 20381 21316
rect 28387 21356 28445 21357
rect 28387 21316 28396 21356
rect 28436 21316 28445 21356
rect 28387 21315 28445 21316
rect 39619 21356 39677 21357
rect 39619 21316 39628 21356
rect 39668 21316 39677 21356
rect 39619 21315 39677 21316
rect 46819 21356 46877 21357
rect 46819 21316 46828 21356
rect 46868 21316 46877 21356
rect 46819 21315 46877 21316
rect 576 21188 99360 21212
rect 576 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 18232 21188
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18600 21148 33352 21188
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33720 21148 48472 21188
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48840 21148 63592 21188
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63960 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 93832 21188
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 94200 21148 99360 21188
rect 576 21124 99360 21148
rect 5827 21020 5885 21021
rect 5827 20980 5836 21020
rect 5876 20980 5885 21020
rect 5827 20979 5885 20980
rect 16003 21020 16061 21021
rect 16003 20980 16012 21020
rect 16052 20980 16061 21020
rect 16003 20979 16061 20980
rect 20043 21020 20085 21029
rect 20043 20980 20044 21020
rect 20084 20980 20085 21020
rect 20043 20971 20085 20980
rect 26475 21020 26517 21029
rect 26475 20980 26476 21020
rect 26516 20980 26517 21020
rect 26475 20971 26517 20980
rect 26859 21020 26901 21029
rect 26859 20980 26860 21020
rect 26900 20980 26901 21020
rect 26859 20971 26901 20980
rect 651 20936 693 20945
rect 651 20896 652 20936
rect 692 20896 693 20936
rect 651 20887 693 20896
rect 26659 20852 26717 20853
rect 26659 20812 26668 20852
rect 26708 20812 26717 20852
rect 26659 20811 26717 20812
rect 27043 20852 27101 20853
rect 27043 20812 27052 20852
rect 27092 20812 27101 20852
rect 27043 20811 27101 20812
rect 52675 20852 52733 20853
rect 52675 20812 52684 20852
rect 52724 20812 52733 20852
rect 52675 20811 52733 20812
rect 5635 20768 5693 20769
rect 5635 20728 5644 20768
rect 5684 20728 5693 20768
rect 5635 20727 5693 20728
rect 11403 20768 11445 20777
rect 11403 20728 11404 20768
rect 11444 20728 11445 20768
rect 11403 20719 11445 20728
rect 11587 20768 11645 20769
rect 11587 20728 11596 20768
rect 11636 20728 11645 20768
rect 11587 20727 11645 20728
rect 11779 20768 11837 20769
rect 11779 20728 11788 20768
rect 11828 20728 11837 20768
rect 11779 20727 11837 20728
rect 12163 20768 12221 20769
rect 12163 20728 12172 20768
rect 12212 20728 12221 20768
rect 12163 20727 12221 20728
rect 12739 20768 12797 20769
rect 12739 20728 12748 20768
rect 12788 20728 12797 20768
rect 12739 20727 12797 20728
rect 13987 20768 14045 20769
rect 13987 20728 13996 20768
rect 14036 20728 14045 20768
rect 13987 20727 14045 20728
rect 14851 20768 14909 20769
rect 14851 20728 14860 20768
rect 14900 20728 14909 20768
rect 14851 20727 14909 20728
rect 20515 20768 20573 20769
rect 20515 20728 20524 20768
rect 20564 20728 20573 20768
rect 20515 20727 20573 20728
rect 20995 20768 21053 20769
rect 20995 20728 21004 20768
rect 21044 20728 21053 20768
rect 20995 20727 21053 20728
rect 21955 20768 22013 20769
rect 21955 20728 21964 20768
rect 22004 20728 22013 20768
rect 21955 20727 22013 20728
rect 39723 20768 39765 20777
rect 39723 20728 39724 20768
rect 39764 20728 39765 20768
rect 39723 20719 39765 20728
rect 39819 20768 39861 20777
rect 39819 20728 39820 20768
rect 39860 20728 39861 20768
rect 39819 20719 39861 20728
rect 39907 20768 39965 20769
rect 39907 20728 39916 20768
rect 39956 20728 39965 20768
rect 39907 20727 39965 20728
rect 40387 20768 40445 20769
rect 40387 20728 40396 20768
rect 40436 20728 40445 20768
rect 40387 20727 40445 20728
rect 40483 20768 40541 20769
rect 40483 20728 40492 20768
rect 40532 20728 40541 20768
rect 40483 20727 40541 20728
rect 45571 20768 45629 20769
rect 45571 20728 45580 20768
rect 45620 20728 45629 20768
rect 45571 20727 45629 20728
rect 46435 20768 46493 20769
rect 46435 20728 46444 20768
rect 46484 20728 46493 20768
rect 46435 20727 46493 20728
rect 46827 20768 46869 20777
rect 46827 20728 46828 20768
rect 46868 20728 46869 20768
rect 46827 20719 46869 20728
rect 11499 20684 11541 20693
rect 11499 20644 11500 20684
rect 11540 20644 11541 20684
rect 11499 20635 11541 20644
rect 12259 20684 12317 20685
rect 12259 20644 12268 20684
rect 12308 20644 12317 20684
rect 12259 20643 12317 20644
rect 13419 20684 13461 20693
rect 13419 20644 13420 20684
rect 13460 20644 13461 20684
rect 13419 20635 13461 20644
rect 13611 20684 13653 20693
rect 13611 20644 13612 20684
rect 13652 20644 13653 20684
rect 13611 20635 13653 20644
rect 5539 20600 5597 20601
rect 5539 20560 5548 20600
rect 5588 20560 5597 20600
rect 5539 20559 5597 20560
rect 40683 20600 40725 20609
rect 40683 20560 40684 20600
rect 40724 20560 40725 20600
rect 40683 20551 40725 20560
rect 44419 20600 44477 20601
rect 44419 20560 44428 20600
rect 44468 20560 44477 20600
rect 44419 20559 44477 20560
rect 52491 20600 52533 20609
rect 52491 20560 52492 20600
rect 52532 20560 52533 20600
rect 52491 20551 52533 20560
rect 576 20432 99360 20456
rect 576 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 19472 20432
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19840 20392 34592 20432
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34960 20392 49712 20432
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 50080 20392 64832 20432
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 65200 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 95072 20432
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95440 20392 99360 20432
rect 576 20368 99360 20392
rect 5347 20180 5405 20181
rect 5347 20140 5356 20180
rect 5396 20140 5405 20180
rect 5347 20139 5405 20140
rect 28395 20180 28437 20189
rect 28395 20140 28396 20180
rect 28436 20140 28437 20180
rect 28395 20131 28437 20140
rect 32035 20180 32093 20181
rect 32035 20140 32044 20180
rect 32084 20140 32093 20180
rect 32035 20139 32093 20140
rect 39139 20180 39197 20181
rect 39139 20140 39148 20180
rect 39188 20140 39197 20180
rect 39139 20139 39197 20140
rect 46059 20180 46101 20189
rect 46059 20140 46060 20180
rect 46100 20140 46101 20180
rect 46059 20131 46101 20140
rect 52107 20180 52149 20189
rect 52107 20140 52108 20180
rect 52148 20140 52149 20180
rect 52107 20131 52149 20140
rect 4491 20096 4533 20105
rect 4491 20056 4492 20096
rect 4532 20056 4533 20096
rect 4491 20047 4533 20056
rect 4675 20096 4733 20097
rect 4675 20056 4684 20096
rect 4724 20056 4733 20096
rect 4675 20055 4733 20056
rect 4867 20096 4925 20097
rect 4867 20056 4876 20096
rect 4916 20056 4925 20096
rect 4867 20055 4925 20056
rect 5155 20096 5213 20097
rect 5155 20056 5164 20096
rect 5204 20056 5213 20096
rect 5155 20055 5213 20056
rect 12075 20096 12117 20105
rect 12075 20056 12076 20096
rect 12116 20056 12117 20096
rect 12075 20047 12117 20056
rect 12163 20096 12221 20097
rect 12163 20056 12172 20096
rect 12212 20056 12221 20096
rect 12163 20055 12221 20056
rect 20619 20096 20661 20105
rect 20619 20056 20620 20096
rect 20660 20056 20661 20096
rect 20619 20047 20661 20056
rect 21003 20096 21045 20105
rect 21003 20056 21004 20096
rect 21044 20056 21045 20096
rect 21003 20047 21045 20056
rect 21379 20096 21437 20097
rect 21379 20056 21388 20096
rect 21428 20056 21437 20096
rect 21379 20055 21437 20056
rect 22243 20096 22301 20097
rect 22243 20056 22252 20096
rect 22292 20056 22301 20096
rect 22243 20055 22301 20056
rect 27915 20096 27957 20105
rect 27915 20056 27916 20096
rect 27956 20056 27957 20096
rect 27915 20047 27957 20056
rect 28099 20096 28157 20097
rect 28099 20056 28108 20096
rect 28148 20056 28157 20096
rect 28099 20055 28157 20056
rect 28299 20096 28341 20105
rect 28299 20056 28300 20096
rect 28340 20056 28341 20096
rect 28299 20047 28341 20056
rect 28483 20096 28541 20097
rect 28483 20056 28492 20096
rect 28532 20056 28541 20096
rect 28483 20055 28541 20056
rect 31171 20096 31229 20097
rect 31171 20056 31180 20096
rect 31220 20056 31229 20096
rect 31171 20055 31229 20056
rect 32419 20096 32477 20097
rect 32419 20056 32428 20096
rect 32468 20056 32477 20096
rect 32419 20055 32477 20056
rect 38659 20096 38717 20097
rect 38659 20056 38668 20096
rect 38708 20056 38717 20096
rect 38659 20055 38717 20056
rect 38947 20096 39005 20097
rect 38947 20056 38956 20096
rect 38996 20056 39005 20096
rect 38947 20055 39005 20056
rect 40099 20096 40157 20097
rect 40099 20056 40108 20096
rect 40148 20056 40157 20096
rect 40099 20055 40157 20056
rect 40771 20096 40829 20097
rect 40771 20056 40780 20096
rect 40820 20056 40829 20096
rect 40771 20055 40829 20056
rect 46723 20096 46781 20097
rect 46723 20056 46732 20096
rect 46772 20056 46781 20096
rect 46723 20055 46781 20056
rect 52483 20096 52541 20097
rect 52483 20056 52492 20096
rect 52532 20056 52541 20096
rect 52483 20055 52541 20056
rect 53347 20096 53405 20097
rect 53347 20056 53356 20096
rect 53396 20056 53405 20096
rect 53347 20055 53405 20056
rect 57475 20096 57533 20097
rect 57475 20056 57484 20096
rect 57524 20056 57533 20096
rect 57475 20055 57533 20056
rect 4587 20012 4629 20021
rect 4587 19972 4588 20012
rect 4628 19972 4629 20012
rect 4587 19963 4629 19972
rect 12451 20012 12509 20013
rect 12451 19972 12460 20012
rect 12500 19972 12509 20012
rect 12451 19971 12509 19972
rect 44995 20012 45053 20013
rect 44995 19972 45004 20012
rect 45044 19972 45053 20012
rect 44995 19971 45053 19972
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 44811 19928 44853 19937
rect 44811 19888 44812 19928
rect 44852 19888 44853 19928
rect 44811 19879 44853 19888
rect 20427 19844 20469 19853
rect 20427 19804 20428 19844
rect 20468 19804 20469 19844
rect 20427 19795 20469 19804
rect 23403 19844 23445 19853
rect 23403 19804 23404 19844
rect 23444 19804 23445 19844
rect 23403 19795 23445 19804
rect 28011 19844 28053 19853
rect 28011 19804 28012 19844
rect 28052 19804 28053 19844
rect 28011 19795 28053 19804
rect 31659 19844 31701 19853
rect 31659 19804 31660 19844
rect 31700 19804 31701 19844
rect 31659 19795 31701 19804
rect 33099 19844 33141 19853
rect 33099 19804 33100 19844
rect 33140 19804 33141 19844
rect 33099 19795 33141 19804
rect 39427 19844 39485 19845
rect 39427 19804 39436 19844
rect 39476 19804 39485 19844
rect 39427 19803 39485 19804
rect 41443 19844 41501 19845
rect 41443 19804 41452 19844
rect 41492 19804 41501 19844
rect 41443 19803 41501 19804
rect 54499 19844 54557 19845
rect 54499 19804 54508 19844
rect 54548 19804 54557 19844
rect 54499 19803 54557 19804
rect 56803 19844 56861 19845
rect 56803 19804 56812 19844
rect 56852 19804 56861 19844
rect 56803 19803 56861 19804
rect 576 19676 99360 19700
rect 576 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 18232 19676
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18600 19636 33352 19676
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33720 19636 48472 19676
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48840 19636 63592 19676
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63960 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 93832 19676
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 94200 19636 99360 19676
rect 576 19612 99360 19636
rect 3723 19508 3765 19517
rect 3723 19468 3724 19508
rect 3764 19468 3765 19508
rect 3723 19459 3765 19468
rect 12163 19508 12221 19509
rect 12163 19468 12172 19508
rect 12212 19468 12221 19508
rect 12163 19467 12221 19468
rect 35403 19508 35445 19517
rect 35403 19468 35404 19508
rect 35444 19468 35445 19508
rect 35403 19459 35445 19468
rect 58051 19508 58109 19509
rect 58051 19468 58060 19508
rect 58100 19468 58109 19508
rect 58051 19467 58109 19468
rect 651 19424 693 19433
rect 651 19384 652 19424
rect 692 19384 693 19424
rect 651 19375 693 19384
rect 3139 19340 3197 19341
rect 3139 19300 3148 19340
rect 3188 19300 3197 19340
rect 3139 19299 3197 19300
rect 5259 19340 5301 19349
rect 5259 19300 5260 19340
rect 5300 19300 5301 19340
rect 5259 19291 5301 19300
rect 55267 19340 55325 19341
rect 55267 19300 55276 19340
rect 55316 19300 55325 19340
rect 55267 19299 55325 19300
rect 3427 19256 3485 19257
rect 3427 19216 3436 19256
rect 3476 19216 3485 19256
rect 3427 19215 3485 19216
rect 4387 19256 4445 19257
rect 4387 19216 4396 19256
rect 4436 19216 4445 19256
rect 4387 19215 4445 19216
rect 4579 19256 4637 19257
rect 4579 19216 4588 19256
rect 4628 19216 4637 19256
rect 4579 19215 4637 19216
rect 7371 19256 7413 19265
rect 7371 19216 7372 19256
rect 7412 19216 7413 19256
rect 7371 19207 7413 19216
rect 7747 19256 7805 19257
rect 7747 19216 7756 19256
rect 7796 19216 7805 19256
rect 7747 19215 7805 19216
rect 8611 19256 8669 19257
rect 8611 19216 8620 19256
rect 8660 19216 8669 19256
rect 8611 19215 8669 19216
rect 12835 19256 12893 19257
rect 12835 19216 12844 19256
rect 12884 19216 12893 19256
rect 12835 19215 12893 19216
rect 19947 19256 19989 19265
rect 19947 19216 19948 19256
rect 19988 19216 19989 19256
rect 19947 19207 19989 19216
rect 20323 19256 20381 19257
rect 20323 19216 20332 19256
rect 20372 19216 20381 19256
rect 20323 19215 20381 19216
rect 21187 19256 21245 19257
rect 21187 19216 21196 19256
rect 21236 19216 21245 19256
rect 21187 19215 21245 19216
rect 22435 19256 22493 19257
rect 22435 19216 22444 19256
rect 22484 19216 22493 19256
rect 22435 19215 22493 19216
rect 28867 19256 28925 19257
rect 28867 19216 28876 19256
rect 28916 19216 28925 19256
rect 28867 19215 28925 19216
rect 29155 19256 29213 19257
rect 29155 19216 29164 19256
rect 29204 19216 29213 19256
rect 29155 19215 29213 19216
rect 31459 19256 31517 19257
rect 31459 19216 31468 19256
rect 31508 19216 31517 19256
rect 31459 19215 31517 19216
rect 32323 19256 32381 19257
rect 32323 19216 32332 19256
rect 32372 19216 32381 19256
rect 32323 19215 32381 19216
rect 35019 19256 35061 19265
rect 35019 19216 35020 19256
rect 35060 19216 35061 19256
rect 35019 19207 35061 19216
rect 35875 19256 35933 19257
rect 35875 19216 35884 19256
rect 35924 19216 35933 19256
rect 35875 19215 35933 19216
rect 54211 19256 54269 19257
rect 54211 19216 54220 19256
rect 54260 19216 54269 19256
rect 54211 19215 54269 19216
rect 56035 19256 56093 19257
rect 56035 19216 56044 19256
rect 56084 19216 56093 19256
rect 56035 19215 56093 19216
rect 56899 19256 56957 19257
rect 56899 19216 56908 19256
rect 56948 19216 56957 19256
rect 56899 19215 56957 19216
rect 29347 19172 29405 19173
rect 29347 19132 29356 19172
rect 29396 19132 29405 19172
rect 29347 19131 29405 19132
rect 31083 19172 31125 19181
rect 31083 19132 31084 19172
rect 31124 19132 31125 19172
rect 31083 19123 31125 19132
rect 55659 19172 55701 19181
rect 55659 19132 55660 19172
rect 55700 19132 55701 19172
rect 55659 19123 55701 19132
rect 2955 19088 2997 19097
rect 2955 19048 2956 19088
rect 2996 19048 2997 19088
rect 2955 19039 2997 19048
rect 9763 19088 9821 19089
rect 9763 19048 9772 19088
rect 9812 19048 9821 19088
rect 9763 19047 9821 19048
rect 33475 19088 33533 19089
rect 33475 19048 33484 19088
rect 33524 19048 33533 19088
rect 33475 19047 33533 19048
rect 53539 19088 53597 19089
rect 53539 19048 53548 19088
rect 53588 19048 53597 19088
rect 53539 19047 53597 19048
rect 55467 19088 55509 19097
rect 55467 19048 55468 19088
rect 55508 19048 55509 19088
rect 55467 19039 55509 19048
rect 576 18920 99360 18944
rect 576 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 19472 18920
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19840 18880 34592 18920
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34960 18880 49712 18920
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 50080 18880 64832 18920
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 65200 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 95072 18920
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95440 18880 99360 18920
rect 576 18856 99360 18880
rect 4675 18752 4733 18753
rect 4675 18712 4684 18752
rect 4724 18712 4733 18752
rect 4675 18711 4733 18712
rect 11211 18752 11253 18761
rect 11211 18712 11212 18752
rect 11252 18712 11253 18752
rect 11211 18703 11253 18712
rect 2283 18668 2325 18677
rect 2283 18628 2284 18668
rect 2324 18628 2325 18668
rect 2283 18619 2325 18628
rect 39435 18668 39477 18677
rect 39435 18628 39436 18668
rect 39476 18628 39477 18668
rect 39435 18619 39477 18628
rect 43083 18668 43125 18677
rect 43083 18628 43084 18668
rect 43124 18628 43125 18668
rect 43083 18619 43125 18628
rect 2659 18584 2717 18585
rect 2659 18544 2668 18584
rect 2708 18544 2717 18584
rect 2659 18543 2717 18544
rect 3523 18584 3581 18585
rect 3523 18544 3532 18584
rect 3572 18544 3581 18584
rect 3523 18543 3581 18544
rect 10723 18584 10781 18585
rect 10723 18544 10732 18584
rect 10772 18544 10781 18584
rect 10723 18543 10781 18544
rect 11011 18584 11069 18585
rect 11011 18544 11020 18584
rect 11060 18544 11069 18584
rect 11011 18543 11069 18544
rect 28291 18584 28349 18585
rect 28291 18544 28300 18584
rect 28340 18544 28349 18584
rect 28291 18543 28349 18544
rect 34051 18584 34109 18585
rect 34051 18544 34060 18584
rect 34100 18544 34109 18584
rect 34051 18543 34109 18544
rect 38179 18584 38237 18585
rect 38179 18544 38188 18584
rect 38228 18544 38237 18584
rect 38179 18543 38237 18544
rect 39043 18584 39101 18585
rect 39043 18544 39052 18584
rect 39092 18544 39101 18584
rect 39043 18543 39101 18544
rect 41827 18584 41885 18585
rect 41827 18544 41836 18584
rect 41876 18544 41885 18584
rect 41827 18543 41885 18544
rect 42691 18584 42749 18585
rect 42691 18544 42700 18584
rect 42740 18544 42749 18584
rect 42691 18543 42749 18544
rect 48747 18584 48789 18593
rect 48747 18544 48748 18584
rect 48788 18544 48789 18584
rect 48747 18535 48789 18544
rect 49123 18584 49181 18585
rect 49123 18544 49132 18584
rect 49172 18544 49181 18584
rect 49123 18543 49181 18544
rect 49987 18584 50045 18585
rect 49987 18544 49996 18584
rect 50036 18544 50045 18584
rect 49987 18543 50045 18544
rect 51331 18584 51389 18585
rect 51331 18544 51340 18584
rect 51380 18544 51389 18584
rect 51331 18543 51389 18544
rect 55179 18584 55221 18593
rect 55179 18544 55180 18584
rect 55220 18544 55221 18584
rect 55179 18535 55221 18544
rect 55363 18584 55421 18585
rect 55363 18544 55372 18584
rect 55412 18544 55421 18584
rect 55363 18543 55421 18544
rect 26851 18500 26909 18501
rect 26851 18460 26860 18500
rect 26900 18460 26909 18500
rect 26851 18459 26909 18460
rect 27235 18500 27293 18501
rect 27235 18460 27244 18500
rect 27284 18460 27293 18500
rect 27235 18459 27293 18460
rect 51147 18500 51189 18509
rect 51147 18460 51148 18500
rect 51188 18460 51189 18500
rect 51147 18451 51189 18460
rect 651 18416 693 18425
rect 651 18376 652 18416
rect 692 18376 693 18416
rect 651 18367 693 18376
rect 26667 18332 26709 18341
rect 26667 18292 26668 18332
rect 26708 18292 26709 18332
rect 26667 18283 26709 18292
rect 27051 18332 27093 18341
rect 27051 18292 27052 18332
rect 27092 18292 27093 18332
rect 27051 18283 27093 18292
rect 27619 18332 27677 18333
rect 27619 18292 27628 18332
rect 27668 18292 27677 18332
rect 27619 18291 27677 18292
rect 33379 18332 33437 18333
rect 33379 18292 33388 18332
rect 33428 18292 33437 18332
rect 33379 18291 33437 18292
rect 37027 18332 37085 18333
rect 37027 18292 37036 18332
rect 37076 18292 37085 18332
rect 37027 18291 37085 18292
rect 40675 18332 40733 18333
rect 40675 18292 40684 18332
rect 40724 18292 40733 18332
rect 40675 18291 40733 18292
rect 52003 18332 52061 18333
rect 52003 18292 52012 18332
rect 52052 18292 52061 18332
rect 52003 18291 52061 18292
rect 55275 18332 55317 18341
rect 55275 18292 55276 18332
rect 55316 18292 55317 18332
rect 55275 18283 55317 18292
rect 576 18164 99360 18188
rect 576 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 18232 18164
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18600 18124 33352 18164
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33720 18124 48472 18164
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48840 18124 63592 18164
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63960 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 93832 18164
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 94200 18124 99360 18164
rect 576 18100 99360 18124
rect 11011 17996 11069 17997
rect 11011 17956 11020 17996
rect 11060 17956 11069 17996
rect 11011 17955 11069 17956
rect 28099 17996 28157 17997
rect 28099 17956 28108 17996
rect 28148 17956 28157 17996
rect 28099 17955 28157 17956
rect 28963 17996 29021 17997
rect 28963 17956 28972 17996
rect 29012 17956 29021 17996
rect 28963 17955 29021 17956
rect 49323 17996 49365 18005
rect 49323 17956 49324 17996
rect 49364 17956 49365 17996
rect 49323 17947 49365 17956
rect 651 17912 693 17921
rect 651 17872 652 17912
rect 692 17872 693 17912
rect 651 17863 693 17872
rect 15819 17912 15861 17921
rect 15819 17872 15820 17912
rect 15860 17872 15861 17912
rect 15819 17863 15861 17872
rect 48843 17912 48885 17921
rect 48843 17872 48844 17912
rect 48884 17872 48885 17912
rect 48843 17863 48885 17872
rect 16003 17828 16061 17829
rect 16003 17788 16012 17828
rect 16052 17788 16061 17828
rect 16003 17787 16061 17788
rect 49027 17828 49085 17829
rect 49027 17788 49036 17828
rect 49076 17788 49085 17828
rect 49027 17787 49085 17788
rect 49507 17828 49565 17829
rect 49507 17788 49516 17828
rect 49556 17788 49565 17828
rect 49507 17787 49565 17788
rect 2563 17744 2621 17745
rect 2563 17704 2572 17744
rect 2612 17704 2621 17744
rect 2563 17703 2621 17704
rect 3427 17744 3485 17745
rect 3427 17704 3436 17744
rect 3476 17704 3485 17744
rect 3427 17703 3485 17704
rect 8995 17744 9053 17745
rect 8995 17704 9004 17744
rect 9044 17704 9053 17744
rect 8995 17703 9053 17704
rect 9859 17744 9917 17745
rect 9859 17704 9868 17744
rect 9908 17704 9917 17744
rect 9859 17703 9917 17704
rect 17443 17744 17501 17745
rect 17443 17704 17452 17744
rect 17492 17704 17501 17744
rect 17443 17703 17501 17704
rect 25707 17744 25749 17753
rect 25707 17704 25708 17744
rect 25748 17704 25749 17744
rect 25707 17695 25749 17704
rect 26083 17744 26141 17745
rect 26083 17704 26092 17744
rect 26132 17704 26141 17744
rect 26083 17703 26141 17704
rect 26947 17744 27005 17745
rect 26947 17704 26956 17744
rect 26996 17704 27005 17744
rect 26947 17703 27005 17704
rect 28291 17744 28349 17745
rect 28291 17704 28300 17744
rect 28340 17704 28349 17744
rect 28291 17703 28349 17704
rect 29251 17744 29309 17745
rect 29251 17704 29260 17744
rect 29300 17704 29309 17744
rect 29251 17703 29309 17704
rect 37891 17744 37949 17745
rect 37891 17704 37900 17744
rect 37940 17704 37949 17744
rect 37891 17703 37949 17704
rect 42691 17744 42749 17745
rect 42691 17704 42700 17744
rect 42740 17704 42749 17744
rect 42691 17703 42749 17704
rect 43563 17744 43605 17753
rect 43563 17704 43564 17744
rect 43604 17704 43605 17744
rect 43563 17695 43605 17704
rect 49707 17744 49749 17753
rect 49707 17704 49708 17744
rect 49748 17704 49749 17744
rect 51147 17744 51189 17753
rect 49707 17695 49749 17704
rect 50371 17711 50429 17712
rect 50371 17671 50380 17711
rect 50420 17671 50429 17711
rect 51147 17704 51148 17744
rect 51188 17704 51189 17744
rect 51147 17695 51189 17704
rect 51331 17744 51389 17745
rect 51331 17704 51340 17744
rect 51380 17704 51389 17744
rect 51331 17703 51389 17704
rect 52387 17744 52445 17745
rect 52387 17704 52396 17744
rect 52436 17704 52445 17744
rect 52387 17703 52445 17704
rect 55171 17744 55229 17745
rect 55171 17704 55180 17744
rect 55220 17704 55229 17744
rect 55171 17703 55229 17704
rect 55459 17744 55517 17745
rect 55459 17704 55468 17744
rect 55508 17704 55517 17744
rect 55459 17703 55517 17704
rect 50371 17670 50429 17671
rect 2187 17660 2229 17669
rect 2187 17620 2188 17660
rect 2228 17620 2229 17660
rect 2187 17611 2229 17620
rect 8619 17660 8661 17669
rect 8619 17620 8620 17660
rect 8660 17620 8661 17660
rect 8619 17611 8661 17620
rect 16779 17660 16821 17669
rect 16779 17620 16780 17660
rect 16820 17620 16821 17660
rect 16779 17611 16821 17620
rect 51243 17660 51285 17669
rect 51243 17620 51244 17660
rect 51284 17620 51285 17660
rect 51243 17611 51285 17620
rect 4579 17576 4637 17577
rect 4579 17536 4588 17576
rect 4628 17536 4637 17576
rect 4579 17535 4637 17536
rect 29155 17576 29213 17577
rect 29155 17536 29164 17576
rect 29204 17536 29213 17576
rect 29155 17535 29213 17536
rect 29443 17576 29501 17577
rect 29443 17536 29452 17576
rect 29492 17536 29501 17576
rect 29443 17535 29501 17536
rect 38563 17576 38621 17577
rect 38563 17536 38572 17576
rect 38612 17536 38621 17576
rect 38563 17535 38621 17536
rect 52291 17576 52349 17577
rect 52291 17536 52300 17576
rect 52340 17536 52349 17576
rect 52291 17535 52349 17536
rect 52579 17576 52637 17577
rect 52579 17536 52588 17576
rect 52628 17536 52637 17576
rect 52579 17535 52637 17536
rect 55659 17576 55701 17585
rect 55659 17536 55660 17576
rect 55700 17536 55701 17576
rect 55659 17527 55701 17536
rect 576 17408 99360 17432
rect 576 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 19472 17408
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19840 17368 34592 17408
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34960 17368 49712 17408
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 50080 17368 64832 17408
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 65200 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 95072 17408
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95440 17368 99360 17408
rect 576 17344 99360 17368
rect 3051 17240 3093 17249
rect 3051 17200 3052 17240
rect 3092 17200 3093 17240
rect 3051 17191 3093 17200
rect 4003 17240 4061 17241
rect 4003 17200 4012 17240
rect 4052 17200 4061 17240
rect 4003 17199 4061 17200
rect 11971 17240 12029 17241
rect 11971 17200 11980 17240
rect 12020 17200 12029 17240
rect 11971 17199 12029 17200
rect 17251 17240 17309 17241
rect 17251 17200 17260 17240
rect 17300 17200 17309 17240
rect 17251 17199 17309 17200
rect 28579 17240 28637 17241
rect 28579 17200 28588 17240
rect 28628 17200 28637 17240
rect 28579 17199 28637 17200
rect 50179 17240 50237 17241
rect 50179 17200 50188 17240
rect 50228 17200 50237 17240
rect 50179 17199 50237 17200
rect 14859 17156 14901 17165
rect 14859 17116 14860 17156
rect 14900 17116 14901 17156
rect 14859 17107 14901 17116
rect 21283 17156 21341 17157
rect 21283 17116 21292 17156
rect 21332 17116 21341 17156
rect 21283 17115 21341 17116
rect 26187 17156 26229 17165
rect 26187 17116 26188 17156
rect 26228 17116 26229 17156
rect 26187 17107 26229 17116
rect 33187 17156 33245 17157
rect 33187 17116 33196 17156
rect 33236 17116 33245 17156
rect 33187 17115 33245 17116
rect 40867 17156 40925 17157
rect 40867 17116 40876 17156
rect 40916 17116 40925 17156
rect 40867 17115 40925 17116
rect 47787 17156 47829 17165
rect 47787 17116 47788 17156
rect 47828 17116 47829 17156
rect 47787 17107 47829 17116
rect 52779 17156 52821 17165
rect 52779 17116 52780 17156
rect 52820 17116 52821 17156
rect 52779 17107 52821 17116
rect 56619 17156 56661 17165
rect 56619 17116 56620 17156
rect 56660 17116 56661 17156
rect 56619 17107 56661 17116
rect 4675 17072 4733 17073
rect 4675 17032 4684 17072
rect 4724 17032 4733 17072
rect 4675 17031 4733 17032
rect 9579 17072 9621 17081
rect 9579 17032 9580 17072
rect 9620 17032 9621 17072
rect 9579 17023 9621 17032
rect 9955 17072 10013 17073
rect 9955 17032 9964 17072
rect 10004 17032 10013 17072
rect 9955 17031 10013 17032
rect 10819 17072 10877 17073
rect 10819 17032 10828 17072
rect 10868 17032 10877 17072
rect 10819 17031 10877 17032
rect 15235 17072 15293 17073
rect 15235 17032 15244 17072
rect 15284 17032 15293 17072
rect 15235 17031 15293 17032
rect 16099 17072 16157 17073
rect 16099 17032 16108 17072
rect 16148 17032 16157 17072
rect 16099 17031 16157 17032
rect 20131 17072 20189 17073
rect 20131 17032 20140 17072
rect 20180 17032 20189 17072
rect 20131 17031 20189 17032
rect 20419 17072 20477 17073
rect 20419 17032 20428 17072
rect 20468 17032 20477 17072
rect 20419 17031 20477 17032
rect 23395 17072 23453 17073
rect 23395 17032 23404 17072
rect 23444 17032 23453 17072
rect 23395 17031 23453 17032
rect 26563 17072 26621 17073
rect 26563 17032 26572 17072
rect 26612 17032 26621 17072
rect 26563 17031 26621 17032
rect 27427 17072 27485 17073
rect 27427 17032 27436 17072
rect 27476 17032 27485 17072
rect 27427 17031 27485 17032
rect 32707 17072 32765 17073
rect 32707 17032 32716 17072
rect 32756 17032 32765 17072
rect 32707 17031 32765 17032
rect 33091 17072 33149 17073
rect 33091 17032 33100 17072
rect 33140 17032 33149 17072
rect 33091 17031 33149 17032
rect 33763 17072 33821 17073
rect 33763 17032 33772 17072
rect 33812 17032 33821 17072
rect 33763 17031 33821 17032
rect 35395 17072 35453 17073
rect 35395 17032 35404 17072
rect 35444 17032 35453 17072
rect 35395 17031 35453 17032
rect 36075 17072 36117 17081
rect 36075 17032 36076 17072
rect 36116 17032 36117 17072
rect 36075 17023 36117 17032
rect 36267 17072 36309 17081
rect 36267 17032 36268 17072
rect 36308 17032 36309 17072
rect 36267 17023 36309 17032
rect 36643 17072 36701 17073
rect 36643 17032 36652 17072
rect 36692 17032 36701 17072
rect 36643 17031 36701 17032
rect 37507 17072 37565 17073
rect 37507 17032 37516 17072
rect 37556 17032 37565 17072
rect 37507 17031 37565 17032
rect 40387 17072 40445 17073
rect 40387 17032 40396 17072
rect 40436 17032 40445 17072
rect 40387 17031 40445 17032
rect 40675 17072 40733 17073
rect 40675 17032 40684 17072
rect 40724 17032 40733 17072
rect 40675 17031 40733 17032
rect 45091 17072 45149 17073
rect 45091 17032 45100 17072
rect 45140 17032 45149 17072
rect 45091 17031 45149 17032
rect 46051 17072 46109 17073
rect 46051 17032 46060 17072
rect 46100 17032 46109 17072
rect 46051 17031 46109 17032
rect 48163 17072 48221 17073
rect 48163 17032 48172 17072
rect 48212 17032 48221 17072
rect 48163 17031 48221 17032
rect 49027 17072 49085 17073
rect 49027 17032 49036 17072
rect 49076 17032 49085 17072
rect 49027 17031 49085 17032
rect 53155 17072 53213 17073
rect 53155 17032 53164 17072
rect 53204 17032 53213 17072
rect 53155 17031 53213 17032
rect 54019 17072 54077 17073
rect 54019 17032 54028 17072
rect 54068 17032 54077 17072
rect 54019 17031 54077 17032
rect 56995 17072 57053 17073
rect 56995 17032 57004 17072
rect 57044 17032 57053 17072
rect 56995 17031 57053 17032
rect 57859 17072 57917 17073
rect 57859 17032 57868 17072
rect 57908 17032 57917 17072
rect 57859 17031 57917 17032
rect 3235 16988 3293 16989
rect 3235 16948 3244 16988
rect 3284 16948 3293 16988
rect 3235 16947 3293 16948
rect 38667 16988 38709 16997
rect 38667 16948 38668 16988
rect 38708 16948 38709 16988
rect 38667 16939 38709 16948
rect 651 16904 693 16913
rect 651 16864 652 16904
rect 692 16864 693 16904
rect 651 16855 693 16864
rect 19459 16820 19517 16821
rect 19459 16780 19468 16820
rect 19508 16780 19517 16820
rect 19459 16779 19517 16780
rect 20715 16820 20757 16829
rect 20715 16780 20716 16820
rect 20756 16780 20757 16820
rect 20715 16771 20757 16780
rect 24067 16820 24125 16821
rect 24067 16780 24076 16820
rect 24116 16780 24125 16820
rect 24067 16779 24125 16780
rect 34435 16820 34493 16821
rect 34435 16780 34444 16820
rect 34484 16780 34493 16820
rect 34435 16779 34493 16780
rect 55171 16820 55229 16821
rect 55171 16780 55180 16820
rect 55220 16780 55229 16820
rect 55171 16779 55229 16780
rect 59011 16820 59069 16821
rect 59011 16780 59020 16820
rect 59060 16780 59069 16820
rect 59011 16779 59069 16780
rect 576 16652 99360 16676
rect 576 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 18232 16652
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18600 16612 33352 16652
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33720 16612 48472 16652
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48840 16612 63592 16652
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63960 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 93832 16652
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 94200 16612 99360 16652
rect 576 16588 99360 16612
rect 10731 16484 10773 16493
rect 10731 16444 10732 16484
rect 10772 16444 10773 16484
rect 10731 16435 10773 16444
rect 651 16400 693 16409
rect 651 16360 652 16400
rect 692 16360 693 16400
rect 651 16351 693 16360
rect 21283 16400 21341 16401
rect 21283 16360 21292 16400
rect 21332 16360 21341 16400
rect 21283 16359 21341 16360
rect 46539 16400 46581 16409
rect 46539 16360 46540 16400
rect 46580 16360 46581 16400
rect 46539 16351 46581 16360
rect 16971 16316 17013 16325
rect 16971 16276 16972 16316
rect 17012 16276 17013 16316
rect 16971 16267 17013 16276
rect 18499 16316 18557 16317
rect 18499 16276 18508 16316
rect 18548 16276 18557 16316
rect 18499 16275 18557 16276
rect 34339 16316 34397 16317
rect 34339 16276 34348 16316
rect 34388 16276 34397 16316
rect 34339 16275 34397 16276
rect 10243 16232 10301 16233
rect 10243 16192 10252 16232
rect 10292 16192 10301 16232
rect 10243 16191 10301 16192
rect 14947 16232 15005 16233
rect 14947 16192 14956 16232
rect 14996 16192 15005 16232
rect 14947 16191 15005 16192
rect 15811 16232 15869 16233
rect 15811 16192 15820 16232
rect 15860 16192 15869 16232
rect 15811 16191 15869 16192
rect 17155 16232 17213 16233
rect 17155 16192 17164 16232
rect 17204 16192 17213 16232
rect 17155 16191 17213 16192
rect 19267 16232 19325 16233
rect 19267 16192 19276 16232
rect 19316 16192 19325 16232
rect 19267 16191 19325 16192
rect 20131 16232 20189 16233
rect 20131 16192 20140 16232
rect 20180 16192 20189 16232
rect 20131 16191 20189 16192
rect 31083 16232 31125 16241
rect 31083 16192 31084 16232
rect 31124 16192 31125 16232
rect 31083 16183 31125 16192
rect 31459 16232 31517 16233
rect 31459 16192 31468 16232
rect 31508 16192 31517 16232
rect 31459 16191 31517 16192
rect 32323 16232 32381 16233
rect 32323 16192 32332 16232
rect 32372 16192 32381 16232
rect 32323 16191 32381 16192
rect 34051 16232 34109 16233
rect 34051 16192 34060 16232
rect 34100 16192 34109 16232
rect 34051 16191 34109 16192
rect 34147 16232 34205 16233
rect 34147 16192 34156 16232
rect 34196 16192 34205 16232
rect 34147 16191 34205 16192
rect 41443 16232 41501 16233
rect 41443 16192 41452 16232
rect 41492 16192 41501 16232
rect 41443 16191 41501 16192
rect 45963 16232 46005 16241
rect 45963 16192 45964 16232
rect 46004 16192 46005 16232
rect 45963 16183 46005 16192
rect 56035 16232 56093 16233
rect 56035 16192 56044 16232
rect 56084 16192 56093 16232
rect 56035 16191 56093 16192
rect 14571 16148 14613 16157
rect 14571 16108 14572 16148
rect 14612 16108 14613 16148
rect 14571 16099 14613 16108
rect 18891 16148 18933 16157
rect 18891 16108 18892 16148
rect 18932 16108 18933 16148
rect 18891 16099 18933 16108
rect 10731 16064 10773 16073
rect 10731 16024 10732 16064
rect 10772 16024 10773 16064
rect 10731 16015 10773 16024
rect 17827 16064 17885 16065
rect 17827 16024 17836 16064
rect 17876 16024 17885 16064
rect 17827 16023 17885 16024
rect 18699 16064 18741 16073
rect 18699 16024 18700 16064
rect 18740 16024 18741 16064
rect 18699 16015 18741 16024
rect 33475 16064 33533 16065
rect 33475 16024 33484 16064
rect 33524 16024 33533 16064
rect 33475 16023 33533 16024
rect 42115 16064 42173 16065
rect 42115 16024 42124 16064
rect 42164 16024 42173 16064
rect 42115 16023 42173 16024
rect 46347 16064 46389 16073
rect 46347 16024 46348 16064
rect 46388 16024 46389 16064
rect 46347 16015 46389 16024
rect 55363 16064 55421 16065
rect 55363 16024 55372 16064
rect 55412 16024 55421 16064
rect 55363 16023 55421 16024
rect 576 15896 99360 15920
rect 576 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 19472 15896
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19840 15856 34592 15896
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34960 15856 49712 15896
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 50080 15856 64832 15896
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 65200 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 95072 15896
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95440 15856 99360 15896
rect 576 15832 99360 15856
rect 643 15728 701 15729
rect 643 15688 652 15728
rect 692 15688 701 15728
rect 643 15687 701 15688
rect 15627 15728 15669 15737
rect 15627 15688 15628 15728
rect 15668 15688 15669 15728
rect 15627 15679 15669 15688
rect 19939 15728 19997 15729
rect 19939 15688 19948 15728
rect 19988 15688 19997 15728
rect 19939 15687 19997 15688
rect 27715 15728 27773 15729
rect 27715 15688 27724 15728
rect 27764 15688 27773 15728
rect 27715 15687 27773 15688
rect 39331 15728 39389 15729
rect 39331 15688 39340 15728
rect 39380 15688 39389 15728
rect 39331 15687 39389 15688
rect 40971 15728 41013 15737
rect 40971 15688 40972 15728
rect 41012 15688 41013 15728
rect 40971 15679 41013 15688
rect 18691 15644 18749 15645
rect 18691 15604 18700 15644
rect 18740 15604 18749 15644
rect 18691 15603 18749 15604
rect 25323 15644 25365 15653
rect 25323 15604 25324 15644
rect 25364 15604 25365 15644
rect 25323 15595 25365 15604
rect 41739 15644 41781 15653
rect 41739 15604 41740 15644
rect 41780 15604 41781 15644
rect 41739 15595 41781 15604
rect 16003 15560 16061 15561
rect 16003 15520 16012 15560
rect 16052 15520 16061 15560
rect 16003 15519 16061 15520
rect 16963 15560 17021 15561
rect 16963 15520 16972 15560
rect 17012 15520 17021 15560
rect 16963 15519 17021 15520
rect 17451 15560 17493 15569
rect 17451 15520 17452 15560
rect 17492 15520 17493 15560
rect 17451 15511 17493 15520
rect 17635 15560 17693 15561
rect 17635 15520 17644 15560
rect 17684 15520 17693 15560
rect 17635 15519 17693 15520
rect 17827 15560 17885 15561
rect 17827 15520 17836 15560
rect 17876 15520 17885 15560
rect 17827 15519 17885 15520
rect 18027 15560 18069 15569
rect 18027 15520 18028 15560
rect 18068 15520 18069 15560
rect 18027 15511 18069 15520
rect 18211 15560 18269 15561
rect 18211 15520 18220 15560
rect 18260 15520 18269 15560
rect 18211 15519 18269 15520
rect 18499 15560 18557 15561
rect 18499 15520 18508 15560
rect 18548 15520 18557 15560
rect 18499 15519 18557 15520
rect 20035 15560 20093 15561
rect 20035 15520 20044 15560
rect 20084 15520 20093 15560
rect 20035 15519 20093 15520
rect 20419 15560 20477 15561
rect 20419 15520 20428 15560
rect 20468 15520 20477 15560
rect 20419 15519 20477 15520
rect 22915 15560 22973 15561
rect 22915 15520 22924 15560
rect 22964 15520 22973 15560
rect 22915 15519 22973 15520
rect 25699 15560 25757 15561
rect 25699 15520 25708 15560
rect 25748 15520 25757 15560
rect 25699 15519 25757 15520
rect 26563 15560 26621 15561
rect 26563 15520 26572 15560
rect 26612 15520 26621 15560
rect 26563 15519 26621 15520
rect 33475 15560 33533 15561
rect 33475 15520 33484 15560
rect 33524 15520 33533 15560
rect 33475 15519 33533 15520
rect 33579 15560 33621 15569
rect 33579 15520 33580 15560
rect 33620 15520 33621 15560
rect 33579 15511 33621 15520
rect 33675 15560 33717 15569
rect 33675 15520 33676 15560
rect 33716 15520 33717 15560
rect 33675 15511 33717 15520
rect 33859 15560 33917 15561
rect 33859 15520 33868 15560
rect 33908 15520 33917 15560
rect 33859 15519 33917 15520
rect 38659 15560 38717 15561
rect 38659 15520 38668 15560
rect 38708 15520 38717 15560
rect 38659 15519 38717 15520
rect 39531 15560 39573 15569
rect 39531 15520 39532 15560
rect 39572 15520 39573 15560
rect 39531 15511 39573 15520
rect 39627 15560 39669 15569
rect 39627 15520 39628 15560
rect 39668 15520 39669 15560
rect 39627 15511 39669 15520
rect 39715 15560 39773 15561
rect 39715 15520 39724 15560
rect 39764 15520 39773 15560
rect 39715 15519 39773 15520
rect 40675 15560 40733 15561
rect 40675 15520 40684 15560
rect 40724 15520 40733 15560
rect 40675 15519 40733 15520
rect 40771 15560 40829 15561
rect 40771 15520 40780 15560
rect 40820 15520 40829 15560
rect 40771 15519 40829 15520
rect 42115 15560 42173 15561
rect 42115 15520 42124 15560
rect 42164 15520 42173 15560
rect 42115 15519 42173 15520
rect 42979 15560 43037 15561
rect 42979 15520 42988 15560
rect 43028 15520 43037 15560
rect 42979 15519 43037 15520
rect 15811 15476 15869 15477
rect 15811 15436 15820 15476
rect 15860 15436 15869 15476
rect 15811 15435 15869 15436
rect 34539 15476 34581 15485
rect 34539 15436 34540 15476
rect 34580 15436 34581 15476
rect 34539 15427 34581 15436
rect 17547 15392 17589 15401
rect 17547 15352 17548 15392
rect 17588 15352 17589 15392
rect 17547 15343 17589 15352
rect 17931 15392 17973 15401
rect 17931 15352 17932 15392
rect 17972 15352 17973 15392
rect 17931 15343 17973 15352
rect 16491 15308 16533 15317
rect 16491 15268 16492 15308
rect 16532 15268 16533 15308
rect 16491 15259 16533 15268
rect 20227 15308 20285 15309
rect 20227 15268 20236 15308
rect 20276 15268 20285 15308
rect 20227 15267 20285 15268
rect 22243 15308 22301 15309
rect 22243 15268 22252 15308
rect 22292 15268 22301 15308
rect 22243 15267 22301 15268
rect 44131 15308 44189 15309
rect 44131 15268 44140 15308
rect 44180 15268 44189 15308
rect 44131 15267 44189 15268
rect 576 15140 99360 15164
rect 576 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 18232 15140
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18600 15100 33352 15140
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33720 15100 48472 15140
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48840 15100 63592 15140
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63960 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 93832 15140
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 94200 15100 99360 15140
rect 576 15076 99360 15100
rect 9091 14972 9149 14973
rect 9091 14932 9100 14972
rect 9140 14932 9149 14972
rect 9091 14931 9149 14932
rect 51531 14888 51573 14897
rect 51531 14848 51532 14888
rect 51572 14848 51573 14888
rect 51531 14839 51573 14848
rect 55467 14888 55509 14897
rect 55467 14848 55468 14888
rect 55508 14848 55509 14888
rect 55467 14839 55509 14848
rect 4003 14804 4061 14805
rect 4003 14764 4012 14804
rect 4052 14764 4061 14804
rect 4003 14763 4061 14764
rect 37803 14804 37845 14813
rect 37803 14764 37804 14804
rect 37844 14764 37845 14804
rect 37803 14755 37845 14764
rect 56523 14804 56565 14813
rect 56523 14764 56524 14804
rect 56564 14764 56565 14804
rect 56523 14755 56565 14764
rect 5155 14720 5213 14721
rect 5155 14680 5164 14720
rect 5204 14680 5213 14720
rect 5155 14679 5213 14680
rect 6307 14720 6365 14721
rect 6307 14680 6316 14720
rect 6356 14680 6365 14720
rect 6307 14679 6365 14680
rect 8035 14720 8093 14721
rect 8035 14680 8044 14720
rect 8084 14680 8093 14720
rect 8035 14679 8093 14680
rect 8419 14720 8477 14721
rect 8419 14680 8428 14720
rect 8468 14680 8477 14720
rect 8419 14679 8477 14680
rect 8899 14720 8957 14721
rect 8899 14680 8908 14720
rect 8948 14680 8957 14720
rect 8899 14679 8957 14680
rect 10635 14720 10677 14729
rect 10635 14680 10636 14720
rect 10676 14680 10677 14720
rect 10635 14671 10677 14680
rect 11299 14720 11357 14721
rect 11299 14680 11308 14720
rect 11348 14680 11357 14720
rect 11299 14679 11357 14680
rect 21291 14720 21333 14729
rect 21291 14680 21292 14720
rect 21332 14680 21333 14720
rect 21291 14671 21333 14680
rect 21667 14720 21725 14721
rect 21667 14680 21676 14720
rect 21716 14680 21725 14720
rect 21667 14679 21725 14680
rect 22531 14720 22589 14721
rect 22531 14680 22540 14720
rect 22580 14680 22589 14720
rect 22531 14679 22589 14680
rect 33667 14720 33725 14721
rect 33667 14680 33676 14720
rect 33716 14680 33725 14720
rect 33667 14679 33725 14680
rect 34051 14720 34109 14721
rect 34051 14680 34060 14720
rect 34100 14680 34109 14720
rect 34051 14679 34109 14680
rect 34531 14720 34589 14721
rect 34531 14680 34540 14720
rect 34580 14680 34589 14720
rect 34531 14679 34589 14680
rect 35779 14720 35837 14721
rect 35779 14680 35788 14720
rect 35828 14680 35837 14720
rect 35779 14679 35837 14680
rect 36643 14720 36701 14721
rect 36643 14680 36652 14720
rect 36692 14680 36701 14720
rect 36643 14679 36701 14680
rect 38275 14720 38333 14721
rect 38275 14680 38284 14720
rect 38324 14680 38333 14720
rect 38275 14679 38333 14680
rect 38659 14720 38717 14721
rect 38659 14680 38668 14720
rect 38708 14680 38717 14720
rect 38659 14679 38717 14680
rect 51235 14720 51293 14721
rect 51235 14680 51244 14720
rect 51284 14680 51293 14720
rect 51235 14679 51293 14680
rect 52195 14720 52253 14721
rect 52195 14680 52204 14720
rect 52244 14680 52253 14720
rect 52195 14679 52253 14680
rect 53635 14720 53693 14721
rect 53635 14680 53644 14720
rect 53684 14680 53693 14720
rect 53635 14679 53693 14680
rect 55371 14720 55413 14729
rect 55371 14680 55372 14720
rect 55412 14680 55413 14720
rect 55371 14671 55413 14680
rect 55555 14720 55613 14721
rect 55555 14680 55564 14720
rect 55604 14680 55613 14720
rect 55555 14679 55613 14680
rect 56035 14720 56093 14721
rect 56035 14680 56044 14720
rect 56084 14680 56093 14720
rect 56035 14679 56093 14680
rect 56131 14720 56189 14721
rect 56131 14680 56140 14720
rect 56180 14680 56189 14720
rect 56131 14679 56189 14680
rect 57187 14720 57245 14721
rect 57187 14680 57196 14720
rect 57236 14680 57245 14720
rect 57187 14679 57245 14680
rect 59395 14720 59453 14721
rect 59395 14680 59404 14720
rect 59444 14680 59453 14720
rect 59395 14679 59453 14680
rect 59779 14720 59837 14721
rect 59779 14680 59788 14720
rect 59828 14680 59837 14720
rect 59779 14679 59837 14680
rect 8515 14636 8573 14637
rect 8515 14596 8524 14636
rect 8564 14596 8573 14636
rect 8515 14595 8573 14596
rect 34147 14636 34205 14637
rect 34147 14596 34156 14636
rect 34196 14596 34205 14636
rect 34147 14595 34205 14596
rect 35211 14636 35253 14645
rect 35211 14596 35212 14636
rect 35252 14596 35253 14636
rect 35211 14587 35253 14596
rect 35403 14636 35445 14645
rect 35403 14596 35404 14636
rect 35444 14596 35445 14636
rect 35403 14587 35445 14596
rect 59299 14636 59357 14637
rect 59299 14596 59308 14636
rect 59348 14596 59357 14636
rect 59299 14595 59357 14596
rect 643 14552 701 14553
rect 643 14512 652 14552
rect 692 14512 701 14552
rect 643 14511 701 14512
rect 3819 14552 3861 14561
rect 3819 14512 3820 14552
rect 3860 14512 3861 14552
rect 3819 14503 3861 14512
rect 4483 14552 4541 14553
rect 4483 14512 4492 14552
rect 4532 14512 4541 14552
rect 4483 14511 4541 14512
rect 5835 14552 5877 14561
rect 5835 14512 5836 14552
rect 5876 14512 5877 14552
rect 5835 14503 5877 14512
rect 8803 14552 8861 14553
rect 8803 14512 8812 14552
rect 8852 14512 8861 14552
rect 8803 14511 8861 14512
rect 23683 14552 23741 14553
rect 23683 14512 23692 14552
rect 23732 14512 23741 14552
rect 23683 14511 23741 14512
rect 38763 14552 38805 14561
rect 38763 14512 38764 14552
rect 38804 14512 38805 14552
rect 38763 14503 38805 14512
rect 52963 14552 53021 14553
rect 52963 14512 52972 14552
rect 53012 14512 53021 14552
rect 52963 14511 53021 14512
rect 56331 14552 56373 14561
rect 56331 14512 56332 14552
rect 56372 14512 56373 14552
rect 56331 14503 56373 14512
rect 576 14384 99360 14408
rect 576 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 19472 14384
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19840 14344 34592 14384
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34960 14344 49712 14384
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 50080 14344 64832 14384
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 65200 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 95072 14384
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95440 14344 99360 14384
rect 576 14320 99360 14344
rect 5347 14216 5405 14217
rect 5347 14176 5356 14216
rect 5396 14176 5405 14216
rect 5347 14175 5405 14176
rect 11875 14216 11933 14217
rect 11875 14176 11884 14216
rect 11924 14176 11933 14216
rect 11875 14175 11933 14176
rect 18499 14216 18557 14217
rect 18499 14176 18508 14216
rect 18548 14176 18557 14216
rect 18499 14175 18557 14176
rect 55179 14216 55221 14225
rect 55179 14176 55180 14216
rect 55220 14176 55221 14216
rect 55179 14167 55221 14176
rect 61411 14216 61469 14217
rect 61411 14176 61420 14216
rect 61460 14176 61469 14216
rect 61411 14175 61469 14176
rect 2955 14132 2997 14141
rect 2955 14092 2956 14132
rect 2996 14092 2997 14132
rect 2955 14083 2997 14092
rect 7179 14132 7221 14141
rect 7179 14092 7180 14132
rect 7220 14092 7221 14132
rect 7179 14083 7221 14092
rect 9195 14132 9237 14141
rect 9195 14092 9196 14132
rect 9236 14092 9237 14132
rect 9195 14083 9237 14092
rect 43555 14132 43613 14133
rect 43555 14092 43564 14132
rect 43604 14092 43613 14132
rect 43555 14091 43613 14092
rect 50571 14132 50613 14141
rect 50571 14092 50572 14132
rect 50612 14092 50613 14132
rect 50571 14083 50613 14092
rect 57859 14132 57917 14133
rect 57859 14092 57868 14132
rect 57908 14092 57917 14132
rect 57859 14091 57917 14092
rect 3331 14048 3389 14049
rect 3331 14008 3340 14048
rect 3380 14008 3389 14048
rect 3331 14007 3389 14008
rect 4195 14048 4253 14049
rect 4195 14008 4204 14048
rect 4244 14008 4253 14048
rect 4195 14007 4253 14008
rect 6211 14048 6269 14049
rect 6211 14008 6220 14048
rect 6260 14008 6269 14048
rect 6211 14007 6269 14008
rect 7083 14048 7125 14057
rect 7083 14008 7084 14048
rect 7124 14008 7125 14048
rect 7083 13999 7125 14008
rect 7267 14048 7325 14049
rect 7267 14008 7276 14048
rect 7316 14008 7325 14048
rect 7267 14007 7325 14008
rect 9091 14048 9149 14049
rect 9091 14008 9100 14048
rect 9140 14008 9149 14048
rect 9091 14007 9149 14008
rect 9291 14048 9333 14057
rect 9291 14008 9292 14048
rect 9332 14008 9333 14048
rect 9291 13999 9333 14008
rect 9483 14048 9525 14057
rect 9483 14008 9484 14048
rect 9524 14008 9525 14048
rect 9483 13999 9525 14008
rect 9859 14048 9917 14049
rect 9859 14008 9868 14048
rect 9908 14008 9917 14048
rect 9859 14007 9917 14008
rect 10723 14048 10781 14049
rect 10723 14008 10732 14048
rect 10772 14008 10781 14048
rect 10723 14007 10781 14008
rect 12075 14048 12117 14057
rect 12075 14008 12076 14048
rect 12116 14008 12117 14048
rect 12075 13999 12117 14008
rect 12739 14048 12797 14049
rect 12739 14008 12748 14048
rect 12788 14008 12797 14048
rect 12739 14007 12797 14008
rect 19171 14048 19229 14049
rect 19171 14008 19180 14048
rect 19220 14008 19229 14048
rect 19171 14007 19229 14008
rect 26851 14048 26909 14049
rect 26851 14008 26860 14048
rect 26900 14008 26909 14048
rect 26851 14007 26909 14008
rect 27723 14048 27765 14057
rect 27723 14008 27724 14048
rect 27764 14008 27765 14048
rect 27723 13999 27765 14008
rect 39139 14048 39197 14049
rect 39139 14008 39148 14048
rect 39188 14008 39197 14048
rect 39139 14007 39197 14008
rect 43747 14048 43805 14049
rect 43747 14008 43756 14048
rect 43796 14008 43805 14048
rect 43747 14007 43805 14008
rect 44035 14048 44093 14049
rect 44035 14008 44044 14048
rect 44084 14008 44093 14048
rect 44035 14007 44093 14008
rect 45379 14048 45437 14049
rect 45379 14008 45388 14048
rect 45428 14008 45437 14048
rect 45379 14007 45437 14008
rect 46243 14048 46301 14049
rect 46243 14008 46252 14048
rect 46292 14008 46301 14048
rect 46243 14007 46301 14008
rect 46635 14048 46677 14057
rect 46635 14008 46636 14048
rect 46676 14008 46677 14048
rect 46635 13999 46677 14008
rect 47307 14048 47349 14057
rect 47307 14008 47308 14048
rect 47348 14008 47349 14048
rect 47307 13999 47349 14008
rect 47971 14048 48029 14049
rect 47971 14008 47980 14048
rect 48020 14008 48029 14048
rect 47971 14007 48029 14008
rect 49315 14048 49373 14049
rect 49315 14008 49324 14048
rect 49364 14008 49373 14048
rect 49315 14007 49373 14008
rect 50179 14048 50237 14049
rect 50179 14008 50188 14048
rect 50228 14008 50237 14048
rect 50179 14007 50237 14008
rect 55363 14048 55421 14049
rect 55363 14008 55372 14048
rect 55412 14008 55421 14048
rect 55363 14007 55421 14008
rect 55651 14048 55709 14049
rect 55651 14008 55660 14048
rect 55700 14008 55709 14048
rect 55651 14007 55709 14008
rect 56707 14048 56765 14049
rect 56707 14008 56716 14048
rect 56756 14008 56765 14048
rect 56707 14007 56765 14008
rect 56995 14048 57053 14049
rect 56995 14008 57004 14048
rect 57044 14008 57053 14048
rect 56995 14007 57053 14008
rect 59019 14048 59061 14057
rect 59019 14008 59020 14048
rect 59060 14008 59061 14048
rect 59019 13999 59061 14008
rect 59395 14048 59453 14049
rect 59395 14008 59404 14048
rect 59444 14008 59453 14048
rect 59395 14007 59453 14008
rect 60259 14048 60317 14049
rect 60259 14008 60268 14048
rect 60308 14008 60317 14048
rect 60259 14007 60317 14008
rect 5731 13964 5789 13965
rect 5731 13924 5740 13964
rect 5780 13924 5789 13964
rect 5731 13923 5789 13924
rect 6891 13964 6933 13973
rect 6891 13924 6892 13964
rect 6932 13924 6933 13964
rect 6891 13915 6933 13924
rect 17539 13964 17597 13965
rect 17539 13924 17548 13964
rect 17588 13924 17597 13964
rect 17539 13923 17597 13924
rect 44235 13964 44277 13973
rect 44235 13924 44236 13964
rect 44276 13924 44277 13964
rect 44235 13915 44277 13924
rect 5547 13880 5589 13889
rect 5547 13840 5548 13880
rect 5588 13840 5589 13880
rect 5547 13831 5589 13840
rect 57291 13880 57333 13889
rect 57291 13840 57292 13880
rect 57332 13840 57333 13880
rect 57291 13831 57333 13840
rect 17355 13796 17397 13805
rect 17355 13756 17356 13796
rect 17396 13756 17397 13796
rect 17355 13747 17397 13756
rect 38467 13796 38525 13797
rect 38467 13756 38476 13796
rect 38516 13756 38525 13796
rect 38467 13755 38525 13756
rect 48163 13796 48221 13797
rect 48163 13756 48172 13796
rect 48212 13756 48221 13796
rect 48163 13755 48221 13756
rect 56035 13796 56093 13797
rect 56035 13756 56044 13796
rect 56084 13756 56093 13796
rect 56035 13755 56093 13756
rect 576 13628 99360 13652
rect 576 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 18232 13628
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18600 13588 33352 13628
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33720 13588 48472 13628
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48840 13588 63592 13628
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63960 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 93832 13628
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 94200 13588 99360 13628
rect 576 13564 99360 13588
rect 6403 13460 6461 13461
rect 6403 13420 6412 13460
rect 6452 13420 6461 13460
rect 6403 13419 6461 13420
rect 9291 13460 9333 13469
rect 9291 13420 9292 13460
rect 9332 13420 9333 13460
rect 9291 13411 9333 13420
rect 12259 13460 12317 13461
rect 12259 13420 12268 13460
rect 12308 13420 12317 13460
rect 12259 13419 12317 13420
rect 19267 13460 19325 13461
rect 19267 13420 19276 13460
rect 19316 13420 19325 13460
rect 19267 13419 19325 13420
rect 49611 13460 49653 13469
rect 49611 13420 49612 13460
rect 49652 13420 49653 13460
rect 49611 13411 49653 13420
rect 23115 13376 23157 13385
rect 23115 13336 23116 13376
rect 23156 13336 23157 13376
rect 23115 13327 23157 13336
rect 9091 13292 9149 13293
rect 9091 13252 9100 13292
rect 9140 13252 9149 13292
rect 9091 13251 9149 13252
rect 9475 13292 9533 13293
rect 9475 13252 9484 13292
rect 9524 13252 9533 13292
rect 9475 13251 9533 13252
rect 4011 13208 4053 13217
rect 4011 13168 4012 13208
rect 4052 13168 4053 13208
rect 4011 13159 4053 13168
rect 4387 13208 4445 13209
rect 4387 13168 4396 13208
rect 4436 13168 4445 13208
rect 4387 13167 4445 13168
rect 5251 13208 5309 13209
rect 5251 13168 5260 13208
rect 5300 13168 5309 13208
rect 5251 13167 5309 13168
rect 10243 13208 10301 13209
rect 10243 13168 10252 13208
rect 10292 13168 10301 13208
rect 10243 13167 10301 13168
rect 11107 13208 11165 13209
rect 11107 13168 11116 13208
rect 11156 13168 11165 13208
rect 11107 13167 11165 13168
rect 16875 13208 16917 13217
rect 16875 13168 16876 13208
rect 16916 13168 16917 13208
rect 16875 13159 16917 13168
rect 17251 13208 17309 13209
rect 17251 13168 17260 13208
rect 17300 13168 17309 13208
rect 17251 13167 17309 13168
rect 18115 13208 18173 13209
rect 18115 13168 18124 13208
rect 18164 13168 18173 13208
rect 18115 13167 18173 13168
rect 23019 13208 23061 13217
rect 23019 13168 23020 13208
rect 23060 13168 23061 13208
rect 23019 13159 23061 13168
rect 23203 13208 23261 13209
rect 23203 13168 23212 13208
rect 23252 13168 23261 13208
rect 23203 13167 23261 13168
rect 23491 13208 23549 13209
rect 23491 13168 23500 13208
rect 23540 13168 23549 13208
rect 23491 13167 23549 13168
rect 26083 13208 26141 13209
rect 26083 13168 26092 13208
rect 26132 13168 26141 13208
rect 26083 13167 26141 13168
rect 38475 13208 38517 13217
rect 38475 13168 38476 13208
rect 38516 13168 38517 13208
rect 38475 13159 38517 13168
rect 38851 13208 38909 13209
rect 38851 13168 38860 13208
rect 38900 13168 38909 13208
rect 38851 13167 38909 13168
rect 39715 13208 39773 13209
rect 39715 13168 39724 13208
rect 39764 13168 39773 13208
rect 39715 13167 39773 13168
rect 41635 13208 41693 13209
rect 41635 13168 41644 13208
rect 41684 13168 41693 13208
rect 41635 13167 41693 13168
rect 48643 13208 48701 13209
rect 48643 13168 48652 13208
rect 48692 13168 48701 13208
rect 48643 13167 48701 13168
rect 49795 13208 49853 13209
rect 49795 13168 49804 13208
rect 49844 13168 49853 13208
rect 49795 13167 49853 13168
rect 49899 13208 49941 13217
rect 49899 13168 49900 13208
rect 49940 13168 49941 13208
rect 49899 13159 49941 13168
rect 54787 13208 54845 13209
rect 54787 13168 54796 13208
rect 54836 13168 54845 13208
rect 54787 13167 54845 13168
rect 55651 13208 55709 13209
rect 55651 13168 55660 13208
rect 55700 13168 55709 13208
rect 55651 13167 55709 13168
rect 56043 13208 56085 13217
rect 56043 13168 56044 13208
rect 56084 13168 56085 13208
rect 56043 13159 56085 13168
rect 56611 13208 56669 13209
rect 56611 13168 56620 13208
rect 56660 13168 56669 13208
rect 56611 13167 56669 13168
rect 9867 13124 9909 13133
rect 9867 13084 9868 13124
rect 9908 13084 9909 13124
rect 9867 13075 9909 13084
rect 643 13040 701 13041
rect 643 13000 652 13040
rect 692 13000 701 13040
rect 643 12999 701 13000
rect 9675 13040 9717 13049
rect 9675 13000 9676 13040
rect 9716 13000 9717 13040
rect 9675 12991 9717 13000
rect 24163 13040 24221 13041
rect 24163 13000 24172 13040
rect 24212 13000 24221 13040
rect 24163 12999 24221 13000
rect 26755 13040 26813 13041
rect 26755 13000 26764 13040
rect 26804 13000 26813 13040
rect 26755 12999 26813 13000
rect 40867 13040 40925 13041
rect 40867 13000 40876 13040
rect 40916 13000 40925 13040
rect 40867 12999 40925 13000
rect 42307 13040 42365 13041
rect 42307 13000 42316 13040
rect 42356 13000 42365 13040
rect 42307 12999 42365 13000
rect 49315 13040 49373 13041
rect 49315 13000 49324 13040
rect 49364 13000 49373 13040
rect 49315 12999 49373 13000
rect 53635 13040 53693 13041
rect 53635 13000 53644 13040
rect 53684 13000 53693 13040
rect 53635 12999 53693 13000
rect 576 12872 99360 12896
rect 576 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 19472 12872
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19840 12832 34592 12872
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34960 12832 49712 12872
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 50080 12832 64832 12872
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 65200 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 95072 12872
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95440 12832 99360 12872
rect 576 12808 99360 12832
rect 643 12704 701 12705
rect 643 12664 652 12704
rect 692 12664 701 12704
rect 643 12663 701 12664
rect 31651 12704 31709 12705
rect 31651 12664 31660 12704
rect 31700 12664 31709 12704
rect 31651 12663 31709 12664
rect 50475 12704 50517 12713
rect 50475 12664 50476 12704
rect 50516 12664 50517 12704
rect 50475 12655 50517 12664
rect 23203 12620 23261 12621
rect 23203 12580 23212 12620
rect 23252 12580 23261 12620
rect 23203 12579 23261 12580
rect 23787 12620 23829 12629
rect 23787 12580 23788 12620
rect 23828 12580 23829 12620
rect 23787 12571 23829 12580
rect 28299 12620 28341 12629
rect 28299 12580 28300 12620
rect 28340 12580 28341 12620
rect 28299 12571 28341 12580
rect 42699 12620 42741 12629
rect 42699 12580 42700 12620
rect 42740 12580 42741 12620
rect 42699 12571 42741 12580
rect 49419 12620 49461 12629
rect 49419 12580 49420 12620
rect 49460 12580 49461 12620
rect 49419 12571 49461 12580
rect 9475 12536 9533 12537
rect 9475 12496 9484 12536
rect 9524 12496 9533 12536
rect 9475 12495 9533 12496
rect 19371 12536 19413 12545
rect 19371 12496 19372 12536
rect 19412 12496 19413 12536
rect 19371 12487 19413 12496
rect 21283 12536 21341 12537
rect 21283 12496 21292 12536
rect 21332 12496 21341 12536
rect 21283 12495 21341 12496
rect 22723 12536 22781 12537
rect 22723 12496 22732 12536
rect 22772 12496 22781 12536
rect 22723 12495 22781 12496
rect 23011 12536 23069 12537
rect 23011 12496 23020 12536
rect 23060 12496 23069 12536
rect 23011 12495 23069 12496
rect 23499 12536 23541 12545
rect 23499 12496 23500 12536
rect 23540 12496 23541 12536
rect 23499 12487 23541 12496
rect 23595 12536 23637 12545
rect 23595 12496 23596 12536
rect 23636 12496 23637 12536
rect 23595 12487 23637 12496
rect 23691 12536 23733 12545
rect 23691 12496 23692 12536
rect 23732 12496 23733 12536
rect 23691 12487 23733 12496
rect 23972 12535 24014 12544
rect 23972 12495 23973 12535
rect 24013 12495 24014 12535
rect 23972 12486 24014 12495
rect 24171 12536 24213 12545
rect 24171 12496 24172 12536
rect 24212 12496 24213 12536
rect 24171 12487 24213 12496
rect 28675 12536 28733 12537
rect 28675 12496 28684 12536
rect 28724 12496 28733 12536
rect 28675 12495 28733 12496
rect 29539 12536 29597 12537
rect 29539 12496 29548 12536
rect 29588 12496 29597 12536
rect 29539 12495 29597 12496
rect 31171 12536 31229 12537
rect 31171 12496 31180 12536
rect 31220 12496 31229 12536
rect 31171 12495 31229 12496
rect 31275 12536 31317 12545
rect 31275 12496 31276 12536
rect 31316 12496 31317 12536
rect 31275 12487 31317 12496
rect 31747 12536 31805 12537
rect 31747 12496 31756 12536
rect 31796 12496 31805 12536
rect 31747 12495 31805 12496
rect 35875 12536 35933 12537
rect 35875 12496 35884 12536
rect 35924 12496 35933 12536
rect 35875 12495 35933 12496
rect 41731 12536 41789 12537
rect 41731 12496 41740 12536
rect 41780 12496 41789 12536
rect 41731 12495 41789 12496
rect 42603 12536 42645 12545
rect 42603 12496 42604 12536
rect 42644 12496 42645 12536
rect 42603 12487 42645 12496
rect 42787 12536 42845 12537
rect 42787 12496 42796 12536
rect 42836 12496 42845 12536
rect 42787 12495 42845 12496
rect 49323 12536 49365 12545
rect 49323 12496 49324 12536
rect 49364 12496 49365 12536
rect 49323 12487 49365 12496
rect 49507 12536 49565 12537
rect 49507 12496 49516 12536
rect 49556 12496 49565 12536
rect 49507 12495 49565 12496
rect 50563 12536 50621 12537
rect 50563 12496 50572 12536
rect 50612 12496 50621 12536
rect 50563 12495 50621 12496
rect 50947 12536 51005 12537
rect 50947 12496 50956 12536
rect 50996 12496 51005 12536
rect 50947 12495 51005 12496
rect 53155 12536 53213 12537
rect 53155 12496 53164 12536
rect 53204 12496 53213 12536
rect 53155 12495 53213 12496
rect 54115 12536 54173 12537
rect 54115 12496 54124 12536
rect 54164 12496 54173 12536
rect 54115 12495 54173 12496
rect 54411 12536 54453 12545
rect 54411 12496 54412 12536
rect 54452 12496 54453 12536
rect 54411 12487 54453 12496
rect 54787 12536 54845 12537
rect 54787 12496 54796 12536
rect 54836 12496 54845 12536
rect 54787 12495 54845 12496
rect 55651 12536 55709 12537
rect 55651 12496 55660 12536
rect 55700 12496 55709 12536
rect 55651 12495 55709 12496
rect 30699 12452 30741 12461
rect 30699 12412 30700 12452
rect 30740 12412 30741 12452
rect 30699 12403 30741 12412
rect 30883 12452 30941 12453
rect 30883 12412 30892 12452
rect 30932 12412 30941 12452
rect 30883 12411 30941 12412
rect 41155 12452 41213 12453
rect 41155 12412 41164 12452
rect 41204 12412 41213 12452
rect 41155 12411 41213 12412
rect 56811 12452 56853 12461
rect 56811 12412 56812 12452
rect 56852 12412 56853 12452
rect 56811 12403 56853 12412
rect 9003 12368 9045 12377
rect 9003 12328 9004 12368
rect 9044 12328 9045 12368
rect 9003 12319 9045 12328
rect 18795 12368 18837 12377
rect 18795 12328 18796 12368
rect 18836 12328 18837 12368
rect 18795 12319 18837 12328
rect 23979 12368 24021 12377
rect 23979 12328 23980 12368
rect 24020 12328 24021 12368
rect 23979 12319 24021 12328
rect 21771 12284 21813 12293
rect 21771 12244 21772 12284
rect 21812 12244 21813 12284
rect 21771 12235 21813 12244
rect 31939 12284 31997 12285
rect 31939 12244 31948 12284
rect 31988 12244 31997 12284
rect 31939 12243 31997 12244
rect 35211 12284 35253 12293
rect 35211 12244 35212 12284
rect 35252 12244 35253 12284
rect 35211 12235 35253 12244
rect 42403 12284 42461 12285
rect 42403 12244 42412 12284
rect 42452 12244 42461 12284
rect 42403 12243 42461 12244
rect 576 12116 99360 12140
rect 576 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 18232 12116
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18600 12076 33352 12116
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33720 12076 48472 12116
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48840 12076 63592 12116
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63960 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 93832 12116
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 94200 12076 99360 12116
rect 576 12052 99360 12076
rect 30307 11948 30365 11949
rect 30307 11908 30316 11948
rect 30356 11908 30365 11948
rect 30307 11907 30365 11908
rect 41931 11948 41973 11957
rect 41931 11908 41932 11948
rect 41972 11908 41973 11948
rect 41931 11899 41973 11908
rect 49507 11948 49565 11949
rect 49507 11908 49516 11948
rect 49556 11908 49565 11948
rect 49507 11907 49565 11908
rect 53835 11948 53877 11957
rect 53835 11908 53836 11948
rect 53876 11908 53877 11948
rect 53835 11899 53877 11908
rect 29931 11864 29973 11873
rect 29931 11824 29932 11864
rect 29972 11824 29973 11864
rect 29931 11815 29973 11824
rect 42891 11864 42933 11873
rect 42891 11824 42892 11864
rect 42932 11824 42933 11864
rect 42891 11815 42933 11824
rect 23683 11780 23741 11781
rect 23683 11740 23692 11780
rect 23732 11740 23741 11780
rect 23683 11739 23741 11740
rect 18115 11696 18173 11697
rect 18115 11656 18124 11696
rect 18164 11656 18173 11696
rect 18115 11655 18173 11656
rect 18987 11696 19029 11705
rect 18987 11656 18988 11696
rect 19028 11656 19029 11696
rect 18987 11647 19029 11656
rect 23307 11696 23349 11705
rect 23307 11656 23308 11696
rect 23348 11656 23349 11696
rect 23307 11647 23349 11656
rect 23395 11696 23453 11697
rect 23395 11656 23404 11696
rect 23444 11656 23453 11696
rect 23395 11655 23453 11656
rect 24163 11696 24221 11697
rect 24163 11656 24172 11696
rect 24212 11656 24221 11696
rect 24163 11655 24221 11656
rect 29931 11696 29973 11705
rect 29931 11656 29932 11696
rect 29972 11656 29973 11696
rect 29931 11647 29973 11656
rect 31459 11696 31517 11697
rect 31459 11656 31468 11696
rect 31508 11656 31517 11696
rect 31459 11655 31517 11656
rect 32323 11696 32381 11697
rect 32323 11656 32332 11696
rect 32372 11656 32381 11696
rect 32323 11655 32381 11656
rect 41347 11696 41405 11697
rect 41347 11656 41356 11696
rect 41396 11656 41405 11696
rect 41347 11655 41405 11656
rect 41635 11696 41693 11697
rect 41635 11656 41644 11696
rect 41684 11656 41693 11696
rect 41635 11655 41693 11656
rect 42595 11696 42653 11697
rect 42595 11656 42604 11696
rect 42644 11656 42653 11696
rect 42595 11655 42653 11656
rect 43075 11696 43133 11697
rect 43075 11656 43084 11696
rect 43124 11656 43133 11696
rect 43075 11655 43133 11656
rect 43179 11696 43221 11705
rect 43179 11656 43180 11696
rect 43220 11656 43221 11696
rect 43179 11647 43221 11656
rect 47299 11696 47357 11697
rect 47299 11656 47308 11696
rect 47348 11656 47357 11696
rect 47299 11655 47357 11656
rect 49027 11696 49085 11697
rect 49027 11656 49036 11696
rect 49076 11656 49085 11696
rect 49027 11655 49085 11656
rect 49315 11696 49373 11697
rect 49315 11656 49324 11696
rect 49364 11656 49373 11696
rect 49315 11655 49373 11656
rect 50179 11696 50237 11697
rect 50179 11656 50188 11696
rect 50228 11656 50237 11696
rect 50179 11655 50237 11656
rect 53539 11696 53597 11697
rect 53539 11656 53548 11696
rect 53588 11656 53597 11696
rect 53539 11655 53597 11656
rect 61795 11696 61853 11697
rect 61795 11656 61804 11696
rect 61844 11656 61853 11696
rect 61795 11655 61853 11656
rect 32715 11612 32757 11621
rect 32715 11572 32716 11612
rect 32756 11572 32757 11612
rect 32715 11563 32757 11572
rect 48835 11612 48893 11613
rect 48835 11572 48844 11612
rect 48884 11572 48893 11612
rect 48835 11571 48893 11572
rect 643 11528 701 11529
rect 643 11488 652 11528
rect 692 11488 701 11528
rect 643 11487 701 11488
rect 24835 11528 24893 11529
rect 24835 11488 24844 11528
rect 24884 11488 24893 11528
rect 24835 11487 24893 11488
rect 30123 11528 30165 11537
rect 30123 11488 30124 11528
rect 30164 11488 30165 11528
rect 30123 11479 30165 11488
rect 40675 11528 40733 11529
rect 40675 11488 40684 11528
rect 40724 11488 40733 11528
rect 40675 11487 40733 11488
rect 46627 11528 46685 11529
rect 46627 11488 46636 11528
rect 46676 11488 46685 11528
rect 46627 11487 46685 11488
rect 61123 11528 61181 11529
rect 61123 11488 61132 11528
rect 61172 11488 61181 11528
rect 61123 11487 61181 11488
rect 576 11360 99360 11384
rect 576 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 19472 11360
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19840 11320 34592 11360
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34960 11320 49712 11360
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 50080 11320 64832 11360
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 65200 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 95072 11360
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95440 11320 99360 11360
rect 576 11296 99360 11320
rect 643 11192 701 11193
rect 643 11152 652 11192
rect 692 11152 701 11192
rect 643 11151 701 11152
rect 18691 11192 18749 11193
rect 18691 11152 18700 11192
rect 18740 11152 18749 11192
rect 18691 11151 18749 11152
rect 32227 11192 32285 11193
rect 32227 11152 32236 11192
rect 32276 11152 32285 11192
rect 32227 11151 32285 11152
rect 33091 11192 33149 11193
rect 33091 11152 33100 11192
rect 33140 11152 33149 11192
rect 33091 11151 33149 11152
rect 41923 11192 41981 11193
rect 41923 11152 41932 11192
rect 41972 11152 41981 11192
rect 41923 11151 41981 11152
rect 59211 11192 59253 11201
rect 59211 11152 59212 11192
rect 59252 11152 59253 11192
rect 59211 11143 59253 11152
rect 61987 11192 62045 11193
rect 61987 11152 61996 11192
rect 62036 11152 62045 11192
rect 61987 11151 62045 11152
rect 24459 11108 24501 11117
rect 24459 11068 24460 11108
rect 24500 11068 24501 11108
rect 24459 11059 24501 11068
rect 44331 11108 44373 11117
rect 44331 11068 44332 11108
rect 44372 11068 44373 11108
rect 44331 11059 44373 11068
rect 10243 11024 10301 11025
rect 10243 10984 10252 11024
rect 10292 10984 10301 11024
rect 10243 10983 10301 10984
rect 13603 11024 13661 11025
rect 13603 10984 13612 11024
rect 13652 10984 13661 11024
rect 13603 10983 13661 10984
rect 15427 11024 15485 11025
rect 15427 10984 15436 11024
rect 15476 10984 15485 11024
rect 15427 10983 15485 10984
rect 16107 11024 16149 11033
rect 16107 10984 16108 11024
rect 16148 10984 16149 11024
rect 16107 10975 16149 10984
rect 16299 11024 16341 11033
rect 16299 10984 16300 11024
rect 16340 10984 16341 11024
rect 16299 10975 16341 10984
rect 16675 11024 16733 11025
rect 16675 10984 16684 11024
rect 16724 10984 16733 11024
rect 16675 10983 16733 10984
rect 17539 11024 17597 11025
rect 17539 10984 17548 11024
rect 17588 10984 17597 11024
rect 17539 10983 17597 10984
rect 20707 11024 20765 11025
rect 20707 10984 20716 11024
rect 20756 10984 20765 11024
rect 20707 10983 20765 10984
rect 21667 11024 21725 11025
rect 21667 10984 21676 11024
rect 21716 10984 21725 11024
rect 21667 10983 21725 10984
rect 24835 11024 24893 11025
rect 24835 10984 24844 11024
rect 24884 10984 24893 11024
rect 24835 10983 24893 10984
rect 25699 11024 25757 11025
rect 25699 10984 25708 11024
rect 25748 10984 25757 11024
rect 25699 10983 25757 10984
rect 31171 11024 31229 11025
rect 31171 10984 31180 11024
rect 31220 10984 31229 11024
rect 31363 11024 31421 11025
rect 31171 10983 31229 10984
rect 31275 10989 31317 10998
rect 31275 10949 31276 10989
rect 31316 10949 31317 10989
rect 31363 10984 31372 11024
rect 31412 10984 31421 11024
rect 31363 10983 31421 10984
rect 31947 11024 31989 11033
rect 31947 10984 31948 11024
rect 31988 10984 31989 11024
rect 31947 10975 31989 10984
rect 32043 11024 32085 11033
rect 32043 10984 32044 11024
rect 32084 10984 32085 11024
rect 32043 10975 32085 10984
rect 33763 11024 33821 11025
rect 33763 10984 33772 11024
rect 33812 10984 33821 11024
rect 33763 10983 33821 10984
rect 37027 11024 37085 11025
rect 37027 10984 37036 11024
rect 37076 10984 37085 11024
rect 37027 10983 37085 10984
rect 37891 11024 37949 11025
rect 37891 10984 37900 11024
rect 37940 10984 37949 11024
rect 37891 10983 37949 10984
rect 38283 11024 38325 11033
rect 38283 10984 38284 11024
rect 38324 10984 38325 11024
rect 38283 10975 38325 10984
rect 41155 11024 41213 11025
rect 41155 10984 41164 11024
rect 41204 10984 41213 11024
rect 41155 10983 41213 10984
rect 43075 11024 43133 11025
rect 43075 10984 43084 11024
rect 43124 10984 43133 11024
rect 43075 10983 43133 10984
rect 43939 11024 43997 11025
rect 43939 10984 43948 11024
rect 43988 10984 43997 11024
rect 43939 10983 43997 10984
rect 52579 11024 52637 11025
rect 52579 10984 52588 11024
rect 52628 10984 52637 11024
rect 52579 10983 52637 10984
rect 58723 11024 58781 11025
rect 58723 10984 58732 11024
rect 58772 10984 58781 11024
rect 58723 10983 58781 10984
rect 59011 11024 59069 11025
rect 59011 10984 59020 11024
rect 59060 10984 59069 11024
rect 59011 10983 59069 10984
rect 59595 11024 59637 11033
rect 59595 10984 59596 11024
rect 59636 10984 59637 11024
rect 59595 10975 59637 10984
rect 59971 11024 60029 11025
rect 59971 10984 59980 11024
rect 60020 10984 60029 11024
rect 59971 10983 60029 10984
rect 60835 11024 60893 11025
rect 60835 10984 60844 11024
rect 60884 10984 60893 11024
rect 60835 10983 60893 10984
rect 31275 10940 31317 10949
rect 51723 10940 51765 10949
rect 51723 10900 51724 10940
rect 51764 10900 51765 10940
rect 51723 10891 51765 10900
rect 9579 10772 9621 10781
rect 9579 10732 9580 10772
rect 9620 10732 9621 10772
rect 9579 10723 9621 10732
rect 12931 10772 12989 10773
rect 12931 10732 12940 10772
rect 12980 10732 12989 10772
rect 12931 10731 12989 10732
rect 26851 10772 26909 10773
rect 26851 10732 26860 10772
rect 26900 10732 26909 10772
rect 26851 10731 26909 10732
rect 30891 10772 30933 10781
rect 30891 10732 30892 10772
rect 30932 10732 30933 10772
rect 30891 10723 30933 10732
rect 35883 10772 35925 10781
rect 35883 10732 35884 10772
rect 35924 10732 35925 10772
rect 35883 10723 35925 10732
rect 40483 10772 40541 10773
rect 40483 10732 40492 10772
rect 40532 10732 40541 10772
rect 40483 10731 40541 10732
rect 576 10604 99360 10628
rect 576 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 18232 10604
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18600 10564 33352 10604
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33720 10564 48472 10604
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48840 10564 63592 10604
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63960 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 93832 10604
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 94200 10564 99360 10604
rect 576 10540 99360 10564
rect 15331 10436 15389 10437
rect 15331 10396 15340 10436
rect 15380 10396 15389 10436
rect 15331 10395 15389 10396
rect 21963 10436 22005 10445
rect 21963 10396 21964 10436
rect 22004 10396 22005 10436
rect 21963 10387 22005 10396
rect 49219 10436 49277 10437
rect 49219 10396 49228 10436
rect 49268 10396 49277 10436
rect 49219 10395 49277 10396
rect 55171 10436 55229 10437
rect 55171 10396 55180 10436
rect 55220 10396 55229 10436
rect 55171 10395 55229 10396
rect 58539 10436 58581 10445
rect 58539 10396 58540 10436
rect 58580 10396 58581 10436
rect 58539 10387 58581 10396
rect 58923 10436 58965 10445
rect 58923 10396 58924 10436
rect 58964 10396 58965 10436
rect 58923 10387 58965 10396
rect 59787 10436 59829 10445
rect 59787 10396 59788 10436
rect 59828 10396 59829 10436
rect 59787 10387 59829 10396
rect 3147 10352 3189 10361
rect 3147 10312 3148 10352
rect 3188 10312 3189 10352
rect 3147 10303 3189 10312
rect 55843 10352 55901 10353
rect 55843 10312 55852 10352
rect 55892 10312 55901 10352
rect 55843 10311 55901 10312
rect 3331 10268 3389 10269
rect 3331 10228 3340 10268
rect 3380 10228 3389 10268
rect 3331 10227 3389 10228
rect 37899 10268 37941 10277
rect 37899 10228 37900 10268
rect 37940 10228 37941 10268
rect 37899 10219 37941 10228
rect 59971 10268 60029 10269
rect 59971 10228 59980 10268
rect 60020 10228 60029 10268
rect 59971 10227 60029 10228
rect 4771 10184 4829 10185
rect 4771 10144 4780 10184
rect 4820 10144 4829 10184
rect 4771 10143 4829 10144
rect 9859 10184 9917 10185
rect 9859 10144 9868 10184
rect 9908 10144 9917 10184
rect 9859 10143 9917 10144
rect 12547 10184 12605 10185
rect 12547 10144 12556 10184
rect 12596 10144 12605 10184
rect 12547 10143 12605 10144
rect 12739 10184 12797 10185
rect 12739 10144 12748 10184
rect 12788 10144 12797 10184
rect 12739 10143 12797 10144
rect 12939 10184 12981 10193
rect 12939 10144 12940 10184
rect 12980 10144 12981 10184
rect 12939 10135 12981 10144
rect 13315 10184 13373 10185
rect 13315 10144 13324 10184
rect 13364 10144 13373 10184
rect 13315 10143 13373 10144
rect 14179 10184 14237 10185
rect 14179 10144 14188 10184
rect 14228 10144 14237 10184
rect 14179 10143 14237 10144
rect 21091 10184 21149 10185
rect 21091 10144 21100 10184
rect 21140 10144 21149 10184
rect 21091 10143 21149 10144
rect 21475 10184 21533 10185
rect 21475 10144 21484 10184
rect 21524 10144 21533 10184
rect 21475 10143 21533 10144
rect 21867 10184 21909 10193
rect 21867 10144 21868 10184
rect 21908 10144 21909 10184
rect 21867 10135 21909 10144
rect 22051 10184 22109 10185
rect 22051 10144 22060 10184
rect 22100 10144 22109 10184
rect 22051 10143 22109 10144
rect 27819 10184 27861 10193
rect 27819 10144 27820 10184
rect 27860 10144 27861 10184
rect 27819 10135 27861 10144
rect 28011 10184 28053 10193
rect 28011 10144 28012 10184
rect 28052 10144 28053 10184
rect 28011 10135 28053 10144
rect 28203 10184 28245 10193
rect 28203 10144 28204 10184
rect 28244 10144 28245 10184
rect 28203 10135 28245 10144
rect 28387 10184 28445 10185
rect 28387 10144 28396 10184
rect 28436 10144 28445 10184
rect 28387 10143 28445 10144
rect 37027 10184 37085 10185
rect 37027 10144 37036 10184
rect 37076 10144 37085 10184
rect 37027 10143 37085 10144
rect 38179 10184 38237 10185
rect 38179 10144 38188 10184
rect 38228 10144 38237 10184
rect 38179 10143 38237 10144
rect 39051 10184 39093 10193
rect 39051 10144 39052 10184
rect 39092 10144 39093 10184
rect 39051 10135 39093 10144
rect 41443 10184 41501 10185
rect 41443 10144 41452 10184
rect 41492 10144 41501 10184
rect 41443 10143 41501 10144
rect 41731 10184 41789 10185
rect 41731 10144 41740 10184
rect 41780 10144 41789 10184
rect 41731 10143 41789 10144
rect 47203 10184 47261 10185
rect 47203 10144 47212 10184
rect 47252 10144 47261 10184
rect 47203 10143 47261 10144
rect 48067 10184 48125 10185
rect 48067 10144 48076 10184
rect 48116 10144 48125 10184
rect 48067 10143 48125 10144
rect 55363 10184 55421 10185
rect 55363 10144 55372 10184
rect 55412 10144 55421 10184
rect 55363 10143 55421 10144
rect 56515 10184 56573 10185
rect 56515 10144 56524 10184
rect 56564 10144 56573 10184
rect 56515 10143 56573 10144
rect 58443 10184 58485 10193
rect 58443 10144 58444 10184
rect 58484 10144 58485 10184
rect 58443 10135 58485 10144
rect 58627 10184 58685 10185
rect 58627 10144 58636 10184
rect 58676 10144 58685 10184
rect 58627 10143 58685 10144
rect 58819 10184 58877 10185
rect 58819 10144 58828 10184
rect 58868 10144 58877 10184
rect 58819 10143 58877 10144
rect 59019 10184 59061 10193
rect 59019 10144 59020 10184
rect 59060 10144 59061 10184
rect 59019 10135 59061 10144
rect 61411 10184 61469 10185
rect 61411 10144 61420 10184
rect 61460 10144 61469 10184
rect 61411 10143 61469 10144
rect 4107 10100 4149 10109
rect 4107 10060 4108 10100
rect 4148 10060 4149 10100
rect 4107 10051 4149 10060
rect 28299 10100 28341 10109
rect 28299 10060 28300 10100
rect 28340 10060 28341 10100
rect 28299 10051 28341 10060
rect 41251 10100 41309 10101
rect 41251 10060 41260 10100
rect 41300 10060 41309 10100
rect 41251 10059 41309 10060
rect 46827 10100 46869 10109
rect 46827 10060 46828 10100
rect 46868 10060 46869 10100
rect 46827 10051 46869 10060
rect 60747 10100 60789 10109
rect 60747 10060 60748 10100
rect 60788 10060 60789 10100
rect 60747 10051 60789 10060
rect 643 10016 701 10017
rect 643 9976 652 10016
rect 692 9976 701 10016
rect 643 9975 701 9976
rect 10531 10016 10589 10017
rect 10531 9976 10540 10016
rect 10580 9976 10589 10016
rect 10531 9975 10589 9976
rect 21579 10016 21621 10025
rect 21579 9976 21580 10016
rect 21620 9976 21621 10016
rect 21579 9967 21621 9976
rect 27915 10016 27957 10025
rect 27915 9976 27916 10016
rect 27956 9976 27957 10016
rect 27915 9967 27957 9976
rect 55459 10016 55517 10017
rect 55459 9976 55468 10016
rect 55508 9976 55517 10016
rect 55459 9975 55517 9976
rect 576 9848 99360 9872
rect 576 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 19472 9848
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19840 9808 34592 9848
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34960 9808 49712 9848
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 50080 9808 64832 9848
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 65200 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 95072 9848
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95440 9808 99360 9848
rect 576 9784 99360 9808
rect 643 9680 701 9681
rect 643 9640 652 9680
rect 692 9640 701 9680
rect 643 9639 701 9640
rect 4675 9680 4733 9681
rect 4675 9640 4684 9680
rect 4724 9640 4733 9680
rect 4675 9639 4733 9640
rect 9187 9680 9245 9681
rect 9187 9640 9196 9680
rect 9236 9640 9245 9680
rect 9187 9639 9245 9640
rect 12739 9680 12797 9681
rect 12739 9640 12748 9680
rect 12788 9640 12797 9680
rect 12739 9639 12797 9640
rect 20995 9680 21053 9681
rect 20995 9640 21004 9680
rect 21044 9640 21053 9680
rect 20995 9639 21053 9640
rect 32995 9680 33053 9681
rect 32995 9640 33004 9680
rect 33044 9640 33053 9680
rect 32995 9639 33053 9640
rect 33475 9680 33533 9681
rect 33475 9640 33484 9680
rect 33524 9640 33533 9680
rect 33475 9639 33533 9640
rect 47011 9680 47069 9681
rect 47011 9640 47020 9680
rect 47060 9640 47069 9680
rect 47011 9639 47069 9640
rect 50467 9680 50525 9681
rect 50467 9640 50476 9680
rect 50516 9640 50525 9680
rect 50467 9639 50525 9640
rect 59403 9680 59445 9689
rect 59403 9640 59404 9680
rect 59444 9640 59445 9680
rect 59403 9631 59445 9640
rect 61987 9680 62045 9681
rect 61987 9640 61996 9680
rect 62036 9640 62045 9680
rect 61987 9639 62045 9640
rect 2283 9596 2325 9605
rect 2283 9556 2284 9596
rect 2324 9556 2325 9596
rect 2283 9547 2325 9556
rect 10347 9596 10389 9605
rect 10347 9556 10348 9596
rect 10388 9556 10389 9596
rect 10347 9547 10389 9556
rect 39531 9596 39573 9605
rect 39531 9556 39532 9596
rect 39572 9556 39573 9596
rect 39531 9547 39573 9556
rect 59595 9596 59637 9605
rect 59595 9556 59596 9596
rect 59636 9556 59637 9596
rect 59595 9547 59637 9556
rect 2659 9512 2717 9513
rect 2659 9472 2668 9512
rect 2708 9472 2717 9512
rect 2659 9471 2717 9472
rect 3523 9512 3581 9513
rect 3523 9472 3532 9512
rect 3572 9472 3581 9512
rect 3523 9471 3581 9472
rect 6795 9512 6837 9521
rect 6795 9472 6796 9512
rect 6836 9472 6837 9512
rect 6795 9463 6837 9472
rect 7171 9512 7229 9513
rect 7171 9472 7180 9512
rect 7220 9472 7229 9512
rect 7171 9471 7229 9472
rect 8035 9512 8093 9513
rect 8035 9472 8044 9512
rect 8084 9472 8093 9512
rect 8035 9471 8093 9472
rect 10723 9512 10781 9513
rect 10723 9472 10732 9512
rect 10772 9472 10781 9512
rect 10723 9471 10781 9472
rect 11587 9512 11645 9513
rect 11587 9472 11596 9512
rect 11636 9472 11645 9512
rect 11587 9471 11645 9472
rect 20323 9512 20381 9513
rect 20323 9472 20332 9512
rect 20372 9472 20381 9512
rect 20323 9471 20381 9472
rect 21859 9512 21917 9513
rect 21859 9472 21868 9512
rect 21908 9472 21917 9512
rect 21859 9471 21917 9472
rect 33099 9512 33141 9521
rect 33099 9472 33100 9512
rect 33140 9472 33141 9512
rect 33099 9463 33141 9472
rect 33195 9512 33237 9521
rect 33195 9472 33196 9512
rect 33236 9472 33237 9512
rect 33195 9463 33237 9472
rect 33291 9512 33333 9521
rect 33291 9472 33292 9512
rect 33332 9472 33333 9512
rect 33291 9463 33333 9472
rect 34147 9512 34205 9513
rect 34147 9472 34156 9512
rect 34196 9472 34205 9512
rect 34147 9471 34205 9472
rect 36355 9512 36413 9513
rect 36355 9472 36364 9512
rect 36404 9472 36413 9512
rect 36355 9471 36413 9472
rect 38275 9512 38333 9513
rect 38275 9472 38284 9512
rect 38324 9472 38333 9512
rect 38275 9471 38333 9472
rect 39139 9512 39197 9513
rect 39139 9472 39148 9512
rect 39188 9472 39197 9512
rect 39139 9471 39197 9472
rect 46339 9512 46397 9513
rect 46339 9472 46348 9512
rect 46388 9472 46397 9512
rect 46339 9471 46397 9472
rect 47203 9512 47261 9513
rect 47203 9472 47212 9512
rect 47252 9472 47261 9512
rect 47203 9471 47261 9472
rect 47883 9512 47925 9521
rect 47883 9472 47884 9512
rect 47924 9472 47925 9512
rect 47883 9463 47925 9472
rect 48075 9512 48117 9521
rect 48075 9472 48076 9512
rect 48116 9472 48117 9512
rect 48075 9463 48117 9472
rect 48451 9512 48509 9513
rect 48451 9472 48460 9512
rect 48500 9472 48509 9512
rect 48451 9471 48509 9472
rect 49315 9512 49373 9513
rect 49315 9472 49324 9512
rect 49364 9472 49373 9512
rect 49315 9471 49373 9472
rect 53451 9512 53493 9521
rect 53451 9472 53452 9512
rect 53492 9472 53493 9512
rect 53451 9463 53493 9472
rect 55275 9512 55317 9521
rect 55275 9472 55276 9512
rect 55316 9472 55317 9512
rect 55275 9463 55317 9472
rect 55651 9512 55709 9513
rect 55651 9472 55660 9512
rect 55700 9472 55709 9512
rect 55651 9471 55709 9472
rect 56515 9512 56573 9513
rect 56515 9472 56524 9512
rect 56564 9472 56573 9512
rect 56515 9471 56573 9472
rect 59971 9512 60029 9513
rect 59971 9472 59980 9512
rect 60020 9472 60029 9512
rect 59971 9471 60029 9472
rect 60835 9512 60893 9513
rect 60835 9472 60844 9512
rect 60884 9472 60893 9512
rect 60835 9471 60893 9472
rect 54883 9428 54941 9429
rect 54883 9388 54892 9428
rect 54932 9388 54941 9428
rect 54883 9387 54941 9388
rect 59203 9428 59261 9429
rect 59203 9388 59212 9428
rect 59252 9388 59261 9428
rect 59203 9387 59261 9388
rect 37123 9344 37181 9345
rect 37123 9304 37132 9344
rect 37172 9304 37181 9344
rect 37123 9303 37181 9304
rect 22531 9260 22589 9261
rect 22531 9220 22540 9260
rect 22580 9220 22589 9260
rect 22531 9219 22589 9220
rect 35683 9260 35741 9261
rect 35683 9220 35692 9260
rect 35732 9220 35741 9260
rect 35683 9219 35741 9220
rect 53259 9260 53301 9269
rect 53259 9220 53260 9260
rect 53300 9220 53301 9260
rect 53259 9211 53301 9220
rect 54699 9260 54741 9269
rect 54699 9220 54700 9260
rect 54740 9220 54741 9260
rect 54699 9211 54741 9220
rect 57667 9260 57725 9261
rect 57667 9220 57676 9260
rect 57716 9220 57725 9260
rect 57667 9219 57725 9220
rect 576 9092 99360 9116
rect 576 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 18232 9092
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18600 9052 33352 9092
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33720 9052 48472 9092
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48840 9052 63592 9092
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63960 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 93832 9092
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 94200 9052 99360 9092
rect 576 9028 99360 9052
rect 19075 8840 19133 8841
rect 19075 8800 19084 8840
rect 19124 8800 19133 8840
rect 19075 8799 19133 8800
rect 33291 8840 33333 8849
rect 33291 8800 33292 8840
rect 33332 8800 33333 8840
rect 33291 8791 33333 8800
rect 56803 8840 56861 8841
rect 56803 8800 56812 8840
rect 56852 8800 56861 8840
rect 56803 8799 56861 8800
rect 34443 8756 34485 8765
rect 34443 8716 34444 8756
rect 34484 8716 34485 8756
rect 34443 8707 34485 8716
rect 44523 8756 44565 8765
rect 44523 8716 44524 8756
rect 44564 8716 44565 8756
rect 44523 8707 44565 8716
rect 3331 8672 3389 8673
rect 3331 8632 3340 8672
rect 3380 8632 3389 8672
rect 3331 8631 3389 8632
rect 4195 8672 4253 8673
rect 4195 8632 4204 8672
rect 4244 8632 4253 8672
rect 4195 8631 4253 8632
rect 17059 8672 17117 8673
rect 17059 8632 17068 8672
rect 17108 8632 17117 8672
rect 17059 8631 17117 8632
rect 17923 8672 17981 8673
rect 17923 8632 17932 8672
rect 17972 8632 17981 8672
rect 17923 8631 17981 8632
rect 23491 8672 23549 8673
rect 23491 8632 23500 8672
rect 23540 8632 23549 8672
rect 23491 8631 23549 8632
rect 24451 8672 24509 8673
rect 24451 8632 24460 8672
rect 24500 8632 24509 8672
rect 24451 8631 24509 8632
rect 25899 8672 25941 8681
rect 25899 8632 25900 8672
rect 25940 8632 25941 8672
rect 25899 8623 25941 8632
rect 26083 8672 26141 8673
rect 26083 8632 26092 8672
rect 26132 8632 26141 8672
rect 26083 8631 26141 8632
rect 27235 8672 27293 8673
rect 27235 8632 27244 8672
rect 27284 8632 27293 8672
rect 27235 8631 27293 8632
rect 27339 8672 27381 8681
rect 27339 8632 27340 8672
rect 27380 8632 27381 8672
rect 27339 8623 27381 8632
rect 28003 8672 28061 8673
rect 28003 8632 28012 8672
rect 28052 8632 28061 8672
rect 28003 8631 28061 8632
rect 28291 8672 28349 8673
rect 28291 8632 28300 8672
rect 28340 8632 28349 8672
rect 28291 8631 28349 8632
rect 29155 8672 29213 8673
rect 29155 8632 29164 8672
rect 29204 8632 29213 8672
rect 29155 8631 29213 8632
rect 29547 8672 29589 8681
rect 29547 8632 29548 8672
rect 29588 8632 29589 8672
rect 29547 8623 29589 8632
rect 29643 8672 29685 8681
rect 29643 8632 29644 8672
rect 29684 8632 29685 8672
rect 29643 8623 29685 8632
rect 29739 8672 29781 8681
rect 29739 8632 29740 8672
rect 29780 8632 29781 8672
rect 29739 8623 29781 8632
rect 29835 8672 29877 8681
rect 29835 8632 29836 8672
rect 29876 8632 29877 8672
rect 29835 8623 29877 8632
rect 32323 8672 32381 8673
rect 32323 8632 32332 8672
rect 32372 8632 32381 8672
rect 32323 8631 32381 8632
rect 33195 8672 33237 8681
rect 33195 8632 33196 8672
rect 33236 8632 33237 8672
rect 33195 8623 33237 8632
rect 33379 8672 33437 8673
rect 33379 8632 33388 8672
rect 33428 8632 33437 8672
rect 33379 8631 33437 8632
rect 33859 8672 33917 8673
rect 33859 8632 33868 8672
rect 33908 8632 33917 8672
rect 33859 8631 33917 8632
rect 34147 8672 34205 8673
rect 34147 8632 34156 8672
rect 34196 8632 34205 8672
rect 34147 8631 34205 8632
rect 34347 8672 34389 8681
rect 34347 8632 34348 8672
rect 34388 8632 34389 8672
rect 34347 8623 34389 8632
rect 34539 8672 34581 8681
rect 34539 8632 34540 8672
rect 34580 8632 34581 8672
rect 34539 8623 34581 8632
rect 38379 8672 38421 8681
rect 38379 8632 38380 8672
rect 38420 8632 38421 8672
rect 38379 8623 38421 8632
rect 42499 8672 42557 8673
rect 42499 8632 42508 8672
rect 42548 8632 42557 8672
rect 42499 8631 42557 8632
rect 43363 8672 43421 8673
rect 43363 8632 43372 8672
rect 43412 8632 43421 8672
rect 43363 8631 43421 8632
rect 45667 8672 45725 8673
rect 45667 8632 45676 8672
rect 45716 8632 45725 8672
rect 45667 8631 45725 8632
rect 46723 8672 46781 8673
rect 46723 8632 46732 8672
rect 46772 8632 46781 8672
rect 46723 8631 46781 8632
rect 47107 8672 47165 8673
rect 47107 8632 47116 8672
rect 47156 8632 47165 8672
rect 47107 8631 47165 8632
rect 54123 8672 54165 8681
rect 54123 8632 54124 8672
rect 54164 8632 54165 8672
rect 54123 8623 54165 8632
rect 54499 8672 54557 8673
rect 54499 8632 54508 8672
rect 54548 8632 54557 8672
rect 54499 8631 54557 8632
rect 55363 8672 55421 8673
rect 55363 8632 55372 8672
rect 55412 8632 55421 8672
rect 55363 8631 55421 8632
rect 57475 8672 57533 8673
rect 57475 8632 57484 8672
rect 57524 8632 57533 8672
rect 57475 8631 57533 8632
rect 2955 8588 2997 8597
rect 2955 8548 2956 8588
rect 2996 8548 2997 8588
rect 2955 8539 2997 8548
rect 16683 8588 16725 8597
rect 16683 8548 16684 8588
rect 16724 8548 16725 8588
rect 16683 8539 16725 8548
rect 25995 8588 26037 8597
rect 25995 8548 25996 8588
rect 26036 8548 26037 8588
rect 25995 8539 26037 8548
rect 27811 8588 27869 8589
rect 27811 8548 27820 8588
rect 27860 8548 27869 8588
rect 27811 8547 27869 8548
rect 42123 8588 42165 8597
rect 42123 8548 42124 8588
rect 42164 8548 42165 8588
rect 42123 8539 42165 8548
rect 46627 8588 46685 8589
rect 46627 8548 46636 8588
rect 46676 8548 46685 8588
rect 46627 8547 46685 8548
rect 643 8504 701 8505
rect 643 8464 652 8504
rect 692 8464 701 8504
rect 643 8463 701 8464
rect 5347 8504 5405 8505
rect 5347 8464 5356 8504
rect 5396 8464 5405 8504
rect 5347 8463 5405 8464
rect 23979 8504 24021 8513
rect 23979 8464 23980 8504
rect 24020 8464 24021 8504
rect 23979 8455 24021 8464
rect 26955 8504 26997 8513
rect 26955 8464 26956 8504
rect 26996 8464 26997 8504
rect 26955 8455 26997 8464
rect 28483 8504 28541 8505
rect 28483 8464 28492 8504
rect 28532 8464 28541 8504
rect 28483 8463 28541 8464
rect 31651 8504 31709 8505
rect 31651 8464 31660 8504
rect 31700 8464 31709 8504
rect 31651 8463 31709 8464
rect 33675 8504 33717 8513
rect 33675 8464 33676 8504
rect 33716 8464 33717 8504
rect 33675 8455 33717 8464
rect 37995 8504 38037 8513
rect 37995 8464 37996 8504
rect 38036 8464 38037 8504
rect 37995 8455 38037 8464
rect 46339 8504 46397 8505
rect 46339 8464 46348 8504
rect 46388 8464 46397 8504
rect 46339 8463 46397 8464
rect 56515 8504 56573 8505
rect 56515 8464 56524 8504
rect 56564 8464 56573 8504
rect 56515 8463 56573 8464
rect 576 8336 99360 8360
rect 576 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 19472 8336
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19840 8296 34592 8336
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34960 8296 49712 8336
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 50080 8296 64832 8336
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 65200 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 95072 8336
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95440 8296 99360 8336
rect 576 8272 99360 8296
rect 643 8168 701 8169
rect 643 8128 652 8168
rect 692 8128 701 8168
rect 643 8127 701 8128
rect 3723 8168 3765 8177
rect 3723 8128 3724 8168
rect 3764 8128 3765 8168
rect 3723 8119 3765 8128
rect 6123 8168 6165 8177
rect 6123 8128 6124 8168
rect 6164 8128 6165 8168
rect 6123 8119 6165 8128
rect 16483 8168 16541 8169
rect 16483 8128 16492 8168
rect 16532 8128 16541 8168
rect 16483 8127 16541 8128
rect 27619 8168 27677 8169
rect 27619 8128 27628 8168
rect 27668 8128 27677 8168
rect 27619 8127 27677 8128
rect 33099 8168 33141 8177
rect 33099 8128 33100 8168
rect 33140 8128 33141 8168
rect 33099 8119 33141 8128
rect 33963 8168 34005 8177
rect 33963 8128 33964 8168
rect 34004 8128 34005 8168
rect 33963 8119 34005 8128
rect 47499 8168 47541 8177
rect 47499 8128 47500 8168
rect 47540 8128 47541 8168
rect 47499 8119 47541 8128
rect 55563 8168 55605 8177
rect 55563 8128 55564 8168
rect 55604 8128 55605 8168
rect 55563 8119 55605 8128
rect 21963 8084 22005 8093
rect 21963 8044 21964 8084
rect 22004 8044 22005 8084
rect 21963 8035 22005 8044
rect 25315 8084 25373 8085
rect 25315 8044 25324 8084
rect 25364 8044 25373 8084
rect 25315 8043 25373 8044
rect 30027 8084 30069 8093
rect 30027 8044 30028 8084
rect 30068 8044 30069 8084
rect 30027 8035 30069 8044
rect 48555 8084 48597 8093
rect 48555 8044 48556 8084
rect 48596 8044 48597 8084
rect 48555 8035 48597 8044
rect 4395 8000 4437 8009
rect 4395 7960 4396 8000
rect 4436 7960 4437 8000
rect 4395 7951 4437 7960
rect 4491 8000 4533 8009
rect 4491 7960 4492 8000
rect 4532 7960 4533 8000
rect 4491 7951 4533 7960
rect 4579 8000 4637 8001
rect 4579 7960 4588 8000
rect 4628 7960 4637 8000
rect 4579 7959 4637 7960
rect 5443 8000 5501 8001
rect 5443 7960 5452 8000
rect 5492 7960 5501 8000
rect 5443 7959 5501 7960
rect 5635 8000 5693 8001
rect 5635 7960 5644 8000
rect 5684 7960 5693 8000
rect 5635 7959 5693 7960
rect 5923 8000 5981 8001
rect 5923 7960 5932 8000
rect 5972 7960 5981 8000
rect 5923 7959 5981 7960
rect 6595 8000 6653 8001
rect 6595 7960 6604 8000
rect 6644 7960 6653 8000
rect 6595 7959 6653 7960
rect 7555 8000 7613 8001
rect 7555 7960 7564 8000
rect 7604 7960 7613 8000
rect 7555 7959 7613 7960
rect 15811 8000 15869 8001
rect 15811 7960 15820 8000
rect 15860 7960 15869 8000
rect 15811 7959 15869 7960
rect 18123 8000 18165 8009
rect 18123 7960 18124 8000
rect 18164 7960 18165 8000
rect 18123 7951 18165 7960
rect 22339 8000 22397 8001
rect 22339 7960 22348 8000
rect 22388 7960 22397 8000
rect 22339 7959 22397 7960
rect 23203 8000 23261 8001
rect 23203 7960 23212 8000
rect 23252 7960 23261 8000
rect 23203 7959 23261 7960
rect 25411 8000 25469 8001
rect 25411 7960 25420 8000
rect 25460 7960 25469 8000
rect 25411 7959 25469 7960
rect 25795 8000 25853 8001
rect 25795 7960 25804 8000
rect 25844 7960 25853 8000
rect 25795 7959 25853 7960
rect 28771 8000 28829 8001
rect 28771 7960 28780 8000
rect 28820 7960 28829 8000
rect 28771 7959 28829 7960
rect 29635 8000 29693 8001
rect 29635 7960 29644 8000
rect 29684 7960 29693 8000
rect 29635 7959 29693 7960
rect 33379 8000 33437 8001
rect 33379 7960 33388 8000
rect 33428 7960 33437 8000
rect 33379 7959 33437 7960
rect 33483 8000 33525 8009
rect 33483 7960 33484 8000
rect 33524 7960 33525 8000
rect 33483 7951 33525 7960
rect 34051 8000 34109 8001
rect 34051 7960 34060 8000
rect 34100 7960 34109 8000
rect 34051 7959 34109 7960
rect 34435 8000 34493 8001
rect 34435 7960 34444 8000
rect 34484 7960 34493 8000
rect 34435 7959 34493 7960
rect 46531 8000 46589 8001
rect 46531 7960 46540 8000
rect 46580 7960 46589 8000
rect 46531 7959 46589 7960
rect 46635 8000 46677 8009
rect 46635 7960 46636 8000
rect 46676 7960 46677 8000
rect 46635 7951 46677 7960
rect 46731 8000 46773 8009
rect 46731 7960 46732 8000
rect 46772 7960 46773 8000
rect 46731 7951 46773 7960
rect 47115 8000 47157 8009
rect 47115 7960 47116 8000
rect 47156 7960 47157 8000
rect 47115 7951 47157 7960
rect 47203 8000 47261 8001
rect 47203 7960 47212 8000
rect 47252 7960 47261 8000
rect 47203 7959 47261 7960
rect 49219 8000 49277 8001
rect 49219 7960 49228 8000
rect 49268 7960 49277 8000
rect 49219 7959 49277 7960
rect 3907 7916 3965 7917
rect 3907 7876 3916 7916
rect 3956 7876 3965 7916
rect 3907 7875 3965 7876
rect 24363 7916 24405 7925
rect 24363 7876 24364 7916
rect 24404 7876 24405 7916
rect 24363 7867 24405 7876
rect 55747 7916 55805 7917
rect 55747 7876 55756 7916
rect 55796 7876 55805 7916
rect 55747 7875 55805 7876
rect 18699 7832 18741 7841
rect 18699 7792 18700 7832
rect 18740 7792 18741 7832
rect 18699 7783 18741 7792
rect 4771 7748 4829 7749
rect 4771 7708 4780 7748
rect 4820 7708 4829 7748
rect 4771 7707 4829 7708
rect 6891 7748 6933 7757
rect 6891 7708 6892 7748
rect 6932 7708 6933 7748
rect 6891 7699 6933 7708
rect 576 7580 99360 7604
rect 576 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 18232 7580
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18600 7540 33352 7580
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33720 7540 48472 7580
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48840 7540 63592 7580
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63960 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 93832 7580
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 94200 7540 99360 7580
rect 576 7516 99360 7540
rect 11499 7412 11541 7421
rect 11499 7372 11500 7412
rect 11540 7372 11541 7412
rect 11499 7363 11541 7372
rect 14755 7412 14813 7413
rect 14755 7372 14764 7412
rect 14804 7372 14813 7412
rect 14755 7371 14813 7372
rect 25411 7412 25469 7413
rect 25411 7372 25420 7412
rect 25460 7372 25469 7412
rect 25411 7371 25469 7372
rect 33291 7412 33333 7421
rect 33291 7372 33292 7412
rect 33332 7372 33333 7412
rect 33291 7363 33333 7372
rect 34243 7412 34301 7413
rect 34243 7372 34252 7412
rect 34292 7372 34301 7412
rect 34243 7371 34301 7372
rect 49323 7412 49365 7421
rect 49323 7372 49324 7412
rect 49364 7372 49365 7412
rect 49323 7363 49365 7372
rect 50371 7412 50429 7413
rect 50371 7372 50380 7412
rect 50420 7372 50429 7412
rect 50371 7371 50429 7372
rect 56715 7412 56757 7421
rect 56715 7372 56716 7412
rect 56756 7372 56757 7412
rect 56715 7363 56757 7372
rect 38851 7244 38909 7245
rect 38851 7204 38860 7244
rect 38900 7204 38909 7244
rect 38851 7203 38909 7204
rect 39723 7244 39765 7253
rect 39723 7204 39724 7244
rect 39764 7204 39765 7244
rect 39723 7195 39765 7204
rect 11203 7160 11261 7161
rect 11203 7120 11212 7160
rect 11252 7120 11261 7160
rect 11203 7119 11261 7120
rect 12163 7160 12221 7161
rect 12163 7120 12172 7160
rect 12212 7120 12221 7160
rect 12163 7119 12221 7120
rect 12739 7160 12797 7161
rect 12739 7120 12748 7160
rect 12788 7120 12797 7160
rect 12739 7119 12797 7120
rect 13603 7160 13661 7161
rect 13603 7120 13612 7160
rect 13652 7120 13661 7160
rect 13603 7119 13661 7120
rect 23395 7160 23453 7161
rect 23395 7120 23404 7160
rect 23444 7120 23453 7160
rect 23395 7119 23453 7120
rect 24259 7160 24317 7161
rect 24259 7120 24268 7160
rect 24308 7120 24317 7160
rect 24259 7119 24317 7120
rect 33187 7160 33245 7161
rect 33187 7120 33196 7160
rect 33236 7120 33245 7160
rect 33187 7119 33245 7120
rect 33387 7160 33429 7169
rect 33387 7120 33388 7160
rect 33428 7120 33429 7160
rect 33387 7111 33429 7120
rect 33571 7160 33629 7161
rect 33571 7120 33580 7160
rect 33620 7120 33629 7160
rect 33571 7119 33629 7120
rect 40387 7160 40445 7161
rect 40387 7120 40396 7160
rect 40436 7120 40445 7160
rect 40387 7119 40445 7120
rect 49795 7160 49853 7161
rect 49795 7120 49804 7160
rect 49844 7120 49853 7160
rect 49795 7119 49853 7120
rect 51523 7160 51581 7161
rect 51523 7120 51532 7160
rect 51572 7120 51581 7160
rect 51523 7119 51581 7120
rect 52387 7160 52445 7161
rect 52387 7120 52396 7160
rect 52436 7120 52445 7160
rect 52387 7119 52445 7120
rect 56419 7160 56477 7161
rect 56419 7120 56428 7160
rect 56468 7120 56477 7160
rect 56419 7119 56477 7120
rect 12363 7076 12405 7085
rect 12363 7036 12364 7076
rect 12404 7036 12405 7076
rect 12363 7027 12405 7036
rect 23019 7076 23061 7085
rect 23019 7036 23020 7076
rect 23060 7036 23061 7076
rect 23019 7027 23061 7036
rect 48931 7076 48989 7077
rect 48931 7036 48940 7076
rect 48980 7036 48989 7076
rect 48931 7035 48989 7036
rect 52779 7076 52821 7085
rect 52779 7036 52780 7076
rect 52820 7036 52821 7076
rect 52779 7027 52821 7036
rect 643 6992 701 6993
rect 643 6952 652 6992
rect 692 6952 701 6992
rect 643 6951 701 6952
rect 38667 6992 38709 7001
rect 38667 6952 38668 6992
rect 38708 6952 38709 6992
rect 38667 6943 38709 6952
rect 576 6824 99360 6848
rect 576 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 19472 6824
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19840 6784 34592 6824
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34960 6784 49712 6824
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 50080 6784 64832 6824
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 65200 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 95072 6824
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95440 6784 99360 6824
rect 576 6760 99360 6784
rect 12651 6656 12693 6665
rect 12651 6616 12652 6656
rect 12692 6616 12693 6656
rect 12651 6607 12693 6616
rect 33475 6656 33533 6657
rect 33475 6616 33484 6656
rect 33524 6616 33533 6656
rect 33475 6615 33533 6616
rect 40291 6656 40349 6657
rect 40291 6616 40300 6656
rect 40340 6616 40349 6656
rect 40291 6615 40349 6616
rect 40675 6656 40733 6657
rect 40675 6616 40684 6656
rect 40724 6616 40733 6656
rect 40675 6615 40733 6616
rect 40963 6656 41021 6657
rect 40963 6616 40972 6656
rect 41012 6616 41021 6656
rect 40963 6615 41021 6616
rect 46923 6656 46965 6665
rect 46923 6616 46924 6656
rect 46964 6616 46965 6656
rect 46923 6607 46965 6616
rect 37899 6572 37941 6581
rect 37899 6532 37900 6572
rect 37940 6532 37941 6572
rect 37899 6523 37941 6532
rect 9667 6488 9725 6489
rect 9667 6448 9676 6488
rect 9716 6448 9725 6488
rect 9667 6447 9725 6448
rect 12163 6488 12221 6489
rect 12163 6448 12172 6488
rect 12212 6448 12221 6488
rect 12163 6447 12221 6448
rect 13123 6488 13181 6489
rect 13123 6448 13132 6488
rect 13172 6448 13181 6488
rect 13123 6447 13181 6448
rect 19171 6488 19229 6489
rect 19171 6448 19180 6488
rect 19220 6448 19229 6488
rect 19171 6447 19229 6448
rect 34147 6488 34205 6489
rect 34147 6448 34156 6488
rect 34196 6448 34205 6488
rect 34147 6447 34205 6448
rect 34339 6488 34397 6489
rect 34339 6448 34348 6488
rect 34388 6448 34397 6488
rect 34339 6447 34397 6448
rect 35299 6488 35357 6489
rect 35299 6448 35308 6488
rect 35348 6448 35357 6488
rect 35299 6447 35357 6448
rect 38275 6488 38333 6489
rect 38275 6448 38284 6488
rect 38324 6448 38333 6488
rect 38275 6447 38333 6448
rect 39139 6488 39197 6489
rect 39139 6448 39148 6488
rect 39188 6448 39197 6488
rect 39139 6447 39197 6448
rect 40771 6488 40829 6489
rect 40771 6448 40780 6488
rect 40820 6448 40829 6488
rect 40771 6447 40829 6448
rect 46435 6488 46493 6489
rect 46435 6448 46444 6488
rect 46484 6448 46493 6488
rect 46435 6447 46493 6448
rect 46723 6488 46781 6489
rect 46723 6448 46732 6488
rect 46772 6448 46781 6488
rect 46723 6447 46781 6448
rect 17635 6404 17693 6405
rect 17635 6364 17644 6404
rect 17684 6364 17693 6404
rect 17635 6363 17693 6364
rect 10339 6320 10397 6321
rect 10339 6280 10348 6320
rect 10388 6280 10397 6320
rect 10339 6279 10397 6280
rect 18499 6320 18557 6321
rect 18499 6280 18508 6320
rect 18548 6280 18557 6320
rect 18499 6279 18557 6280
rect 17451 6236 17493 6245
rect 17451 6196 17452 6236
rect 17492 6196 17493 6236
rect 17451 6187 17493 6196
rect 576 6068 99360 6092
rect 576 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 18232 6068
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18600 6028 33352 6068
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33720 6028 48472 6068
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48840 6028 63592 6068
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63960 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 93832 6068
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 94200 6028 99360 6068
rect 576 6004 99360 6028
rect 4587 5900 4629 5909
rect 4587 5860 4588 5900
rect 4628 5860 4629 5900
rect 4587 5851 4629 5860
rect 12355 5900 12413 5901
rect 12355 5860 12364 5900
rect 12404 5860 12413 5900
rect 12355 5859 12413 5860
rect 19075 5900 19133 5901
rect 19075 5860 19084 5900
rect 19124 5860 19133 5900
rect 19075 5859 19133 5860
rect 33475 5900 33533 5901
rect 33475 5860 33484 5900
rect 33524 5860 33533 5900
rect 33475 5859 33533 5860
rect 44611 5900 44669 5901
rect 44611 5860 44620 5900
rect 44660 5860 44669 5900
rect 44611 5859 44669 5860
rect 46339 5900 46397 5901
rect 46339 5860 46348 5900
rect 46388 5860 46397 5900
rect 46339 5859 46397 5860
rect 2947 5732 3005 5733
rect 2947 5692 2956 5732
rect 2996 5692 3005 5732
rect 2947 5691 3005 5692
rect 12171 5732 12213 5741
rect 12171 5692 12172 5732
rect 12212 5692 12213 5732
rect 12171 5683 12213 5692
rect 37411 5732 37469 5733
rect 37411 5692 37420 5732
rect 37460 5692 37469 5732
rect 37411 5691 37469 5692
rect 2083 5648 2141 5649
rect 2083 5608 2092 5648
rect 2132 5608 2141 5648
rect 2083 5607 2141 5608
rect 2763 5648 2805 5657
rect 2763 5608 2764 5648
rect 2804 5608 2805 5648
rect 2763 5599 2805 5608
rect 4491 5648 4533 5657
rect 4491 5608 4492 5648
rect 4532 5608 4533 5648
rect 4491 5599 4533 5608
rect 4675 5648 4733 5649
rect 4675 5608 4684 5648
rect 4724 5608 4733 5648
rect 4675 5607 4733 5608
rect 5155 5648 5213 5649
rect 5155 5608 5164 5648
rect 5204 5608 5213 5648
rect 5155 5607 5213 5608
rect 6211 5648 6269 5649
rect 6211 5608 6220 5648
rect 6260 5608 6269 5648
rect 6211 5607 6269 5608
rect 9771 5648 9813 5657
rect 9771 5608 9772 5648
rect 9812 5608 9813 5648
rect 9771 5599 9813 5608
rect 10147 5648 10205 5649
rect 10147 5608 10156 5648
rect 10196 5608 10205 5648
rect 10147 5607 10205 5608
rect 11011 5648 11069 5649
rect 11011 5608 11020 5648
rect 11060 5608 11069 5648
rect 11011 5607 11069 5608
rect 13027 5648 13085 5649
rect 13027 5608 13036 5648
rect 13076 5608 13085 5648
rect 13027 5607 13085 5608
rect 16683 5648 16725 5657
rect 16683 5608 16684 5648
rect 16724 5608 16725 5648
rect 16683 5599 16725 5608
rect 17059 5648 17117 5649
rect 17059 5608 17068 5648
rect 17108 5608 17117 5648
rect 17059 5607 17117 5608
rect 17923 5648 17981 5649
rect 17923 5608 17932 5648
rect 17972 5608 17981 5648
rect 17923 5607 17981 5608
rect 19651 5648 19709 5649
rect 19651 5608 19660 5648
rect 19700 5608 19709 5648
rect 19651 5607 19709 5608
rect 20611 5648 20669 5649
rect 20611 5608 20620 5648
rect 20660 5608 20669 5648
rect 20611 5607 20669 5608
rect 30211 5648 30269 5649
rect 30211 5608 30220 5648
rect 30260 5608 30269 5648
rect 30211 5607 30269 5608
rect 31459 5648 31517 5649
rect 31459 5608 31468 5648
rect 31508 5608 31517 5648
rect 31459 5607 31517 5608
rect 32323 5648 32381 5649
rect 32323 5608 32332 5648
rect 32372 5608 32381 5648
rect 32323 5607 32381 5608
rect 36547 5648 36605 5649
rect 36547 5608 36556 5648
rect 36596 5608 36605 5648
rect 36547 5607 36605 5608
rect 37227 5648 37269 5657
rect 37227 5608 37228 5648
rect 37268 5608 37269 5648
rect 37227 5599 37269 5608
rect 39331 5648 39389 5649
rect 39331 5608 39340 5648
rect 39380 5608 39389 5648
rect 39331 5607 39389 5608
rect 39531 5648 39573 5657
rect 39531 5608 39532 5648
rect 39572 5608 39573 5648
rect 39531 5599 39573 5608
rect 42595 5648 42653 5649
rect 42595 5608 42604 5648
rect 42644 5608 42653 5648
rect 42595 5607 42653 5608
rect 43459 5648 43517 5649
rect 43459 5608 43468 5648
rect 43508 5608 43517 5648
rect 43459 5607 43517 5608
rect 47491 5648 47549 5649
rect 47491 5608 47500 5648
rect 47540 5608 47549 5648
rect 47491 5607 47549 5608
rect 48355 5648 48413 5649
rect 48355 5608 48364 5648
rect 48404 5608 48413 5648
rect 48355 5607 48413 5608
rect 54019 5648 54077 5649
rect 54019 5608 54028 5648
rect 54068 5608 54077 5648
rect 54019 5607 54077 5608
rect 30891 5564 30933 5573
rect 30891 5524 30892 5564
rect 30932 5524 30933 5564
rect 30891 5515 30933 5524
rect 31083 5564 31125 5573
rect 31083 5524 31084 5564
rect 31124 5524 31125 5564
rect 31083 5515 31125 5524
rect 39435 5564 39477 5573
rect 39435 5524 39436 5564
rect 39476 5524 39477 5564
rect 39435 5515 39477 5524
rect 42219 5564 42261 5573
rect 42219 5524 42220 5564
rect 42260 5524 42261 5564
rect 42219 5515 42261 5524
rect 48747 5564 48789 5573
rect 48747 5524 48748 5564
rect 48788 5524 48789 5564
rect 48747 5515 48789 5524
rect 643 5480 701 5481
rect 643 5440 652 5480
rect 692 5440 701 5480
rect 643 5439 701 5440
rect 3147 5480 3189 5489
rect 3147 5440 3148 5480
rect 3188 5440 3189 5480
rect 3147 5431 3189 5440
rect 5059 5480 5117 5481
rect 5059 5440 5068 5480
rect 5108 5440 5117 5480
rect 5059 5439 5117 5440
rect 5347 5480 5405 5481
rect 5347 5440 5356 5480
rect 5396 5440 5405 5480
rect 5347 5439 5405 5440
rect 5539 5480 5597 5481
rect 5539 5440 5548 5480
rect 5588 5440 5597 5480
rect 5539 5439 5597 5440
rect 37611 5480 37653 5489
rect 37611 5440 37612 5480
rect 37652 5440 37653 5480
rect 37611 5431 37653 5440
rect 53347 5480 53405 5481
rect 53347 5440 53356 5480
rect 53396 5440 53405 5480
rect 53347 5439 53405 5440
rect 576 5312 99360 5336
rect 576 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 95072 5312
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95440 5272 99360 5312
rect 576 5248 99360 5272
rect 1315 5144 1373 5145
rect 1315 5104 1324 5144
rect 1364 5104 1373 5144
rect 1315 5103 1373 5104
rect 41547 5144 41589 5153
rect 41547 5104 41548 5144
rect 41588 5104 41589 5144
rect 41547 5095 41589 5104
rect 50083 5144 50141 5145
rect 50083 5104 50092 5144
rect 50132 5104 50141 5144
rect 50083 5103 50141 5104
rect 3723 5060 3765 5069
rect 3723 5020 3724 5060
rect 3764 5020 3765 5060
rect 3723 5011 3765 5020
rect 6987 5060 7029 5069
rect 6987 5020 6988 5060
rect 7028 5020 7029 5060
rect 6987 5011 7029 5020
rect 38379 5060 38421 5069
rect 38379 5020 38380 5060
rect 38420 5020 38421 5060
rect 38379 5011 38421 5020
rect 50371 5060 50429 5061
rect 50371 5020 50380 5060
rect 50420 5020 50429 5060
rect 50371 5019 50429 5020
rect 2467 4976 2525 4977
rect 2467 4936 2476 4976
rect 2516 4936 2525 4976
rect 2467 4935 2525 4936
rect 3331 4976 3389 4977
rect 3331 4936 3340 4976
rect 3380 4936 3389 4976
rect 3331 4935 3389 4936
rect 3915 4976 3957 4985
rect 3915 4936 3916 4976
rect 3956 4936 3957 4976
rect 3915 4927 3957 4936
rect 4291 4976 4349 4977
rect 4291 4936 4300 4976
rect 4340 4936 4349 4976
rect 4291 4935 4349 4936
rect 5155 4976 5213 4977
rect 5155 4936 5164 4976
rect 5204 4936 5213 4976
rect 5155 4935 5213 4936
rect 7363 4976 7421 4977
rect 7363 4936 7372 4976
rect 7412 4936 7421 4976
rect 7363 4935 7421 4936
rect 8227 4976 8285 4977
rect 8227 4936 8236 4976
rect 8276 4936 8285 4976
rect 8227 4935 8285 4936
rect 26851 4976 26909 4977
rect 26851 4936 26860 4976
rect 26900 4936 26909 4976
rect 26851 4935 26909 4936
rect 27531 4976 27573 4985
rect 27531 4936 27532 4976
rect 27572 4936 27573 4976
rect 27531 4927 27573 4936
rect 27723 4976 27765 4985
rect 27723 4936 27724 4976
rect 27764 4936 27765 4976
rect 27723 4927 27765 4936
rect 28099 4976 28157 4977
rect 28099 4936 28108 4976
rect 28148 4936 28157 4976
rect 28099 4935 28157 4936
rect 28963 4976 29021 4977
rect 28963 4936 28972 4976
rect 29012 4936 29021 4976
rect 28963 4935 29021 4936
rect 37123 4976 37181 4977
rect 37123 4936 37132 4976
rect 37172 4936 37181 4976
rect 37123 4935 37181 4936
rect 37987 4976 38045 4977
rect 37987 4936 37996 4976
rect 38036 4936 38045 4976
rect 37987 4935 38045 4936
rect 39907 4976 39965 4977
rect 39907 4936 39916 4976
rect 39956 4936 39965 4976
rect 39907 4935 39965 4936
rect 41059 4976 41117 4977
rect 41059 4936 41068 4976
rect 41108 4936 41117 4976
rect 41059 4935 41117 4936
rect 41347 4976 41405 4977
rect 41347 4936 41356 4976
rect 41396 4936 41405 4976
rect 41347 4935 41405 4936
rect 50179 4976 50237 4977
rect 50179 4936 50188 4976
rect 50228 4936 50237 4976
rect 50179 4935 50237 4936
rect 51915 4976 51957 4985
rect 51915 4936 51916 4976
rect 51956 4936 51957 4976
rect 51915 4927 51957 4936
rect 52291 4976 52349 4977
rect 52291 4936 52300 4976
rect 52340 4936 52349 4976
rect 52291 4935 52349 4936
rect 53155 4976 53213 4977
rect 53155 4936 53164 4976
rect 53204 4936 53213 4976
rect 53155 4935 53213 4936
rect 835 4892 893 4893
rect 835 4852 844 4892
rect 884 4852 893 4892
rect 835 4851 893 4852
rect 6315 4892 6357 4901
rect 6315 4852 6316 4892
rect 6356 4852 6357 4892
rect 6315 4843 6357 4852
rect 9387 4892 9429 4901
rect 9387 4852 9388 4892
rect 9428 4852 9429 4892
rect 9387 4843 9429 4852
rect 30123 4892 30165 4901
rect 30123 4852 30124 4892
rect 30164 4852 30165 4892
rect 30123 4843 30165 4852
rect 35979 4892 36021 4901
rect 35979 4852 35980 4892
rect 36020 4852 36021 4892
rect 35979 4843 36021 4852
rect 39427 4892 39485 4893
rect 39427 4852 39436 4892
rect 39476 4852 39485 4892
rect 39427 4851 39485 4852
rect 54315 4892 54357 4901
rect 54315 4852 54316 4892
rect 54356 4852 54357 4892
rect 54315 4843 54357 4852
rect 651 4808 693 4817
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 40203 4724 40245 4733
rect 40203 4684 40204 4724
rect 40244 4684 40245 4724
rect 40203 4675 40245 4684
rect 576 4556 99360 4580
rect 576 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 93832 4556
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 94200 4516 99360 4556
rect 576 4492 99360 4516
rect 4395 4388 4437 4397
rect 4395 4348 4396 4388
rect 4436 4348 4437 4388
rect 4395 4339 4437 4348
rect 26179 4388 26237 4389
rect 26179 4348 26188 4388
rect 26228 4348 26237 4388
rect 26179 4347 26237 4348
rect 41163 4388 41205 4397
rect 41163 4348 41164 4388
rect 41204 4348 41205 4388
rect 41163 4339 41205 4348
rect 51915 4388 51957 4397
rect 51915 4348 51916 4388
rect 51956 4348 51957 4388
rect 51915 4339 51957 4348
rect 835 4220 893 4221
rect 835 4180 844 4220
rect 884 4180 893 4220
rect 835 4179 893 4180
rect 4579 4220 4637 4221
rect 4579 4180 4588 4220
rect 4628 4180 4637 4220
rect 4579 4179 4637 4180
rect 12931 4220 12989 4221
rect 12931 4180 12940 4220
rect 12980 4180 12989 4220
rect 12931 4179 12989 4180
rect 16971 4220 17013 4229
rect 16971 4180 16972 4220
rect 17012 4180 17013 4220
rect 16971 4171 17013 4180
rect 52099 4220 52157 4221
rect 52099 4180 52108 4220
rect 52148 4180 52157 4220
rect 52099 4179 52157 4180
rect 16291 4136 16349 4137
rect 16291 4096 16300 4136
rect 16340 4096 16349 4136
rect 16291 4095 16349 4096
rect 17635 4136 17693 4137
rect 17635 4096 17644 4136
rect 17684 4096 17693 4136
rect 17635 4095 17693 4096
rect 18691 4136 18749 4137
rect 18691 4096 18700 4136
rect 18740 4096 18749 4136
rect 18691 4095 18749 4096
rect 22915 4136 22973 4137
rect 22915 4096 22924 4136
rect 22964 4096 22973 4136
rect 22915 4095 22973 4096
rect 24163 4136 24221 4137
rect 24163 4096 24172 4136
rect 24212 4096 24221 4136
rect 24163 4095 24221 4096
rect 25027 4136 25085 4137
rect 25027 4096 25036 4136
rect 25076 4096 25085 4136
rect 25027 4095 25085 4096
rect 30979 4136 31037 4137
rect 30979 4096 30988 4136
rect 31028 4096 31037 4136
rect 30979 4095 31037 4096
rect 41059 4136 41117 4137
rect 41059 4096 41068 4136
rect 41108 4096 41117 4136
rect 41059 4095 41117 4096
rect 41259 4136 41301 4145
rect 41259 4096 41260 4136
rect 41300 4096 41301 4136
rect 41259 4087 41301 4096
rect 49219 4136 49277 4137
rect 49219 4096 49228 4136
rect 49268 4096 49277 4136
rect 49219 4095 49277 4096
rect 49603 4136 49661 4137
rect 49603 4096 49612 4136
rect 49652 4096 49661 4136
rect 49603 4095 49661 4096
rect 18027 4052 18069 4061
rect 18027 4012 18028 4052
rect 18068 4012 18069 4052
rect 18027 4003 18069 4012
rect 23595 4052 23637 4061
rect 23595 4012 23596 4052
rect 23636 4012 23637 4052
rect 23595 4003 23637 4012
rect 23787 4052 23829 4061
rect 23787 4012 23788 4052
rect 23828 4012 23829 4052
rect 23787 4003 23829 4012
rect 49123 4052 49181 4053
rect 49123 4012 49132 4052
rect 49172 4012 49181 4052
rect 49123 4011 49181 4012
rect 651 3968 693 3977
rect 651 3928 652 3968
rect 692 3928 693 3968
rect 651 3919 693 3928
rect 12747 3968 12789 3977
rect 12747 3928 12748 3968
rect 12788 3928 12789 3968
rect 17827 3968 17885 3969
rect 12747 3919 12789 3928
rect 17539 3963 17597 3964
rect 17539 3923 17548 3963
rect 17588 3923 17597 3963
rect 17827 3928 17836 3968
rect 17876 3928 17885 3968
rect 17827 3927 17885 3928
rect 31651 3968 31709 3969
rect 31651 3928 31660 3968
rect 31700 3928 31709 3968
rect 31651 3927 31709 3928
rect 17539 3922 17597 3923
rect 576 3800 99360 3824
rect 576 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 95072 3800
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95440 3760 99360 3800
rect 576 3736 99360 3760
rect 14179 3632 14237 3633
rect 14179 3592 14188 3632
rect 14228 3592 14237 3632
rect 14179 3591 14237 3592
rect 18691 3632 18749 3633
rect 18691 3592 18700 3632
rect 18740 3592 18749 3632
rect 18691 3591 18749 3592
rect 21763 3632 21821 3633
rect 21763 3592 21772 3632
rect 21812 3592 21821 3632
rect 21763 3591 21821 3592
rect 40099 3632 40157 3633
rect 40099 3592 40108 3632
rect 40148 3592 40157 3632
rect 40099 3591 40157 3592
rect 41635 3632 41693 3633
rect 41635 3592 41644 3632
rect 41684 3592 41693 3632
rect 41635 3591 41693 3592
rect 49507 3632 49565 3633
rect 49507 3592 49516 3632
rect 49556 3592 49565 3632
rect 49507 3591 49565 3592
rect 11787 3548 11829 3557
rect 11787 3508 11788 3548
rect 11828 3508 11829 3548
rect 11787 3499 11829 3508
rect 19371 3548 19413 3557
rect 19371 3508 19372 3548
rect 19412 3508 19413 3548
rect 19371 3499 19413 3508
rect 49227 3548 49269 3557
rect 49227 3508 49228 3548
rect 49268 3508 49269 3548
rect 49227 3499 49269 3508
rect 50475 3548 50517 3557
rect 50475 3508 50476 3548
rect 50516 3508 50517 3548
rect 50475 3499 50517 3508
rect 50370 3485 50428 3486
rect 12163 3464 12221 3465
rect 12163 3424 12172 3464
rect 12212 3424 12221 3464
rect 12163 3423 12221 3424
rect 13027 3464 13085 3465
rect 13027 3424 13036 3464
rect 13076 3424 13085 3464
rect 13027 3423 13085 3424
rect 16299 3464 16341 3473
rect 16299 3424 16300 3464
rect 16340 3424 16341 3464
rect 16299 3415 16341 3424
rect 16675 3464 16733 3465
rect 16675 3424 16684 3464
rect 16724 3424 16733 3464
rect 16675 3423 16733 3424
rect 17539 3464 17597 3465
rect 17539 3424 17548 3464
rect 17588 3424 17597 3464
rect 17539 3423 17597 3424
rect 19747 3464 19805 3465
rect 19747 3424 19756 3464
rect 19796 3424 19805 3464
rect 19747 3423 19805 3424
rect 20611 3464 20669 3465
rect 20611 3424 20620 3464
rect 20660 3424 20669 3464
rect 20611 3423 20669 3424
rect 31083 3464 31125 3473
rect 31083 3424 31084 3464
rect 31124 3424 31125 3464
rect 31083 3415 31125 3424
rect 31459 3464 31517 3465
rect 31459 3424 31468 3464
rect 31508 3424 31517 3464
rect 31459 3423 31517 3424
rect 32323 3464 32381 3465
rect 32323 3424 32332 3464
rect 32372 3424 32381 3464
rect 32323 3423 32381 3424
rect 33571 3464 33629 3465
rect 33571 3424 33580 3464
rect 33620 3424 33629 3464
rect 33571 3423 33629 3424
rect 40771 3464 40829 3465
rect 40771 3424 40780 3464
rect 40820 3424 40829 3464
rect 40771 3423 40829 3424
rect 40963 3464 41021 3465
rect 40963 3424 40972 3464
rect 41012 3424 41021 3464
rect 40963 3423 41021 3424
rect 45763 3464 45821 3465
rect 45763 3424 45772 3464
rect 45812 3424 45821 3464
rect 45763 3423 45821 3424
rect 46443 3464 46485 3473
rect 46443 3424 46444 3464
rect 46484 3424 46485 3464
rect 46443 3415 46485 3424
rect 49131 3464 49173 3473
rect 49131 3424 49132 3464
rect 49172 3424 49173 3464
rect 49131 3415 49173 3424
rect 49315 3464 49373 3465
rect 49315 3424 49324 3464
rect 49364 3424 49373 3464
rect 49315 3423 49373 3424
rect 50179 3464 50237 3465
rect 50179 3424 50188 3464
rect 50228 3424 50237 3464
rect 50370 3445 50379 3485
rect 50419 3445 50428 3485
rect 50370 3444 50428 3445
rect 50563 3464 50621 3465
rect 50179 3423 50237 3424
rect 50563 3424 50572 3464
rect 50612 3424 50621 3464
rect 50563 3423 50621 3424
rect 54019 3464 54077 3465
rect 54019 3424 54028 3464
rect 54068 3424 54077 3464
rect 54019 3423 54077 3424
rect 835 3380 893 3381
rect 835 3340 844 3380
rect 884 3340 893 3380
rect 835 3339 893 3340
rect 39427 3380 39485 3381
rect 39427 3340 39436 3380
rect 39476 3340 39485 3380
rect 39427 3339 39485 3340
rect 41827 3380 41885 3381
rect 41827 3340 41836 3380
rect 41876 3340 41885 3380
rect 41827 3339 41885 3340
rect 46627 3380 46685 3381
rect 46627 3340 46636 3380
rect 46676 3340 46685 3380
rect 46627 3339 46685 3340
rect 48739 3380 48797 3381
rect 48739 3340 48748 3380
rect 48788 3340 48797 3380
rect 48739 3339 48797 3340
rect 651 3212 693 3221
rect 651 3172 652 3212
rect 692 3172 693 3212
rect 651 3163 693 3172
rect 39243 3212 39285 3221
rect 39243 3172 39244 3212
rect 39284 3172 39285 3212
rect 39243 3163 39285 3172
rect 42027 3212 42069 3221
rect 42027 3172 42028 3212
rect 42068 3172 42069 3212
rect 42027 3163 42069 3172
rect 46827 3212 46869 3221
rect 46827 3172 46828 3212
rect 46868 3172 46869 3212
rect 46827 3163 46869 3172
rect 48555 3212 48597 3221
rect 48555 3172 48556 3212
rect 48596 3172 48597 3212
rect 48555 3163 48597 3172
rect 53347 3212 53405 3213
rect 53347 3172 53356 3212
rect 53396 3172 53405 3212
rect 53347 3171 53405 3172
rect 576 3044 99360 3068
rect 576 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 93832 3044
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 94200 3004 99360 3044
rect 576 2980 99360 3004
rect 16875 2876 16917 2885
rect 16875 2836 16876 2876
rect 16916 2836 16917 2876
rect 16875 2827 16917 2836
rect 18123 2876 18165 2885
rect 18123 2836 18124 2876
rect 18164 2836 18165 2876
rect 18123 2827 18165 2836
rect 30595 2876 30653 2877
rect 30595 2836 30604 2876
rect 30644 2836 30653 2876
rect 30595 2835 30653 2836
rect 40483 2876 40541 2877
rect 40483 2836 40492 2876
rect 40532 2836 40541 2876
rect 40483 2835 40541 2836
rect 40675 2876 40733 2877
rect 40675 2836 40684 2876
rect 40724 2836 40733 2876
rect 40675 2835 40733 2836
rect 44995 2876 45053 2877
rect 44995 2836 45004 2876
rect 45044 2836 45053 2876
rect 44995 2835 45053 2836
rect 49987 2876 50045 2877
rect 49987 2836 49996 2876
rect 50036 2836 50045 2876
rect 49987 2835 50045 2836
rect 54595 2876 54653 2877
rect 54595 2836 54604 2876
rect 54644 2836 54653 2876
rect 54595 2835 54653 2836
rect 17547 2792 17589 2801
rect 17547 2752 17548 2792
rect 17588 2752 17589 2792
rect 17547 2743 17589 2752
rect 52011 2792 52053 2801
rect 52011 2752 52012 2792
rect 52052 2752 52053 2792
rect 52011 2743 52053 2752
rect 835 2708 893 2709
rect 835 2668 844 2708
rect 884 2668 893 2708
rect 835 2667 893 2668
rect 14667 2708 14709 2717
rect 14667 2668 14668 2708
rect 14708 2668 14709 2708
rect 14667 2659 14709 2668
rect 17059 2708 17117 2709
rect 17059 2668 17068 2708
rect 17108 2668 17117 2708
rect 17059 2667 17117 2668
rect 23307 2708 23349 2717
rect 23307 2668 23308 2708
rect 23348 2668 23349 2708
rect 23307 2659 23349 2668
rect 27051 2708 27093 2717
rect 27051 2668 27052 2708
rect 27092 2668 27093 2708
rect 27051 2659 27093 2668
rect 51811 2708 51869 2709
rect 51811 2668 51820 2708
rect 51860 2668 51869 2708
rect 51811 2667 51869 2668
rect 12643 2624 12701 2625
rect 12643 2584 12652 2624
rect 12692 2584 12701 2624
rect 12643 2583 12701 2584
rect 13507 2624 13565 2625
rect 13507 2584 13516 2624
rect 13556 2584 13565 2624
rect 13507 2583 13565 2584
rect 14851 2624 14909 2625
rect 14851 2584 14860 2624
rect 14900 2584 14909 2624
rect 14851 2583 14909 2584
rect 15531 2624 15573 2633
rect 15531 2584 15532 2624
rect 15572 2584 15573 2624
rect 15531 2575 15573 2584
rect 17451 2624 17493 2633
rect 17451 2584 17452 2624
rect 17492 2584 17493 2624
rect 17451 2575 17493 2584
rect 17635 2624 17693 2625
rect 17635 2584 17644 2624
rect 17684 2584 17693 2624
rect 18211 2624 18269 2625
rect 17635 2583 17693 2584
rect 18018 2611 18060 2620
rect 18018 2571 18019 2611
rect 18059 2571 18060 2611
rect 18211 2584 18220 2624
rect 18260 2584 18269 2624
rect 18211 2583 18269 2584
rect 18691 2624 18749 2625
rect 18691 2584 18700 2624
rect 18740 2584 18749 2624
rect 18691 2583 18749 2584
rect 18979 2624 19037 2625
rect 18979 2584 18988 2624
rect 19028 2584 19037 2624
rect 18979 2583 19037 2584
rect 21283 2624 21341 2625
rect 21283 2584 21292 2624
rect 21332 2584 21341 2624
rect 21283 2583 21341 2584
rect 22147 2624 22205 2625
rect 22147 2584 22156 2624
rect 22196 2584 22205 2624
rect 22147 2583 22205 2584
rect 23779 2624 23837 2625
rect 23779 2584 23788 2624
rect 23828 2584 23837 2624
rect 23779 2583 23837 2584
rect 25027 2624 25085 2625
rect 25027 2584 25036 2624
rect 25076 2584 25085 2624
rect 25027 2583 25085 2584
rect 25891 2624 25949 2625
rect 25891 2584 25900 2624
rect 25940 2584 25949 2624
rect 25891 2583 25949 2584
rect 27331 2624 27389 2625
rect 27331 2584 27340 2624
rect 27380 2584 27389 2624
rect 27331 2583 27389 2584
rect 28579 2624 28637 2625
rect 28579 2584 28588 2624
rect 28628 2584 28637 2624
rect 28579 2583 28637 2584
rect 29443 2624 29501 2625
rect 29443 2584 29452 2624
rect 29492 2584 29501 2624
rect 29443 2583 29501 2584
rect 38091 2624 38133 2633
rect 38091 2584 38092 2624
rect 38132 2584 38133 2624
rect 38091 2575 38133 2584
rect 38467 2624 38525 2625
rect 38467 2584 38476 2624
rect 38516 2584 38525 2624
rect 38467 2583 38525 2584
rect 39331 2624 39389 2625
rect 39331 2584 39340 2624
rect 39380 2584 39389 2624
rect 39331 2583 39389 2584
rect 41827 2624 41885 2625
rect 41827 2584 41836 2624
rect 41876 2584 41885 2624
rect 41827 2583 41885 2584
rect 42691 2624 42749 2625
rect 42691 2584 42700 2624
rect 42740 2584 42749 2624
rect 42691 2583 42749 2584
rect 43083 2624 43125 2633
rect 43083 2584 43084 2624
rect 43124 2584 43125 2624
rect 43083 2575 43125 2584
rect 46147 2624 46205 2625
rect 46147 2584 46156 2624
rect 46196 2584 46205 2624
rect 46147 2583 46205 2584
rect 47011 2624 47069 2625
rect 47011 2584 47020 2624
rect 47060 2584 47069 2624
rect 47011 2583 47069 2584
rect 47403 2624 47445 2633
rect 47403 2584 47404 2624
rect 47444 2584 47445 2624
rect 47403 2575 47445 2584
rect 47595 2624 47637 2633
rect 47595 2584 47596 2624
rect 47636 2584 47637 2624
rect 47595 2575 47637 2584
rect 47971 2624 48029 2625
rect 47971 2584 47980 2624
rect 48020 2584 48029 2624
rect 47971 2583 48029 2584
rect 48835 2624 48893 2625
rect 48835 2584 48844 2624
rect 48884 2584 48893 2624
rect 48835 2583 48893 2584
rect 52203 2624 52245 2633
rect 52203 2584 52204 2624
rect 52244 2584 52245 2624
rect 52203 2575 52245 2584
rect 52579 2624 52637 2625
rect 52579 2584 52588 2624
rect 52628 2584 52637 2624
rect 52579 2583 52637 2584
rect 53443 2624 53501 2625
rect 53443 2584 53452 2624
rect 53492 2584 53501 2624
rect 53443 2583 53501 2584
rect 18018 2562 18060 2571
rect 12267 2540 12309 2549
rect 12267 2500 12268 2540
rect 12308 2500 12309 2540
rect 12267 2491 12309 2500
rect 19171 2540 19229 2541
rect 19171 2500 19180 2540
rect 19220 2500 19229 2540
rect 19171 2499 19229 2500
rect 20907 2540 20949 2549
rect 20907 2500 20908 2540
rect 20948 2500 20949 2540
rect 20907 2491 20949 2500
rect 24459 2540 24501 2549
rect 24459 2500 24460 2540
rect 24500 2500 24501 2540
rect 24459 2491 24501 2500
rect 24651 2540 24693 2549
rect 24651 2500 24652 2540
rect 24692 2500 24693 2540
rect 24651 2491 24693 2500
rect 28011 2540 28053 2549
rect 28011 2500 28012 2540
rect 28052 2500 28053 2540
rect 28011 2491 28053 2500
rect 28203 2540 28245 2549
rect 28203 2500 28204 2540
rect 28244 2500 28245 2540
rect 28203 2491 28245 2500
rect 651 2456 693 2465
rect 651 2416 652 2456
rect 692 2416 693 2456
rect 651 2407 693 2416
rect 576 2288 99360 2312
rect 576 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 95072 2288
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95440 2248 99360 2288
rect 576 2224 99360 2248
rect 13323 2120 13365 2129
rect 13323 2080 13324 2120
rect 13364 2080 13365 2120
rect 13323 2071 13365 2080
rect 13507 1868 13565 1869
rect 13507 1828 13516 1868
rect 13556 1828 13565 1868
rect 13507 1827 13565 1828
rect 576 1532 99360 1556
rect 576 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 93832 1532
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 94200 1492 99360 1532
rect 576 1468 99360 1492
rect 576 776 99360 800
rect 576 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 95072 776
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95440 736 99360 776
rect 576 712 99360 736
<< via1 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 37324 38200 37364 38240
rect 36652 37948 36692 37988
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 37612 37612 37652 37652
rect 9484 37444 9524 37484
rect 20716 37444 20756 37484
rect 10348 37360 10388 37400
rect 18700 37360 18740 37400
rect 19564 37360 19604 37400
rect 20908 37360 20948 37400
rect 25420 37360 25460 37400
rect 35596 37360 35636 37400
rect 36460 37360 36500 37400
rect 18316 37276 18356 37316
rect 35212 37276 35252 37316
rect 9292 37192 9332 37232
rect 9676 37192 9716 37232
rect 21580 37192 21620 37232
rect 24748 37192 24788 37232
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 11788 36856 11828 36896
rect 9388 36772 9428 36812
rect 7276 36688 7316 36728
rect 9772 36688 9812 36728
rect 10636 36688 10676 36728
rect 18796 36688 18836 36728
rect 19180 36688 19220 36728
rect 20044 36688 20084 36728
rect 21388 36688 21428 36728
rect 24556 36688 24596 36728
rect 24940 36688 24980 36728
rect 25804 36688 25844 36728
rect 32812 36688 32852 36728
rect 36556 36688 36596 36728
rect 36940 36688 36980 36728
rect 37804 36688 37844 36728
rect 5836 36604 5876 36644
rect 21196 36604 21236 36644
rect 31372 36604 31412 36644
rect 5644 36520 5684 36560
rect 6604 36520 6644 36560
rect 31180 36520 31220 36560
rect 32140 36520 32180 36560
rect 38956 36520 38996 36560
rect 22060 36436 22100 36476
rect 26956 36436 26996 36476
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 7084 36100 7124 36140
rect 19276 36100 19316 36140
rect 19852 36100 19892 36140
rect 25996 36100 26036 36140
rect 32620 36100 32660 36140
rect 35212 36100 35252 36140
rect 36460 36100 36500 36140
rect 19468 35932 19508 35972
rect 20044 35932 20084 35972
rect 23212 35932 23252 35972
rect 35404 35932 35444 35972
rect 36651 35932 36691 35972
rect 36844 35932 36884 35972
rect 4684 35848 4724 35888
rect 5068 35848 5108 35888
rect 5932 35848 5972 35888
rect 9196 35848 9236 35888
rect 9388 35848 9428 35888
rect 9964 35848 10004 35888
rect 10828 35848 10868 35888
rect 22156 35848 22196 35888
rect 22348 35848 22388 35888
rect 23980 35848 24020 35888
rect 24844 35848 24884 35888
rect 26860 35848 26900 35888
rect 30220 35848 30260 35888
rect 30604 35848 30644 35888
rect 31468 35848 31508 35888
rect 36076 35848 36116 35888
rect 36268 35848 36308 35888
rect 37516 35848 37556 35888
rect 9292 35764 9332 35804
rect 9580 35764 9620 35804
rect 22252 35764 22292 35804
rect 23596 35764 23636 35804
rect 36172 35764 36212 35804
rect 11980 35680 12020 35720
rect 23404 35680 23444 35720
rect 26188 35680 26228 35720
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 9484 35344 9524 35384
rect 25228 35344 25268 35384
rect 7372 35260 7412 35300
rect 22156 35260 22196 35300
rect 36268 35260 36308 35300
rect 5836 35176 5876 35216
rect 6508 35176 6548 35216
rect 7276 35176 7316 35216
rect 7468 35176 7508 35216
rect 10348 35176 10388 35216
rect 21292 35176 21332 35216
rect 21484 35176 21524 35216
rect 21676 35176 21716 35216
rect 22060 35176 22100 35216
rect 25324 35176 25364 35216
rect 32908 35176 32948 35216
rect 33100 35176 33140 35216
rect 33196 35176 33236 35216
rect 33292 35176 33332 35216
rect 35788 35176 35828 35216
rect 36172 35176 36212 35216
rect 5068 35092 5108 35132
rect 9292 35092 9332 35132
rect 9676 35092 9716 35132
rect 24844 35092 24884 35132
rect 31468 35092 31508 35132
rect 32236 35092 32276 35132
rect 21388 35008 21428 35048
rect 24652 35008 24692 35048
rect 4876 34924 4916 34964
rect 25516 34924 25556 34964
rect 31276 34924 31316 34964
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 6316 34588 6356 34628
rect 20332 34588 20372 34628
rect 32716 34588 32756 34628
rect 16876 34420 16916 34460
rect 3916 34336 3956 34376
rect 4300 34336 4340 34376
rect 5164 34336 5204 34376
rect 8044 34336 8084 34376
rect 8428 34336 8468 34376
rect 8716 34336 8756 34376
rect 14860 34336 14900 34376
rect 15724 34336 15764 34376
rect 17740 34336 17780 34376
rect 20812 34336 20852 34376
rect 30316 34336 30356 34376
rect 30700 34336 30740 34376
rect 31564 34336 31604 34376
rect 33868 34336 33908 34376
rect 37324 34336 37364 34376
rect 37708 34336 37748 34376
rect 38572 34336 38612 34376
rect 14476 34252 14516 34292
rect 7948 34168 7988 34208
rect 8236 34168 8276 34208
rect 8908 34168 8948 34208
rect 17068 34168 17108 34208
rect 20332 34168 20372 34208
rect 33772 34168 33812 34208
rect 34060 34168 34100 34208
rect 39724 34168 39764 34208
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 10732 33664 10772 33704
rect 11116 33664 11156 33704
rect 12076 33664 12116 33704
rect 14956 33664 14996 33704
rect 15340 33664 15380 33704
rect 16204 33664 16244 33704
rect 17548 33664 17588 33704
rect 24268 33664 24308 33704
rect 24556 33664 24596 33704
rect 47500 33664 47540 33704
rect 17356 33580 17396 33620
rect 11404 33496 11444 33536
rect 18220 33412 18260 33452
rect 25036 33412 25076 33452
rect 46828 33412 46868 33452
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 15436 33076 15476 33116
rect 15916 33076 15956 33116
rect 47788 33076 47828 33116
rect 43372 32992 43412 33032
rect 15628 32908 15668 32948
rect 16108 32908 16148 32948
rect 43564 32908 43604 32948
rect 44332 32908 44372 32948
rect 6508 32824 6548 32864
rect 7468 32824 7508 32864
rect 8812 32824 8852 32864
rect 9196 32824 9236 32864
rect 10060 32824 10100 32864
rect 21772 32824 21812 32864
rect 22156 32824 22196 32864
rect 23020 32824 23060 32864
rect 25612 32824 25652 32864
rect 25996 32824 26036 32864
rect 26860 32824 26900 32864
rect 36940 32824 36980 32864
rect 45004 32824 45044 32864
rect 45772 32824 45812 32864
rect 46636 32824 46676 32864
rect 45388 32740 45428 32780
rect 6988 32656 7028 32696
rect 11212 32656 11252 32696
rect 24172 32656 24212 32696
rect 28012 32656 28052 32696
rect 37612 32656 37652 32696
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 44908 32320 44948 32360
rect 45484 32320 45524 32360
rect 8812 32236 8852 32276
rect 33868 32236 33908 32276
rect 38092 32236 38132 32276
rect 39916 32236 39956 32276
rect 42508 32236 42548 32276
rect 9196 32152 9236 32192
rect 10060 32152 10100 32192
rect 16972 32152 17012 32192
rect 17164 32152 17204 32192
rect 34252 32152 34292 32192
rect 35116 32152 35156 32192
rect 37228 32152 37268 32192
rect 37420 32152 37460 32192
rect 37612 32152 37652 32192
rect 37996 32152 38036 32192
rect 40012 32152 40052 32192
rect 40396 32152 40436 32192
rect 42892 32152 42932 32192
rect 43756 32152 43796 32192
rect 36268 32068 36308 32108
rect 45676 32068 45716 32108
rect 11212 31900 11252 31940
rect 17068 31900 17108 31940
rect 37324 31900 37364 31940
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 38284 31564 38324 31604
rect 22348 31480 22388 31520
rect 33772 31480 33812 31520
rect 37132 31480 37172 31520
rect 38476 31396 38516 31436
rect 3916 31312 3956 31352
rect 4876 31312 4916 31352
rect 11788 31312 11828 31352
rect 22636 31312 22676 31352
rect 23884 31312 23924 31352
rect 24172 31312 24212 31352
rect 27628 31312 27668 31352
rect 31180 31312 31220 31352
rect 33100 31312 33140 31352
rect 34060 31312 34100 31352
rect 36172 31312 36212 31352
rect 36460 31312 36500 31352
rect 37420 31312 37460 31352
rect 37612 31312 37652 31352
rect 38764 31312 38804 31352
rect 38860 31312 38900 31352
rect 44524 31312 44564 31352
rect 11116 31144 11156 31184
rect 24364 31144 24404 31184
rect 26956 31144 26996 31184
rect 30508 31144 30548 31184
rect 35500 31144 35540 31184
rect 44332 31144 44372 31184
rect 44620 31144 44660 31184
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 18220 30808 18260 30848
rect 22540 30808 22580 30848
rect 30412 30808 30452 30848
rect 34636 30808 34676 30848
rect 35980 30808 36020 30848
rect 39436 30808 39476 30848
rect 17932 30724 17972 30764
rect 20140 30724 20180 30764
rect 32812 30724 32852 30764
rect 41836 30724 41876 30764
rect 45484 30724 45524 30764
rect 2860 30640 2900 30680
rect 3244 30640 3284 30680
rect 4108 30640 4148 30680
rect 6124 30640 6164 30680
rect 16204 30640 16244 30680
rect 16876 30640 16916 30680
rect 17068 30640 17108 30680
rect 17260 30640 17300 30680
rect 17452 30640 17492 30680
rect 17740 30640 17780 30680
rect 18316 30640 18356 30680
rect 20524 30640 20564 30680
rect 21388 30640 21428 30680
rect 24268 30640 24308 30680
rect 24940 30640 24980 30680
rect 25132 30640 25172 30680
rect 25228 30640 25268 30680
rect 25324 30640 25364 30680
rect 25708 30640 25748 30680
rect 25804 30640 25844 30680
rect 26764 30640 26804 30680
rect 31564 30640 31604 30680
rect 32428 30640 32468 30680
rect 34156 30640 34196 30680
rect 35116 30640 35156 30680
rect 35788 30640 35828 30680
rect 37132 30640 37172 30680
rect 37996 30640 38036 30680
rect 38380 30640 38420 30680
rect 40588 30640 40628 30680
rect 41452 30640 41492 30680
rect 45004 30640 45044 30680
rect 45388 30640 45428 30680
rect 46444 30640 46484 30680
rect 46540 30640 46580 30680
rect 46636 30640 46676 30680
rect 49228 30640 49268 30680
rect 5260 30556 5300 30596
rect 15436 30556 15476 30596
rect 26092 30556 26132 30596
rect 47500 30556 47540 30596
rect 48556 30556 48596 30596
rect 17164 30472 17204 30512
rect 5452 30388 5492 30428
rect 15244 30388 15284 30428
rect 18508 30388 18548 30428
rect 27436 30388 27476 30428
rect 47308 30388 47348 30428
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 3916 30052 3956 30092
rect 9676 30052 9716 30092
rect 16780 30052 16820 30092
rect 17260 30052 17300 30092
rect 23212 30052 23252 30092
rect 44908 30052 44948 30092
rect 49324 30052 49364 30092
rect 45580 29968 45620 30008
rect 3724 29884 3764 29924
rect 4108 29884 4148 29924
rect 4588 29884 4628 29924
rect 29740 29884 29780 29924
rect 5260 29800 5300 29840
rect 10156 29800 10196 29840
rect 10540 29800 10580 29840
rect 10924 29800 10964 29840
rect 14380 29800 14420 29840
rect 14764 29800 14804 29840
rect 15628 29800 15668 29840
rect 17932 29800 17972 29840
rect 20812 29800 20852 29840
rect 21196 29800 21236 29840
rect 22060 29800 22100 29840
rect 25324 29800 25364 29840
rect 25612 29800 25652 29840
rect 26092 29800 26132 29840
rect 27052 29800 27092 29840
rect 27340 29800 27380 29840
rect 27724 29800 27764 29840
rect 28588 29800 28628 29840
rect 30028 29800 30068 29840
rect 30412 29800 30452 29840
rect 39628 29800 39668 29840
rect 44524 29800 44564 29840
rect 44812 29800 44852 29840
rect 45004 29800 45044 29840
rect 45292 29800 45332 29840
rect 46924 29800 46964 29840
rect 47308 29800 47348 29840
rect 48172 29800 48212 29840
rect 3532 29632 3572 29672
rect 11020 29632 11060 29672
rect 25804 29632 25844 29672
rect 30508 29632 30548 29672
rect 40300 29632 40340 29672
rect 45772 29632 45812 29672
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 5164 29296 5204 29336
rect 10252 29296 10292 29336
rect 15052 29296 15092 29336
rect 17836 29296 17876 29336
rect 44812 29296 44852 29336
rect 2764 29212 2804 29252
rect 3148 29128 3188 29168
rect 4012 29128 4052 29168
rect 7852 29128 7892 29168
rect 8236 29128 8276 29168
rect 9100 29128 9140 29168
rect 11884 29128 11924 29168
rect 15436 29128 15476 29168
rect 15820 29128 15860 29168
rect 16684 29128 16724 29168
rect 22156 29128 22196 29168
rect 23116 29128 23156 29168
rect 26092 29128 26132 29168
rect 30604 29128 30644 29168
rect 39916 29128 39956 29168
rect 40876 29128 40916 29168
rect 45484 29128 45524 29168
rect 15244 29044 15284 29084
rect 44620 29044 44660 29084
rect 22636 28960 22676 29000
rect 40396 28960 40436 29000
rect 11212 28876 11252 28916
rect 26764 28876 26804 28916
rect 29932 28876 29972 28916
rect 44428 28876 44468 28916
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 16204 28540 16244 28580
rect 40492 28540 40532 28580
rect 46924 28540 46964 28580
rect 19948 28456 19988 28496
rect 40300 28456 40340 28496
rect 16396 28372 16436 28412
rect 19276 28372 19316 28412
rect 28780 28372 28820 28412
rect 19660 28288 19700 28328
rect 20620 28288 20660 28328
rect 27148 28288 27188 28328
rect 29068 28288 29108 28328
rect 29164 28288 29204 28328
rect 32908 28288 32948 28328
rect 33868 28288 33908 28328
rect 40972 28288 41012 28328
rect 44524 28288 44564 28328
rect 44908 28288 44948 28328
rect 45772 28288 45812 28328
rect 26476 28120 26516 28160
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 4972 27784 5012 27824
rect 4300 27700 4340 27740
rect 4684 27700 4724 27740
rect 5932 27700 5972 27740
rect 26188 27700 26228 27740
rect 4204 27616 4244 27656
rect 4396 27616 4436 27656
rect 4588 27616 4628 27656
rect 4780 27616 4820 27656
rect 5068 27616 5108 27656
rect 5452 27616 5492 27656
rect 5740 27616 5780 27656
rect 9772 27616 9812 27656
rect 11116 27616 11156 27656
rect 11212 27616 11252 27656
rect 11596 27616 11636 27656
rect 26572 27616 26612 27656
rect 27436 27616 27476 27656
rect 28780 27616 28820 27656
rect 33676 27616 33716 27656
rect 34540 27616 34580 27656
rect 34924 27616 34964 27656
rect 39628 27616 39668 27656
rect 40492 27616 40532 27656
rect 40876 27616 40916 27656
rect 11404 27532 11444 27572
rect 28588 27532 28628 27572
rect 5260 27364 5300 27404
rect 9484 27364 9524 27404
rect 12268 27364 12308 27404
rect 29452 27364 29492 27404
rect 32524 27364 32564 27404
rect 38476 27364 38516 27404
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 4204 27028 4244 27068
rect 5068 27028 5108 27068
rect 11116 27028 11156 27068
rect 28780 27028 28820 27068
rect 3436 26860 3476 26900
rect 3820 26860 3860 26900
rect 42700 26860 42740 26900
rect 4876 26776 4916 26816
rect 5740 26776 5780 26816
rect 10156 26776 10196 26816
rect 11020 26776 11060 26816
rect 11212 26776 11252 26816
rect 28684 26776 28724 26816
rect 28876 26776 28916 26816
rect 33196 26776 33236 26816
rect 34444 26776 34484 26816
rect 35308 26776 35348 26816
rect 40684 26776 40724 26816
rect 41548 26776 41588 26816
rect 42892 26776 42932 26816
rect 34060 26692 34100 26732
rect 40300 26692 40340 26732
rect 3244 26608 3284 26648
rect 3628 26608 3668 26648
rect 10828 26608 10868 26648
rect 33868 26608 33908 26648
rect 36460 26608 36500 26648
rect 43564 26608 43604 26648
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 4876 26272 4916 26312
rect 9484 26272 9524 26312
rect 33580 26272 33620 26312
rect 34060 26272 34100 26312
rect 41452 26272 41492 26312
rect 43948 26272 43988 26312
rect 2476 26188 2516 26228
rect 7084 26188 7124 26228
rect 10540 26188 10580 26228
rect 11692 26188 11732 26228
rect 23980 26188 24020 26228
rect 28684 26188 28724 26228
rect 2860 26104 2900 26144
rect 3724 26104 3764 26144
rect 7468 26104 7508 26144
rect 8332 26104 8372 26144
rect 10060 26104 10100 26144
rect 10444 26104 10484 26144
rect 10828 26104 10868 26144
rect 12076 26104 12116 26144
rect 12940 26104 12980 26144
rect 17836 26104 17876 26144
rect 18508 26104 18548 26144
rect 18700 26104 18740 26144
rect 19084 26104 19124 26144
rect 19948 26104 19988 26144
rect 22732 26104 22772 26144
rect 23596 26104 23636 26144
rect 28396 26104 28436 26144
rect 28780 26104 28820 26144
rect 29164 26104 29204 26144
rect 35116 26104 35156 26144
rect 35596 26104 35636 26144
rect 36556 26104 36596 26144
rect 44428 26104 44468 26144
rect 47020 26104 47060 26144
rect 33388 26020 33428 26060
rect 34252 26020 34292 26060
rect 41644 26020 41684 26060
rect 11500 25852 11540 25892
rect 14092 25852 14132 25892
rect 21100 25852 21140 25892
rect 21580 25852 21620 25892
rect 27724 25852 27764 25892
rect 34444 25852 34484 25892
rect 46348 25852 46388 25892
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 4780 25516 4820 25556
rect 6124 25516 6164 25556
rect 16876 25516 16916 25556
rect 28972 25516 29012 25556
rect 47596 25516 47636 25556
rect 24556 25432 24596 25472
rect 2380 25264 2420 25304
rect 2764 25264 2804 25304
rect 3628 25264 3668 25304
rect 5836 25264 5876 25304
rect 6796 25264 6836 25304
rect 11404 25264 11444 25304
rect 11788 25264 11828 25304
rect 12652 25264 12692 25304
rect 16588 25264 16628 25304
rect 16684 25264 16724 25304
rect 21772 25264 21812 25304
rect 22060 25264 22100 25304
rect 24268 25264 24308 25304
rect 28780 25264 28820 25304
rect 29644 25264 29684 25304
rect 45580 25264 45620 25304
rect 46444 25264 46484 25304
rect 25132 25180 25172 25220
rect 45196 25180 45236 25220
rect 13804 25096 13844 25136
rect 22252 25096 22292 25136
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 16588 24760 16628 24800
rect 45100 24760 45140 24800
rect 12748 24676 12788 24716
rect 16972 24676 17012 24716
rect 22924 24676 22964 24716
rect 27148 24676 27188 24716
rect 11884 24592 11924 24632
rect 15244 24592 15284 24632
rect 16108 24592 16148 24632
rect 16396 24592 16436 24632
rect 16876 24592 16916 24632
rect 17068 24592 17108 24632
rect 20908 24592 20948 24632
rect 21100 24592 21140 24632
rect 23596 24592 23636 24632
rect 25900 24592 25940 24632
rect 26764 24592 26804 24632
rect 33868 24592 33908 24632
rect 34060 24592 34100 24632
rect 35116 24592 35156 24632
rect 43372 24592 43412 24632
rect 43564 24592 43604 24632
rect 46156 24592 46196 24632
rect 46540 24592 46580 24632
rect 46924 24592 46964 24632
rect 47788 24592 47828 24632
rect 24748 24508 24788 24548
rect 31468 24508 31508 24548
rect 44908 24508 44948 24548
rect 12172 24424 12212 24464
rect 15916 24424 15956 24464
rect 21004 24340 21044 24380
rect 31276 24340 31316 24380
rect 33964 24340 34004 24380
rect 34924 24340 34964 24380
rect 43468 24340 43508 24380
rect 45964 24340 46004 24380
rect 48940 24340 48980 24380
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 16876 24004 16916 24044
rect 46348 24004 46388 24044
rect 21484 23920 21524 23960
rect 20332 23836 20372 23876
rect 46156 23836 46196 23876
rect 47692 23836 47732 23876
rect 15436 23752 15476 23792
rect 15820 23752 15860 23792
rect 16204 23752 16244 23792
rect 17068 23752 17108 23792
rect 18316 23752 18356 23792
rect 19180 23752 19220 23792
rect 20812 23752 20852 23792
rect 21964 23752 22004 23792
rect 22060 23752 22100 23792
rect 30220 23752 30260 23792
rect 30604 23752 30644 23792
rect 31468 23752 31508 23792
rect 34828 23752 34868 23792
rect 34924 23752 34964 23792
rect 35020 23752 35060 23792
rect 35212 23752 35252 23792
rect 35500 23752 35540 23792
rect 39916 23752 39956 23792
rect 42028 23752 42068 23792
rect 42892 23752 42932 23792
rect 43468 23752 43508 23792
rect 43852 23752 43892 23792
rect 45484 23752 45524 23792
rect 45580 23752 45620 23792
rect 45676 23752 45716 23792
rect 48364 23752 48404 23792
rect 15916 23668 15956 23708
rect 17740 23668 17780 23708
rect 17932 23668 17972 23708
rect 43276 23668 43316 23708
rect 21676 23584 21716 23624
rect 32620 23584 32660 23624
rect 35692 23584 35732 23624
rect 40588 23584 40628 23624
rect 40876 23584 40916 23624
rect 43948 23584 43988 23624
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 34444 23248 34484 23288
rect 39244 23248 39284 23288
rect 20716 23164 20756 23204
rect 36844 23164 36884 23204
rect 40300 23164 40340 23204
rect 2092 23080 2132 23120
rect 6124 23080 6164 23120
rect 20908 23080 20948 23120
rect 21196 23080 21236 23120
rect 28204 23080 28244 23120
rect 33772 23080 33812 23120
rect 37228 23080 37268 23120
rect 38092 23080 38132 23120
rect 40492 23080 40532 23120
rect 40780 23080 40820 23120
rect 2956 22996 2996 23036
rect 4492 22996 4532 23036
rect 2764 22828 2804 22868
rect 3148 22828 3188 22868
rect 4300 22828 4340 22868
rect 5452 22828 5492 22868
rect 27532 22828 27572 22868
rect 34444 22828 34484 22868
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 1228 22492 1268 22532
rect 6220 22492 6260 22532
rect 16012 22492 16052 22532
rect 28108 22492 28148 22532
rect 49612 22492 49652 22532
rect 652 22408 692 22448
rect 34252 22408 34292 22448
rect 33484 22324 33524 22364
rect 2380 22240 2420 22280
rect 3244 22240 3284 22280
rect 3628 22240 3668 22280
rect 3820 22240 3860 22280
rect 4204 22240 4244 22280
rect 5068 22240 5108 22280
rect 9964 22240 10004 22280
rect 13996 22240 14036 22280
rect 14860 22240 14900 22280
rect 21964 22240 22004 22280
rect 26092 22240 26132 22280
rect 26956 22240 26996 22280
rect 34924 22240 34964 22280
rect 35212 22240 35252 22280
rect 41068 22240 41108 22280
rect 45004 22240 45044 22280
rect 49324 22240 49364 22280
rect 50284 22240 50324 22280
rect 13612 22156 13652 22196
rect 25708 22156 25748 22196
rect 9484 22072 9524 22112
rect 21292 22072 21332 22112
rect 33292 22072 33332 22112
rect 35116 22072 35156 22112
rect 35404 22072 35444 22112
rect 40396 22072 40436 22112
rect 44908 22072 44948 22112
rect 45196 22072 45236 22112
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 13708 21736 13748 21776
rect 34828 21736 34868 21776
rect 32428 21652 32468 21692
rect 36268 21652 36308 21692
rect 4492 21568 4532 21608
rect 4684 21568 4724 21608
rect 8044 21568 8084 21608
rect 8428 21568 8468 21608
rect 9292 21568 9332 21608
rect 11020 21568 11060 21608
rect 13036 21568 13076 21608
rect 14764 21568 14804 21608
rect 15724 21568 15764 21608
rect 21004 21568 21044 21608
rect 25804 21568 25844 21608
rect 26188 21568 26228 21608
rect 27052 21568 27092 21608
rect 29068 21568 29108 21608
rect 31180 21568 31220 21608
rect 32140 21568 32180 21608
rect 32812 21568 32852 21608
rect 33676 21568 33716 21608
rect 36652 21568 36692 21608
rect 37516 21568 37556 21608
rect 38956 21568 38996 21608
rect 43084 21568 43124 21608
rect 44044 21568 44084 21608
rect 44428 21568 44468 21608
rect 44812 21568 44852 21608
rect 45676 21568 45716 21608
rect 10444 21484 10484 21524
rect 28204 21484 28244 21524
rect 38668 21484 38708 21524
rect 15244 21400 15284 21440
rect 31468 21400 31508 21440
rect 43756 21400 43796 21440
rect 4588 21316 4628 21356
rect 11692 21316 11732 21356
rect 20332 21316 20372 21356
rect 28396 21316 28436 21356
rect 39628 21316 39668 21356
rect 46828 21316 46868 21356
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 5836 20980 5876 21020
rect 16012 20980 16052 21020
rect 20044 20980 20084 21020
rect 26476 20980 26516 21020
rect 26860 20980 26900 21020
rect 652 20896 692 20936
rect 26668 20812 26708 20852
rect 27052 20812 27092 20852
rect 52684 20812 52724 20852
rect 5644 20728 5684 20768
rect 11404 20728 11444 20768
rect 11596 20728 11636 20768
rect 11788 20728 11828 20768
rect 12172 20728 12212 20768
rect 12748 20728 12788 20768
rect 13996 20728 14036 20768
rect 14860 20728 14900 20768
rect 20524 20728 20564 20768
rect 21004 20728 21044 20768
rect 21964 20728 22004 20768
rect 39724 20728 39764 20768
rect 39820 20728 39860 20768
rect 39916 20728 39956 20768
rect 40396 20728 40436 20768
rect 40492 20728 40532 20768
rect 45580 20728 45620 20768
rect 46444 20728 46484 20768
rect 46828 20728 46868 20768
rect 11500 20644 11540 20684
rect 12268 20644 12308 20684
rect 13420 20644 13460 20684
rect 13612 20644 13652 20684
rect 5548 20560 5588 20600
rect 40684 20560 40724 20600
rect 44428 20560 44468 20600
rect 52492 20560 52532 20600
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 5356 20140 5396 20180
rect 28396 20140 28436 20180
rect 32044 20140 32084 20180
rect 39148 20140 39188 20180
rect 46060 20140 46100 20180
rect 52108 20140 52148 20180
rect 4492 20056 4532 20096
rect 4684 20056 4724 20096
rect 4876 20056 4916 20096
rect 5164 20056 5204 20096
rect 12076 20056 12116 20096
rect 12172 20056 12212 20096
rect 20620 20056 20660 20096
rect 21004 20056 21044 20096
rect 21388 20056 21428 20096
rect 22252 20056 22292 20096
rect 27916 20056 27956 20096
rect 28108 20056 28148 20096
rect 28300 20056 28340 20096
rect 28492 20056 28532 20096
rect 31180 20056 31220 20096
rect 32428 20056 32468 20096
rect 38668 20056 38708 20096
rect 38956 20056 38996 20096
rect 40108 20056 40148 20096
rect 40780 20056 40820 20096
rect 46732 20056 46772 20096
rect 52492 20056 52532 20096
rect 53356 20056 53396 20096
rect 57484 20056 57524 20096
rect 4588 19972 4628 20012
rect 12460 19972 12500 20012
rect 45004 19972 45044 20012
rect 652 19888 692 19928
rect 44812 19888 44852 19928
rect 20428 19804 20468 19844
rect 23404 19804 23444 19844
rect 28012 19804 28052 19844
rect 31660 19804 31700 19844
rect 33100 19804 33140 19844
rect 39436 19804 39476 19844
rect 41452 19804 41492 19844
rect 54508 19804 54548 19844
rect 56812 19804 56852 19844
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 3724 19468 3764 19508
rect 12172 19468 12212 19508
rect 35404 19468 35444 19508
rect 58060 19468 58100 19508
rect 652 19384 692 19424
rect 3148 19300 3188 19340
rect 5260 19300 5300 19340
rect 55276 19300 55316 19340
rect 3436 19216 3476 19256
rect 4396 19216 4436 19256
rect 4588 19216 4628 19256
rect 7372 19216 7412 19256
rect 7756 19216 7796 19256
rect 8620 19216 8660 19256
rect 12844 19216 12884 19256
rect 19948 19216 19988 19256
rect 20332 19216 20372 19256
rect 21196 19216 21236 19256
rect 22444 19216 22484 19256
rect 28876 19216 28916 19256
rect 29164 19216 29204 19256
rect 31468 19216 31508 19256
rect 32332 19216 32372 19256
rect 35020 19216 35060 19256
rect 35884 19216 35924 19256
rect 54220 19216 54260 19256
rect 56044 19216 56084 19256
rect 56908 19216 56948 19256
rect 29356 19132 29396 19172
rect 31084 19132 31124 19172
rect 55660 19132 55700 19172
rect 2956 19048 2996 19088
rect 9772 19048 9812 19088
rect 33484 19048 33524 19088
rect 53548 19048 53588 19088
rect 55468 19048 55508 19088
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 4684 18712 4724 18752
rect 11212 18712 11252 18752
rect 2284 18628 2324 18668
rect 39436 18628 39476 18668
rect 43084 18628 43124 18668
rect 2668 18544 2708 18584
rect 3532 18544 3572 18584
rect 10732 18544 10772 18584
rect 11020 18544 11060 18584
rect 28300 18544 28340 18584
rect 34060 18544 34100 18584
rect 38188 18544 38228 18584
rect 39052 18544 39092 18584
rect 41836 18544 41876 18584
rect 42700 18544 42740 18584
rect 48748 18544 48788 18584
rect 49132 18544 49172 18584
rect 49996 18544 50036 18584
rect 51340 18544 51380 18584
rect 55180 18544 55220 18584
rect 55372 18544 55412 18584
rect 26860 18460 26900 18500
rect 27244 18460 27284 18500
rect 51148 18460 51188 18500
rect 652 18376 692 18416
rect 26668 18292 26708 18332
rect 27052 18292 27092 18332
rect 27628 18292 27668 18332
rect 33388 18292 33428 18332
rect 37036 18292 37076 18332
rect 40684 18292 40724 18332
rect 52012 18292 52052 18332
rect 55276 18292 55316 18332
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 11020 17956 11060 17996
rect 28108 17956 28148 17996
rect 28972 17956 29012 17996
rect 49324 17956 49364 17996
rect 652 17872 692 17912
rect 15820 17872 15860 17912
rect 48844 17872 48884 17912
rect 16012 17788 16052 17828
rect 49036 17788 49076 17828
rect 49516 17788 49556 17828
rect 2572 17704 2612 17744
rect 3436 17704 3476 17744
rect 9004 17704 9044 17744
rect 9868 17704 9908 17744
rect 17452 17704 17492 17744
rect 25708 17704 25748 17744
rect 26092 17704 26132 17744
rect 26956 17704 26996 17744
rect 28300 17704 28340 17744
rect 29260 17704 29300 17744
rect 37900 17704 37940 17744
rect 42700 17704 42740 17744
rect 43564 17704 43604 17744
rect 49708 17704 49748 17744
rect 50380 17671 50420 17711
rect 51148 17704 51188 17744
rect 51340 17704 51380 17744
rect 52396 17704 52436 17744
rect 55180 17704 55220 17744
rect 55468 17704 55508 17744
rect 2188 17620 2228 17660
rect 8620 17620 8660 17660
rect 16780 17620 16820 17660
rect 51244 17620 51284 17660
rect 4588 17536 4628 17576
rect 29164 17536 29204 17576
rect 29452 17536 29492 17576
rect 38572 17536 38612 17576
rect 52300 17536 52340 17576
rect 52588 17536 52628 17576
rect 55660 17536 55700 17576
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 3052 17200 3092 17240
rect 4012 17200 4052 17240
rect 11980 17200 12020 17240
rect 17260 17200 17300 17240
rect 28588 17200 28628 17240
rect 50188 17200 50228 17240
rect 14860 17116 14900 17156
rect 21292 17116 21332 17156
rect 26188 17116 26228 17156
rect 33196 17116 33236 17156
rect 40876 17116 40916 17156
rect 47788 17116 47828 17156
rect 52780 17116 52820 17156
rect 56620 17116 56660 17156
rect 4684 17032 4724 17072
rect 9580 17032 9620 17072
rect 9964 17032 10004 17072
rect 10828 17032 10868 17072
rect 15244 17032 15284 17072
rect 16108 17032 16148 17072
rect 20140 17032 20180 17072
rect 20428 17032 20468 17072
rect 23404 17032 23444 17072
rect 26572 17032 26612 17072
rect 27436 17032 27476 17072
rect 32716 17032 32756 17072
rect 33100 17032 33140 17072
rect 33772 17032 33812 17072
rect 35404 17032 35444 17072
rect 36076 17032 36116 17072
rect 36268 17032 36308 17072
rect 36652 17032 36692 17072
rect 37516 17032 37556 17072
rect 40396 17032 40436 17072
rect 40684 17032 40724 17072
rect 45100 17032 45140 17072
rect 46060 17032 46100 17072
rect 48172 17032 48212 17072
rect 49036 17032 49076 17072
rect 53164 17032 53204 17072
rect 54028 17032 54068 17072
rect 57004 17032 57044 17072
rect 57868 17032 57908 17072
rect 3244 16948 3284 16988
rect 38668 16948 38708 16988
rect 652 16864 692 16904
rect 19468 16780 19508 16820
rect 20716 16780 20756 16820
rect 24076 16780 24116 16820
rect 34444 16780 34484 16820
rect 55180 16780 55220 16820
rect 59020 16780 59060 16820
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 10732 16444 10772 16484
rect 652 16360 692 16400
rect 21292 16360 21332 16400
rect 46540 16360 46580 16400
rect 16972 16276 17012 16316
rect 18508 16276 18548 16316
rect 34348 16276 34388 16316
rect 10252 16192 10292 16232
rect 14956 16192 14996 16232
rect 15820 16192 15860 16232
rect 17164 16192 17204 16232
rect 19276 16192 19316 16232
rect 20140 16192 20180 16232
rect 31084 16192 31124 16232
rect 31468 16192 31508 16232
rect 32332 16192 32372 16232
rect 34060 16192 34100 16232
rect 34156 16192 34196 16232
rect 41452 16192 41492 16232
rect 45964 16192 46004 16232
rect 56044 16192 56084 16232
rect 14572 16108 14612 16148
rect 18892 16108 18932 16148
rect 10732 16024 10772 16064
rect 17836 16024 17876 16064
rect 18700 16024 18740 16064
rect 33484 16024 33524 16064
rect 42124 16024 42164 16064
rect 46348 16024 46388 16064
rect 55372 16024 55412 16064
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 652 15688 692 15728
rect 15628 15688 15668 15728
rect 19948 15688 19988 15728
rect 27724 15688 27764 15728
rect 39340 15688 39380 15728
rect 40972 15688 41012 15728
rect 18700 15604 18740 15644
rect 25324 15604 25364 15644
rect 41740 15604 41780 15644
rect 16012 15520 16052 15560
rect 16972 15520 17012 15560
rect 17452 15520 17492 15560
rect 17644 15520 17684 15560
rect 17836 15520 17876 15560
rect 18028 15520 18068 15560
rect 18220 15520 18260 15560
rect 18508 15520 18548 15560
rect 20044 15520 20084 15560
rect 20428 15520 20468 15560
rect 22924 15520 22964 15560
rect 25708 15520 25748 15560
rect 26572 15520 26612 15560
rect 33484 15520 33524 15560
rect 33580 15520 33620 15560
rect 33676 15520 33716 15560
rect 33868 15520 33908 15560
rect 38668 15520 38708 15560
rect 39532 15520 39572 15560
rect 39628 15520 39668 15560
rect 39724 15520 39764 15560
rect 40684 15520 40724 15560
rect 40780 15520 40820 15560
rect 42124 15520 42164 15560
rect 42988 15520 43028 15560
rect 15820 15436 15860 15476
rect 34540 15436 34580 15476
rect 17548 15352 17588 15392
rect 17932 15352 17972 15392
rect 16492 15268 16532 15308
rect 20236 15268 20276 15308
rect 22252 15268 22292 15308
rect 44140 15268 44180 15308
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 9100 14932 9140 14972
rect 51532 14848 51572 14888
rect 55468 14848 55508 14888
rect 4012 14764 4052 14804
rect 37804 14764 37844 14804
rect 56524 14764 56564 14804
rect 5164 14680 5204 14720
rect 6316 14680 6356 14720
rect 8044 14680 8084 14720
rect 8428 14680 8468 14720
rect 8908 14680 8948 14720
rect 10636 14680 10676 14720
rect 11308 14680 11348 14720
rect 21292 14680 21332 14720
rect 21676 14680 21716 14720
rect 22540 14680 22580 14720
rect 33676 14680 33716 14720
rect 34060 14680 34100 14720
rect 34540 14680 34580 14720
rect 35788 14680 35828 14720
rect 36652 14680 36692 14720
rect 38284 14680 38324 14720
rect 38668 14680 38708 14720
rect 51244 14680 51284 14720
rect 52204 14680 52244 14720
rect 53644 14680 53684 14720
rect 55372 14680 55412 14720
rect 55564 14680 55604 14720
rect 56044 14680 56084 14720
rect 56140 14680 56180 14720
rect 57196 14680 57236 14720
rect 59404 14680 59444 14720
rect 59788 14680 59828 14720
rect 8524 14596 8564 14636
rect 34156 14596 34196 14636
rect 35212 14596 35252 14636
rect 35404 14596 35444 14636
rect 59308 14596 59348 14636
rect 652 14512 692 14552
rect 3820 14512 3860 14552
rect 4492 14512 4532 14552
rect 5836 14512 5876 14552
rect 8812 14512 8852 14552
rect 23692 14512 23732 14552
rect 38764 14512 38804 14552
rect 52972 14512 53012 14552
rect 56332 14512 56372 14552
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 5356 14176 5396 14216
rect 11884 14176 11924 14216
rect 18508 14176 18548 14216
rect 55180 14176 55220 14216
rect 61420 14176 61460 14216
rect 2956 14092 2996 14132
rect 7180 14092 7220 14132
rect 9196 14092 9236 14132
rect 43564 14092 43604 14132
rect 50572 14092 50612 14132
rect 57868 14092 57908 14132
rect 3340 14008 3380 14048
rect 4204 14008 4244 14048
rect 6220 14008 6260 14048
rect 7084 14008 7124 14048
rect 7276 14008 7316 14048
rect 9100 14008 9140 14048
rect 9292 14008 9332 14048
rect 9484 14008 9524 14048
rect 9868 14008 9908 14048
rect 10732 14008 10772 14048
rect 12076 14008 12116 14048
rect 12748 14008 12788 14048
rect 19180 14008 19220 14048
rect 26860 14008 26900 14048
rect 27724 14008 27764 14048
rect 39148 14008 39188 14048
rect 43756 14008 43796 14048
rect 44044 14008 44084 14048
rect 45388 14008 45428 14048
rect 46252 14008 46292 14048
rect 46636 14008 46676 14048
rect 47308 14008 47348 14048
rect 47980 14008 48020 14048
rect 49324 14008 49364 14048
rect 50188 14008 50228 14048
rect 55372 14008 55412 14048
rect 55660 14008 55700 14048
rect 56716 14008 56756 14048
rect 57004 14008 57044 14048
rect 59020 14008 59060 14048
rect 59404 14008 59444 14048
rect 60268 14008 60308 14048
rect 5740 13924 5780 13964
rect 6892 13924 6932 13964
rect 17548 13924 17588 13964
rect 44236 13924 44276 13964
rect 5548 13840 5588 13880
rect 57292 13840 57332 13880
rect 17356 13756 17396 13796
rect 38476 13756 38516 13796
rect 48172 13756 48212 13796
rect 56044 13756 56084 13796
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 6412 13420 6452 13460
rect 9292 13420 9332 13460
rect 12268 13420 12308 13460
rect 19276 13420 19316 13460
rect 49612 13420 49652 13460
rect 23116 13336 23156 13376
rect 9100 13252 9140 13292
rect 9484 13252 9524 13292
rect 4012 13168 4052 13208
rect 4396 13168 4436 13208
rect 5260 13168 5300 13208
rect 10252 13168 10292 13208
rect 11116 13168 11156 13208
rect 16876 13168 16916 13208
rect 17260 13168 17300 13208
rect 18124 13168 18164 13208
rect 23020 13168 23060 13208
rect 23212 13168 23252 13208
rect 23500 13168 23540 13208
rect 26092 13168 26132 13208
rect 38476 13168 38516 13208
rect 38860 13168 38900 13208
rect 39724 13168 39764 13208
rect 41644 13168 41684 13208
rect 48652 13168 48692 13208
rect 49804 13168 49844 13208
rect 49900 13168 49940 13208
rect 54796 13168 54836 13208
rect 55660 13168 55700 13208
rect 56044 13168 56084 13208
rect 56620 13168 56660 13208
rect 9868 13084 9908 13124
rect 652 13000 692 13040
rect 9676 13000 9716 13040
rect 24172 13000 24212 13040
rect 26764 13000 26804 13040
rect 40876 13000 40916 13040
rect 42316 13000 42356 13040
rect 49324 13000 49364 13040
rect 53644 13000 53684 13040
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 652 12664 692 12704
rect 31660 12664 31700 12704
rect 50476 12664 50516 12704
rect 23212 12580 23252 12620
rect 23788 12580 23828 12620
rect 28300 12580 28340 12620
rect 42700 12580 42740 12620
rect 49420 12580 49460 12620
rect 9484 12496 9524 12536
rect 19372 12496 19412 12536
rect 21292 12496 21332 12536
rect 22732 12496 22772 12536
rect 23020 12496 23060 12536
rect 23500 12496 23540 12536
rect 23596 12496 23636 12536
rect 23692 12496 23732 12536
rect 23973 12495 24013 12535
rect 24172 12496 24212 12536
rect 28684 12496 28724 12536
rect 29548 12496 29588 12536
rect 31180 12496 31220 12536
rect 31276 12496 31316 12536
rect 31756 12496 31796 12536
rect 35884 12496 35924 12536
rect 41740 12496 41780 12536
rect 42604 12496 42644 12536
rect 42796 12496 42836 12536
rect 49324 12496 49364 12536
rect 49516 12496 49556 12536
rect 50572 12496 50612 12536
rect 50956 12496 50996 12536
rect 53164 12496 53204 12536
rect 54124 12496 54164 12536
rect 54412 12496 54452 12536
rect 54796 12496 54836 12536
rect 55660 12496 55700 12536
rect 30700 12412 30740 12452
rect 30892 12412 30932 12452
rect 41164 12412 41204 12452
rect 56812 12412 56852 12452
rect 9004 12328 9044 12368
rect 18796 12328 18836 12368
rect 23980 12328 24020 12368
rect 21772 12244 21812 12284
rect 31948 12244 31988 12284
rect 35212 12244 35252 12284
rect 42412 12244 42452 12284
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 30316 11908 30356 11948
rect 41932 11908 41972 11948
rect 49516 11908 49556 11948
rect 53836 11908 53876 11948
rect 29932 11824 29972 11864
rect 42892 11824 42932 11864
rect 23692 11740 23732 11780
rect 18124 11656 18164 11696
rect 18988 11656 19028 11696
rect 23308 11656 23348 11696
rect 23404 11656 23444 11696
rect 24172 11656 24212 11696
rect 29932 11656 29972 11696
rect 31468 11656 31508 11696
rect 32332 11656 32372 11696
rect 41356 11656 41396 11696
rect 41644 11656 41684 11696
rect 42604 11656 42644 11696
rect 43084 11656 43124 11696
rect 43180 11656 43220 11696
rect 47308 11656 47348 11696
rect 49036 11656 49076 11696
rect 49324 11656 49364 11696
rect 50188 11656 50228 11696
rect 53548 11656 53588 11696
rect 61804 11656 61844 11696
rect 32716 11572 32756 11612
rect 48844 11572 48884 11612
rect 652 11488 692 11528
rect 24844 11488 24884 11528
rect 30124 11488 30164 11528
rect 40684 11488 40724 11528
rect 46636 11488 46676 11528
rect 61132 11488 61172 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 652 11152 692 11192
rect 18700 11152 18740 11192
rect 32236 11152 32276 11192
rect 33100 11152 33140 11192
rect 41932 11152 41972 11192
rect 59212 11152 59252 11192
rect 61996 11152 62036 11192
rect 24460 11068 24500 11108
rect 44332 11068 44372 11108
rect 10252 10984 10292 11024
rect 13612 10984 13652 11024
rect 15436 10984 15476 11024
rect 16108 10984 16148 11024
rect 16300 10984 16340 11024
rect 16684 10984 16724 11024
rect 17548 10984 17588 11024
rect 20716 10984 20756 11024
rect 21676 10984 21716 11024
rect 24844 10984 24884 11024
rect 25708 10984 25748 11024
rect 31180 10984 31220 11024
rect 31276 10949 31316 10989
rect 31372 10984 31412 11024
rect 31948 10984 31988 11024
rect 32044 10984 32084 11024
rect 33772 10984 33812 11024
rect 37036 10984 37076 11024
rect 37900 10984 37940 11024
rect 38284 10984 38324 11024
rect 41164 10984 41204 11024
rect 43084 10984 43124 11024
rect 43948 10984 43988 11024
rect 52588 10984 52628 11024
rect 58732 10984 58772 11024
rect 59020 10984 59060 11024
rect 59596 10984 59636 11024
rect 59980 10984 60020 11024
rect 60844 10984 60884 11024
rect 51724 10900 51764 10940
rect 9580 10732 9620 10772
rect 12940 10732 12980 10772
rect 26860 10732 26900 10772
rect 30892 10732 30932 10772
rect 35884 10732 35924 10772
rect 40492 10732 40532 10772
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 15340 10396 15380 10436
rect 21964 10396 22004 10436
rect 49228 10396 49268 10436
rect 55180 10396 55220 10436
rect 58540 10396 58580 10436
rect 58924 10396 58964 10436
rect 59788 10396 59828 10436
rect 3148 10312 3188 10352
rect 55852 10312 55892 10352
rect 3340 10228 3380 10268
rect 37900 10228 37940 10268
rect 59980 10228 60020 10268
rect 4780 10144 4820 10184
rect 9868 10144 9908 10184
rect 12556 10144 12596 10184
rect 12748 10144 12788 10184
rect 12940 10144 12980 10184
rect 13324 10144 13364 10184
rect 14188 10144 14228 10184
rect 21100 10144 21140 10184
rect 21484 10144 21524 10184
rect 21868 10144 21908 10184
rect 22060 10144 22100 10184
rect 27820 10144 27860 10184
rect 28012 10144 28052 10184
rect 28204 10144 28244 10184
rect 28396 10144 28436 10184
rect 37036 10144 37076 10184
rect 38188 10144 38228 10184
rect 39052 10144 39092 10184
rect 41452 10144 41492 10184
rect 41740 10144 41780 10184
rect 47212 10144 47252 10184
rect 48076 10144 48116 10184
rect 55372 10144 55412 10184
rect 56524 10144 56564 10184
rect 58444 10144 58484 10184
rect 58636 10144 58676 10184
rect 58828 10144 58868 10184
rect 59020 10144 59060 10184
rect 61420 10144 61460 10184
rect 4108 10060 4148 10100
rect 28300 10060 28340 10100
rect 41260 10060 41300 10100
rect 46828 10060 46868 10100
rect 60748 10060 60788 10100
rect 652 9976 692 10016
rect 10540 9976 10580 10016
rect 21580 9976 21620 10016
rect 27916 9976 27956 10016
rect 55468 9976 55508 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 652 9640 692 9680
rect 4684 9640 4724 9680
rect 9196 9640 9236 9680
rect 12748 9640 12788 9680
rect 21004 9640 21044 9680
rect 33004 9640 33044 9680
rect 33484 9640 33524 9680
rect 47020 9640 47060 9680
rect 50476 9640 50516 9680
rect 59404 9640 59444 9680
rect 61996 9640 62036 9680
rect 2284 9556 2324 9596
rect 10348 9556 10388 9596
rect 39532 9556 39572 9596
rect 59596 9556 59636 9596
rect 2668 9472 2708 9512
rect 3532 9472 3572 9512
rect 6796 9472 6836 9512
rect 7180 9472 7220 9512
rect 8044 9472 8084 9512
rect 10732 9472 10772 9512
rect 11596 9472 11636 9512
rect 20332 9472 20372 9512
rect 21868 9472 21908 9512
rect 33100 9472 33140 9512
rect 33196 9472 33236 9512
rect 33292 9472 33332 9512
rect 34156 9472 34196 9512
rect 36364 9472 36404 9512
rect 38284 9472 38324 9512
rect 39148 9472 39188 9512
rect 46348 9472 46388 9512
rect 47212 9472 47252 9512
rect 47884 9472 47924 9512
rect 48076 9472 48116 9512
rect 48460 9472 48500 9512
rect 49324 9472 49364 9512
rect 53452 9472 53492 9512
rect 55276 9472 55316 9512
rect 55660 9472 55700 9512
rect 56524 9472 56564 9512
rect 59980 9472 60020 9512
rect 60844 9472 60884 9512
rect 54892 9388 54932 9428
rect 59212 9388 59252 9428
rect 37132 9304 37172 9344
rect 22540 9220 22580 9260
rect 35692 9220 35732 9260
rect 53260 9220 53300 9260
rect 54700 9220 54740 9260
rect 57676 9220 57716 9260
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 19084 8800 19124 8840
rect 33292 8800 33332 8840
rect 56812 8800 56852 8840
rect 34444 8716 34484 8756
rect 44524 8716 44564 8756
rect 3340 8632 3380 8672
rect 4204 8632 4244 8672
rect 17068 8632 17108 8672
rect 17932 8632 17972 8672
rect 23500 8632 23540 8672
rect 24460 8632 24500 8672
rect 25900 8632 25940 8672
rect 26092 8632 26132 8672
rect 27244 8632 27284 8672
rect 27340 8632 27380 8672
rect 28012 8632 28052 8672
rect 28300 8632 28340 8672
rect 29164 8632 29204 8672
rect 29548 8632 29588 8672
rect 29644 8632 29684 8672
rect 29740 8632 29780 8672
rect 29836 8632 29876 8672
rect 32332 8632 32372 8672
rect 33196 8632 33236 8672
rect 33388 8632 33428 8672
rect 33868 8632 33908 8672
rect 34156 8632 34196 8672
rect 34348 8632 34388 8672
rect 34540 8632 34580 8672
rect 38380 8632 38420 8672
rect 42508 8632 42548 8672
rect 43372 8632 43412 8672
rect 45676 8632 45716 8672
rect 46732 8632 46772 8672
rect 47116 8632 47156 8672
rect 54124 8632 54164 8672
rect 54508 8632 54548 8672
rect 55372 8632 55412 8672
rect 57484 8632 57524 8672
rect 2956 8548 2996 8588
rect 16684 8548 16724 8588
rect 25996 8548 26036 8588
rect 27820 8548 27860 8588
rect 42124 8548 42164 8588
rect 46636 8548 46676 8588
rect 652 8464 692 8504
rect 5356 8464 5396 8504
rect 23980 8464 24020 8504
rect 26956 8464 26996 8504
rect 28492 8464 28532 8504
rect 31660 8464 31700 8504
rect 33676 8464 33716 8504
rect 37996 8464 38036 8504
rect 46348 8464 46388 8504
rect 56524 8464 56564 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 652 8128 692 8168
rect 3724 8128 3764 8168
rect 6124 8128 6164 8168
rect 16492 8128 16532 8168
rect 27628 8128 27668 8168
rect 33100 8128 33140 8168
rect 33964 8128 34004 8168
rect 47500 8128 47540 8168
rect 55564 8128 55604 8168
rect 21964 8044 22004 8084
rect 25324 8044 25364 8084
rect 30028 8044 30068 8084
rect 48556 8044 48596 8084
rect 4396 7960 4436 8000
rect 4492 7960 4532 8000
rect 4588 7960 4628 8000
rect 5452 7960 5492 8000
rect 5644 7960 5684 8000
rect 5932 7960 5972 8000
rect 6604 7960 6644 8000
rect 7564 7960 7604 8000
rect 15820 7960 15860 8000
rect 18124 7960 18164 8000
rect 22348 7960 22388 8000
rect 23212 7960 23252 8000
rect 25420 7960 25460 8000
rect 25804 7960 25844 8000
rect 28780 7960 28820 8000
rect 29644 7960 29684 8000
rect 33388 7960 33428 8000
rect 33484 7960 33524 8000
rect 34060 7960 34100 8000
rect 34444 7960 34484 8000
rect 46540 7960 46580 8000
rect 46636 7960 46676 8000
rect 46732 7960 46772 8000
rect 47116 7960 47156 8000
rect 47212 7960 47252 8000
rect 49228 7960 49268 8000
rect 3916 7876 3956 7916
rect 24364 7876 24404 7916
rect 55756 7876 55796 7916
rect 18700 7792 18740 7832
rect 4780 7708 4820 7748
rect 6892 7708 6932 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 11500 7372 11540 7412
rect 14764 7372 14804 7412
rect 25420 7372 25460 7412
rect 33292 7372 33332 7412
rect 34252 7372 34292 7412
rect 49324 7372 49364 7412
rect 50380 7372 50420 7412
rect 56716 7372 56756 7412
rect 38860 7204 38900 7244
rect 39724 7204 39764 7244
rect 11212 7120 11252 7160
rect 12172 7120 12212 7160
rect 12748 7120 12788 7160
rect 13612 7120 13652 7160
rect 23404 7120 23444 7160
rect 24268 7120 24308 7160
rect 33196 7120 33236 7160
rect 33388 7120 33428 7160
rect 33580 7120 33620 7160
rect 40396 7120 40436 7160
rect 49804 7120 49844 7160
rect 51532 7120 51572 7160
rect 52396 7120 52436 7160
rect 56428 7120 56468 7160
rect 12364 7036 12404 7076
rect 23020 7036 23060 7076
rect 48940 7036 48980 7076
rect 52780 7036 52820 7076
rect 652 6952 692 6992
rect 38668 6952 38708 6992
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 12652 6616 12692 6656
rect 33484 6616 33524 6656
rect 40300 6616 40340 6656
rect 40684 6616 40724 6656
rect 40972 6616 41012 6656
rect 46924 6616 46964 6656
rect 37900 6532 37940 6572
rect 9676 6448 9716 6488
rect 12172 6448 12212 6488
rect 13132 6448 13172 6488
rect 19180 6448 19220 6488
rect 34156 6448 34196 6488
rect 34348 6448 34388 6488
rect 35308 6448 35348 6488
rect 38284 6448 38324 6488
rect 39148 6448 39188 6488
rect 40780 6448 40820 6488
rect 46444 6448 46484 6488
rect 46732 6448 46772 6488
rect 17644 6364 17684 6404
rect 10348 6280 10388 6320
rect 18508 6280 18548 6320
rect 17452 6196 17492 6236
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 4588 5860 4628 5900
rect 12364 5860 12404 5900
rect 19084 5860 19124 5900
rect 33484 5860 33524 5900
rect 44620 5860 44660 5900
rect 46348 5860 46388 5900
rect 2956 5692 2996 5732
rect 12172 5692 12212 5732
rect 37420 5692 37460 5732
rect 2092 5608 2132 5648
rect 2764 5608 2804 5648
rect 4492 5608 4532 5648
rect 4684 5608 4724 5648
rect 5164 5608 5204 5648
rect 6220 5608 6260 5648
rect 9772 5608 9812 5648
rect 10156 5608 10196 5648
rect 11020 5608 11060 5648
rect 13036 5608 13076 5648
rect 16684 5608 16724 5648
rect 17068 5608 17108 5648
rect 17932 5608 17972 5648
rect 19660 5608 19700 5648
rect 20620 5608 20660 5648
rect 30220 5608 30260 5648
rect 31468 5608 31508 5648
rect 32332 5608 32372 5648
rect 36556 5608 36596 5648
rect 37228 5608 37268 5648
rect 39340 5608 39380 5648
rect 39532 5608 39572 5648
rect 42604 5608 42644 5648
rect 43468 5608 43508 5648
rect 47500 5608 47540 5648
rect 48364 5608 48404 5648
rect 54028 5608 54068 5648
rect 30892 5524 30932 5564
rect 31084 5524 31124 5564
rect 39436 5524 39476 5564
rect 42220 5524 42260 5564
rect 48748 5524 48788 5564
rect 652 5440 692 5480
rect 3148 5440 3188 5480
rect 5068 5440 5108 5480
rect 5356 5440 5396 5480
rect 5548 5440 5588 5480
rect 37612 5440 37652 5480
rect 53356 5440 53396 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 1324 5104 1364 5144
rect 41548 5104 41588 5144
rect 50092 5104 50132 5144
rect 3724 5020 3764 5060
rect 6988 5020 7028 5060
rect 38380 5020 38420 5060
rect 50380 5020 50420 5060
rect 2476 4936 2516 4976
rect 3340 4936 3380 4976
rect 3916 4936 3956 4976
rect 4300 4936 4340 4976
rect 5164 4936 5204 4976
rect 7372 4936 7412 4976
rect 8236 4936 8276 4976
rect 26860 4936 26900 4976
rect 27532 4936 27572 4976
rect 27724 4936 27764 4976
rect 28108 4936 28148 4976
rect 28972 4936 29012 4976
rect 37132 4936 37172 4976
rect 37996 4936 38036 4976
rect 39916 4936 39956 4976
rect 41068 4936 41108 4976
rect 41356 4936 41396 4976
rect 50188 4936 50228 4976
rect 51916 4936 51956 4976
rect 52300 4936 52340 4976
rect 53164 4936 53204 4976
rect 844 4852 884 4892
rect 6316 4852 6356 4892
rect 9388 4852 9428 4892
rect 30124 4852 30164 4892
rect 35980 4852 36020 4892
rect 39436 4852 39476 4892
rect 54316 4852 54356 4892
rect 652 4768 692 4808
rect 40204 4684 40244 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 4396 4348 4436 4388
rect 26188 4348 26228 4388
rect 41164 4348 41204 4388
rect 51916 4348 51956 4388
rect 844 4180 884 4220
rect 4588 4180 4628 4220
rect 12940 4180 12980 4220
rect 16972 4180 17012 4220
rect 52108 4180 52148 4220
rect 16300 4096 16340 4136
rect 17644 4096 17684 4136
rect 18700 4096 18740 4136
rect 22924 4096 22964 4136
rect 24172 4096 24212 4136
rect 25036 4096 25076 4136
rect 30988 4096 31028 4136
rect 41068 4096 41108 4136
rect 41260 4096 41300 4136
rect 49228 4096 49268 4136
rect 49612 4096 49652 4136
rect 18028 4012 18068 4052
rect 23596 4012 23636 4052
rect 23788 4012 23828 4052
rect 49132 4012 49172 4052
rect 652 3928 692 3968
rect 12748 3928 12788 3968
rect 17548 3923 17588 3963
rect 17836 3928 17876 3968
rect 31660 3928 31700 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 14188 3592 14228 3632
rect 18700 3592 18740 3632
rect 21772 3592 21812 3632
rect 40108 3592 40148 3632
rect 41644 3592 41684 3632
rect 49516 3592 49556 3632
rect 11788 3508 11828 3548
rect 19372 3508 19412 3548
rect 49228 3508 49268 3548
rect 50476 3508 50516 3548
rect 12172 3424 12212 3464
rect 13036 3424 13076 3464
rect 16300 3424 16340 3464
rect 16684 3424 16724 3464
rect 17548 3424 17588 3464
rect 19756 3424 19796 3464
rect 20620 3424 20660 3464
rect 31084 3424 31124 3464
rect 31468 3424 31508 3464
rect 32332 3424 32372 3464
rect 33580 3424 33620 3464
rect 40780 3424 40820 3464
rect 40972 3424 41012 3464
rect 45772 3424 45812 3464
rect 46444 3424 46484 3464
rect 49132 3424 49172 3464
rect 49324 3424 49364 3464
rect 50188 3424 50228 3464
rect 50379 3445 50419 3485
rect 50572 3424 50612 3464
rect 54028 3424 54068 3464
rect 844 3340 884 3380
rect 39436 3340 39476 3380
rect 41836 3340 41876 3380
rect 46636 3340 46676 3380
rect 48748 3340 48788 3380
rect 652 3172 692 3212
rect 39244 3172 39284 3212
rect 42028 3172 42068 3212
rect 46828 3172 46868 3212
rect 48556 3172 48596 3212
rect 53356 3172 53396 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 16876 2836 16916 2876
rect 18124 2836 18164 2876
rect 30604 2836 30644 2876
rect 40492 2836 40532 2876
rect 40684 2836 40724 2876
rect 45004 2836 45044 2876
rect 49996 2836 50036 2876
rect 54604 2836 54644 2876
rect 17548 2752 17588 2792
rect 52012 2752 52052 2792
rect 844 2668 884 2708
rect 14668 2668 14708 2708
rect 17068 2668 17108 2708
rect 23308 2668 23348 2708
rect 27052 2668 27092 2708
rect 51820 2668 51860 2708
rect 12652 2584 12692 2624
rect 13516 2584 13556 2624
rect 14860 2584 14900 2624
rect 15532 2584 15572 2624
rect 17452 2584 17492 2624
rect 17644 2584 17684 2624
rect 18019 2571 18059 2611
rect 18220 2584 18260 2624
rect 18700 2584 18740 2624
rect 18988 2584 19028 2624
rect 21292 2584 21332 2624
rect 22156 2584 22196 2624
rect 23788 2584 23828 2624
rect 25036 2584 25076 2624
rect 25900 2584 25940 2624
rect 27340 2584 27380 2624
rect 28588 2584 28628 2624
rect 29452 2584 29492 2624
rect 38092 2584 38132 2624
rect 38476 2584 38516 2624
rect 39340 2584 39380 2624
rect 41836 2584 41876 2624
rect 42700 2584 42740 2624
rect 43084 2584 43124 2624
rect 46156 2584 46196 2624
rect 47020 2584 47060 2624
rect 47404 2584 47444 2624
rect 47596 2584 47636 2624
rect 47980 2584 48020 2624
rect 48844 2584 48884 2624
rect 52204 2584 52244 2624
rect 52588 2584 52628 2624
rect 53452 2584 53492 2624
rect 12268 2500 12308 2540
rect 19180 2500 19220 2540
rect 20908 2500 20948 2540
rect 24460 2500 24500 2540
rect 24652 2500 24692 2540
rect 28012 2500 28052 2540
rect 28204 2500 28244 2540
rect 652 2416 692 2456
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 13324 2080 13364 2120
rect 13516 1828 13556 1868
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal2 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 95072 38576 95440 38585
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95072 38527 95440 38536
rect 37324 38240 37364 38249
rect 37364 38200 37652 38240
rect 37324 38191 37364 38200
rect 36652 37988 36692 37997
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 20619 37568 20661 37577
rect 20619 37528 20620 37568
rect 20660 37528 20661 37568
rect 20619 37519 20661 37528
rect 9484 37484 9524 37493
rect 9292 37232 9332 37241
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 9292 36812 9332 37192
rect 9484 37232 9524 37444
rect 10348 37400 10388 37409
rect 9676 37232 9716 37241
rect 9484 37192 9676 37232
rect 9388 36812 9428 36821
rect 9292 36772 9388 36812
rect 9388 36763 9428 36772
rect 75 36728 117 36737
rect 75 36688 76 36728
rect 116 36688 117 36728
rect 75 36679 117 36688
rect 7276 36728 7316 36737
rect 76 20105 116 36679
rect 5835 36644 5877 36653
rect 5835 36604 5836 36644
rect 5876 36604 5877 36644
rect 5835 36595 5877 36604
rect 4683 36560 4725 36569
rect 4683 36520 4684 36560
rect 4724 36520 4725 36560
rect 4683 36511 4725 36520
rect 5643 36560 5685 36569
rect 5643 36520 5644 36560
rect 5684 36520 5685 36560
rect 5643 36511 5685 36520
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 4684 35888 4724 36511
rect 5644 36426 5684 36511
rect 5836 36510 5876 36595
rect 6603 36560 6645 36569
rect 6603 36520 6604 36560
rect 6644 36520 6645 36560
rect 6603 36511 6645 36520
rect 6604 36426 6644 36511
rect 7084 36140 7124 36149
rect 7276 36140 7316 36688
rect 7371 36560 7413 36569
rect 7371 36520 7372 36560
rect 7412 36520 7413 36560
rect 7371 36511 7413 36520
rect 7124 36100 7316 36140
rect 7084 36091 7124 36100
rect 7372 36056 7412 36511
rect 7276 36016 7412 36056
rect 4684 35839 4724 35848
rect 5067 35888 5109 35897
rect 5932 35888 5972 35897
rect 5067 35848 5068 35888
rect 5108 35848 5109 35888
rect 5067 35839 5109 35848
rect 5164 35848 5932 35888
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 5068 35384 5108 35839
rect 4972 35344 5108 35384
rect 4876 34964 4916 34973
rect 3916 34924 4876 34964
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 3916 34376 3956 34924
rect 4876 34915 4916 34924
rect 4972 34385 5012 35344
rect 5067 35216 5109 35225
rect 5067 35176 5068 35216
rect 5108 35176 5109 35216
rect 5067 35167 5109 35176
rect 5068 35132 5108 35167
rect 5068 35081 5108 35092
rect 3916 34327 3956 34336
rect 4299 34376 4341 34385
rect 4299 34336 4300 34376
rect 4340 34336 4341 34376
rect 4299 34327 4341 34336
rect 4971 34376 5013 34385
rect 4971 34336 4972 34376
rect 5012 34336 5013 34376
rect 4971 34327 5013 34336
rect 5164 34376 5204 35848
rect 5835 35216 5877 35225
rect 5835 35176 5836 35216
rect 5876 35176 5877 35216
rect 5835 35167 5877 35176
rect 5836 35082 5876 35167
rect 5164 34327 5204 34336
rect 4300 34242 4340 34327
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 5932 32789 5972 35848
rect 6508 35216 6548 35225
rect 6316 35176 6508 35216
rect 6316 34628 6356 35176
rect 6508 35167 6548 35176
rect 7276 35216 7316 36016
rect 9099 35888 9141 35897
rect 9099 35848 9100 35888
rect 9140 35848 9141 35888
rect 9099 35839 9141 35848
rect 9196 35888 9236 35897
rect 8715 35804 8757 35813
rect 8715 35764 8716 35804
rect 8756 35764 8757 35804
rect 8715 35755 8757 35764
rect 7371 35300 7413 35309
rect 7371 35260 7372 35300
rect 7412 35260 7413 35300
rect 7371 35251 7413 35260
rect 8427 35300 8469 35309
rect 8427 35260 8428 35300
rect 8468 35260 8469 35300
rect 8427 35251 8469 35260
rect 7276 35167 7316 35176
rect 7372 35166 7412 35251
rect 7467 35216 7509 35225
rect 7467 35176 7468 35216
rect 7508 35176 7509 35216
rect 7467 35167 7509 35176
rect 7947 35216 7989 35225
rect 7947 35176 7948 35216
rect 7988 35176 7989 35216
rect 7947 35167 7989 35176
rect 7468 35082 7508 35167
rect 6316 34579 6356 34588
rect 7948 34208 7988 35167
rect 8043 35132 8085 35141
rect 8043 35092 8044 35132
rect 8084 35092 8085 35132
rect 8043 35083 8085 35092
rect 8044 34376 8084 35083
rect 8044 34327 8084 34336
rect 8428 34376 8468 35251
rect 8428 34327 8468 34336
rect 8716 34376 8756 35755
rect 8716 34327 8756 34336
rect 7948 34159 7988 34168
rect 8235 34208 8277 34217
rect 8235 34168 8236 34208
rect 8276 34168 8277 34208
rect 8235 34159 8277 34168
rect 8811 34208 8853 34217
rect 8811 34168 8812 34208
rect 8852 34168 8853 34208
rect 8811 34159 8853 34168
rect 8908 34208 8948 34217
rect 8236 34074 8276 34159
rect 7468 32873 7508 32958
rect 6508 32864 6548 32873
rect 4107 32780 4149 32789
rect 4107 32740 4108 32780
rect 4148 32740 4149 32780
rect 4107 32731 4149 32740
rect 5931 32780 5973 32789
rect 5931 32740 5932 32780
rect 5972 32740 5973 32780
rect 5931 32731 5973 32740
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 3916 31352 3956 31361
rect 3820 31312 3916 31352
rect 2859 30680 2901 30689
rect 2859 30640 2860 30680
rect 2900 30640 2901 30680
rect 2859 30631 2901 30640
rect 3244 30680 3284 30691
rect 2860 30546 2900 30631
rect 3244 30605 3284 30640
rect 3820 30605 3860 31312
rect 3916 31303 3956 31312
rect 3915 30680 3957 30689
rect 4108 30680 4148 32731
rect 6508 32705 6548 32824
rect 7467 32864 7509 32873
rect 7467 32824 7468 32864
rect 7508 32824 7509 32864
rect 7467 32815 7509 32824
rect 8812 32864 8852 34159
rect 8812 32815 8852 32824
rect 6507 32696 6549 32705
rect 6507 32656 6508 32696
rect 6548 32656 6549 32696
rect 6507 32647 6549 32656
rect 6988 32696 7028 32705
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 6988 32201 7028 32656
rect 8812 32276 8852 32285
rect 8908 32276 8948 34168
rect 9100 32864 9140 35839
rect 9196 35132 9236 35848
rect 9388 35888 9428 35897
rect 9484 35888 9524 37192
rect 9676 37183 9716 37192
rect 10348 36905 10388 37360
rect 18700 37400 18740 37409
rect 18315 37316 18357 37325
rect 18315 37276 18316 37316
rect 18356 37276 18357 37316
rect 18315 37267 18357 37276
rect 18316 37182 18356 37267
rect 10347 36896 10389 36905
rect 10347 36856 10348 36896
rect 10388 36856 10389 36896
rect 10347 36847 10389 36856
rect 11787 36896 11829 36905
rect 11787 36856 11788 36896
rect 11828 36856 11829 36896
rect 11787 36847 11829 36856
rect 11788 36762 11828 36847
rect 9772 36728 9812 36737
rect 9772 35897 9812 36688
rect 10636 36728 10676 36737
rect 9428 35848 9524 35888
rect 9771 35888 9813 35897
rect 9771 35848 9772 35888
rect 9812 35848 9813 35888
rect 9388 35839 9428 35848
rect 9771 35839 9813 35848
rect 9963 35888 10005 35897
rect 9963 35848 9964 35888
rect 10004 35848 10005 35888
rect 10636 35888 10676 36688
rect 18700 36569 18740 37360
rect 19564 37400 19604 37409
rect 19604 37360 19988 37400
rect 19564 37351 19604 37360
rect 19275 37316 19317 37325
rect 19275 37276 19276 37316
rect 19316 37276 19317 37316
rect 19275 37267 19317 37276
rect 18795 36728 18837 36737
rect 18795 36688 18796 36728
rect 18836 36688 18837 36728
rect 18795 36679 18837 36688
rect 19180 36728 19220 36737
rect 18796 36594 18836 36679
rect 19180 36569 19220 36688
rect 18699 36560 18741 36569
rect 18699 36520 18700 36560
rect 18740 36520 18741 36560
rect 18699 36511 18741 36520
rect 19179 36560 19221 36569
rect 19179 36520 19180 36560
rect 19220 36520 19221 36560
rect 19179 36511 19221 36520
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 19276 36140 19316 37267
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 19851 36728 19893 36737
rect 19851 36688 19852 36728
rect 19892 36688 19893 36728
rect 19948 36728 19988 37360
rect 20044 36728 20084 36737
rect 19948 36688 20044 36728
rect 20084 36688 20276 36728
rect 19851 36679 19893 36688
rect 20044 36679 20084 36688
rect 19276 36091 19316 36100
rect 19852 36140 19892 36679
rect 19852 36091 19892 36100
rect 19468 35972 19508 35983
rect 19468 35897 19508 35932
rect 20043 35972 20085 35981
rect 20043 35932 20044 35972
rect 20084 35932 20085 35972
rect 20043 35923 20085 35932
rect 10828 35888 10868 35897
rect 10636 35848 10828 35888
rect 9963 35839 10005 35848
rect 9291 35804 9333 35813
rect 9291 35764 9292 35804
rect 9332 35764 9333 35804
rect 9291 35755 9333 35764
rect 9580 35804 9620 35813
rect 9292 35670 9332 35755
rect 9484 35384 9524 35393
rect 9580 35384 9620 35764
rect 9964 35754 10004 35839
rect 10347 35720 10389 35729
rect 10347 35680 10348 35720
rect 10388 35680 10389 35720
rect 10347 35671 10389 35680
rect 9524 35344 9620 35384
rect 9484 35335 9524 35344
rect 10348 35216 10388 35671
rect 10348 35167 10388 35176
rect 9291 35132 9333 35141
rect 9196 35092 9292 35132
rect 9332 35092 9333 35132
rect 9291 35083 9333 35092
rect 9675 35132 9717 35141
rect 9675 35092 9676 35132
rect 9716 35092 9717 35132
rect 9675 35083 9717 35092
rect 9292 34998 9332 35083
rect 9676 34998 9716 35083
rect 9675 33704 9717 33713
rect 9675 33664 9676 33704
rect 9716 33664 9717 33704
rect 9675 33655 9717 33664
rect 10732 33704 10772 35848
rect 10828 35839 10868 35848
rect 19467 35888 19509 35897
rect 19467 35848 19468 35888
rect 19508 35848 19509 35888
rect 19467 35839 19509 35848
rect 20044 35838 20084 35923
rect 11979 35720 12021 35729
rect 11979 35680 11980 35720
rect 12020 35680 12021 35720
rect 11979 35671 12021 35680
rect 11980 35586 12020 35671
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 20236 34628 20276 36688
rect 20332 34628 20372 34637
rect 20236 34588 20332 34628
rect 20332 34579 20372 34588
rect 16875 34460 16917 34469
rect 16875 34420 16876 34460
rect 16916 34420 16917 34460
rect 16875 34411 16917 34420
rect 17739 34460 17781 34469
rect 17739 34420 17740 34460
rect 17780 34420 17781 34460
rect 17739 34411 17781 34420
rect 14860 34376 14900 34385
rect 15724 34376 15764 34385
rect 14900 34336 15092 34376
rect 14860 34327 14900 34336
rect 14475 34292 14517 34301
rect 14475 34252 14476 34292
rect 14516 34252 14517 34292
rect 14475 34243 14517 34252
rect 14476 34158 14516 34243
rect 9676 32873 9716 33655
rect 10732 33545 10772 33664
rect 11115 33704 11157 33713
rect 11115 33664 11116 33704
rect 11156 33664 11157 33704
rect 11115 33655 11157 33664
rect 12076 33704 12116 33713
rect 11116 33570 11156 33655
rect 10059 33536 10101 33545
rect 10059 33496 10060 33536
rect 10100 33496 10101 33536
rect 10059 33487 10101 33496
rect 10731 33536 10773 33545
rect 10731 33496 10732 33536
rect 10772 33496 10773 33536
rect 10731 33487 10773 33496
rect 11403 33536 11445 33545
rect 11403 33496 11404 33536
rect 11444 33496 11445 33536
rect 11403 33487 11445 33496
rect 9196 32864 9236 32873
rect 9100 32824 9196 32864
rect 8852 32236 8948 32276
rect 8812 32227 8852 32236
rect 6987 32192 7029 32201
rect 6987 32152 6988 32192
rect 7028 32152 7029 32192
rect 6987 32143 7029 32152
rect 9196 32192 9236 32824
rect 9675 32864 9717 32873
rect 9675 32824 9676 32864
rect 9716 32824 9717 32864
rect 9675 32815 9717 32824
rect 10060 32864 10100 33487
rect 11404 33402 11444 33487
rect 12076 32873 12116 33664
rect 14956 33704 14996 33713
rect 14956 33125 14996 33664
rect 15052 33704 15092 34336
rect 15435 34292 15477 34301
rect 15435 34252 15436 34292
rect 15476 34252 15477 34292
rect 15435 34243 15477 34252
rect 15340 33704 15380 33713
rect 15052 33664 15340 33704
rect 14955 33116 14997 33125
rect 14955 33076 14956 33116
rect 14996 33076 14997 33116
rect 14955 33067 14997 33076
rect 10060 32815 10100 32824
rect 12075 32864 12117 32873
rect 12075 32824 12076 32864
rect 12116 32824 12117 32864
rect 12075 32815 12117 32824
rect 9196 31529 9236 32152
rect 9195 31520 9237 31529
rect 9195 31480 9196 31520
rect 9236 31480 9237 31520
rect 9195 31471 9237 31480
rect 4876 31352 4916 31361
rect 4876 31193 4916 31312
rect 4875 31184 4917 31193
rect 4875 31144 4876 31184
rect 4916 31144 4917 31184
rect 4875 31135 4917 31144
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 3915 30640 3916 30680
rect 3956 30640 3957 30680
rect 3915 30631 3957 30640
rect 4012 30640 4108 30680
rect 3243 30596 3285 30605
rect 3243 30556 3244 30596
rect 3284 30556 3285 30596
rect 3243 30547 3285 30556
rect 3627 30596 3669 30605
rect 3627 30556 3628 30596
rect 3668 30556 3669 30596
rect 3627 30547 3669 30556
rect 3819 30596 3861 30605
rect 3819 30556 3820 30596
rect 3860 30556 3861 30596
rect 3819 30547 3861 30556
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 3532 29672 3572 29681
rect 2764 29632 3532 29672
rect 2764 29252 2804 29632
rect 3532 29623 3572 29632
rect 2764 29203 2804 29212
rect 3148 29168 3188 29177
rect 3628 29168 3668 30547
rect 3916 30092 3956 30631
rect 3916 30043 3956 30052
rect 3723 29924 3765 29933
rect 3723 29884 3724 29924
rect 3764 29884 3765 29924
rect 3723 29875 3765 29884
rect 3724 29790 3764 29875
rect 3188 29128 3668 29168
rect 4012 29168 4052 30640
rect 4108 30631 4148 30640
rect 6124 30680 6164 30689
rect 5260 30596 5300 30605
rect 6124 30596 6164 30640
rect 5300 30556 6164 30596
rect 8235 30596 8277 30605
rect 8235 30556 8236 30596
rect 8276 30556 8277 30596
rect 5260 30547 5300 30556
rect 8235 30547 8277 30556
rect 5452 30428 5492 30437
rect 5452 30017 5492 30388
rect 4107 30008 4149 30017
rect 4107 29968 4108 30008
rect 4148 29968 4149 30008
rect 4107 29959 4149 29968
rect 5067 30008 5109 30017
rect 5067 29968 5068 30008
rect 5108 29968 5109 30008
rect 5067 29959 5109 29968
rect 5451 30008 5493 30017
rect 5451 29968 5452 30008
rect 5492 29968 5493 30008
rect 5451 29959 5493 29968
rect 4108 29924 4148 29959
rect 4108 29873 4148 29884
rect 4587 29924 4629 29933
rect 4587 29884 4588 29924
rect 4628 29884 4629 29924
rect 4587 29875 4629 29884
rect 4971 29924 5013 29933
rect 4971 29884 4972 29924
rect 5012 29884 5013 29924
rect 4971 29875 5013 29884
rect 4588 29790 4628 29875
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 3148 29119 3188 29128
rect 4012 29119 4052 29128
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 4972 27917 5012 29875
rect 4971 27908 5013 27917
rect 4971 27868 4972 27908
rect 5012 27868 5013 27908
rect 4971 27859 5013 27868
rect 4395 27824 4437 27833
rect 4395 27784 4396 27824
rect 4436 27784 4437 27824
rect 4395 27775 4437 27784
rect 4683 27824 4725 27833
rect 4683 27784 4684 27824
rect 4724 27784 4725 27824
rect 4683 27775 4725 27784
rect 4972 27824 5012 27859
rect 4299 27740 4341 27749
rect 4299 27700 4300 27740
rect 4340 27700 4341 27740
rect 4299 27691 4341 27700
rect 3819 27656 3861 27665
rect 3819 27616 3820 27656
rect 3860 27616 3861 27656
rect 3819 27607 3861 27616
rect 4204 27656 4244 27665
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 3435 26900 3477 26909
rect 3435 26860 3436 26900
rect 3476 26860 3477 26900
rect 3435 26851 3477 26860
rect 3820 26900 3860 27607
rect 4204 27068 4244 27616
rect 4300 27606 4340 27691
rect 4396 27656 4436 27775
rect 4588 27665 4628 27750
rect 4684 27740 4724 27775
rect 4972 27774 5012 27784
rect 4684 27689 4724 27700
rect 4396 27607 4436 27616
rect 4587 27656 4629 27665
rect 4587 27616 4588 27656
rect 4628 27616 4629 27656
rect 4587 27607 4629 27616
rect 4780 27656 4820 27665
rect 5068 27656 5108 29959
rect 5260 29840 5300 29849
rect 5164 29336 5204 29345
rect 5260 29336 5300 29800
rect 5204 29296 5300 29336
rect 5164 29287 5204 29296
rect 5931 29168 5973 29177
rect 5931 29128 5932 29168
rect 5972 29128 5973 29168
rect 5931 29119 5973 29128
rect 7851 29168 7893 29177
rect 7851 29128 7852 29168
rect 7892 29128 7893 29168
rect 7851 29119 7893 29128
rect 8236 29168 8276 30547
rect 9676 30092 9716 32815
rect 15052 32780 15092 33664
rect 15340 33655 15380 33664
rect 15436 33116 15476 34243
rect 15724 34217 15764 34336
rect 16876 34326 16916 34411
rect 17740 34376 17780 34411
rect 17740 34325 17780 34336
rect 15723 34208 15765 34217
rect 15723 34168 15724 34208
rect 15764 34168 15765 34208
rect 15723 34159 15765 34168
rect 16203 34208 16245 34217
rect 16203 34168 16204 34208
rect 16244 34168 16245 34208
rect 16203 34159 16245 34168
rect 17068 34208 17108 34217
rect 16204 33704 16244 34159
rect 16204 33655 16244 33664
rect 15436 33067 15476 33076
rect 15915 33116 15957 33125
rect 15915 33076 15916 33116
rect 15956 33076 15957 33116
rect 15915 33067 15957 33076
rect 15628 32957 15668 33042
rect 15916 32982 15956 33067
rect 17068 32957 17108 34168
rect 20331 34208 20373 34217
rect 20331 34168 20332 34208
rect 20372 34168 20373 34208
rect 20331 34159 20373 34168
rect 20332 34074 20372 34159
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 17548 33704 17588 33713
rect 17356 33620 17396 33629
rect 17548 33620 17588 33664
rect 17396 33580 17588 33620
rect 17356 33571 17396 33580
rect 18220 33452 18260 33461
rect 18124 33412 18220 33452
rect 15627 32948 15669 32957
rect 15627 32908 15628 32948
rect 15668 32908 15669 32948
rect 15627 32899 15669 32908
rect 16108 32948 16148 32957
rect 14764 32740 15092 32780
rect 15627 32780 15669 32789
rect 15627 32740 15628 32780
rect 15668 32740 15669 32780
rect 11212 32696 11252 32705
rect 11252 32656 11348 32696
rect 11212 32647 11252 32656
rect 10059 32192 10101 32201
rect 10059 32152 10060 32192
rect 10100 32152 10101 32192
rect 10059 32143 10101 32152
rect 10060 32058 10100 32143
rect 11211 31940 11253 31949
rect 11211 31900 11212 31940
rect 11252 31900 11253 31940
rect 11211 31891 11253 31900
rect 11212 31806 11252 31891
rect 11116 31184 11156 31193
rect 9676 30043 9716 30052
rect 10924 31144 11116 31184
rect 10155 29840 10197 29849
rect 10540 29840 10580 29849
rect 10155 29800 10156 29840
rect 10196 29800 10197 29840
rect 10155 29791 10197 29800
rect 10252 29800 10540 29840
rect 5739 27824 5781 27833
rect 5739 27784 5740 27824
rect 5780 27784 5781 27824
rect 5739 27775 5781 27784
rect 5451 27740 5493 27749
rect 5451 27700 5452 27740
rect 5492 27700 5493 27740
rect 5451 27691 5493 27700
rect 4820 27616 5068 27656
rect 4780 27607 4820 27616
rect 5068 27607 5108 27616
rect 5452 27656 5492 27691
rect 5452 27605 5492 27616
rect 5740 27656 5780 27775
rect 5932 27740 5972 29119
rect 7852 29034 7892 29119
rect 8236 29093 8276 29128
rect 9100 29168 9140 29177
rect 8235 29084 8277 29093
rect 8235 29044 8236 29084
rect 8276 29044 8277 29084
rect 8235 29035 8277 29044
rect 5932 27691 5972 27700
rect 5740 27607 5780 27616
rect 5067 27488 5109 27497
rect 5067 27448 5068 27488
rect 5108 27448 5109 27488
rect 5067 27439 5109 27448
rect 4204 26909 4244 27028
rect 5068 27068 5108 27439
rect 5259 27404 5301 27413
rect 5259 27364 5260 27404
rect 5300 27364 5301 27404
rect 5259 27355 5301 27364
rect 7083 27404 7125 27413
rect 7083 27364 7084 27404
rect 7124 27364 7125 27404
rect 7083 27355 7125 27364
rect 5260 27270 5300 27355
rect 5068 27019 5108 27028
rect 3820 26851 3860 26860
rect 4203 26900 4245 26909
rect 4203 26860 4204 26900
rect 4244 26860 4245 26900
rect 4203 26851 4245 26860
rect 3436 26766 3476 26851
rect 4876 26816 4916 26825
rect 4780 26776 4876 26816
rect 2475 26648 2517 26657
rect 2475 26608 2476 26648
rect 2516 26608 2517 26648
rect 2475 26599 2517 26608
rect 3244 26648 3284 26657
rect 2379 26480 2421 26489
rect 2379 26440 2380 26480
rect 2420 26440 2421 26480
rect 2379 26431 2421 26440
rect 2380 25304 2420 26431
rect 2476 26228 2516 26599
rect 3244 26489 3284 26608
rect 3627 26648 3669 26657
rect 3627 26608 3628 26648
rect 3668 26608 3669 26648
rect 3627 26599 3669 26608
rect 3628 26514 3668 26599
rect 3243 26480 3285 26489
rect 3243 26440 3244 26480
rect 3284 26440 3285 26480
rect 3243 26431 3285 26440
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 2476 26179 2516 26188
rect 2859 26144 2901 26153
rect 2859 26104 2860 26144
rect 2900 26104 2901 26144
rect 2859 26095 2901 26104
rect 3724 26144 3764 26153
rect 2380 25255 2420 25264
rect 2764 25304 2804 25313
rect 2860 25304 2900 26095
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 3724 25313 3764 26104
rect 4780 25556 4820 26776
rect 4876 26767 4916 26776
rect 5740 26816 5780 26825
rect 5740 26489 5780 26776
rect 4875 26480 4917 26489
rect 4875 26440 4876 26480
rect 4916 26440 4917 26480
rect 4875 26431 4917 26440
rect 5739 26480 5781 26489
rect 5739 26440 5740 26480
rect 5780 26440 5781 26480
rect 5739 26431 5781 26440
rect 6795 26480 6837 26489
rect 6795 26440 6796 26480
rect 6836 26440 6837 26480
rect 6795 26431 6837 26440
rect 4876 26312 4916 26431
rect 4876 26263 4916 26272
rect 4780 25507 4820 25516
rect 6123 25556 6165 25565
rect 6123 25516 6124 25556
rect 6164 25516 6165 25556
rect 6123 25507 6165 25516
rect 6124 25422 6164 25507
rect 2804 25264 2900 25304
rect 3628 25304 3668 25313
rect 3723 25304 3765 25313
rect 3668 25264 3724 25304
rect 3764 25264 3765 25304
rect 2764 23960 2804 25264
rect 3628 25255 3668 25264
rect 3723 25255 3765 25264
rect 5067 25304 5109 25313
rect 5067 25264 5068 25304
rect 5108 25264 5109 25304
rect 5067 25255 5109 25264
rect 5835 25304 5877 25313
rect 5835 25264 5836 25304
rect 5876 25264 5877 25304
rect 5835 25255 5877 25264
rect 6796 25304 6836 26431
rect 7084 26228 7124 27355
rect 7084 26179 7124 26188
rect 7467 26144 7509 26153
rect 7467 26104 7468 26144
rect 7508 26104 7509 26144
rect 7467 26095 7509 26104
rect 8332 26144 8372 26153
rect 7468 26010 7508 26095
rect 8332 25565 8372 26104
rect 8331 25556 8373 25565
rect 8331 25516 8332 25556
rect 8372 25516 8373 25556
rect 8331 25507 8373 25516
rect 6796 25255 6836 25264
rect 3724 25170 3764 25255
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 2668 23920 2804 23960
rect 1227 23120 1269 23129
rect 1227 23080 1228 23120
rect 1268 23080 1269 23120
rect 1227 23071 1269 23080
rect 2091 23120 2133 23129
rect 2091 23080 2092 23120
rect 2132 23080 2133 23120
rect 2091 23071 2133 23080
rect 1228 22532 1268 23071
rect 2092 22986 2132 23071
rect 1228 22483 1268 22492
rect 652 22448 692 22457
rect 652 21617 692 22408
rect 2668 22373 2708 23920
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 2956 23036 2996 23045
rect 2956 22877 2996 22996
rect 4491 23036 4533 23045
rect 4491 22996 4492 23036
rect 4532 22996 4533 23036
rect 4491 22987 4533 22996
rect 4492 22902 4532 22987
rect 2763 22868 2805 22877
rect 2763 22828 2764 22868
rect 2804 22828 2805 22868
rect 2763 22819 2805 22828
rect 2955 22868 2997 22877
rect 2955 22828 2956 22868
rect 2996 22828 2997 22868
rect 2955 22819 2997 22828
rect 3148 22868 3188 22877
rect 4300 22868 4340 22877
rect 3188 22828 3668 22868
rect 3148 22819 3188 22828
rect 2764 22734 2804 22819
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 2667 22364 2709 22373
rect 2667 22324 2668 22364
rect 2708 22324 2709 22364
rect 2667 22315 2709 22324
rect 3243 22364 3285 22373
rect 3243 22324 3244 22364
rect 3284 22324 3285 22364
rect 3243 22315 3285 22324
rect 2379 22280 2421 22289
rect 2379 22240 2380 22280
rect 2420 22240 2421 22280
rect 2379 22231 2421 22240
rect 3244 22280 3284 22315
rect 2380 22146 2420 22231
rect 3244 22229 3284 22240
rect 3628 22280 3668 22828
rect 3820 22828 4300 22868
rect 3723 22364 3765 22373
rect 3723 22324 3724 22364
rect 3764 22324 3765 22364
rect 3723 22315 3765 22324
rect 3628 22231 3668 22240
rect 651 21608 693 21617
rect 651 21568 652 21608
rect 692 21568 693 21608
rect 651 21559 693 21568
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 652 20936 692 20945
rect 652 20777 692 20896
rect 651 20768 693 20777
rect 651 20728 652 20768
rect 692 20728 693 20768
rect 651 20719 693 20728
rect 75 20096 117 20105
rect 75 20056 76 20096
rect 116 20056 117 20096
rect 75 20047 117 20056
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 652 19794 692 19879
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 3724 19517 3764 22315
rect 3820 22280 3860 22828
rect 4300 22819 4340 22828
rect 4107 22700 4149 22709
rect 4107 22660 4108 22700
rect 4148 22660 4149 22700
rect 4107 22651 4149 22660
rect 3820 22231 3860 22240
rect 4108 21608 4148 22651
rect 4203 22364 4245 22373
rect 4203 22324 4204 22364
rect 4244 22324 4245 22364
rect 4203 22315 4245 22324
rect 4204 22280 4244 22315
rect 5068 22289 5108 25255
rect 5836 25170 5876 25255
rect 9100 24473 9140 29128
rect 10156 27665 10196 29791
rect 10252 29336 10292 29800
rect 10540 29791 10580 29800
rect 10924 29840 10964 31144
rect 11116 31135 11156 31144
rect 10924 29791 10964 29800
rect 10252 29287 10292 29296
rect 11020 29672 11060 29681
rect 11020 29177 11060 29632
rect 11019 29168 11061 29177
rect 11019 29128 11020 29168
rect 11060 29128 11061 29168
rect 11019 29119 11061 29128
rect 11212 28916 11252 28925
rect 9771 27656 9813 27665
rect 9771 27616 9772 27656
rect 9812 27616 9813 27656
rect 9771 27607 9813 27616
rect 10155 27656 10197 27665
rect 10155 27616 10156 27656
rect 10196 27616 10197 27656
rect 10155 27607 10197 27616
rect 11116 27656 11156 27665
rect 9772 27522 9812 27607
rect 9484 27404 9524 27413
rect 9484 26489 9524 27364
rect 11116 27068 11156 27616
rect 11212 27656 11252 28876
rect 11212 27607 11252 27616
rect 11116 27019 11156 27028
rect 9579 26816 9621 26825
rect 9579 26776 9580 26816
rect 9620 26776 9621 26816
rect 9579 26767 9621 26776
rect 10155 26816 10197 26825
rect 10155 26776 10156 26816
rect 10196 26776 10197 26816
rect 10155 26767 10197 26776
rect 11020 26816 11060 26825
rect 11212 26816 11252 26825
rect 11308 26816 11348 32656
rect 11787 31940 11829 31949
rect 11787 31900 11788 31940
rect 11828 31900 11829 31940
rect 11787 31891 11829 31900
rect 11788 31352 11828 31891
rect 12075 31520 12117 31529
rect 12075 31480 12076 31520
rect 12116 31480 12117 31520
rect 12075 31471 12117 31480
rect 11788 31303 11828 31312
rect 11883 29168 11925 29177
rect 11883 29128 11884 29168
rect 11924 29128 11925 29168
rect 11883 29119 11925 29128
rect 11884 29034 11924 29119
rect 11596 27656 11636 27665
rect 11404 27572 11444 27581
rect 11596 27572 11636 27616
rect 11444 27532 11636 27572
rect 11404 27523 11444 27532
rect 9483 26480 9525 26489
rect 9483 26440 9484 26480
rect 9524 26440 9525 26480
rect 9483 26431 9525 26440
rect 9484 26312 9524 26321
rect 9580 26312 9620 26767
rect 10156 26682 10196 26767
rect 10828 26648 10868 26657
rect 11020 26648 11060 26776
rect 9524 26272 9620 26312
rect 10252 26608 10828 26648
rect 10868 26608 11060 26648
rect 11116 26776 11212 26816
rect 11252 26776 11348 26816
rect 9484 26263 9524 26272
rect 10060 26144 10100 26153
rect 10252 26144 10292 26608
rect 10828 26599 10868 26608
rect 11116 26480 11156 26776
rect 11212 26767 11252 26776
rect 10100 26104 10292 26144
rect 10444 26440 11156 26480
rect 11883 26480 11925 26489
rect 11883 26440 11884 26480
rect 11924 26440 11925 26480
rect 10444 26144 10484 26440
rect 11883 26431 11925 26440
rect 10540 26228 10580 26237
rect 11691 26228 11733 26237
rect 10580 26188 10868 26228
rect 10540 26179 10580 26188
rect 10060 26095 10100 26104
rect 10444 26095 10484 26104
rect 10828 26144 10868 26188
rect 11691 26188 11692 26228
rect 11732 26188 11733 26228
rect 11691 26179 11733 26188
rect 10828 26095 10868 26104
rect 11692 26094 11732 26179
rect 11500 25892 11540 25901
rect 11404 25304 11444 25313
rect 11500 25304 11540 25852
rect 11444 25264 11540 25304
rect 11787 25304 11829 25313
rect 11787 25264 11788 25304
rect 11828 25264 11829 25304
rect 11404 25255 11444 25264
rect 11787 25255 11829 25264
rect 11788 25170 11828 25255
rect 11884 24632 11924 26431
rect 12076 26144 12116 31471
rect 14379 30428 14421 30437
rect 14379 30388 14380 30428
rect 14420 30388 14421 30428
rect 14379 30379 14421 30388
rect 14380 29840 14420 30379
rect 14380 29791 14420 29800
rect 14764 29840 14804 32740
rect 15627 32731 15669 32740
rect 15435 30680 15477 30689
rect 15435 30640 15436 30680
rect 15476 30640 15477 30680
rect 15435 30631 15477 30640
rect 15436 30596 15476 30631
rect 15436 30545 15476 30556
rect 15243 30428 15285 30437
rect 15243 30388 15244 30428
rect 15284 30388 15285 30428
rect 15243 30379 15285 30388
rect 15244 30294 15284 30379
rect 15628 29840 15668 32731
rect 16108 32201 16148 32908
rect 17067 32948 17109 32957
rect 17067 32908 17068 32948
rect 17108 32908 17109 32948
rect 17067 32899 17109 32908
rect 17068 32780 17108 32899
rect 16972 32740 17108 32780
rect 16107 32192 16149 32201
rect 16107 32152 16108 32192
rect 16148 32152 16149 32192
rect 16107 32143 16149 32152
rect 16972 32192 17012 32740
rect 16972 32143 17012 32152
rect 17163 32192 17205 32201
rect 17163 32152 17164 32192
rect 17204 32152 17205 32192
rect 17163 32143 17205 32152
rect 17067 31940 17109 31949
rect 17067 31900 17068 31940
rect 17108 31900 17109 31940
rect 17067 31891 17109 31900
rect 17068 31806 17108 31891
rect 17164 31613 17204 32143
rect 17739 31940 17781 31949
rect 17739 31900 17740 31940
rect 17780 31900 17781 31940
rect 17739 31891 17781 31900
rect 17163 31604 17205 31613
rect 17163 31564 17164 31604
rect 17204 31564 17205 31604
rect 17163 31555 17205 31564
rect 17260 30689 17300 30774
rect 16203 30680 16245 30689
rect 16203 30640 16204 30680
rect 16244 30640 16245 30680
rect 16203 30631 16245 30640
rect 16876 30680 16916 30689
rect 16204 30546 16244 30631
rect 16395 30260 16437 30269
rect 16395 30220 16396 30260
rect 16436 30220 16437 30260
rect 16395 30211 16437 30220
rect 14804 29800 15092 29840
rect 14764 29791 14804 29800
rect 15052 29336 15092 29800
rect 15628 29791 15668 29800
rect 15052 29177 15092 29296
rect 15051 29168 15093 29177
rect 15051 29128 15052 29168
rect 15092 29128 15093 29168
rect 15051 29119 15093 29128
rect 15436 29168 15476 29177
rect 15819 29168 15861 29177
rect 15476 29128 15764 29168
rect 15436 29119 15476 29128
rect 15243 29084 15285 29093
rect 15243 29044 15244 29084
rect 15284 29044 15380 29084
rect 15243 29035 15285 29044
rect 15244 28950 15284 29035
rect 12268 27404 12308 27413
rect 12268 26237 12308 27364
rect 12267 26228 12309 26237
rect 12267 26188 12268 26228
rect 12308 26188 12309 26228
rect 12267 26179 12309 26188
rect 12076 25313 12116 26104
rect 12940 26144 12980 26153
rect 12075 25304 12117 25313
rect 12075 25264 12076 25304
rect 12116 25264 12117 25304
rect 12075 25255 12117 25264
rect 12652 25304 12692 25313
rect 12940 25304 12980 26104
rect 12692 25264 12980 25304
rect 14092 25892 14132 25901
rect 12652 25255 12692 25264
rect 12748 24716 12788 25264
rect 12748 24667 12788 24676
rect 13804 25136 13844 25145
rect 13804 24641 13844 25096
rect 14092 24725 14132 25852
rect 14091 24716 14133 24725
rect 14091 24676 14092 24716
rect 14132 24676 14133 24716
rect 14091 24667 14133 24676
rect 11884 24583 11924 24592
rect 13803 24632 13845 24641
rect 13803 24592 13804 24632
rect 13844 24592 13845 24632
rect 13803 24583 13845 24592
rect 15243 24632 15285 24641
rect 15243 24592 15244 24632
rect 15284 24592 15285 24632
rect 15243 24583 15285 24592
rect 15244 24498 15284 24583
rect 9099 24464 9141 24473
rect 9099 24424 9100 24464
rect 9140 24424 9141 24464
rect 9099 24415 9141 24424
rect 12171 24464 12213 24473
rect 12171 24424 12172 24464
rect 12212 24424 12213 24464
rect 12171 24415 12213 24424
rect 14859 24464 14901 24473
rect 14859 24424 14860 24464
rect 14900 24424 14901 24464
rect 14859 24415 14901 24424
rect 9100 23960 9140 24415
rect 12172 24330 12212 24415
rect 9100 23920 9332 23960
rect 6124 23120 6164 23129
rect 5451 23036 5493 23045
rect 5451 22996 5452 23036
rect 5492 22996 5493 23036
rect 5451 22987 5493 22996
rect 5452 22868 5492 22987
rect 4204 22229 4244 22240
rect 5067 22280 5109 22289
rect 5067 22240 5068 22280
rect 5108 22240 5109 22280
rect 5067 22231 5109 22240
rect 5068 22146 5108 22231
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 4492 21608 4532 21617
rect 4108 21568 4492 21608
rect 4492 21559 4532 21568
rect 4684 21608 4724 21617
rect 4684 21524 4724 21568
rect 4684 21484 5108 21524
rect 4588 21356 4628 21365
rect 4628 21316 4820 21356
rect 4588 21307 4628 21316
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 4780 20189 4820 21316
rect 5068 20768 5108 21484
rect 5452 20768 5492 22828
rect 6124 22532 6164 23080
rect 6220 22532 6260 22541
rect 6124 22492 6220 22532
rect 6220 22483 6260 22492
rect 8044 21608 8084 21617
rect 8044 21029 8084 21568
rect 8427 21608 8469 21617
rect 8427 21568 8428 21608
rect 8468 21568 8469 21608
rect 8427 21559 8469 21568
rect 9292 21608 9332 23920
rect 9963 22280 10005 22289
rect 9963 22240 9964 22280
rect 10004 22240 10005 22280
rect 9963 22231 10005 22240
rect 13996 22280 14036 22289
rect 9964 22146 10004 22231
rect 13612 22196 13652 22205
rect 9484 22112 9524 22121
rect 9484 21617 9524 22072
rect 13612 21776 13652 22156
rect 13708 21776 13748 21785
rect 13612 21736 13708 21776
rect 13708 21727 13748 21736
rect 9292 21559 9332 21568
rect 9483 21608 9525 21617
rect 9483 21568 9484 21608
rect 9524 21568 9525 21608
rect 9483 21559 9525 21568
rect 10443 21608 10485 21617
rect 10443 21568 10444 21608
rect 10484 21568 10485 21608
rect 10443 21559 10485 21568
rect 11019 21608 11061 21617
rect 11019 21568 11020 21608
rect 11060 21568 11061 21608
rect 11019 21559 11061 21568
rect 11787 21608 11829 21617
rect 11787 21568 11788 21608
rect 11828 21568 11829 21608
rect 11787 21559 11829 21568
rect 12267 21608 12309 21617
rect 12267 21568 12268 21608
rect 12308 21568 12309 21608
rect 12267 21559 12309 21568
rect 13035 21608 13077 21617
rect 13035 21568 13036 21608
rect 13076 21568 13077 21608
rect 13035 21559 13077 21568
rect 8428 21474 8468 21559
rect 5835 21020 5877 21029
rect 5835 20980 5836 21020
rect 5876 20980 5877 21020
rect 5835 20971 5877 20980
rect 8043 21020 8085 21029
rect 8043 20980 8044 21020
rect 8084 20980 8085 21020
rect 8043 20971 8085 20980
rect 5836 20886 5876 20971
rect 5644 20768 5684 20777
rect 5068 20728 5644 20768
rect 5644 20719 5684 20728
rect 5548 20600 5588 20609
rect 4779 20180 4821 20189
rect 4779 20140 4780 20180
rect 4820 20140 4821 20180
rect 4779 20131 4821 20140
rect 5163 20180 5205 20189
rect 5163 20140 5164 20180
rect 5204 20140 5205 20180
rect 5163 20131 5205 20140
rect 5356 20180 5396 20189
rect 4492 20096 4532 20105
rect 4012 20056 4492 20096
rect 2667 19508 2709 19517
rect 2667 19468 2668 19508
rect 2708 19468 2709 19508
rect 2667 19459 2709 19468
rect 3723 19508 3765 19517
rect 3723 19468 3724 19508
rect 3764 19468 3765 19508
rect 3723 19459 3765 19468
rect 652 19424 692 19433
rect 652 19097 692 19384
rect 651 19088 693 19097
rect 651 19048 652 19088
rect 692 19048 693 19088
rect 651 19039 693 19048
rect 2283 19088 2325 19097
rect 2283 19048 2284 19088
rect 2324 19048 2325 19088
rect 2283 19039 2325 19048
rect 2284 18668 2324 19039
rect 2284 18619 2324 18628
rect 2668 18584 2708 19459
rect 3724 19374 3764 19459
rect 3147 19340 3189 19349
rect 3147 19300 3148 19340
rect 3188 19300 3189 19340
rect 3147 19291 3189 19300
rect 2763 19256 2805 19265
rect 2763 19216 2764 19256
rect 2804 19216 2805 19256
rect 2763 19207 2805 19216
rect 652 18416 692 18425
rect 652 18257 692 18376
rect 651 18248 693 18257
rect 651 18208 652 18248
rect 692 18208 693 18248
rect 651 18199 693 18208
rect 652 17912 692 17921
rect 652 17417 692 17872
rect 2572 17744 2612 17753
rect 2668 17744 2708 18544
rect 2612 17704 2708 17744
rect 2572 17695 2612 17704
rect 2188 17660 2228 17669
rect 651 17408 693 17417
rect 651 17368 652 17408
rect 692 17368 693 17408
rect 651 17359 693 17368
rect 2188 17249 2228 17620
rect 2187 17240 2229 17249
rect 2187 17200 2188 17240
rect 2228 17200 2229 17240
rect 2187 17191 2229 17200
rect 652 16904 692 16913
rect 652 16577 692 16864
rect 651 16568 693 16577
rect 651 16528 652 16568
rect 692 16528 693 16568
rect 651 16519 693 16528
rect 652 16400 692 16409
rect 556 16360 652 16400
rect 556 15737 596 16360
rect 652 16351 692 16360
rect 555 15728 597 15737
rect 555 15688 556 15728
rect 596 15688 597 15728
rect 555 15679 597 15688
rect 652 15728 692 15737
rect 652 14897 692 15688
rect 651 14888 693 14897
rect 651 14848 652 14888
rect 692 14848 693 14888
rect 651 14839 693 14848
rect 652 14552 692 14561
rect 652 14057 692 14512
rect 2764 14057 2804 19207
rect 3148 19206 3188 19291
rect 3435 19256 3477 19265
rect 3435 19216 3436 19256
rect 3476 19216 3477 19256
rect 3435 19207 3477 19216
rect 3436 19122 3476 19207
rect 2955 19088 2997 19097
rect 2955 19048 2956 19088
rect 2996 19048 2997 19088
rect 2955 19039 2997 19048
rect 2956 18954 2996 19039
rect 3532 18584 3572 18593
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 3435 17744 3477 17753
rect 3532 17744 3572 18544
rect 3435 17704 3436 17744
rect 3476 17704 3572 17744
rect 3435 17695 3477 17704
rect 3436 17610 3476 17695
rect 3051 17240 3093 17249
rect 3051 17200 3052 17240
rect 3092 17200 3093 17240
rect 3051 17191 3093 17200
rect 4012 17240 4052 20056
rect 4492 20047 4532 20056
rect 4684 20096 4724 20105
rect 4587 20012 4629 20021
rect 4587 19972 4588 20012
rect 4628 19972 4629 20012
rect 4587 19963 4629 19972
rect 4588 19878 4628 19963
rect 4684 19433 4724 20056
rect 4876 20096 4916 20107
rect 4876 20021 4916 20056
rect 5164 20096 5204 20131
rect 5164 20045 5204 20056
rect 4875 20012 4917 20021
rect 4875 19972 4876 20012
rect 4916 19972 4917 20012
rect 4875 19963 4917 19972
rect 4683 19424 4725 19433
rect 4683 19384 4684 19424
rect 4724 19384 4725 19424
rect 4683 19375 4725 19384
rect 5259 19340 5301 19349
rect 5259 19300 5260 19340
rect 5300 19300 5301 19340
rect 5259 19291 5301 19300
rect 4396 19256 4436 19265
rect 4396 19097 4436 19216
rect 4588 19256 4628 19265
rect 4628 19216 4820 19256
rect 4588 19207 4628 19216
rect 4395 19088 4437 19097
rect 4395 19048 4396 19088
rect 4436 19048 4437 19088
rect 4395 19039 4437 19048
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 4684 18752 4724 18761
rect 4780 18752 4820 19216
rect 5260 19206 5300 19291
rect 5356 19265 5396 20140
rect 5548 19349 5588 20560
rect 5547 19340 5589 19349
rect 5547 19300 5548 19340
rect 5588 19300 5589 19340
rect 5547 19291 5589 19300
rect 5355 19256 5397 19265
rect 5355 19216 5356 19256
rect 5396 19216 5397 19256
rect 5355 19207 5397 19216
rect 7371 19256 7413 19265
rect 7371 19216 7372 19256
rect 7412 19216 7413 19256
rect 7371 19207 7413 19216
rect 7756 19256 7796 19265
rect 7372 19122 7412 19207
rect 7756 19097 7796 19216
rect 8620 19256 8660 19265
rect 7755 19088 7797 19097
rect 7755 19048 7756 19088
rect 7796 19048 7797 19088
rect 7755 19039 7797 19048
rect 4724 18712 4820 18752
rect 4684 18703 4724 18712
rect 8620 17837 8660 19216
rect 9484 19181 9524 21559
rect 10444 21524 10484 21559
rect 10444 21473 10484 21484
rect 11020 21474 11060 21559
rect 11692 21356 11732 21365
rect 11403 20768 11445 20777
rect 11403 20728 11404 20768
rect 11444 20728 11445 20768
rect 11403 20719 11445 20728
rect 11596 20768 11636 20777
rect 11692 20768 11732 21316
rect 11636 20728 11732 20768
rect 11788 20768 11828 21559
rect 11596 20719 11636 20728
rect 11788 20719 11828 20728
rect 12171 20768 12213 20777
rect 12171 20728 12172 20768
rect 12212 20728 12213 20768
rect 12171 20719 12213 20728
rect 11404 20634 11444 20719
rect 11500 20684 11540 20693
rect 11500 20432 11540 20644
rect 12172 20516 12212 20719
rect 12268 20684 12308 21559
rect 13036 21474 13076 21559
rect 13996 21449 14036 22240
rect 14763 22280 14805 22289
rect 14763 22240 14764 22280
rect 14804 22240 14805 22280
rect 14763 22231 14805 22240
rect 14860 22280 14900 24415
rect 14860 22231 14900 22240
rect 14764 22037 14804 22231
rect 15340 22037 15380 29044
rect 15724 28664 15764 29128
rect 15819 29128 15820 29168
rect 15860 29128 15861 29168
rect 15819 29119 15861 29128
rect 15820 29034 15860 29119
rect 15724 28624 16244 28664
rect 16204 28580 16244 28624
rect 16204 28531 16244 28540
rect 16396 28412 16436 30211
rect 16780 30092 16820 30101
rect 16876 30092 16916 30640
rect 17067 30680 17109 30689
rect 17067 30640 17068 30680
rect 17108 30640 17109 30680
rect 17067 30631 17109 30640
rect 17259 30680 17301 30689
rect 17259 30640 17260 30680
rect 17300 30640 17301 30680
rect 17259 30631 17301 30640
rect 17452 30680 17492 30689
rect 17068 30546 17108 30631
rect 17164 30512 17204 30521
rect 17452 30512 17492 30640
rect 17740 30680 17780 31891
rect 18124 31613 18164 33412
rect 18220 33403 18260 33412
rect 18232 33284 18600 33293
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18232 33235 18600 33244
rect 20523 32864 20565 32873
rect 20523 32824 20524 32864
rect 20564 32824 20565 32864
rect 20523 32815 20565 32824
rect 19472 32528 19840 32537
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19472 32479 19840 32488
rect 18232 31772 18600 31781
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18232 31723 18600 31732
rect 18123 31604 18165 31613
rect 18123 31564 18124 31604
rect 18164 31564 18165 31604
rect 18123 31555 18165 31564
rect 18315 31604 18357 31613
rect 18315 31564 18316 31604
rect 18356 31564 18357 31604
rect 18315 31555 18357 31564
rect 18220 30848 18260 30857
rect 17931 30764 17973 30773
rect 17931 30724 17932 30764
rect 17972 30724 17973 30764
rect 17931 30715 17973 30724
rect 17740 30631 17780 30640
rect 17932 30630 17972 30715
rect 18220 30689 18260 30808
rect 18219 30680 18261 30689
rect 18219 30640 18220 30680
rect 18260 30640 18261 30680
rect 18219 30631 18261 30640
rect 18316 30680 18356 31555
rect 19472 31016 19840 31025
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19472 30967 19840 30976
rect 20139 30764 20181 30773
rect 20139 30724 20140 30764
rect 20180 30724 20181 30764
rect 20139 30715 20181 30724
rect 18316 30631 18356 30640
rect 20140 30630 20180 30715
rect 20524 30680 20564 32815
rect 17204 30472 17492 30512
rect 17164 30463 17204 30472
rect 18508 30428 18548 30437
rect 18548 30388 18740 30428
rect 18508 30379 18548 30388
rect 17259 30260 17301 30269
rect 17259 30220 17260 30260
rect 17300 30220 17301 30260
rect 17259 30211 17301 30220
rect 18232 30260 18600 30269
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18232 30211 18600 30220
rect 16820 30052 16916 30092
rect 17260 30092 17300 30211
rect 16780 30043 16820 30052
rect 17260 30043 17300 30052
rect 18700 29933 18740 30388
rect 20524 30017 20564 30640
rect 20523 30008 20565 30017
rect 20523 29968 20524 30008
rect 20564 29968 20565 30008
rect 20523 29959 20565 29968
rect 18699 29924 18741 29933
rect 18699 29884 18700 29924
rect 18740 29884 18741 29924
rect 18699 29875 18741 29884
rect 17932 29840 17972 29849
rect 17836 29336 17876 29345
rect 17932 29336 17972 29800
rect 19472 29504 19840 29513
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19472 29455 19840 29464
rect 17876 29296 17972 29336
rect 17836 29287 17876 29296
rect 16683 29168 16725 29177
rect 16683 29128 16684 29168
rect 16724 29128 16725 29168
rect 16683 29119 16725 29128
rect 19275 29168 19317 29177
rect 19275 29128 19276 29168
rect 19316 29128 19317 29168
rect 19275 29119 19317 29128
rect 16684 29034 16724 29119
rect 18232 28748 18600 28757
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18232 28699 18600 28708
rect 16396 28363 16436 28372
rect 19276 28412 19316 29119
rect 20620 29000 20660 37519
rect 20716 37484 20756 37493
rect 20756 37444 20948 37484
rect 20716 37435 20756 37444
rect 20908 37400 20948 37444
rect 20908 37351 20948 37360
rect 25420 37400 25460 37409
rect 35595 37400 35637 37409
rect 25460 37360 26036 37400
rect 25420 37351 25460 37360
rect 21580 37232 21620 37241
rect 21484 37192 21580 37232
rect 21388 36728 21428 36737
rect 21196 36644 21236 36653
rect 21388 36644 21428 36688
rect 21236 36604 21428 36644
rect 21196 36595 21236 36604
rect 21484 36140 21524 37192
rect 21580 37183 21620 37192
rect 24748 37232 24788 37241
rect 24556 36728 24596 36737
rect 23979 36560 24021 36569
rect 23979 36520 23980 36560
rect 24020 36520 24021 36560
rect 23979 36511 24021 36520
rect 22060 36476 22100 36485
rect 22100 36436 22196 36476
rect 22060 36427 22100 36436
rect 21292 36100 21524 36140
rect 21292 35897 21332 36100
rect 22156 35981 22196 36436
rect 22155 35972 22197 35981
rect 22155 35932 22156 35972
rect 22196 35932 22197 35972
rect 22155 35923 22197 35932
rect 23212 35972 23252 35983
rect 21291 35888 21333 35897
rect 21291 35848 21292 35888
rect 21332 35848 21333 35888
rect 21291 35839 21333 35848
rect 21483 35888 21525 35897
rect 21483 35848 21484 35888
rect 21524 35848 21525 35888
rect 21483 35839 21525 35848
rect 22156 35888 22196 35923
rect 23212 35897 23252 35932
rect 21292 35216 21332 35839
rect 21292 35167 21332 35176
rect 21484 35216 21524 35839
rect 22156 35837 22196 35848
rect 22348 35888 22388 35897
rect 22252 35804 22292 35813
rect 22252 35468 22292 35764
rect 22060 35428 22292 35468
rect 21484 35167 21524 35176
rect 21676 35216 21716 35225
rect 21388 35048 21428 35057
rect 21676 35048 21716 35176
rect 22060 35216 22100 35428
rect 22348 35309 22388 35848
rect 23211 35888 23253 35897
rect 23211 35848 23212 35888
rect 23252 35848 23253 35888
rect 23211 35839 23253 35848
rect 23980 35888 24020 36511
rect 23596 35804 23636 35813
rect 23404 35720 23444 35729
rect 23596 35720 23636 35764
rect 23444 35680 23636 35720
rect 23404 35671 23444 35680
rect 22060 35167 22100 35176
rect 22156 35300 22196 35309
rect 21428 35008 21716 35048
rect 21388 34999 21428 35008
rect 20812 34376 20852 34385
rect 20812 34049 20852 34336
rect 20811 34040 20853 34049
rect 22156 34040 22196 35260
rect 22347 35300 22389 35309
rect 22347 35260 22348 35300
rect 22388 35260 22389 35300
rect 22347 35251 22389 35260
rect 23019 34208 23061 34217
rect 23019 34168 23020 34208
rect 23060 34168 23061 34208
rect 23019 34159 23061 34168
rect 20811 34000 20812 34040
rect 20852 34000 20853 34040
rect 20811 33991 20853 34000
rect 21772 34000 22196 34040
rect 22347 34040 22389 34049
rect 22347 34000 22348 34040
rect 22388 34000 22389 34040
rect 21772 32864 21812 34000
rect 22347 33991 22389 34000
rect 21772 32815 21812 32824
rect 22155 32864 22197 32873
rect 22155 32824 22156 32864
rect 22196 32824 22197 32864
rect 22155 32815 22197 32824
rect 22156 32730 22196 32815
rect 22348 31520 22388 33991
rect 23020 32864 23060 34159
rect 23980 32873 24020 35848
rect 24556 35048 24596 36688
rect 24748 35897 24788 37192
rect 24940 36737 24980 36822
rect 24939 36728 24981 36737
rect 24939 36688 24940 36728
rect 24980 36688 24981 36728
rect 24939 36679 24981 36688
rect 25804 36728 25844 36737
rect 25804 36569 25844 36688
rect 24939 36560 24981 36569
rect 24939 36520 24940 36560
rect 24980 36520 24981 36560
rect 24939 36511 24981 36520
rect 25803 36560 25845 36569
rect 25803 36520 25804 36560
rect 25844 36520 25845 36560
rect 25803 36511 25845 36520
rect 24747 35888 24789 35897
rect 24747 35848 24748 35888
rect 24788 35848 24789 35888
rect 24747 35839 24789 35848
rect 24844 35888 24884 35897
rect 24940 35888 24980 36511
rect 25996 36140 26036 37360
rect 35595 37360 35596 37400
rect 35636 37360 35637 37400
rect 35595 37351 35637 37360
rect 36460 37400 36500 37409
rect 35212 37316 35252 37325
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 32812 36728 32852 36737
rect 32620 36688 32812 36728
rect 31372 36644 31412 36655
rect 31372 36569 31412 36604
rect 30219 36560 30261 36569
rect 30219 36520 30220 36560
rect 30260 36520 30261 36560
rect 30219 36511 30261 36520
rect 31179 36560 31221 36569
rect 31179 36520 31180 36560
rect 31220 36520 31221 36560
rect 31179 36511 31221 36520
rect 31371 36560 31413 36569
rect 31371 36520 31372 36560
rect 31412 36520 31413 36560
rect 31371 36511 31413 36520
rect 32139 36560 32181 36569
rect 32139 36520 32140 36560
rect 32180 36520 32181 36560
rect 32139 36511 32181 36520
rect 25996 36091 26036 36100
rect 26956 36476 26996 36485
rect 24884 35848 24980 35888
rect 24844 35839 24884 35848
rect 24843 35300 24885 35309
rect 24843 35260 24844 35300
rect 24884 35260 24885 35300
rect 24843 35251 24885 35260
rect 24844 35132 24884 35251
rect 24844 35083 24884 35092
rect 24652 35048 24692 35057
rect 24556 35008 24652 35048
rect 24652 34999 24692 35008
rect 24555 34040 24597 34049
rect 24555 34000 24556 34040
rect 24596 34000 24597 34040
rect 24555 33991 24597 34000
rect 24267 33704 24309 33713
rect 24267 33664 24268 33704
rect 24308 33664 24309 33704
rect 24267 33655 24309 33664
rect 24556 33704 24596 33991
rect 24940 33704 24980 35848
rect 25227 35888 25269 35897
rect 25227 35848 25228 35888
rect 25268 35848 25269 35888
rect 25227 35839 25269 35848
rect 26860 35888 26900 35897
rect 26956 35888 26996 36436
rect 26900 35848 26996 35888
rect 30220 35888 30260 36511
rect 31180 36426 31220 36511
rect 32140 36426 32180 36511
rect 32620 36140 32660 36688
rect 32812 36679 32852 36688
rect 33099 36560 33141 36569
rect 33099 36520 33100 36560
rect 33140 36520 33141 36560
rect 33099 36511 33141 36520
rect 32620 36091 32660 36100
rect 26860 35839 26900 35848
rect 30220 35839 30260 35848
rect 30604 35888 30644 35897
rect 31468 35888 31508 35897
rect 30644 35848 30740 35888
rect 30604 35839 30644 35848
rect 25228 35384 25268 35839
rect 25228 35335 25268 35344
rect 26188 35720 26228 35729
rect 26188 35309 26228 35680
rect 25323 35300 25365 35309
rect 25323 35260 25324 35300
rect 25364 35260 25365 35300
rect 25323 35251 25365 35260
rect 26187 35300 26229 35309
rect 26187 35260 26188 35300
rect 26228 35260 26229 35300
rect 26187 35251 26229 35260
rect 25324 35216 25364 35251
rect 25324 35165 25364 35176
rect 25516 34964 25556 34973
rect 25035 33704 25077 33713
rect 24940 33664 25036 33704
rect 25076 33664 25077 33704
rect 24556 33655 24596 33664
rect 25035 33655 25077 33664
rect 24268 33570 24308 33655
rect 25036 33452 25076 33655
rect 25036 32873 25076 33412
rect 23020 32815 23060 32824
rect 23979 32864 24021 32873
rect 23979 32824 23980 32864
rect 24020 32824 24021 32864
rect 23979 32815 24021 32824
rect 25035 32864 25077 32873
rect 25035 32824 25036 32864
rect 25076 32824 25077 32864
rect 25516 32864 25556 34924
rect 30315 34964 30357 34973
rect 30315 34924 30316 34964
rect 30356 34924 30357 34964
rect 30315 34915 30357 34924
rect 30316 34376 30356 34915
rect 30700 34385 30740 35848
rect 31508 35848 31604 35888
rect 31468 35839 31508 35848
rect 31467 35132 31509 35141
rect 31467 35092 31468 35132
rect 31508 35092 31509 35132
rect 31467 35083 31509 35092
rect 31468 34998 31508 35083
rect 31275 34964 31317 34973
rect 31275 34924 31276 34964
rect 31316 34924 31317 34964
rect 31275 34915 31317 34924
rect 31276 34830 31316 34915
rect 30316 34327 30356 34336
rect 30699 34376 30741 34385
rect 30699 34336 30700 34376
rect 30740 34336 30741 34376
rect 30699 34327 30741 34336
rect 31564 34376 31604 35848
rect 32908 35216 32948 35225
rect 32716 35176 32908 35216
rect 32235 35132 32277 35141
rect 32235 35092 32236 35132
rect 32276 35092 32277 35132
rect 32235 35083 32277 35092
rect 32236 34998 32276 35083
rect 32716 34628 32756 35176
rect 32908 35167 32948 35176
rect 33100 35216 33140 36511
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 35212 36140 35252 37276
rect 35596 37266 35636 37351
rect 36460 36737 36500 37360
rect 36459 36728 36501 36737
rect 36459 36688 36460 36728
rect 36500 36688 36501 36728
rect 36459 36679 36501 36688
rect 36556 36728 36596 36737
rect 36556 36560 36596 36688
rect 36460 36520 36596 36560
rect 35403 36224 35445 36233
rect 35403 36184 35404 36224
rect 35444 36184 35445 36224
rect 35403 36175 35445 36184
rect 36075 36224 36117 36233
rect 36075 36184 36076 36224
rect 36116 36184 36117 36224
rect 36075 36175 36117 36184
rect 35212 36091 35252 36100
rect 35404 35972 35444 36175
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 33100 35167 33140 35176
rect 33195 35216 33237 35225
rect 33195 35176 33196 35216
rect 33236 35176 33237 35216
rect 33195 35167 33237 35176
rect 33292 35216 33332 35227
rect 33196 35082 33236 35167
rect 33292 35141 33332 35176
rect 33291 35132 33333 35141
rect 33291 35092 33292 35132
rect 33332 35092 33333 35132
rect 33291 35083 33333 35092
rect 33771 35132 33813 35141
rect 33771 35092 33772 35132
rect 33812 35092 33813 35132
rect 33771 35083 33813 35092
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 32716 34579 32756 34588
rect 30700 34242 30740 34327
rect 25995 32948 26037 32957
rect 25995 32908 25996 32948
rect 26036 32908 26037 32948
rect 25995 32899 26037 32908
rect 25612 32864 25652 32873
rect 25516 32824 25612 32864
rect 25035 32815 25077 32824
rect 25612 32815 25652 32824
rect 25996 32864 26036 32899
rect 22348 31471 22388 31480
rect 24172 32696 24212 32705
rect 22636 31352 22676 31361
rect 22539 30848 22581 30857
rect 22539 30808 22540 30848
rect 22580 30808 22581 30848
rect 22539 30799 22581 30808
rect 22540 30714 22580 30799
rect 21388 30680 21428 30689
rect 21195 30008 21237 30017
rect 21195 29968 21196 30008
rect 21236 29968 21237 30008
rect 21195 29959 21237 29968
rect 20811 29924 20853 29933
rect 20811 29884 20812 29924
rect 20852 29884 20853 29924
rect 20811 29875 20853 29884
rect 20812 29840 20852 29875
rect 20812 29789 20852 29800
rect 21196 29840 21236 29959
rect 21196 29791 21236 29800
rect 21388 29177 21428 30640
rect 22636 29849 22676 31312
rect 23884 31352 23924 31361
rect 23884 30857 23924 31312
rect 24172 31352 24212 32656
rect 24172 31303 24212 31312
rect 24363 31184 24405 31193
rect 24363 31144 24364 31184
rect 24404 31144 24405 31184
rect 24363 31135 24405 31144
rect 25707 31184 25749 31193
rect 25707 31144 25708 31184
rect 25748 31144 25749 31184
rect 25707 31135 25749 31144
rect 24364 31050 24404 31135
rect 23883 30848 23925 30857
rect 23883 30808 23884 30848
rect 23924 30808 23925 30848
rect 23883 30799 23925 30808
rect 25323 30764 25365 30773
rect 25323 30724 25324 30764
rect 25364 30724 25365 30764
rect 25323 30715 25365 30724
rect 25611 30764 25653 30773
rect 25611 30724 25612 30764
rect 25652 30724 25653 30764
rect 25611 30715 25653 30724
rect 24268 30680 24308 30689
rect 24268 30101 24308 30640
rect 24940 30680 24980 30689
rect 25132 30680 25172 30689
rect 24980 30640 25132 30680
rect 24940 30631 24980 30640
rect 25132 30631 25172 30640
rect 25227 30680 25269 30689
rect 25227 30640 25228 30680
rect 25268 30640 25269 30680
rect 25227 30631 25269 30640
rect 25324 30680 25364 30715
rect 25228 30546 25268 30631
rect 25324 30629 25364 30640
rect 23211 30092 23253 30101
rect 23211 30052 23212 30092
rect 23252 30052 23253 30092
rect 23211 30043 23253 30052
rect 24267 30092 24309 30101
rect 24267 30052 24268 30092
rect 24308 30052 24309 30092
rect 24267 30043 24309 30052
rect 25323 30092 25365 30101
rect 25323 30052 25324 30092
rect 25364 30052 25365 30092
rect 25323 30043 25365 30052
rect 23212 29958 23252 30043
rect 22060 29840 22100 29849
rect 22060 29177 22100 29800
rect 22635 29840 22677 29849
rect 22635 29800 22636 29840
rect 22676 29800 22677 29840
rect 22635 29791 22677 29800
rect 25324 29840 25364 30043
rect 25324 29791 25364 29800
rect 25612 29840 25652 30715
rect 25708 30680 25748 31135
rect 25708 30631 25748 30640
rect 25803 30680 25845 30689
rect 25803 30640 25804 30680
rect 25844 30640 25845 30680
rect 25803 30631 25845 30640
rect 25804 30546 25844 30631
rect 25996 29840 26036 32824
rect 26859 32864 26901 32873
rect 26859 32824 26860 32864
rect 26900 32824 26901 32864
rect 26859 32815 26901 32824
rect 28587 32864 28629 32873
rect 28587 32824 28588 32864
rect 28628 32824 28629 32864
rect 28587 32815 28629 32824
rect 26860 32730 26900 32815
rect 27627 32696 27669 32705
rect 27627 32656 27628 32696
rect 27668 32656 27669 32696
rect 27627 32647 27669 32656
rect 28011 32696 28053 32705
rect 28011 32656 28012 32696
rect 28052 32656 28053 32696
rect 28011 32647 28053 32656
rect 27628 31352 27668 32647
rect 28012 32562 28052 32647
rect 27628 31303 27668 31312
rect 26956 31184 26996 31193
rect 26956 30773 26996 31144
rect 26955 30764 26997 30773
rect 26955 30724 26956 30764
rect 26996 30724 26997 30764
rect 26955 30715 26997 30724
rect 26764 30680 26804 30691
rect 26764 30605 26804 30640
rect 26091 30596 26133 30605
rect 26091 30556 26092 30596
rect 26132 30556 26133 30596
rect 26091 30547 26133 30556
rect 26763 30596 26805 30605
rect 26763 30556 26764 30596
rect 26804 30556 26805 30596
rect 26763 30547 26805 30556
rect 26092 30462 26132 30547
rect 27436 30428 27476 30437
rect 26092 29840 26132 29849
rect 25996 29800 26092 29840
rect 25612 29791 25652 29800
rect 26092 29791 26132 29800
rect 27051 29840 27093 29849
rect 27051 29800 27052 29840
rect 27092 29800 27093 29840
rect 27051 29791 27093 29800
rect 27340 29840 27380 29849
rect 27436 29840 27476 30388
rect 27380 29800 27476 29840
rect 27723 29840 27765 29849
rect 27723 29800 27724 29840
rect 27764 29800 27765 29840
rect 27340 29791 27380 29800
rect 27723 29791 27765 29800
rect 28588 29840 28628 32815
rect 31180 31352 31220 31361
rect 30412 31312 31180 31352
rect 30412 30848 30452 31312
rect 31180 31303 31220 31312
rect 30412 30799 30452 30808
rect 30508 31184 30548 31193
rect 29740 29924 29780 29933
rect 29780 29884 30068 29924
rect 29740 29875 29780 29884
rect 28588 29791 28628 29800
rect 28971 29840 29013 29849
rect 28971 29800 28972 29840
rect 29012 29800 29013 29840
rect 28971 29791 29013 29800
rect 30028 29840 30068 29884
rect 30028 29791 30068 29800
rect 30412 29840 30452 29849
rect 30508 29840 30548 31144
rect 31564 30689 31604 34336
rect 32427 34376 32469 34385
rect 32427 34336 32428 34376
rect 32468 34336 32469 34376
rect 32427 34327 32469 34336
rect 32428 31361 32468 34327
rect 33772 34208 33812 35083
rect 35404 34385 35444 35932
rect 36076 35888 36116 36175
rect 36460 36140 36500 36520
rect 36652 36233 36692 37948
rect 37612 37652 37652 38200
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 93832 37820 94200 37829
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 93832 37771 94200 37780
rect 37612 37603 37652 37612
rect 36939 37400 36981 37409
rect 36939 37360 36940 37400
rect 36980 37360 36981 37400
rect 36939 37351 36981 37360
rect 36940 36728 36980 37351
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 95072 37064 95440 37073
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95072 37015 95440 37024
rect 36940 36653 36980 36688
rect 37803 36728 37845 36737
rect 37803 36688 37804 36728
rect 37844 36688 37845 36728
rect 37803 36679 37845 36688
rect 38571 36728 38613 36737
rect 38571 36688 38572 36728
rect 38612 36688 38613 36728
rect 38571 36679 38613 36688
rect 36939 36644 36981 36653
rect 36939 36604 36940 36644
rect 36980 36604 36981 36644
rect 36939 36595 36981 36604
rect 37707 36644 37749 36653
rect 37707 36604 37708 36644
rect 37748 36604 37749 36644
rect 37707 36595 37749 36604
rect 36940 36564 36980 36595
rect 37515 36560 37557 36569
rect 37515 36520 37516 36560
rect 37556 36520 37557 36560
rect 37515 36511 37557 36520
rect 36651 36224 36693 36233
rect 36651 36184 36652 36224
rect 36692 36184 36693 36224
rect 36651 36175 36693 36184
rect 36460 36091 36500 36100
rect 36651 35981 36691 36066
rect 36267 35972 36309 35981
rect 36267 35932 36268 35972
rect 36308 35932 36309 35972
rect 36267 35923 36309 35932
rect 36651 35972 36693 35981
rect 36692 35932 36693 35972
rect 36651 35923 36693 35932
rect 36843 35972 36885 35981
rect 36843 35932 36844 35972
rect 36884 35932 36885 35972
rect 36843 35923 36885 35932
rect 36076 35839 36116 35848
rect 36268 35888 36308 35923
rect 36268 35837 36308 35848
rect 36844 35838 36884 35923
rect 37516 35888 37556 36511
rect 37516 35839 37556 35848
rect 36172 35804 36212 35813
rect 35787 35216 35829 35225
rect 35787 35176 35788 35216
rect 35828 35176 35829 35216
rect 35787 35167 35829 35176
rect 36172 35216 36212 35764
rect 36172 35167 36212 35176
rect 36268 35300 36308 35309
rect 35788 35082 35828 35167
rect 36268 34385 36308 35260
rect 33867 34376 33909 34385
rect 33867 34336 33868 34376
rect 33908 34336 33909 34376
rect 33867 34327 33909 34336
rect 35403 34376 35445 34385
rect 35403 34336 35404 34376
rect 35444 34336 35445 34376
rect 35403 34327 35445 34336
rect 36267 34376 36309 34385
rect 36267 34336 36268 34376
rect 36308 34336 36309 34376
rect 36267 34327 36309 34336
rect 37323 34376 37365 34385
rect 37323 34336 37324 34376
rect 37364 34336 37365 34376
rect 37323 34327 37365 34336
rect 37708 34376 37748 36595
rect 37804 36594 37844 36679
rect 33868 34242 33908 34327
rect 37324 34242 37364 34327
rect 33772 34159 33812 34168
rect 34060 34208 34100 34217
rect 33352 33284 33720 33293
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33352 33235 33720 33244
rect 34060 32780 34100 34168
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 33868 32740 34100 32780
rect 36940 32864 36980 32873
rect 33868 32276 33908 32740
rect 34592 32528 34960 32537
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34592 32479 34960 32488
rect 33868 32227 33908 32236
rect 34251 32276 34293 32285
rect 34251 32236 34252 32276
rect 34292 32236 34293 32276
rect 34251 32227 34293 32236
rect 34252 32192 34292 32227
rect 33352 31772 33720 31781
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33352 31723 33720 31732
rect 34252 31529 34292 32152
rect 35116 32192 35156 32201
rect 33771 31520 33813 31529
rect 33771 31480 33772 31520
rect 33812 31480 33813 31520
rect 33771 31471 33813 31480
rect 34251 31520 34293 31529
rect 34251 31480 34252 31520
rect 34292 31480 34293 31520
rect 34251 31471 34293 31480
rect 33772 31386 33812 31471
rect 32427 31352 32469 31361
rect 32427 31312 32428 31352
rect 32468 31312 32469 31352
rect 32427 31303 32469 31312
rect 33099 31352 33141 31361
rect 33099 31312 33100 31352
rect 33140 31312 33141 31352
rect 33099 31303 33141 31312
rect 34060 31352 34100 31361
rect 31563 30680 31605 30689
rect 31563 30640 31564 30680
rect 31604 30640 31605 30680
rect 31563 30631 31605 30640
rect 32428 30680 32468 31303
rect 33100 31218 33140 31303
rect 32811 30764 32853 30773
rect 32811 30724 32812 30764
rect 32852 30724 32853 30764
rect 32811 30715 32853 30724
rect 32428 30631 32468 30640
rect 31564 30546 31604 30631
rect 32812 30630 32852 30715
rect 33771 30680 33813 30689
rect 33771 30640 33772 30680
rect 33812 30640 33813 30680
rect 33771 30631 33813 30640
rect 33352 30260 33720 30269
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33352 30211 33720 30220
rect 30452 29800 30548 29840
rect 30412 29791 30452 29800
rect 22636 29261 22676 29791
rect 27052 29706 27092 29791
rect 27724 29706 27764 29791
rect 25804 29672 25844 29681
rect 25844 29632 26132 29672
rect 25804 29623 25844 29632
rect 22635 29252 22677 29261
rect 22635 29212 22636 29252
rect 22676 29212 22677 29252
rect 22635 29203 22677 29212
rect 21387 29168 21429 29177
rect 21387 29128 21388 29168
rect 21428 29128 21429 29168
rect 21387 29119 21429 29128
rect 22059 29168 22101 29177
rect 22059 29128 22060 29168
rect 22100 29128 22101 29168
rect 22059 29119 22101 29128
rect 22156 29168 22196 29177
rect 20620 28960 20756 29000
rect 19276 28328 19316 28372
rect 19948 28496 19988 28505
rect 19660 28328 19700 28337
rect 19276 28288 19660 28328
rect 19660 28279 19700 28288
rect 19472 27992 19840 28001
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19472 27943 19840 27952
rect 18232 27236 18600 27245
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18232 27187 18600 27196
rect 19472 26480 19840 26489
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19472 26431 19840 26440
rect 17836 26144 17876 26153
rect 17836 25565 17876 26104
rect 18508 26144 18548 26153
rect 18700 26144 18740 26153
rect 18548 26104 18700 26144
rect 18508 26095 18548 26104
rect 18700 26095 18740 26104
rect 19083 26144 19125 26153
rect 19083 26104 19084 26144
rect 19124 26104 19125 26144
rect 19083 26095 19125 26104
rect 19948 26144 19988 28456
rect 20619 28328 20661 28337
rect 20619 28288 20620 28328
rect 20660 28288 20661 28328
rect 20619 28279 20661 28288
rect 20620 28194 20660 28279
rect 18232 25724 18600 25733
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18232 25675 18600 25684
rect 16875 25556 16917 25565
rect 16875 25516 16876 25556
rect 16916 25516 16917 25556
rect 16875 25507 16917 25516
rect 17835 25556 17877 25565
rect 17835 25516 17836 25556
rect 17876 25516 17877 25556
rect 17835 25507 17877 25516
rect 16876 25422 16916 25507
rect 16588 25304 16628 25313
rect 16588 24800 16628 25264
rect 16684 25304 16724 25313
rect 16724 25264 17012 25304
rect 16684 25255 16724 25264
rect 16588 24751 16628 24760
rect 16972 24716 17012 25264
rect 16972 24667 17012 24676
rect 16108 24632 16148 24641
rect 15915 24464 15957 24473
rect 15915 24424 15916 24464
rect 15956 24424 15957 24464
rect 15915 24415 15957 24424
rect 15916 23960 15956 24415
rect 15820 23920 15956 23960
rect 15436 23792 15476 23803
rect 15436 23717 15476 23752
rect 15820 23792 15860 23920
rect 15820 23743 15860 23752
rect 15915 23792 15957 23801
rect 15915 23752 15916 23792
rect 15956 23752 15957 23792
rect 15915 23743 15957 23752
rect 15435 23708 15477 23717
rect 15435 23668 15436 23708
rect 15476 23668 15477 23708
rect 15435 23659 15477 23668
rect 15916 23708 15956 23743
rect 15916 23657 15956 23668
rect 16011 22532 16053 22541
rect 16011 22492 16012 22532
rect 16052 22492 16053 22532
rect 16011 22483 16053 22492
rect 16012 22398 16052 22483
rect 14763 22028 14805 22037
rect 14763 21988 14764 22028
rect 14804 21988 14805 22028
rect 14763 21979 14805 21988
rect 15339 22028 15381 22037
rect 15339 21988 15340 22028
rect 15380 21988 15381 22028
rect 15339 21979 15381 21988
rect 14764 21608 14804 21979
rect 14764 21559 14804 21568
rect 15723 21608 15765 21617
rect 15723 21568 15724 21608
rect 15764 21568 15765 21608
rect 15723 21559 15765 21568
rect 15724 21474 15764 21559
rect 13995 21440 14037 21449
rect 13995 21400 13996 21440
rect 14036 21400 14037 21440
rect 13995 21391 14037 21400
rect 15243 21440 15285 21449
rect 15243 21400 15244 21440
rect 15284 21400 15285 21440
rect 15243 21391 15285 21400
rect 12748 20768 12788 20777
rect 12268 20635 12308 20644
rect 12460 20728 12748 20768
rect 12172 20476 12308 20516
rect 11500 20392 12212 20432
rect 12076 20096 12116 20105
rect 11404 20056 12076 20096
rect 9483 19172 9525 19181
rect 9483 19132 9484 19172
rect 9524 19132 9525 19172
rect 9483 19123 9525 19132
rect 8619 17828 8661 17837
rect 8619 17788 8620 17828
rect 8660 17788 8661 17828
rect 8619 17779 8661 17788
rect 4203 17744 4245 17753
rect 4203 17704 4204 17744
rect 4244 17704 4245 17744
rect 4203 17695 4245 17704
rect 9004 17744 9044 17753
rect 9484 17744 9524 19123
rect 9771 19088 9813 19097
rect 9771 19048 9772 19088
rect 9812 19048 9813 19088
rect 9771 19039 9813 19048
rect 10731 19088 10773 19097
rect 10731 19048 10732 19088
rect 10772 19048 10773 19088
rect 10731 19039 10773 19048
rect 9772 18954 9812 19039
rect 10732 18584 10772 19039
rect 11212 18752 11252 18761
rect 11404 18752 11444 20056
rect 12076 20047 12116 20056
rect 12172 20096 12212 20392
rect 12172 20047 12212 20056
rect 12172 19508 12212 19517
rect 12268 19508 12308 20476
rect 12460 20012 12500 20728
rect 12748 20719 12788 20728
rect 13996 20768 14036 21391
rect 15244 21306 15284 21391
rect 16012 21020 16052 21029
rect 16108 21020 16148 24592
rect 16395 24632 16437 24641
rect 16395 24592 16396 24632
rect 16436 24592 16437 24632
rect 16395 24583 16437 24592
rect 16876 24632 16916 24641
rect 16396 24498 16436 24583
rect 16876 24044 16916 24592
rect 17068 24632 17108 24641
rect 17068 24473 17108 24592
rect 17067 24464 17109 24473
rect 17067 24424 17068 24464
rect 17108 24424 17109 24464
rect 17067 24415 17109 24424
rect 18232 24212 18600 24221
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18232 24163 18600 24172
rect 16876 23995 16916 24004
rect 19084 23801 19124 26095
rect 19472 24968 19840 24977
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19472 24919 19840 24928
rect 19948 23960 19988 26104
rect 20716 23960 20756 28960
rect 22156 28337 22196 29128
rect 23115 29168 23157 29177
rect 23115 29128 23116 29168
rect 23156 29128 23157 29168
rect 23115 29119 23157 29128
rect 26092 29168 26132 29632
rect 26092 29119 26132 29128
rect 22636 29093 22676 29095
rect 22635 29084 22677 29093
rect 22635 29044 22636 29084
rect 22676 29044 22677 29084
rect 22635 29035 22677 29044
rect 22636 29000 22676 29035
rect 23116 29034 23156 29119
rect 22636 28951 22676 28960
rect 24267 29000 24309 29009
rect 24267 28960 24268 29000
rect 24308 28960 24309 29000
rect 24267 28951 24309 28960
rect 22155 28328 22197 28337
rect 22155 28288 22156 28328
rect 22196 28288 22197 28328
rect 22155 28279 22197 28288
rect 23979 28160 24021 28169
rect 23979 28120 23980 28160
rect 24020 28120 24021 28160
rect 23979 28111 24021 28120
rect 23980 26228 24020 28111
rect 23980 26179 24020 26188
rect 22732 26144 22772 26153
rect 21100 25892 21140 25901
rect 21100 25313 21140 25852
rect 21580 25892 21620 25901
rect 21620 25852 22100 25892
rect 21580 25843 21620 25852
rect 21099 25304 21141 25313
rect 21099 25264 21100 25304
rect 21140 25264 21141 25304
rect 21099 25255 21141 25264
rect 21771 25304 21813 25313
rect 21771 25264 21772 25304
rect 21812 25264 21813 25304
rect 21771 25255 21813 25264
rect 22060 25304 22100 25852
rect 22732 25481 22772 26104
rect 23595 26144 23637 26153
rect 23595 26104 23596 26144
rect 23636 26104 23637 26144
rect 23595 26095 23637 26104
rect 23596 26010 23636 26095
rect 22731 25472 22773 25481
rect 22731 25432 22732 25472
rect 22772 25432 22773 25472
rect 22731 25423 22773 25432
rect 22060 25255 22100 25264
rect 21772 25170 21812 25255
rect 22252 25136 22292 25145
rect 20907 24716 20949 24725
rect 20907 24676 20908 24716
rect 20948 24676 20949 24716
rect 20907 24667 20949 24676
rect 19180 23920 19988 23960
rect 20524 23920 20756 23960
rect 20908 24632 20948 24667
rect 16204 23792 16244 23801
rect 16204 23717 16244 23752
rect 17067 23792 17109 23801
rect 17067 23752 17068 23792
rect 17108 23752 17109 23792
rect 17067 23743 17109 23752
rect 17643 23792 17685 23801
rect 17643 23752 17644 23792
rect 17684 23752 17685 23792
rect 17643 23743 17685 23752
rect 18315 23792 18357 23801
rect 18315 23752 18316 23792
rect 18356 23752 18357 23792
rect 18315 23743 18357 23752
rect 19083 23792 19125 23801
rect 19083 23752 19084 23792
rect 19124 23752 19125 23792
rect 19083 23743 19125 23752
rect 19180 23792 19220 23920
rect 20331 23876 20373 23885
rect 20331 23836 20332 23876
rect 20372 23836 20373 23876
rect 20331 23827 20373 23836
rect 19180 23743 19220 23752
rect 16203 23708 16245 23717
rect 16203 23668 16204 23708
rect 16244 23668 16245 23708
rect 16203 23659 16245 23668
rect 16204 22541 16244 23659
rect 17068 23658 17108 23743
rect 16203 22532 16245 22541
rect 16203 22492 16204 22532
rect 16244 22492 16245 22532
rect 16203 22483 16245 22492
rect 17644 21617 17684 23743
rect 17740 23708 17780 23717
rect 17932 23708 17972 23717
rect 17780 23668 17932 23708
rect 17740 23659 17780 23668
rect 17932 23659 17972 23668
rect 18316 23658 18356 23743
rect 20332 23742 20372 23827
rect 19472 23456 19840 23465
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19472 23407 19840 23416
rect 18232 22700 18600 22709
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18232 22651 18600 22660
rect 20043 22028 20085 22037
rect 20043 21988 20044 22028
rect 20084 21988 20085 22028
rect 20043 21979 20085 21988
rect 19472 21944 19840 21953
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19472 21895 19840 21904
rect 17643 21608 17685 21617
rect 17643 21568 17644 21608
rect 17684 21568 17685 21608
rect 17643 21559 17685 21568
rect 19947 21356 19989 21365
rect 19947 21316 19948 21356
rect 19988 21316 19989 21356
rect 19947 21307 19989 21316
rect 18232 21188 18600 21197
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18232 21139 18600 21148
rect 16052 20980 16148 21020
rect 16012 20971 16052 20980
rect 13996 20719 14036 20728
rect 14860 20768 14900 20777
rect 14900 20728 14996 20768
rect 14860 20719 14900 20728
rect 13420 20684 13460 20693
rect 13612 20684 13652 20693
rect 13460 20644 13612 20684
rect 13420 20635 13460 20644
rect 13612 20635 13652 20644
rect 12460 19963 12500 19972
rect 12212 19468 12308 19508
rect 12172 19459 12212 19468
rect 11252 18712 11444 18752
rect 12844 19256 12884 19265
rect 11212 18703 11252 18712
rect 10732 18535 10772 18544
rect 11020 18584 11060 18593
rect 11020 17996 11060 18544
rect 11020 17947 11060 17956
rect 9867 17828 9909 17837
rect 9867 17788 9868 17828
rect 9908 17788 9909 17828
rect 9867 17779 9909 17788
rect 10827 17828 10869 17837
rect 10827 17788 10828 17828
rect 10868 17788 10869 17828
rect 10827 17779 10869 17788
rect 9868 17744 9908 17779
rect 9044 17704 9716 17744
rect 9004 17695 9044 17704
rect 3052 17106 3092 17191
rect 4012 16997 4052 17200
rect 3243 16988 3285 16997
rect 3243 16948 3244 16988
rect 3284 16948 3285 16988
rect 3243 16939 3285 16948
rect 4011 16988 4053 16997
rect 4011 16948 4012 16988
rect 4052 16948 4053 16988
rect 4011 16939 4053 16948
rect 3244 16854 3284 16939
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 4012 14804 4052 14813
rect 4012 14561 4052 14764
rect 3820 14552 3860 14561
rect 3820 14141 3860 14512
rect 4011 14552 4053 14561
rect 4011 14512 4012 14552
rect 4052 14512 4053 14552
rect 4011 14503 4053 14512
rect 2955 14132 2997 14141
rect 2955 14092 2956 14132
rect 2996 14092 2997 14132
rect 2955 14083 2997 14092
rect 3819 14132 3861 14141
rect 3819 14092 3820 14132
rect 3860 14092 3861 14132
rect 3819 14083 3861 14092
rect 651 14048 693 14057
rect 651 14008 652 14048
rect 692 14008 693 14048
rect 651 13999 693 14008
rect 2763 14048 2805 14057
rect 2763 14008 2764 14048
rect 2804 14008 2805 14048
rect 2763 13999 2805 14008
rect 2956 13998 2996 14083
rect 4204 14057 4244 17695
rect 8620 17660 8660 17669
rect 4588 17576 4628 17585
rect 4628 17536 4820 17576
rect 4588 17527 4628 17536
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 4684 17072 4724 17081
rect 4780 17072 4820 17536
rect 4724 17032 4820 17072
rect 4684 17023 4724 17032
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 5164 14720 5204 14729
rect 4492 14561 4532 14646
rect 4491 14552 4533 14561
rect 4491 14512 4492 14552
rect 4532 14512 4533 14552
rect 4491 14503 4533 14512
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 5164 14216 5204 14680
rect 6316 14720 6356 14729
rect 8044 14720 8084 14729
rect 6356 14680 6452 14720
rect 6316 14671 6356 14680
rect 5836 14552 5876 14561
rect 5356 14216 5396 14225
rect 5164 14176 5356 14216
rect 5356 14167 5396 14176
rect 5836 14057 5876 14512
rect 3339 14048 3381 14057
rect 3339 14008 3340 14048
rect 3380 14008 3381 14048
rect 3339 13999 3381 14008
rect 4203 14048 4245 14057
rect 4203 14008 4204 14048
rect 4244 14008 4245 14048
rect 4203 13999 4245 14008
rect 5835 14048 5877 14057
rect 5835 14008 5836 14048
rect 5876 14008 5877 14048
rect 5835 13999 5877 14008
rect 6220 14048 6260 14057
rect 6260 14008 6356 14048
rect 6220 13999 6260 14008
rect 3340 13914 3380 13999
rect 4204 13914 4244 13999
rect 4395 13964 4437 13973
rect 4395 13924 4396 13964
rect 4436 13924 4437 13964
rect 4395 13915 4437 13924
rect 5739 13964 5781 13973
rect 5739 13924 5740 13964
rect 5780 13924 5781 13964
rect 5739 13915 5781 13924
rect 4011 13880 4053 13889
rect 4011 13840 4012 13880
rect 4052 13840 4053 13880
rect 4011 13831 4053 13840
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 651 13208 693 13217
rect 651 13168 652 13208
rect 692 13168 693 13208
rect 651 13159 693 13168
rect 4012 13208 4052 13831
rect 4012 13159 4052 13168
rect 4396 13208 4436 13915
rect 5547 13880 5589 13889
rect 5547 13840 5548 13880
rect 5588 13840 5589 13880
rect 5547 13831 5589 13840
rect 5548 13746 5588 13831
rect 5740 13830 5780 13915
rect 5836 13217 5876 13999
rect 6316 13460 6356 14008
rect 6412 13889 6452 14680
rect 7275 14552 7317 14561
rect 7275 14512 7276 14552
rect 7316 14512 7317 14552
rect 7275 14503 7317 14512
rect 7179 14132 7221 14141
rect 7179 14092 7180 14132
rect 7220 14092 7221 14132
rect 7179 14083 7221 14092
rect 7084 14048 7124 14059
rect 7084 13973 7124 14008
rect 7180 13998 7220 14083
rect 7276 14048 7316 14503
rect 8044 14141 8084 14680
rect 8428 14720 8468 14729
rect 8428 14141 8468 14680
rect 8524 14636 8564 14645
rect 8620 14636 8660 17620
rect 9580 17072 9620 17081
rect 9676 17072 9716 17704
rect 9868 17693 9908 17704
rect 9964 17072 10004 17081
rect 10828 17072 10868 17779
rect 12844 17669 12884 19216
rect 14859 17912 14901 17921
rect 14859 17872 14860 17912
rect 14900 17872 14901 17912
rect 14859 17863 14901 17872
rect 11979 17660 12021 17669
rect 11979 17620 11980 17660
rect 12020 17620 12021 17660
rect 11979 17611 12021 17620
rect 12843 17660 12885 17669
rect 12843 17620 12844 17660
rect 12884 17620 12885 17660
rect 12843 17611 12885 17620
rect 11980 17240 12020 17611
rect 11980 17191 12020 17200
rect 14860 17156 14900 17863
rect 14860 17107 14900 17116
rect 9676 17032 9964 17072
rect 9580 15140 9620 17032
rect 9100 15100 9620 15140
rect 9100 14972 9140 15100
rect 9100 14923 9140 14932
rect 8907 14720 8949 14729
rect 8907 14680 8908 14720
rect 8948 14680 8949 14720
rect 8907 14671 8949 14680
rect 9099 14720 9141 14729
rect 9099 14680 9100 14720
rect 9140 14680 9141 14720
rect 9099 14671 9141 14680
rect 8564 14596 8660 14636
rect 8524 14587 8564 14596
rect 8908 14586 8948 14671
rect 8811 14552 8853 14561
rect 8811 14512 8812 14552
rect 8852 14512 8853 14552
rect 8811 14503 8853 14512
rect 8812 14418 8852 14503
rect 8043 14132 8085 14141
rect 8043 14092 8044 14132
rect 8084 14092 8085 14132
rect 8043 14083 8085 14092
rect 8427 14132 8469 14141
rect 8427 14092 8428 14132
rect 8468 14092 8469 14132
rect 8427 14083 8469 14092
rect 7276 13999 7316 14008
rect 9100 14048 9140 14671
rect 9195 14132 9237 14141
rect 9195 14092 9196 14132
rect 9236 14092 9237 14132
rect 9195 14083 9237 14092
rect 6891 13964 6933 13973
rect 6891 13924 6892 13964
rect 6932 13924 6933 13964
rect 6891 13915 6933 13924
rect 7083 13964 7125 13973
rect 7083 13924 7084 13964
rect 7124 13924 7125 13964
rect 7083 13915 7125 13924
rect 6411 13880 6453 13889
rect 6411 13840 6412 13880
rect 6452 13840 6453 13880
rect 6411 13831 6453 13840
rect 6892 13830 6932 13915
rect 9003 13880 9045 13889
rect 9003 13840 9004 13880
rect 9044 13840 9045 13880
rect 9003 13831 9045 13840
rect 6412 13460 6452 13469
rect 6316 13420 6412 13460
rect 6412 13411 6452 13420
rect 4396 13159 4436 13168
rect 5259 13208 5301 13217
rect 5259 13168 5260 13208
rect 5300 13168 5301 13208
rect 5259 13159 5301 13168
rect 5835 13208 5877 13217
rect 5835 13168 5836 13208
rect 5876 13168 5877 13208
rect 5835 13159 5877 13168
rect 8043 13208 8085 13217
rect 8043 13168 8044 13208
rect 8084 13168 8085 13208
rect 8043 13159 8085 13168
rect 652 13040 692 13159
rect 5260 13074 5300 13159
rect 652 12991 692 13000
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 652 12704 692 12713
rect 652 12377 692 12664
rect 651 12368 693 12377
rect 651 12328 652 12368
rect 692 12328 693 12368
rect 651 12319 693 12328
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 651 11528 693 11537
rect 651 11488 652 11528
rect 692 11488 693 11528
rect 651 11479 693 11488
rect 652 11394 692 11479
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 652 11192 692 11201
rect 652 10697 692 11152
rect 651 10688 693 10697
rect 651 10648 652 10688
rect 692 10648 693 10688
rect 651 10639 693 10648
rect 843 10688 885 10697
rect 843 10648 844 10688
rect 884 10648 885 10688
rect 843 10639 885 10648
rect 652 10016 692 10025
rect 652 9857 692 9976
rect 651 9848 693 9857
rect 651 9808 652 9848
rect 692 9808 693 9848
rect 651 9799 693 9808
rect 652 9680 692 9689
rect 652 9017 692 9640
rect 651 9008 693 9017
rect 651 8968 652 9008
rect 692 8968 693 9008
rect 651 8959 693 8968
rect 652 8504 692 8513
rect 556 8464 652 8504
rect 556 8177 596 8464
rect 652 8455 692 8464
rect 555 8168 597 8177
rect 555 8128 556 8168
rect 596 8128 597 8168
rect 555 8119 597 8128
rect 652 8168 692 8177
rect 652 7337 692 8128
rect 651 7328 693 7337
rect 651 7288 652 7328
rect 692 7288 693 7328
rect 651 7279 693 7288
rect 652 6992 692 7001
rect 652 6497 692 6952
rect 651 6488 693 6497
rect 651 6448 652 6488
rect 692 6448 693 6488
rect 651 6439 693 6448
rect 651 5648 693 5657
rect 651 5608 652 5648
rect 692 5608 693 5648
rect 651 5599 693 5608
rect 652 5480 692 5599
rect 652 5431 692 5440
rect 844 4892 884 10639
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 2283 10352 2325 10361
rect 2283 10312 2284 10352
rect 2324 10312 2325 10352
rect 2283 10303 2325 10312
rect 3147 10352 3189 10361
rect 3147 10312 3148 10352
rect 3188 10312 3189 10352
rect 3147 10303 3189 10312
rect 2284 9596 2324 10303
rect 3148 10218 3188 10303
rect 3339 10268 3381 10277
rect 3339 10228 3340 10268
rect 3380 10228 3381 10268
rect 3339 10219 3381 10228
rect 4107 10268 4149 10277
rect 4107 10228 4108 10268
rect 4148 10228 4149 10268
rect 4107 10219 4149 10228
rect 3340 10134 3380 10219
rect 2284 9547 2324 9556
rect 4108 10100 4148 10219
rect 2668 9512 2708 9521
rect 2668 8756 2708 9472
rect 3532 9512 3572 9521
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 2668 8716 3380 8756
rect 2092 5648 2132 5657
rect 1324 5608 2092 5648
rect 1324 5144 1364 5608
rect 2092 5599 2132 5608
rect 2763 5648 2805 5657
rect 2763 5608 2764 5648
rect 2804 5608 2805 5648
rect 2763 5599 2805 5608
rect 2764 5514 2804 5599
rect 1324 5095 1364 5104
rect 2475 4976 2517 4985
rect 2475 4936 2476 4976
rect 2516 4936 2517 4976
rect 2475 4927 2517 4936
rect 844 4843 884 4852
rect 2476 4842 2516 4927
rect 2860 4901 2900 8716
rect 3340 8672 3380 8716
rect 3532 8681 3572 9472
rect 3340 8623 3380 8632
rect 3531 8672 3573 8681
rect 3531 8632 3532 8672
rect 3572 8632 3573 8672
rect 3531 8623 3573 8632
rect 2956 8588 2996 8597
rect 2996 8548 3284 8588
rect 2956 8539 2996 8548
rect 3244 8252 3284 8548
rect 3244 8212 3764 8252
rect 3724 8168 3764 8212
rect 3724 8119 3764 8128
rect 4108 8000 4148 10060
rect 4780 10184 4820 10193
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 4684 9680 4724 9689
rect 4780 9680 4820 10144
rect 4724 9640 4820 9680
rect 4684 9631 4724 9640
rect 6123 9512 6165 9521
rect 6123 9472 6124 9512
rect 6164 9472 6165 9512
rect 6123 9463 6165 9472
rect 6795 9512 6837 9521
rect 6795 9472 6796 9512
rect 6836 9472 6837 9512
rect 6795 9463 6837 9472
rect 7180 9512 7220 9521
rect 4203 8672 4245 8681
rect 4203 8632 4204 8672
rect 4244 8632 4245 8672
rect 4203 8623 4245 8632
rect 4204 8538 4244 8623
rect 5356 8504 5396 8513
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 4396 8000 4436 8009
rect 4108 7960 4396 8000
rect 4396 7951 4436 7960
rect 4491 8000 4533 8009
rect 4491 7960 4492 8000
rect 4532 7960 4533 8000
rect 4491 7951 4533 7960
rect 4588 8000 4628 8009
rect 5356 8000 5396 8464
rect 6124 8168 6164 9463
rect 6796 9378 6836 9463
rect 6603 8672 6645 8681
rect 6603 8632 6604 8672
rect 6644 8632 6645 8672
rect 6603 8623 6645 8632
rect 6124 8119 6164 8128
rect 5452 8000 5492 8009
rect 5356 7960 5452 8000
rect 3916 7916 3956 7925
rect 3916 7748 3956 7876
rect 4492 7866 4532 7951
rect 4588 7748 4628 7960
rect 5452 7951 5492 7960
rect 5644 8000 5684 8009
rect 4780 7748 4820 7757
rect 3916 7708 4780 7748
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 4587 6656 4629 6665
rect 4587 6616 4588 6656
rect 4628 6616 4629 6656
rect 4587 6607 4629 6616
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 4588 5900 4628 6607
rect 4588 5851 4628 5860
rect 2956 5732 2996 5743
rect 2956 5657 2996 5692
rect 4780 5657 4820 7708
rect 5644 6665 5684 7960
rect 5931 8000 5973 8009
rect 5931 7960 5932 8000
rect 5972 7960 5973 8000
rect 5931 7951 5973 7960
rect 6604 8000 6644 8623
rect 6604 7951 6644 7960
rect 5932 7866 5972 7951
rect 6892 7748 6932 7757
rect 5643 6656 5685 6665
rect 5643 6616 5644 6656
rect 5684 6616 5685 6656
rect 5643 6607 5685 6616
rect 2955 5648 2997 5657
rect 2955 5608 2956 5648
rect 2996 5608 2997 5648
rect 2955 5599 2997 5608
rect 4491 5648 4533 5657
rect 4491 5608 4492 5648
rect 4532 5608 4533 5648
rect 4491 5599 4533 5608
rect 4684 5648 4724 5657
rect 4492 5514 4532 5599
rect 3148 5480 3188 5489
rect 4684 5480 4724 5608
rect 4779 5648 4821 5657
rect 4779 5608 4780 5648
rect 4820 5608 4821 5648
rect 4779 5599 4821 5608
rect 5163 5648 5205 5657
rect 5163 5608 5164 5648
rect 5204 5608 5205 5648
rect 5163 5599 5205 5608
rect 6220 5648 6260 5657
rect 6260 5608 6356 5648
rect 5164 5514 5204 5599
rect 6220 5580 6260 5608
rect 5067 5480 5109 5489
rect 3188 5440 3764 5480
rect 4684 5440 5068 5480
rect 5108 5440 5109 5480
rect 3148 5431 3188 5440
rect 3724 5060 3764 5440
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 3724 5011 3764 5020
rect 3340 4976 3380 4987
rect 3340 4901 3380 4936
rect 3916 4976 3956 4985
rect 4300 4976 4340 4987
rect 3956 4936 4244 4976
rect 3916 4927 3956 4936
rect 2859 4892 2901 4901
rect 2859 4852 2860 4892
rect 2900 4852 2901 4892
rect 2859 4843 2901 4852
rect 3339 4892 3381 4901
rect 3339 4852 3340 4892
rect 3380 4852 3381 4892
rect 3339 4843 3381 4852
rect 651 4808 693 4817
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 652 4674 692 4759
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 4204 4388 4244 4936
rect 4300 4901 4340 4936
rect 4299 4892 4341 4901
rect 4299 4852 4300 4892
rect 4340 4852 4341 4892
rect 4299 4843 4341 4852
rect 4396 4388 4436 4397
rect 4204 4348 4396 4388
rect 4396 4339 4436 4348
rect 843 4220 885 4229
rect 843 4180 844 4220
rect 884 4180 885 4220
rect 843 4171 885 4180
rect 4588 4220 4628 4229
rect 4780 4220 4820 5440
rect 5067 5431 5109 5440
rect 5356 5480 5396 5489
rect 5068 5346 5108 5431
rect 5356 5069 5396 5440
rect 5547 5480 5589 5489
rect 5547 5440 5548 5480
rect 5588 5440 5589 5480
rect 5547 5431 5589 5440
rect 5548 5346 5588 5431
rect 5355 5060 5397 5069
rect 5355 5020 5356 5060
rect 5396 5020 5397 5060
rect 5355 5011 5397 5020
rect 5163 4976 5205 4985
rect 5163 4936 5164 4976
rect 5204 4936 5205 4976
rect 5163 4927 5205 4936
rect 5164 4842 5204 4927
rect 6316 4892 6356 5608
rect 6892 4985 6932 7708
rect 7180 6413 7220 9472
rect 8044 9512 8084 13159
rect 9004 12368 9044 13831
rect 9100 13292 9140 14008
rect 9196 13998 9236 14083
rect 9291 14048 9333 14057
rect 9484 14048 9524 14057
rect 9291 14008 9292 14048
rect 9332 14008 9333 14048
rect 9291 13999 9333 14008
rect 9388 14008 9484 14048
rect 9292 13914 9332 13999
rect 9292 13460 9332 13469
rect 9388 13460 9428 14008
rect 9484 13999 9524 14008
rect 9579 14048 9621 14057
rect 9579 14008 9580 14048
rect 9620 14008 9621 14048
rect 9579 13999 9621 14008
rect 9868 14048 9908 17032
rect 9964 17023 10004 17032
rect 10732 17032 10828 17072
rect 10732 16484 10772 17032
rect 10828 17023 10868 17032
rect 10732 16435 10772 16444
rect 14956 16409 14996 20728
rect 19472 20432 19840 20441
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19472 20383 19840 20392
rect 18232 19676 18600 19685
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18232 19627 18600 19636
rect 19948 19256 19988 21307
rect 20044 21020 20084 21979
rect 20331 21356 20373 21365
rect 20331 21316 20332 21356
rect 20372 21316 20373 21356
rect 20331 21307 20373 21316
rect 20332 21222 20372 21307
rect 20044 20971 20084 20980
rect 20524 20768 20564 23920
rect 20811 23876 20853 23885
rect 20811 23836 20812 23876
rect 20852 23836 20853 23876
rect 20811 23827 20853 23836
rect 20812 23792 20852 23827
rect 20812 23741 20852 23752
rect 20716 23204 20756 23213
rect 20756 23164 20852 23204
rect 20716 23155 20756 23164
rect 20812 21608 20852 23164
rect 20908 23120 20948 24592
rect 21099 24632 21141 24641
rect 21099 24592 21100 24632
rect 21140 24592 21141 24632
rect 21099 24583 21141 24592
rect 21483 24632 21525 24641
rect 21483 24592 21484 24632
rect 21524 24592 21525 24632
rect 21483 24583 21525 24592
rect 21100 24498 21140 24583
rect 21003 24380 21045 24389
rect 21003 24340 21004 24380
rect 21044 24340 21045 24380
rect 21003 24331 21045 24340
rect 21004 24246 21044 24331
rect 21484 23960 21524 24583
rect 21963 24380 22005 24389
rect 21963 24340 21964 24380
rect 22004 24340 22005 24380
rect 21963 24331 22005 24340
rect 21484 23911 21524 23920
rect 21003 23876 21045 23885
rect 21003 23836 21004 23876
rect 21044 23836 21236 23876
rect 21003 23827 21045 23836
rect 20908 23071 20948 23080
rect 21196 23120 21236 23836
rect 21964 23792 22004 24331
rect 22252 23960 22292 25096
rect 21964 23743 22004 23752
rect 22060 23920 22292 23960
rect 22060 23792 22100 23920
rect 22060 23743 22100 23752
rect 21676 23624 21716 23633
rect 21716 23584 22004 23624
rect 21676 23575 21716 23584
rect 21196 23071 21236 23080
rect 21964 22280 22004 23584
rect 21964 22231 22004 22240
rect 21292 22112 21332 22121
rect 21100 22072 21292 22112
rect 21004 21608 21044 21617
rect 20812 21568 21004 21608
rect 21004 21559 21044 21568
rect 21004 20768 21044 20777
rect 20564 20728 21004 20768
rect 20524 20719 20564 20728
rect 20620 20096 20660 20728
rect 21004 20719 21044 20728
rect 20620 20047 20660 20056
rect 21004 20096 21044 20105
rect 21100 20096 21140 22072
rect 21292 22063 21332 22072
rect 21964 20768 22004 20777
rect 21964 20609 22004 20728
rect 21963 20600 22005 20609
rect 21963 20560 21964 20600
rect 22004 20560 22005 20600
rect 21963 20551 22005 20560
rect 21044 20056 21140 20096
rect 21388 20096 21428 20107
rect 22732 20105 22772 25423
rect 24268 25304 24308 28951
rect 26764 28916 26804 28925
rect 26475 28160 26517 28169
rect 26475 28120 26476 28160
rect 26516 28120 26517 28160
rect 26475 28111 26517 28120
rect 26476 28026 26516 28111
rect 26764 27749 26804 28876
rect 27147 28412 27189 28421
rect 27147 28372 27148 28412
rect 27188 28372 27189 28412
rect 27147 28363 27189 28372
rect 28779 28412 28821 28421
rect 28779 28372 28780 28412
rect 28820 28372 28821 28412
rect 28779 28363 28821 28372
rect 27148 28328 27188 28363
rect 27148 28277 27188 28288
rect 28780 28278 28820 28363
rect 28875 28328 28917 28337
rect 28875 28288 28876 28328
rect 28916 28288 28917 28328
rect 28875 28279 28917 28288
rect 26187 27740 26229 27749
rect 26187 27700 26188 27740
rect 26228 27700 26229 27740
rect 26187 27691 26229 27700
rect 26763 27740 26805 27749
rect 26763 27700 26764 27740
rect 26804 27700 26805 27740
rect 26763 27691 26805 27700
rect 26188 27606 26228 27691
rect 26572 27656 26612 27665
rect 26572 26573 26612 27616
rect 27436 27656 27476 27665
rect 26571 26564 26613 26573
rect 26571 26524 26572 26564
rect 26612 26524 26613 26564
rect 26571 26515 26613 26524
rect 26091 26144 26133 26153
rect 26091 26104 26092 26144
rect 26132 26104 26133 26144
rect 26091 26095 26133 26104
rect 24555 25472 24597 25481
rect 24555 25432 24556 25472
rect 24596 25432 24597 25472
rect 24555 25423 24597 25432
rect 24556 25338 24596 25423
rect 24268 25255 24308 25264
rect 25132 25220 25172 25229
rect 25172 25180 25268 25220
rect 25132 25171 25172 25180
rect 22923 24716 22965 24725
rect 22923 24676 22924 24716
rect 22964 24676 22965 24716
rect 22923 24667 22965 24676
rect 22924 24582 22964 24667
rect 25228 24641 25268 25180
rect 26092 24725 26132 26095
rect 27147 25892 27189 25901
rect 27147 25852 27148 25892
rect 27188 25852 27189 25892
rect 27147 25843 27189 25852
rect 26091 24716 26133 24725
rect 26091 24676 26092 24716
rect 26132 24676 26133 24716
rect 26091 24667 26133 24676
rect 26763 24716 26805 24725
rect 26763 24676 26764 24716
rect 26804 24676 26805 24716
rect 26763 24667 26805 24676
rect 27148 24716 27188 25843
rect 27148 24667 27188 24676
rect 23595 24632 23637 24641
rect 23595 24592 23596 24632
rect 23636 24592 23637 24632
rect 23595 24583 23637 24592
rect 25227 24632 25269 24641
rect 25227 24592 25228 24632
rect 25268 24592 25269 24632
rect 25227 24583 25269 24592
rect 25899 24632 25941 24641
rect 25899 24592 25900 24632
rect 25940 24592 25941 24632
rect 25899 24583 25941 24592
rect 23596 24498 23636 24583
rect 24747 24548 24789 24557
rect 24747 24508 24748 24548
rect 24788 24508 24789 24548
rect 24747 24499 24789 24508
rect 24748 24414 24788 24499
rect 25900 24498 25940 24583
rect 26092 22280 26132 24667
rect 26764 24632 26804 24667
rect 27436 24641 27476 27616
rect 28780 27656 28820 27665
rect 28588 27572 28628 27581
rect 28780 27572 28820 27616
rect 28628 27532 28820 27572
rect 28588 27523 28628 27532
rect 28780 27068 28820 27077
rect 28876 27068 28916 28279
rect 28820 27028 28916 27068
rect 28780 27019 28820 27028
rect 28684 26816 28724 26827
rect 28684 26741 28724 26776
rect 28875 26816 28917 26825
rect 28875 26776 28876 26816
rect 28916 26776 28917 26816
rect 28875 26767 28917 26776
rect 28683 26732 28725 26741
rect 28683 26692 28684 26732
rect 28724 26692 28820 26732
rect 28683 26683 28725 26692
rect 28684 26228 28724 26237
rect 28396 26188 28684 26228
rect 28396 26144 28436 26188
rect 28684 26179 28724 26188
rect 28396 26095 28436 26104
rect 28780 26144 28820 26692
rect 28876 26682 28916 26767
rect 28875 26564 28917 26573
rect 28875 26524 28876 26564
rect 28916 26524 28917 26564
rect 28875 26515 28917 26524
rect 28780 26095 28820 26104
rect 27723 25892 27765 25901
rect 27723 25852 27724 25892
rect 27764 25852 27765 25892
rect 27723 25843 27765 25852
rect 27724 25758 27764 25843
rect 28780 25304 28820 25313
rect 28876 25304 28916 26515
rect 28972 25556 29012 29791
rect 30508 29672 30548 29681
rect 30508 29168 30548 29632
rect 30604 29168 30644 29177
rect 30508 29128 30604 29168
rect 30604 29119 30644 29128
rect 31563 29168 31605 29177
rect 31563 29128 31564 29168
rect 31604 29128 31605 29168
rect 31563 29119 31605 29128
rect 29932 28916 29972 28925
rect 29164 28876 29932 28916
rect 29067 28328 29109 28337
rect 29067 28288 29068 28328
rect 29108 28288 29109 28328
rect 29067 28279 29109 28288
rect 29164 28328 29204 28876
rect 29932 28867 29972 28876
rect 29164 28279 29204 28288
rect 29068 28194 29108 28279
rect 29452 27404 29492 27413
rect 29164 27364 29452 27404
rect 29164 26825 29204 27364
rect 29452 27355 29492 27364
rect 29163 26816 29205 26825
rect 29163 26776 29164 26816
rect 29204 26776 29205 26816
rect 29163 26767 29205 26776
rect 29164 26144 29204 26767
rect 30603 26648 30645 26657
rect 30603 26608 30604 26648
rect 30644 26608 30645 26648
rect 30603 26599 30645 26608
rect 29164 26095 29204 26104
rect 28972 25507 29012 25516
rect 30604 25313 30644 26599
rect 28820 25264 28916 25304
rect 29643 25304 29685 25313
rect 29643 25264 29644 25304
rect 29684 25264 29685 25304
rect 26764 24581 26804 24592
rect 26955 24632 26997 24641
rect 26955 24592 26956 24632
rect 26996 24592 26997 24632
rect 26955 24583 26997 24592
rect 27435 24632 27477 24641
rect 27435 24592 27436 24632
rect 27476 24592 27477 24632
rect 27435 24583 27477 24592
rect 25707 22196 25749 22205
rect 25707 22156 25708 22196
rect 25748 22156 25749 22196
rect 25707 22147 25749 22156
rect 25708 22062 25748 22147
rect 25803 21608 25845 21617
rect 25803 21568 25804 21608
rect 25844 21568 25845 21608
rect 26092 21608 26132 22240
rect 26956 22280 26996 24583
rect 28204 23120 28244 23129
rect 27532 22868 27572 22877
rect 26956 22231 26996 22240
rect 27052 22828 27532 22868
rect 26475 22196 26517 22205
rect 26475 22156 26476 22196
rect 26516 22156 26517 22196
rect 26475 22147 26517 22156
rect 26188 21608 26228 21617
rect 26092 21568 26188 21608
rect 25803 21559 25845 21568
rect 26188 21559 26228 21568
rect 25804 21474 25844 21559
rect 26476 21020 26516 22147
rect 27052 21776 27092 22828
rect 27532 22819 27572 22828
rect 28108 22532 28148 22541
rect 28204 22532 28244 23080
rect 28148 22492 28244 22532
rect 28108 22483 28148 22492
rect 26476 20971 26516 20980
rect 26668 21736 27092 21776
rect 26668 20852 26708 21736
rect 26859 21608 26901 21617
rect 27051 21608 27093 21617
rect 26859 21568 26860 21608
rect 26900 21568 26901 21608
rect 26859 21559 26901 21568
rect 26956 21568 27052 21608
rect 27092 21568 27093 21608
rect 26860 21020 26900 21559
rect 26860 20971 26900 20980
rect 21004 20047 21044 20056
rect 21388 20021 21428 20056
rect 22251 20096 22293 20105
rect 22251 20056 22252 20096
rect 22292 20056 22293 20096
rect 22251 20047 22293 20056
rect 22731 20096 22773 20105
rect 22731 20056 22732 20096
rect 22772 20056 22773 20096
rect 22731 20047 22773 20056
rect 20331 20012 20373 20021
rect 20331 19972 20332 20012
rect 20372 19972 20373 20012
rect 20331 19963 20373 19972
rect 21387 20012 21429 20021
rect 21387 19972 21388 20012
rect 21428 19972 21429 20012
rect 21387 19963 21429 19972
rect 19948 19207 19988 19216
rect 20332 19256 20372 19963
rect 22252 19962 22292 20047
rect 26668 20021 26708 20812
rect 25227 20012 25269 20021
rect 25227 19972 25228 20012
rect 25268 19972 25269 20012
rect 25227 19963 25269 19972
rect 26667 20012 26709 20021
rect 26667 19972 26668 20012
rect 26708 19972 26709 20012
rect 26667 19963 26709 19972
rect 20427 19844 20469 19853
rect 20427 19804 20428 19844
rect 20468 19804 20469 19844
rect 20427 19795 20469 19804
rect 20811 19844 20853 19853
rect 20811 19804 20812 19844
rect 20852 19804 20853 19844
rect 20811 19795 20853 19804
rect 23404 19844 23444 19853
rect 20428 19710 20468 19795
rect 20332 19207 20372 19216
rect 19472 18920 19840 18929
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19472 18871 19840 18880
rect 18232 18164 18600 18173
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18232 18115 18600 18124
rect 15819 17912 15861 17921
rect 15819 17872 15820 17912
rect 15860 17872 15861 17912
rect 15819 17863 15861 17872
rect 15820 17778 15860 17863
rect 16012 17828 16052 17837
rect 16012 17669 16052 17788
rect 17452 17744 17492 17753
rect 17260 17704 17452 17744
rect 16011 17660 16053 17669
rect 16011 17620 16012 17660
rect 16052 17620 16053 17660
rect 16011 17611 16053 17620
rect 16779 17660 16821 17669
rect 16779 17620 16780 17660
rect 16820 17620 16821 17660
rect 16779 17611 16821 17620
rect 16780 17526 16820 17611
rect 17260 17240 17300 17704
rect 17452 17695 17492 17704
rect 17547 17660 17589 17669
rect 17547 17620 17548 17660
rect 17588 17620 17589 17660
rect 17547 17611 17589 17620
rect 17260 17191 17300 17200
rect 15244 17072 15284 17081
rect 14955 16400 14997 16409
rect 14955 16360 14956 16400
rect 14996 16360 14997 16400
rect 14955 16351 14997 16360
rect 15244 16241 15284 17032
rect 16108 17072 16148 17081
rect 15819 16400 15861 16409
rect 15819 16360 15820 16400
rect 15860 16360 15861 16400
rect 15819 16351 15861 16360
rect 10252 16232 10292 16241
rect 9908 14008 10196 14048
rect 9868 13999 9908 14008
rect 9332 13420 9428 13460
rect 9292 13411 9332 13420
rect 9100 13243 9140 13252
rect 9484 13292 9524 13301
rect 9580 13292 9620 13999
rect 9524 13252 9620 13292
rect 9484 13243 9524 13252
rect 10156 13208 10196 14008
rect 10252 13889 10292 16192
rect 14955 16232 14997 16241
rect 14955 16192 14956 16232
rect 14996 16192 14997 16232
rect 14955 16183 14997 16192
rect 15243 16232 15285 16241
rect 15243 16192 15244 16232
rect 15284 16192 15285 16232
rect 15243 16183 15285 16192
rect 15820 16232 15860 16351
rect 16108 16232 16148 17032
rect 16972 16316 17012 16325
rect 17012 16276 17204 16316
rect 16972 16267 17012 16276
rect 15860 16192 16148 16232
rect 17164 16232 17204 16276
rect 15820 16183 15860 16192
rect 14572 16148 14612 16157
rect 10732 16064 10772 16073
rect 10635 14720 10677 14729
rect 10635 14680 10636 14720
rect 10676 14680 10677 14720
rect 10635 14671 10677 14680
rect 10636 14586 10676 14671
rect 10732 14048 10772 16024
rect 14572 15737 14612 16108
rect 14956 16098 14996 16183
rect 14571 15728 14613 15737
rect 14571 15688 14572 15728
rect 14612 15688 14613 15728
rect 14571 15679 14613 15688
rect 15627 15728 15669 15737
rect 15627 15688 15628 15728
rect 15668 15688 15669 15728
rect 15627 15679 15669 15688
rect 15628 15594 15668 15679
rect 15916 15560 15956 16192
rect 17164 16183 17204 16192
rect 16012 15560 16052 15569
rect 15916 15520 16012 15560
rect 16012 15511 16052 15520
rect 16971 15560 17013 15569
rect 16971 15520 16972 15560
rect 17012 15520 17013 15560
rect 16971 15511 17013 15520
rect 17452 15560 17492 15569
rect 17548 15560 17588 17611
rect 19472 17408 19840 17417
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19472 17359 19840 17368
rect 20140 17072 20180 17081
rect 20428 17072 20468 17081
rect 19468 16820 19508 16829
rect 18232 16652 18600 16661
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18232 16603 18600 16612
rect 19468 16325 19508 16780
rect 20140 16409 20180 17032
rect 20332 17032 20428 17072
rect 20139 16400 20181 16409
rect 20139 16360 20140 16400
rect 20180 16360 20181 16400
rect 20139 16351 20181 16360
rect 18027 16316 18069 16325
rect 18027 16276 18028 16316
rect 18068 16276 18069 16316
rect 18027 16267 18069 16276
rect 18507 16316 18549 16325
rect 18507 16276 18508 16316
rect 18548 16276 18549 16316
rect 18507 16267 18549 16276
rect 19467 16316 19509 16325
rect 19467 16276 19468 16316
rect 19508 16276 19509 16316
rect 19467 16267 19509 16276
rect 20043 16316 20085 16325
rect 20043 16276 20044 16316
rect 20084 16276 20085 16316
rect 20043 16267 20085 16276
rect 17836 16064 17876 16073
rect 17492 15520 17588 15560
rect 17644 15560 17684 15569
rect 17452 15511 17492 15520
rect 15819 15476 15861 15485
rect 15819 15436 15820 15476
rect 15860 15436 15861 15476
rect 15819 15427 15861 15436
rect 15820 15342 15860 15427
rect 16972 15426 17012 15511
rect 17547 15392 17589 15401
rect 17547 15352 17548 15392
rect 17588 15352 17589 15392
rect 17547 15343 17589 15352
rect 16492 15308 16532 15317
rect 11308 14720 11348 14729
rect 11308 14225 11348 14680
rect 11307 14216 11349 14225
rect 11307 14176 11308 14216
rect 11348 14176 11349 14216
rect 11307 14167 11349 14176
rect 11883 14216 11925 14225
rect 11883 14176 11884 14216
rect 11924 14176 11925 14216
rect 11883 14167 11925 14176
rect 11884 14082 11924 14167
rect 12075 14048 12117 14057
rect 10772 14008 11156 14048
rect 10732 13999 10772 14008
rect 10251 13880 10293 13889
rect 10251 13840 10252 13880
rect 10292 13840 10293 13880
rect 10251 13831 10293 13840
rect 10252 13208 10292 13217
rect 10156 13168 10252 13208
rect 10252 13159 10292 13168
rect 11116 13208 11156 14008
rect 12075 14008 12076 14048
rect 12116 14008 12117 14048
rect 12075 13999 12117 14008
rect 12267 14048 12309 14057
rect 12267 14008 12268 14048
rect 12308 14008 12309 14048
rect 12267 13999 12309 14008
rect 12747 14048 12789 14057
rect 12747 14008 12748 14048
rect 12788 14008 12789 14048
rect 12747 13999 12789 14008
rect 12076 13914 12116 13999
rect 12268 13460 12308 13999
rect 12748 13914 12788 13999
rect 12268 13411 12308 13420
rect 11116 13159 11156 13168
rect 9868 13124 9908 13133
rect 9676 13040 9716 13049
rect 9868 13040 9908 13084
rect 9716 13000 9908 13040
rect 9676 12991 9716 13000
rect 9483 12536 9525 12545
rect 9483 12496 9484 12536
rect 9524 12496 9525 12536
rect 9483 12487 9525 12496
rect 10251 12536 10293 12545
rect 10251 12496 10252 12536
rect 10292 12496 10293 12536
rect 10251 12487 10293 12496
rect 9484 12402 9524 12487
rect 9004 12319 9044 12328
rect 10252 11024 10292 12487
rect 16492 11033 16532 15268
rect 17548 15258 17588 15343
rect 17644 15317 17684 15520
rect 17836 15560 17876 16024
rect 17836 15485 17876 15520
rect 18028 15560 18068 16267
rect 18508 16182 18548 16267
rect 19275 16232 19317 16241
rect 19275 16192 19276 16232
rect 19316 16192 19317 16232
rect 19275 16183 19317 16192
rect 18892 16148 18932 16157
rect 18700 16108 18892 16148
rect 18700 16064 18740 16108
rect 18892 16099 18932 16108
rect 19276 16098 19316 16183
rect 18700 16015 18740 16024
rect 18795 15980 18837 15989
rect 18795 15940 18796 15980
rect 18836 15940 18837 15980
rect 18795 15931 18837 15940
rect 18699 15644 18741 15653
rect 18699 15604 18700 15644
rect 18740 15604 18741 15644
rect 18699 15595 18741 15604
rect 18028 15511 18068 15520
rect 18220 15560 18260 15569
rect 17835 15476 17877 15485
rect 17835 15436 17836 15476
rect 17876 15436 17877 15476
rect 17835 15427 17877 15436
rect 17932 15392 17972 15401
rect 18220 15392 18260 15520
rect 18508 15560 18548 15569
rect 18508 15401 18548 15520
rect 18700 15510 18740 15595
rect 18796 15569 18836 15931
rect 19472 15896 19840 15905
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19472 15847 19840 15856
rect 19948 15728 19988 15737
rect 18795 15560 18837 15569
rect 18795 15520 18796 15560
rect 18836 15520 18837 15560
rect 18795 15511 18837 15520
rect 17972 15352 18260 15392
rect 18507 15392 18549 15401
rect 18507 15352 18508 15392
rect 18548 15352 18549 15392
rect 17932 15343 17972 15352
rect 18507 15343 18549 15352
rect 18699 15392 18741 15401
rect 18699 15352 18700 15392
rect 18740 15352 18741 15392
rect 18699 15343 18741 15352
rect 17643 15308 17685 15317
rect 17643 15268 17644 15308
rect 17684 15268 17685 15308
rect 17643 15259 17685 15268
rect 18232 15140 18600 15149
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18232 15091 18600 15100
rect 18123 14552 18165 14561
rect 18123 14512 18124 14552
rect 18164 14512 18165 14552
rect 18123 14503 18165 14512
rect 17547 13964 17589 13973
rect 17547 13924 17548 13964
rect 17588 13924 17589 13964
rect 17547 13915 17589 13924
rect 17548 13830 17588 13915
rect 17356 13796 17396 13805
rect 16876 13756 17356 13796
rect 16876 13208 16916 13756
rect 17356 13747 17396 13756
rect 16876 13159 16916 13168
rect 17259 13208 17301 13217
rect 17259 13168 17260 13208
rect 17300 13168 17301 13208
rect 17259 13159 17301 13168
rect 18124 13208 18164 14503
rect 18508 14216 18548 14225
rect 18700 14216 18740 15343
rect 18548 14176 18740 14216
rect 18508 13973 18548 14176
rect 18507 13964 18549 13973
rect 18507 13924 18508 13964
rect 18548 13924 18549 13964
rect 18507 13915 18549 13924
rect 18232 13628 18600 13637
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18232 13579 18600 13588
rect 18124 13159 18164 13168
rect 17260 13074 17300 13159
rect 18699 12452 18741 12461
rect 18699 12412 18700 12452
rect 18740 12412 18741 12452
rect 18699 12403 18741 12412
rect 18232 12116 18600 12125
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18232 12067 18600 12076
rect 18124 11696 18164 11705
rect 13612 11024 13652 11033
rect 10252 10975 10292 10984
rect 12844 10984 13612 11024
rect 9580 10772 9620 10781
rect 9195 9680 9237 9689
rect 9195 9640 9196 9680
rect 9236 9640 9237 9680
rect 9195 9631 9237 9640
rect 9196 9546 9236 9631
rect 8044 9463 8084 9472
rect 9580 8009 9620 10732
rect 12747 10268 12789 10277
rect 12747 10228 12748 10268
rect 12788 10228 12789 10268
rect 12747 10219 12789 10228
rect 9868 10184 9908 10193
rect 9868 9689 9908 10144
rect 12556 10184 12596 10193
rect 10731 10100 10773 10109
rect 10731 10060 10732 10100
rect 10772 10060 10773 10100
rect 12556 10100 12596 10144
rect 12748 10184 12788 10219
rect 12748 10133 12788 10144
rect 12651 10100 12693 10109
rect 12556 10060 12652 10100
rect 12692 10060 12693 10100
rect 10731 10051 10773 10060
rect 12651 10051 12693 10060
rect 10540 10016 10580 10025
rect 10348 9976 10540 10016
rect 9867 9680 9909 9689
rect 9867 9640 9868 9680
rect 9908 9640 9909 9680
rect 9867 9631 9909 9640
rect 10348 9596 10388 9976
rect 10540 9967 10580 9976
rect 10348 9547 10388 9556
rect 10732 9512 10772 10051
rect 12748 9680 12788 9689
rect 12844 9680 12884 10984
rect 13612 10975 13652 10984
rect 15436 11024 15476 11033
rect 12940 10772 12980 10781
rect 12940 10184 12980 10732
rect 15340 10436 15380 10445
rect 15436 10436 15476 10984
rect 16108 11024 16148 11033
rect 16300 11024 16340 11033
rect 16148 10984 16300 11024
rect 16108 10975 16148 10984
rect 16300 10975 16340 10984
rect 16491 11024 16533 11033
rect 16491 10984 16492 11024
rect 16532 10984 16533 11024
rect 16491 10975 16533 10984
rect 16684 11024 16724 11033
rect 15380 10396 15476 10436
rect 15340 10387 15380 10396
rect 13131 10268 13173 10277
rect 13131 10228 13132 10268
rect 13172 10228 13173 10268
rect 13131 10219 13173 10228
rect 12940 10135 12980 10144
rect 12788 9640 12884 9680
rect 12748 9631 12788 9640
rect 11596 9512 11636 9521
rect 10732 9463 10772 9472
rect 11500 9472 11596 9512
rect 7563 8000 7605 8009
rect 7563 7960 7564 8000
rect 7604 7960 7605 8000
rect 7563 7951 7605 7960
rect 9579 8000 9621 8009
rect 9579 7960 9580 8000
rect 9620 7960 9621 8000
rect 9579 7951 9621 7960
rect 11211 8000 11253 8009
rect 11211 7960 11212 8000
rect 11252 7960 11253 8000
rect 11211 7951 11253 7960
rect 7564 7866 7604 7951
rect 11019 7412 11061 7421
rect 11019 7372 11020 7412
rect 11060 7372 11061 7412
rect 11019 7363 11061 7372
rect 9676 6488 9716 6497
rect 7179 6404 7221 6413
rect 7179 6364 7180 6404
rect 7220 6364 7221 6404
rect 7179 6355 7221 6364
rect 7371 6320 7413 6329
rect 9676 6320 9716 6448
rect 10155 6404 10197 6413
rect 10155 6364 10156 6404
rect 10196 6364 10197 6404
rect 10155 6355 10197 6364
rect 7371 6280 7372 6320
rect 7412 6280 7413 6320
rect 7371 6271 7413 6280
rect 9388 6280 9716 6320
rect 6987 5060 7029 5069
rect 6987 5020 6988 5060
rect 7028 5020 7029 5060
rect 6987 5011 7029 5020
rect 6891 4976 6933 4985
rect 6891 4936 6892 4976
rect 6932 4936 6933 4976
rect 6891 4927 6933 4936
rect 6988 4926 7028 5011
rect 7372 4976 7412 6271
rect 7372 4901 7412 4936
rect 8235 4976 8277 4985
rect 8235 4936 8236 4976
rect 8276 4936 8277 4976
rect 8235 4927 8277 4936
rect 6316 4843 6356 4852
rect 7371 4892 7413 4901
rect 7371 4852 7372 4892
rect 7412 4852 7413 4892
rect 7371 4843 7413 4852
rect 8236 4842 8276 4927
rect 9388 4892 9428 6280
rect 9771 6236 9813 6245
rect 9771 6196 9772 6236
rect 9812 6196 9813 6236
rect 9771 6187 9813 6196
rect 9772 5648 9812 6187
rect 9772 5599 9812 5608
rect 10156 5648 10196 6355
rect 10348 6329 10388 6414
rect 10347 6320 10389 6329
rect 10347 6280 10348 6320
rect 10388 6280 10389 6320
rect 10347 6271 10389 6280
rect 10156 5599 10196 5608
rect 11020 5648 11060 7363
rect 11212 7160 11252 7951
rect 11500 7421 11540 9472
rect 11596 9463 11636 9472
rect 11499 7412 11541 7421
rect 11499 7372 11500 7412
rect 11540 7372 11541 7412
rect 11499 7363 11541 7372
rect 11500 7278 11540 7363
rect 11212 7111 11252 7120
rect 12171 7160 12213 7169
rect 12748 7160 12788 7169
rect 12171 7120 12172 7160
rect 12212 7120 12213 7160
rect 12171 7111 12213 7120
rect 12652 7120 12748 7160
rect 12172 7026 12212 7111
rect 12364 7076 12404 7085
rect 12172 6488 12212 6499
rect 12172 6413 12212 6448
rect 12171 6404 12213 6413
rect 12171 6364 12172 6404
rect 12212 6364 12213 6404
rect 12171 6355 12213 6364
rect 12364 5900 12404 7036
rect 12652 6656 12692 7120
rect 12748 7111 12788 7120
rect 12652 6607 12692 6616
rect 12364 5851 12404 5860
rect 13132 6488 13172 10219
rect 13324 10184 13364 10195
rect 16492 10193 16532 10975
rect 13324 10109 13364 10144
rect 14187 10184 14229 10193
rect 14187 10144 14188 10184
rect 14228 10144 14229 10184
rect 14187 10135 14229 10144
rect 16491 10184 16533 10193
rect 16491 10144 16492 10184
rect 16532 10144 16533 10184
rect 16491 10135 16533 10144
rect 13323 10100 13365 10109
rect 13323 10060 13324 10100
rect 13364 10060 13365 10100
rect 13323 10051 13365 10060
rect 14188 10050 14228 10135
rect 16684 10109 16724 10984
rect 17547 11024 17589 11033
rect 17547 10984 17548 11024
rect 17588 10984 17589 11024
rect 17547 10975 17589 10984
rect 17548 10890 17588 10975
rect 18124 10277 18164 11656
rect 18700 11192 18740 12403
rect 18796 12368 18836 15511
rect 19948 15401 19988 15688
rect 20044 15560 20084 16267
rect 20044 15511 20084 15520
rect 20140 16232 20180 16241
rect 19947 15392 19989 15401
rect 19947 15352 19948 15392
rect 19988 15352 19989 15392
rect 19947 15343 19989 15352
rect 20140 15065 20180 16192
rect 20332 15989 20372 17032
rect 20428 17023 20468 17032
rect 20716 16820 20756 16829
rect 20428 16780 20716 16820
rect 20331 15980 20373 15989
rect 20331 15940 20332 15980
rect 20372 15940 20373 15980
rect 20331 15931 20373 15940
rect 20428 15560 20468 16780
rect 20716 16771 20756 16780
rect 20236 15308 20276 15317
rect 20139 15056 20181 15065
rect 20139 15016 20140 15056
rect 20180 15016 20181 15056
rect 20139 15007 20181 15016
rect 20140 14561 20180 15007
rect 20236 14729 20276 15268
rect 20428 15065 20468 15520
rect 20427 15056 20469 15065
rect 20427 15016 20428 15056
rect 20468 15016 20469 15056
rect 20427 15007 20469 15016
rect 20235 14720 20277 14729
rect 20235 14680 20236 14720
rect 20276 14680 20277 14720
rect 20235 14671 20277 14680
rect 20139 14552 20181 14561
rect 20139 14512 20140 14552
rect 20180 14512 20181 14552
rect 20139 14503 20181 14512
rect 20812 14477 20852 19795
rect 21196 19256 21236 19265
rect 21196 17156 21236 19216
rect 22444 19256 22484 19265
rect 21292 17156 21332 17165
rect 21196 17116 21292 17156
rect 21292 17107 21332 17116
rect 21291 16400 21333 16409
rect 21291 16360 21292 16400
rect 21332 16360 21333 16400
rect 21291 16351 21333 16360
rect 21292 16266 21332 16351
rect 22444 15569 22484 19216
rect 23404 17072 23444 19804
rect 25228 17669 25268 19963
rect 26860 18500 26900 18511
rect 26860 18425 26900 18460
rect 26859 18416 26901 18425
rect 26859 18376 26860 18416
rect 26900 18376 26901 18416
rect 26859 18367 26901 18376
rect 26187 18332 26229 18341
rect 26187 18292 26188 18332
rect 26228 18292 26229 18332
rect 26187 18283 26229 18292
rect 26668 18332 26708 18341
rect 25707 17744 25749 17753
rect 25707 17704 25708 17744
rect 25748 17704 25749 17744
rect 25707 17695 25749 17704
rect 26092 17744 26132 17755
rect 25227 17660 25269 17669
rect 25227 17620 25228 17660
rect 25268 17620 25269 17660
rect 25227 17611 25269 17620
rect 23404 17023 23444 17032
rect 24076 16820 24116 16829
rect 22443 15560 22485 15569
rect 22443 15520 22444 15560
rect 22484 15520 22485 15560
rect 22443 15511 22485 15520
rect 22635 15560 22677 15569
rect 22635 15520 22636 15560
rect 22676 15520 22677 15560
rect 22635 15511 22677 15520
rect 22923 15560 22965 15569
rect 22923 15520 22924 15560
rect 22964 15520 22965 15560
rect 22923 15511 22965 15520
rect 22252 15308 22292 15317
rect 22252 15140 22292 15268
rect 22060 15100 22292 15140
rect 21291 14720 21333 14729
rect 21291 14680 21292 14720
rect 21332 14680 21333 14720
rect 21291 14671 21333 14680
rect 21676 14720 21716 14729
rect 21292 14586 21332 14671
rect 21676 14477 21716 14680
rect 20811 14468 20853 14477
rect 20811 14428 20812 14468
rect 20852 14428 20853 14468
rect 20811 14419 20853 14428
rect 21291 14468 21333 14477
rect 21291 14428 21292 14468
rect 21332 14428 21333 14468
rect 21291 14419 21333 14428
rect 21675 14468 21717 14477
rect 21675 14428 21676 14468
rect 21716 14428 21717 14468
rect 21675 14419 21717 14428
rect 19472 14384 19840 14393
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19472 14335 19840 14344
rect 19180 14048 19220 14057
rect 19180 13460 19220 14008
rect 19276 13460 19316 13469
rect 19180 13420 19276 13460
rect 19276 13411 19316 13420
rect 18987 13208 19029 13217
rect 18987 13168 18988 13208
rect 19028 13168 19029 13208
rect 18987 13159 19029 13168
rect 18988 12629 19028 13159
rect 19472 12872 19840 12881
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19472 12823 19840 12832
rect 21292 12629 21332 14419
rect 18987 12620 19029 12629
rect 18987 12580 18988 12620
rect 19028 12580 19029 12620
rect 18987 12571 19029 12580
rect 21291 12620 21333 12629
rect 21291 12580 21292 12620
rect 21332 12580 21333 12620
rect 21291 12571 21333 12580
rect 18796 12319 18836 12328
rect 18988 11696 19028 12571
rect 19371 12536 19413 12545
rect 19371 12496 19372 12536
rect 19412 12496 19413 12536
rect 19371 12487 19413 12496
rect 21292 12536 21332 12571
rect 19372 12402 19412 12487
rect 21292 12485 21332 12496
rect 21675 12536 21717 12545
rect 21675 12496 21676 12536
rect 21716 12496 21717 12536
rect 21675 12487 21717 12496
rect 18988 11647 19028 11656
rect 19472 11360 19840 11369
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19472 11311 19840 11320
rect 21099 11360 21141 11369
rect 21099 11320 21100 11360
rect 21140 11320 21141 11360
rect 21099 11311 21141 11320
rect 18700 11143 18740 11152
rect 20716 11024 20756 11033
rect 20620 10984 20716 11024
rect 18232 10604 18600 10613
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18232 10555 18600 10564
rect 18123 10268 18165 10277
rect 18123 10228 18124 10268
rect 18164 10228 18165 10268
rect 18123 10219 18165 10228
rect 16683 10100 16725 10109
rect 16683 10060 16684 10100
rect 16724 10060 16725 10100
rect 16683 10051 16725 10060
rect 17067 10100 17109 10109
rect 17067 10060 17068 10100
rect 17108 10060 17109 10100
rect 17067 10051 17109 10060
rect 17068 8672 17108 10051
rect 17068 8623 17108 8632
rect 17932 8672 17972 8681
rect 16684 8588 16724 8597
rect 16492 8548 16684 8588
rect 16492 8168 16532 8548
rect 16684 8539 16724 8548
rect 16492 8119 16532 8128
rect 14763 8000 14805 8009
rect 14763 7960 14764 8000
rect 14804 7960 14805 8000
rect 14763 7951 14805 7960
rect 15819 8000 15861 8009
rect 15819 7960 15820 8000
rect 15860 7960 15861 8000
rect 15819 7951 15861 7960
rect 14764 7412 14804 7951
rect 15820 7866 15860 7951
rect 14764 7363 14804 7372
rect 13515 7160 13557 7169
rect 13612 7160 13652 7169
rect 13515 7120 13516 7160
rect 13556 7120 13612 7160
rect 13515 7111 13557 7120
rect 13612 7111 13652 7120
rect 12171 5732 12213 5741
rect 12171 5692 12172 5732
rect 12212 5692 12213 5732
rect 12171 5683 12213 5692
rect 13035 5732 13077 5741
rect 13035 5692 13036 5732
rect 13076 5692 13077 5732
rect 13035 5683 13077 5692
rect 11020 5599 11060 5608
rect 12172 5598 12212 5683
rect 13036 5648 13076 5683
rect 13036 5597 13076 5608
rect 9388 4843 9428 4852
rect 4628 4180 4820 4220
rect 12939 4220 12981 4229
rect 12939 4180 12940 4220
rect 12980 4180 12981 4220
rect 4588 4171 4628 4180
rect 12939 4171 12981 4180
rect 844 4086 884 4171
rect 12940 4086 12980 4171
rect 651 3968 693 3977
rect 651 3928 652 3968
rect 692 3928 693 3968
rect 651 3919 693 3928
rect 11787 3968 11829 3977
rect 11787 3928 11788 3968
rect 11828 3928 11829 3968
rect 11787 3919 11829 3928
rect 12747 3968 12789 3977
rect 12747 3928 12748 3968
rect 12788 3928 12789 3968
rect 12747 3919 12789 3928
rect 652 3834 692 3919
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 11788 3548 11828 3919
rect 12748 3834 12788 3919
rect 11788 3499 11828 3508
rect 13132 3473 13172 6448
rect 12171 3464 12213 3473
rect 12171 3424 12172 3464
rect 12212 3424 12213 3464
rect 12171 3415 12213 3424
rect 12651 3464 12693 3473
rect 12651 3424 12652 3464
rect 12692 3424 12693 3464
rect 12651 3415 12693 3424
rect 13036 3464 13076 3473
rect 843 3380 885 3389
rect 843 3340 844 3380
rect 884 3340 885 3380
rect 843 3331 885 3340
rect 844 3246 884 3331
rect 12172 3330 12212 3415
rect 651 3212 693 3221
rect 651 3172 652 3212
rect 692 3172 693 3212
rect 651 3163 693 3172
rect 652 3078 692 3163
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 843 2708 885 2717
rect 843 2668 844 2708
rect 884 2668 885 2708
rect 843 2659 885 2668
rect 844 2574 884 2659
rect 12652 2624 12692 3415
rect 13036 2624 13076 3424
rect 13131 3464 13173 3473
rect 13131 3424 13132 3464
rect 13172 3424 13173 3464
rect 13131 3415 13173 3424
rect 13516 2624 13556 7111
rect 17644 6404 17684 6413
rect 17644 6245 17684 6364
rect 17452 6236 17492 6245
rect 16684 6196 17452 6236
rect 16684 5648 16724 6196
rect 17452 6187 17492 6196
rect 17643 6236 17685 6245
rect 17643 6196 17644 6236
rect 17684 6196 17685 6236
rect 17643 6187 17685 6196
rect 16779 5732 16821 5741
rect 16779 5692 16780 5732
rect 16820 5692 16821 5732
rect 16779 5683 16821 5692
rect 17067 5732 17109 5741
rect 17067 5692 17068 5732
rect 17108 5692 17109 5732
rect 17067 5683 17109 5692
rect 16684 5599 16724 5608
rect 14187 4136 14229 4145
rect 14187 4096 14188 4136
rect 14228 4096 14229 4136
rect 14187 4087 14229 4096
rect 16299 4136 16341 4145
rect 16299 4096 16300 4136
rect 16340 4096 16341 4136
rect 16299 4087 16341 4096
rect 14188 3632 14228 4087
rect 16300 4002 16340 4087
rect 14188 3583 14228 3592
rect 16300 3464 16340 3473
rect 16300 2885 16340 3424
rect 16684 3464 16724 3473
rect 16780 3464 16820 5683
rect 17068 5648 17108 5683
rect 17932 5657 17972 8632
rect 18124 8000 18164 10219
rect 19472 9848 19840 9857
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19472 9799 19840 9808
rect 20332 9512 20372 9521
rect 18232 9092 18600 9101
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18232 9043 18600 9052
rect 20332 8849 20372 9472
rect 19083 8840 19125 8849
rect 19083 8800 19084 8840
rect 19124 8800 19125 8840
rect 19083 8791 19125 8800
rect 20331 8840 20373 8849
rect 20331 8800 20332 8840
rect 20372 8800 20373 8840
rect 20331 8791 20373 8800
rect 19084 8706 19124 8791
rect 20620 8681 20660 10984
rect 20716 10975 20756 10984
rect 21003 10184 21045 10193
rect 21003 10144 21004 10184
rect 21044 10144 21045 10184
rect 21003 10135 21045 10144
rect 21100 10184 21140 11311
rect 21676 11033 21716 12487
rect 21771 12284 21813 12293
rect 21771 12244 21772 12284
rect 21812 12244 21813 12284
rect 21771 12235 21813 12244
rect 21675 11024 21717 11033
rect 21675 10984 21676 11024
rect 21716 10984 21717 11024
rect 21675 10975 21717 10984
rect 21676 10890 21716 10975
rect 21100 10135 21140 10144
rect 21483 10184 21525 10193
rect 21483 10144 21484 10184
rect 21524 10144 21525 10184
rect 21483 10135 21525 10144
rect 21004 9680 21044 10135
rect 21484 10050 21524 10135
rect 21004 9631 21044 9640
rect 21580 10016 21620 10025
rect 21580 9521 21620 9976
rect 21579 9512 21621 9521
rect 21579 9472 21580 9512
rect 21620 9472 21621 9512
rect 21579 9463 21621 9472
rect 20619 8672 20661 8681
rect 20619 8632 20620 8672
rect 20660 8632 20661 8672
rect 20619 8623 20661 8632
rect 19472 8336 19840 8345
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19472 8287 19840 8296
rect 18124 7673 18164 7960
rect 18699 8000 18741 8009
rect 18699 7960 18700 8000
rect 18740 7960 18741 8000
rect 18699 7951 18741 7960
rect 18700 7832 18740 7951
rect 18123 7664 18165 7673
rect 18123 7624 18124 7664
rect 18164 7624 18165 7664
rect 18123 7615 18165 7624
rect 18232 7580 18600 7589
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18232 7531 18600 7540
rect 18508 6320 18548 6329
rect 18123 6236 18165 6245
rect 18508 6236 18548 6280
rect 18123 6196 18124 6236
rect 18164 6196 18548 6236
rect 18123 6187 18165 6196
rect 17068 5597 17108 5608
rect 17931 5648 17973 5657
rect 17931 5608 17932 5648
rect 17972 5608 17973 5648
rect 17931 5599 17973 5608
rect 16971 4220 17013 4229
rect 16971 4180 16972 4220
rect 17012 4180 17013 4220
rect 16971 4171 17013 4180
rect 16972 4086 17012 4171
rect 17643 4136 17685 4145
rect 17643 4096 17644 4136
rect 17684 4096 17780 4136
rect 17643 4087 17685 4096
rect 17548 3977 17588 4058
rect 17644 4002 17684 4087
rect 17547 3968 17589 3977
rect 17547 3923 17548 3968
rect 17588 3923 17589 3968
rect 17547 3919 17589 3923
rect 17548 3914 17588 3919
rect 17643 3884 17685 3893
rect 17643 3844 17644 3884
rect 17684 3844 17685 3884
rect 17643 3835 17685 3844
rect 17547 3800 17589 3809
rect 17547 3760 17548 3800
rect 17588 3760 17589 3800
rect 17547 3751 17589 3760
rect 17548 3473 17588 3751
rect 16724 3424 16820 3464
rect 17547 3464 17589 3473
rect 17547 3424 17548 3464
rect 17588 3424 17589 3464
rect 16684 3415 16724 3424
rect 17547 3415 17589 3424
rect 17548 3330 17588 3415
rect 17644 2960 17684 3835
rect 17068 2920 17684 2960
rect 16299 2876 16341 2885
rect 16299 2836 16300 2876
rect 16340 2836 16341 2876
rect 16299 2827 16341 2836
rect 16875 2876 16917 2885
rect 16875 2836 16876 2876
rect 16916 2836 16917 2876
rect 16875 2827 16917 2836
rect 16876 2742 16916 2827
rect 14668 2708 14708 2717
rect 14708 2668 14900 2708
rect 14668 2659 14708 2668
rect 13036 2584 13516 2624
rect 12652 2575 12692 2584
rect 13516 2575 13556 2584
rect 13611 2624 13653 2633
rect 13611 2584 13612 2624
rect 13652 2584 13653 2624
rect 13611 2575 13653 2584
rect 14860 2624 14900 2668
rect 15532 2633 15572 2718
rect 17068 2708 17108 2920
rect 17547 2792 17589 2801
rect 17547 2752 17548 2792
rect 17588 2752 17589 2792
rect 17547 2743 17589 2752
rect 17068 2659 17108 2668
rect 17452 2633 17492 2718
rect 17548 2658 17588 2743
rect 14860 2575 14900 2584
rect 15531 2624 15573 2633
rect 15531 2584 15532 2624
rect 15572 2584 15573 2624
rect 15531 2575 15573 2584
rect 17451 2624 17493 2633
rect 17451 2584 17452 2624
rect 17492 2584 17493 2624
rect 17451 2575 17493 2584
rect 17644 2624 17684 2920
rect 17740 2624 17780 4096
rect 17835 3968 17877 3977
rect 17835 3928 17836 3968
rect 17876 3928 17877 3968
rect 17835 3919 17877 3928
rect 17836 3834 17876 3919
rect 17932 3809 17972 5599
rect 18027 4052 18069 4061
rect 18027 4012 18028 4052
rect 18068 4012 18069 4052
rect 18027 4003 18069 4012
rect 18028 3918 18068 4003
rect 17931 3800 17973 3809
rect 18124 3800 18164 6187
rect 18232 6068 18600 6077
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18232 6019 18600 6028
rect 18700 5741 18740 7792
rect 19947 7664 19989 7673
rect 19947 7624 19948 7664
rect 19988 7624 19989 7664
rect 19947 7615 19989 7624
rect 19472 6824 19840 6833
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19472 6775 19840 6784
rect 19180 6488 19220 6497
rect 19084 5900 19124 5909
rect 19180 5900 19220 6448
rect 19124 5860 19220 5900
rect 19084 5851 19124 5860
rect 18699 5732 18741 5741
rect 18699 5692 18700 5732
rect 18740 5692 18741 5732
rect 18699 5683 18741 5692
rect 19659 5648 19701 5657
rect 19659 5608 19660 5648
rect 19700 5608 19701 5648
rect 19659 5599 19701 5608
rect 19660 5514 19700 5599
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 17931 3760 17932 3800
rect 17972 3760 17973 3800
rect 17931 3751 17973 3760
rect 18028 3760 18164 3800
rect 18700 4136 18740 4145
rect 18028 2708 18068 3760
rect 18700 3632 18740 4096
rect 19371 3968 19413 3977
rect 19371 3928 19372 3968
rect 19412 3928 19413 3968
rect 19371 3919 19413 3928
rect 18700 3583 18740 3592
rect 19372 3548 19412 3919
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 19372 3499 19412 3508
rect 19756 3464 19796 3473
rect 19948 3464 19988 7615
rect 20620 5648 20660 8623
rect 21772 6320 21812 12235
rect 21963 10436 22005 10445
rect 21963 10396 21964 10436
rect 22004 10396 22005 10436
rect 21963 10387 22005 10396
rect 21964 10302 22004 10387
rect 21868 10193 21908 10278
rect 21867 10184 21909 10193
rect 21867 10144 21868 10184
rect 21908 10144 21909 10184
rect 21867 10135 21909 10144
rect 22060 10184 22100 15100
rect 22539 15056 22581 15065
rect 22539 15016 22540 15056
rect 22580 15016 22581 15056
rect 22539 15007 22581 15016
rect 22540 14720 22580 15007
rect 22540 14671 22580 14680
rect 22636 11369 22676 15511
rect 22924 15426 22964 15511
rect 23691 14552 23733 14561
rect 23691 14512 23692 14552
rect 23732 14512 23733 14552
rect 23691 14503 23733 14512
rect 23692 14418 23732 14503
rect 23116 13376 23156 13385
rect 23156 13336 23540 13376
rect 23116 13327 23156 13336
rect 23020 13208 23060 13217
rect 23020 12629 23060 13168
rect 23212 13208 23252 13217
rect 23500 13208 23540 13336
rect 23252 13168 23348 13208
rect 23212 13159 23252 13168
rect 23019 12620 23061 12629
rect 23019 12580 23020 12620
rect 23060 12580 23061 12620
rect 23019 12571 23061 12580
rect 23212 12620 23252 12629
rect 22731 12536 22773 12545
rect 22731 12496 22732 12536
rect 22772 12496 22773 12536
rect 22731 12487 22773 12496
rect 23020 12536 23060 12571
rect 22732 12402 22772 12487
rect 23020 12461 23060 12496
rect 23019 12452 23061 12461
rect 23019 12412 23020 12452
rect 23060 12412 23061 12452
rect 23019 12403 23061 12412
rect 23212 11696 23252 12580
rect 23308 12545 23348 13168
rect 23500 13159 23540 13168
rect 23691 13040 23733 13049
rect 23691 13000 23692 13040
rect 23732 13000 23733 13040
rect 23691 12991 23733 13000
rect 23307 12536 23349 12545
rect 23500 12536 23540 12545
rect 23307 12496 23308 12536
rect 23348 12496 23349 12536
rect 23307 12487 23349 12496
rect 23404 12496 23500 12536
rect 23308 11696 23348 11705
rect 23212 11656 23308 11696
rect 23308 11647 23348 11656
rect 23404 11696 23444 12496
rect 23500 12487 23540 12496
rect 23596 12536 23636 12545
rect 23596 12377 23636 12496
rect 23692 12536 23732 12991
rect 23883 12704 23925 12713
rect 23883 12664 23884 12704
rect 23924 12664 23925 12704
rect 23883 12655 23925 12664
rect 23787 12620 23829 12629
rect 23787 12580 23788 12620
rect 23828 12580 23829 12620
rect 23787 12571 23829 12580
rect 23692 12487 23732 12496
rect 23788 12486 23828 12571
rect 23884 12536 23924 12655
rect 24076 12545 24116 16780
rect 25228 16241 25268 17611
rect 25708 17610 25748 17695
rect 26092 17669 26132 17704
rect 26091 17660 26133 17669
rect 26091 17620 26092 17660
rect 26132 17620 26133 17660
rect 26091 17611 26133 17620
rect 26188 17156 26228 18283
rect 26668 17753 26708 18292
rect 26667 17744 26709 17753
rect 26956 17744 26996 21568
rect 27051 21559 27093 21568
rect 27052 21474 27092 21559
rect 28203 21524 28245 21533
rect 28203 21484 28204 21524
rect 28244 21484 28245 21524
rect 28203 21475 28245 21484
rect 28204 21390 28244 21475
rect 28780 21449 28820 25264
rect 29643 25255 29685 25264
rect 30603 25304 30645 25313
rect 30603 25264 30604 25304
rect 30644 25264 30645 25304
rect 30603 25255 30645 25264
rect 29644 25170 29684 25255
rect 30219 24380 30261 24389
rect 30219 24340 30220 24380
rect 30260 24340 30261 24380
rect 30219 24331 30261 24340
rect 30220 23792 30260 24331
rect 30604 23801 30644 25255
rect 31564 24641 31604 29119
rect 33352 28748 33720 28757
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33352 28699 33720 28708
rect 32908 28328 32948 28337
rect 32524 27404 32564 27413
rect 32524 26825 32564 27364
rect 32523 26816 32565 26825
rect 32523 26776 32524 26816
rect 32564 26776 32565 26816
rect 32523 26767 32565 26776
rect 32908 26573 32948 28288
rect 33676 27656 33716 27665
rect 33772 27656 33812 30631
rect 34060 30269 34100 31312
rect 34592 31016 34960 31025
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34592 30967 34960 30976
rect 35116 30857 35156 32152
rect 36940 32117 36980 32824
rect 37612 32696 37652 32705
rect 37420 32656 37612 32696
rect 37227 32192 37269 32201
rect 37227 32152 37228 32192
rect 37268 32152 37269 32192
rect 37227 32143 37269 32152
rect 37420 32192 37460 32656
rect 37612 32647 37652 32656
rect 37708 32285 37748 34336
rect 38572 34376 38612 36679
rect 38955 36560 38997 36569
rect 38955 36520 38956 36560
rect 38996 36520 38997 36560
rect 38955 36511 38997 36520
rect 38956 36426 38996 36511
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 93832 36308 94200 36317
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 93832 36259 94200 36268
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 95072 35552 95440 35561
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95072 35503 95440 35512
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 93832 34796 94200 34805
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 93832 34747 94200 34756
rect 37707 32276 37749 32285
rect 37707 32236 37708 32276
rect 37748 32236 37749 32276
rect 37707 32227 37749 32236
rect 38092 32276 38132 32285
rect 37420 32143 37460 32152
rect 37612 32192 37652 32203
rect 36267 32108 36309 32117
rect 36267 32068 36268 32108
rect 36308 32068 36309 32108
rect 36267 32059 36309 32068
rect 36939 32108 36981 32117
rect 36939 32068 36940 32108
rect 36980 32068 36981 32108
rect 36939 32059 36981 32068
rect 36268 31974 36308 32059
rect 37228 32058 37268 32143
rect 37612 32117 37652 32152
rect 37611 32108 37653 32117
rect 37611 32068 37612 32108
rect 37652 32068 37653 32108
rect 37611 32059 37653 32068
rect 37323 31940 37365 31949
rect 37323 31900 37324 31940
rect 37364 31900 37365 31940
rect 37323 31891 37365 31900
rect 37324 31806 37364 31891
rect 37132 31520 37172 31529
rect 37708 31520 37748 32227
rect 37995 32192 38037 32201
rect 37995 32152 37996 32192
rect 38036 32152 38037 32192
rect 37995 32143 38037 32152
rect 37996 32058 38036 32143
rect 37708 31480 37844 31520
rect 36171 31436 36213 31445
rect 36171 31396 36172 31436
rect 36212 31396 36213 31436
rect 36171 31387 36213 31396
rect 36172 31352 36212 31387
rect 36172 31301 36212 31312
rect 36460 31352 36500 31361
rect 35500 31184 35540 31193
rect 34635 30848 34677 30857
rect 34635 30808 34636 30848
rect 34676 30808 34677 30848
rect 34635 30799 34677 30808
rect 35115 30848 35157 30857
rect 35115 30808 35116 30848
rect 35156 30808 35157 30848
rect 35115 30799 35157 30808
rect 34636 30714 34676 30799
rect 35500 30773 35540 31144
rect 35979 30848 36021 30857
rect 35979 30808 35980 30848
rect 36020 30808 36021 30848
rect 35979 30799 36021 30808
rect 35499 30764 35541 30773
rect 35499 30724 35500 30764
rect 35540 30724 35541 30764
rect 35499 30715 35541 30724
rect 35787 30764 35829 30773
rect 35787 30724 35788 30764
rect 35828 30724 35829 30764
rect 35787 30715 35829 30724
rect 34155 30680 34197 30689
rect 34155 30640 34156 30680
rect 34196 30640 34197 30680
rect 34155 30631 34197 30640
rect 35115 30680 35157 30689
rect 35115 30640 35116 30680
rect 35156 30640 35157 30680
rect 35115 30631 35157 30640
rect 35595 30680 35637 30689
rect 35595 30640 35596 30680
rect 35636 30640 35637 30680
rect 35595 30631 35637 30640
rect 35788 30680 35828 30715
rect 35980 30714 36020 30799
rect 36460 30689 36500 31312
rect 37132 30773 37172 31480
rect 37419 31352 37461 31361
rect 37419 31312 37420 31352
rect 37460 31312 37461 31352
rect 37419 31303 37461 31312
rect 37612 31352 37652 31361
rect 37420 31218 37460 31303
rect 37612 30857 37652 31312
rect 37611 30848 37653 30857
rect 37611 30808 37612 30848
rect 37652 30808 37653 30848
rect 37611 30799 37653 30808
rect 37131 30764 37173 30773
rect 37131 30724 37132 30764
rect 37172 30724 37173 30764
rect 37131 30715 37173 30724
rect 34156 30546 34196 30631
rect 35116 30546 35156 30631
rect 34059 30260 34101 30269
rect 34059 30220 34060 30260
rect 34100 30220 34101 30260
rect 34059 30211 34101 30220
rect 34060 29000 34100 30211
rect 34592 29504 34960 29513
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34592 29455 34960 29464
rect 33868 28960 34100 29000
rect 33868 28328 33908 28960
rect 33868 28279 33908 28288
rect 34592 27992 34960 28001
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34592 27943 34960 27952
rect 33716 27616 33812 27656
rect 34540 27656 34580 27665
rect 33676 27607 33716 27616
rect 33352 27236 33720 27245
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33352 27187 33720 27196
rect 33195 26816 33237 26825
rect 33195 26776 33196 26816
rect 33236 26776 33237 26816
rect 33195 26767 33237 26776
rect 34444 26816 34484 26825
rect 34540 26816 34580 27616
rect 34484 26776 34580 26816
rect 34924 27656 34964 27665
rect 33196 26682 33236 26767
rect 34060 26732 34100 26741
rect 33868 26648 33908 26657
rect 33388 26608 33868 26648
rect 32907 26564 32949 26573
rect 32907 26524 32908 26564
rect 32948 26524 32949 26564
rect 32907 26515 32949 26524
rect 33388 26060 33428 26608
rect 33579 26480 33621 26489
rect 33579 26440 33580 26480
rect 33620 26440 33621 26480
rect 33579 26431 33621 26440
rect 33580 26312 33620 26431
rect 33580 26263 33620 26272
rect 33388 26011 33428 26020
rect 33352 25724 33720 25733
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33352 25675 33720 25684
rect 31563 24632 31605 24641
rect 31563 24592 31564 24632
rect 31604 24592 31605 24632
rect 31563 24583 31605 24592
rect 32043 24632 32085 24641
rect 32043 24592 32044 24632
rect 32084 24592 32085 24632
rect 32043 24583 32085 24592
rect 33868 24632 33908 26608
rect 34060 26312 34100 26692
rect 34444 26657 34484 26776
rect 34924 26657 34964 27616
rect 35307 26816 35349 26825
rect 35307 26776 35308 26816
rect 35348 26776 35349 26816
rect 35307 26767 35349 26776
rect 35308 26682 35348 26767
rect 34443 26648 34485 26657
rect 34443 26608 34444 26648
rect 34484 26608 34485 26648
rect 34443 26599 34485 26608
rect 34923 26648 34965 26657
rect 34923 26608 34924 26648
rect 34964 26608 34965 26648
rect 34923 26599 34965 26608
rect 35115 26648 35157 26657
rect 35115 26608 35116 26648
rect 35156 26608 35157 26648
rect 35115 26599 35157 26608
rect 34592 26480 34960 26489
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34592 26431 34960 26440
rect 34060 26263 34100 26272
rect 35116 26144 35156 26599
rect 35116 26095 35156 26104
rect 35596 26144 35636 30631
rect 35788 30629 35828 30640
rect 36459 30680 36501 30689
rect 36459 30640 36460 30680
rect 36500 30640 36501 30680
rect 36459 30631 36501 30640
rect 37132 30680 37172 30715
rect 37804 30680 37844 31480
rect 37996 30680 38036 30689
rect 37804 30640 37996 30680
rect 37132 30630 37172 30640
rect 37996 30631 38036 30640
rect 38092 29849 38132 32236
rect 38283 32192 38325 32201
rect 38283 32152 38284 32192
rect 38324 32152 38325 32192
rect 38283 32143 38325 32152
rect 38284 31604 38324 32143
rect 38284 31555 38324 31564
rect 38475 31436 38517 31445
rect 38475 31396 38476 31436
rect 38516 31396 38517 31436
rect 38475 31387 38517 31396
rect 38476 31302 38516 31387
rect 38572 31361 38612 34336
rect 39724 34208 39764 34217
rect 38859 32276 38901 32285
rect 38859 32236 38860 32276
rect 38900 32236 38901 32276
rect 38859 32227 38901 32236
rect 38763 31940 38805 31949
rect 38763 31900 38764 31940
rect 38804 31900 38805 31940
rect 38763 31891 38805 31900
rect 38571 31352 38613 31361
rect 38571 31312 38572 31352
rect 38612 31312 38613 31352
rect 38571 31303 38613 31312
rect 38764 31352 38804 31891
rect 38764 31303 38804 31312
rect 38860 31352 38900 32227
rect 39724 32201 39764 34168
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 95072 34040 95440 34049
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95072 33991 95440 34000
rect 47500 33704 47540 33713
rect 47540 33664 47828 33704
rect 47500 33655 47540 33664
rect 45675 33452 45717 33461
rect 45675 33412 45676 33452
rect 45716 33412 45717 33452
rect 45675 33403 45717 33412
rect 46827 33452 46869 33461
rect 46827 33412 46828 33452
rect 46868 33412 46869 33452
rect 46827 33403 46869 33412
rect 42507 33032 42549 33041
rect 42507 32992 42508 33032
rect 42548 32992 42549 33032
rect 42507 32983 42549 32992
rect 43371 33032 43413 33041
rect 43371 32992 43372 33032
rect 43412 32992 43413 33032
rect 43371 32983 43413 32992
rect 39915 32276 39957 32285
rect 39915 32236 39916 32276
rect 39956 32236 39957 32276
rect 39915 32227 39957 32236
rect 42508 32276 42548 32983
rect 43372 32898 43412 32983
rect 43563 32948 43605 32957
rect 43563 32908 43564 32948
rect 43604 32908 43605 32948
rect 43563 32899 43605 32908
rect 44331 32948 44373 32957
rect 44331 32908 44332 32948
rect 44372 32908 44373 32948
rect 44331 32899 44373 32908
rect 43564 32814 43604 32899
rect 44332 32780 44372 32899
rect 45004 32864 45044 32873
rect 44332 32740 44660 32780
rect 42508 32227 42548 32236
rect 39723 32192 39765 32201
rect 39723 32152 39724 32192
rect 39764 32152 39765 32192
rect 39723 32143 39765 32152
rect 39916 32142 39956 32227
rect 40012 32192 40052 32201
rect 38860 31303 38900 31312
rect 39436 30848 39476 30857
rect 40012 30848 40052 32152
rect 40395 32192 40437 32201
rect 40395 32152 40396 32192
rect 40436 32152 40437 32192
rect 40395 32143 40437 32152
rect 42892 32192 42932 32201
rect 40396 32058 40436 32143
rect 42892 31613 42932 32152
rect 43756 32192 43796 32201
rect 42891 31604 42933 31613
rect 42891 31564 42892 31604
rect 42932 31564 42933 31604
rect 42891 31555 42933 31564
rect 39476 30808 40052 30848
rect 39436 30799 39476 30808
rect 41835 30764 41877 30773
rect 41835 30724 41836 30764
rect 41876 30724 41877 30764
rect 41835 30715 41877 30724
rect 38379 30680 38421 30689
rect 38379 30640 38380 30680
rect 38420 30640 38421 30680
rect 38379 30631 38421 30640
rect 40588 30680 40628 30689
rect 38380 30546 38420 30631
rect 39915 30260 39957 30269
rect 39915 30220 39916 30260
rect 39956 30220 39957 30260
rect 39915 30211 39957 30220
rect 38091 29840 38133 29849
rect 38091 29800 38092 29840
rect 38132 29800 38133 29840
rect 38091 29791 38133 29800
rect 39627 29840 39669 29849
rect 39627 29800 39628 29840
rect 39668 29800 39669 29840
rect 39627 29791 39669 29800
rect 39628 29706 39668 29791
rect 39916 29168 39956 30211
rect 39916 29119 39956 29128
rect 40300 29672 40340 29681
rect 40300 28664 40340 29632
rect 40204 28624 40340 28664
rect 40396 29000 40436 29009
rect 40204 27749 40244 28624
rect 40300 28496 40340 28505
rect 40203 27740 40245 27749
rect 40203 27700 40204 27740
rect 40244 27700 40245 27740
rect 40203 27691 40245 27700
rect 40300 27665 40340 28456
rect 39627 27656 39669 27665
rect 39627 27616 39628 27656
rect 39668 27616 39669 27656
rect 39627 27607 39669 27616
rect 40299 27656 40341 27665
rect 40299 27616 40300 27656
rect 40340 27616 40341 27656
rect 40396 27656 40436 28960
rect 40492 28580 40532 28589
rect 40588 28580 40628 30640
rect 41452 30680 41492 30689
rect 41452 30269 41492 30640
rect 41836 30630 41876 30715
rect 40683 30260 40725 30269
rect 40683 30220 40684 30260
rect 40724 30220 40725 30260
rect 40683 30211 40725 30220
rect 41451 30260 41493 30269
rect 41451 30220 41452 30260
rect 41492 30220 41493 30260
rect 41451 30211 41493 30220
rect 40532 28540 40628 28580
rect 40492 28531 40532 28540
rect 40492 27656 40532 27665
rect 40396 27616 40492 27656
rect 40299 27607 40341 27616
rect 38476 27404 38516 27413
rect 38476 26741 38516 27364
rect 39628 26825 39668 27607
rect 39627 26816 39669 26825
rect 39627 26776 39628 26816
rect 39668 26776 39669 26816
rect 39627 26767 39669 26776
rect 38475 26732 38517 26741
rect 38475 26692 38476 26732
rect 38516 26692 38517 26732
rect 38475 26683 38517 26692
rect 40299 26732 40341 26741
rect 40299 26692 40300 26732
rect 40340 26692 40341 26732
rect 40299 26683 40341 26692
rect 36459 26648 36501 26657
rect 36459 26608 36460 26648
rect 36500 26608 36501 26648
rect 36459 26599 36501 26608
rect 36460 26514 36500 26599
rect 40300 26598 40340 26683
rect 40492 26657 40532 27616
rect 40684 26816 40724 30211
rect 42892 29597 42932 31555
rect 43756 29849 43796 32152
rect 44523 31520 44565 31529
rect 44523 31480 44524 31520
rect 44564 31480 44565 31520
rect 44523 31471 44565 31480
rect 44524 31352 44564 31471
rect 44524 31303 44564 31312
rect 44332 31184 44372 31193
rect 44332 30689 44372 31144
rect 44620 31184 44660 32740
rect 44908 32360 44948 32369
rect 45004 32360 45044 32824
rect 44948 32320 45044 32360
rect 45388 32780 45428 32789
rect 45388 32360 45428 32740
rect 45484 32360 45524 32369
rect 45388 32320 45484 32360
rect 44908 32311 44948 32320
rect 45484 32311 45524 32320
rect 45676 32108 45716 33403
rect 46828 33318 46868 33403
rect 47788 33116 47828 33664
rect 48472 33284 48840 33293
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48472 33235 48840 33244
rect 63592 33284 63960 33293
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63592 33235 63960 33244
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 93832 33284 94200 33293
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 93832 33235 94200 33244
rect 47788 33067 47828 33076
rect 45195 31604 45237 31613
rect 45195 31564 45196 31604
rect 45236 31564 45237 31604
rect 45195 31555 45237 31564
rect 44660 31144 45140 31184
rect 44620 31135 44660 31144
rect 44331 30680 44373 30689
rect 44331 30640 44332 30680
rect 44372 30640 44373 30680
rect 44331 30631 44373 30640
rect 45004 30680 45044 30689
rect 44908 30092 44948 30101
rect 45004 30092 45044 30640
rect 44948 30052 45044 30092
rect 44908 30043 44948 30052
rect 43755 29840 43797 29849
rect 43755 29800 43756 29840
rect 43796 29800 43797 29840
rect 43755 29791 43797 29800
rect 44523 29840 44565 29849
rect 44523 29800 44524 29840
rect 44564 29800 44565 29840
rect 44523 29791 44565 29800
rect 44812 29840 44852 29849
rect 44524 29706 44564 29791
rect 40875 29588 40917 29597
rect 40875 29548 40876 29588
rect 40916 29548 40917 29588
rect 40875 29539 40917 29548
rect 42891 29588 42933 29597
rect 42891 29548 42892 29588
rect 42932 29548 42933 29588
rect 42891 29539 42933 29548
rect 40876 29168 40916 29539
rect 44812 29336 44852 29800
rect 45004 29840 45044 29849
rect 45100 29840 45140 31144
rect 45044 29800 45140 29840
rect 45004 29791 45044 29800
rect 40876 29119 40916 29128
rect 44620 29296 44812 29336
rect 44620 29084 44660 29296
rect 44812 29287 44852 29296
rect 44620 29035 44660 29044
rect 44428 28916 44468 28925
rect 40971 28328 41013 28337
rect 40971 28288 40972 28328
rect 41012 28288 41013 28328
rect 40971 28279 41013 28288
rect 43947 28328 43989 28337
rect 43947 28288 43948 28328
rect 43988 28288 43989 28328
rect 44428 28328 44468 28876
rect 45196 28337 45236 31555
rect 45676 31529 45716 32068
rect 45772 32864 45812 32873
rect 45772 31613 45812 32824
rect 46636 32864 46676 32873
rect 46636 32780 46676 32824
rect 46636 32740 46772 32780
rect 45771 31604 45813 31613
rect 45771 31564 45772 31604
rect 45812 31564 45813 31604
rect 45771 31555 45813 31564
rect 45675 31520 45717 31529
rect 45675 31480 45676 31520
rect 45716 31480 45717 31520
rect 45675 31471 45717 31480
rect 46443 31520 46485 31529
rect 46443 31480 46444 31520
rect 46484 31480 46485 31520
rect 46443 31471 46485 31480
rect 45483 30764 45525 30773
rect 45483 30724 45484 30764
rect 45524 30724 45525 30764
rect 45483 30715 45525 30724
rect 45387 30680 45429 30689
rect 45387 30640 45388 30680
rect 45428 30640 45429 30680
rect 45387 30631 45429 30640
rect 45388 30546 45428 30631
rect 45484 30630 45524 30715
rect 46444 30680 46484 31471
rect 46444 30631 46484 30640
rect 46539 30680 46581 30689
rect 46539 30640 46540 30680
rect 46580 30640 46581 30680
rect 46539 30631 46581 30640
rect 46636 30680 46676 30691
rect 46540 30546 46580 30631
rect 46636 30605 46676 30640
rect 46635 30596 46677 30605
rect 46635 30556 46636 30596
rect 46676 30556 46677 30596
rect 46635 30547 46677 30556
rect 45580 30008 45620 30017
rect 45580 29849 45620 29968
rect 46732 29849 46772 32740
rect 49712 32528 50080 32537
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 49712 32479 50080 32488
rect 64832 32528 65200 32537
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 64832 32479 65200 32488
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 95072 32528 95440 32537
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95072 32479 95440 32488
rect 48472 31772 48840 31781
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48472 31723 48840 31732
rect 63592 31772 63960 31781
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63592 31723 63960 31732
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 93832 31772 94200 31781
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 93832 31723 94200 31732
rect 49712 31016 50080 31025
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 49712 30967 50080 30976
rect 64832 31016 65200 31025
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 64832 30967 65200 30976
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 95072 31016 95440 31025
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95072 30967 95440 30976
rect 49228 30680 49268 30689
rect 47499 30596 47541 30605
rect 47499 30556 47500 30596
rect 47540 30556 47541 30596
rect 47499 30547 47541 30556
rect 48555 30596 48597 30605
rect 48555 30556 48556 30596
rect 48596 30556 48597 30596
rect 48555 30547 48597 30556
rect 47500 30462 47540 30547
rect 48556 30462 48596 30547
rect 47308 30428 47348 30437
rect 46924 30388 47308 30428
rect 45292 29840 45332 29849
rect 44524 28328 44564 28337
rect 44428 28288 44524 28328
rect 43947 28279 43989 28288
rect 44524 28279 44564 28288
rect 44907 28328 44949 28337
rect 44907 28288 44908 28328
rect 44948 28288 44949 28328
rect 44907 28279 44949 28288
rect 45195 28328 45237 28337
rect 45195 28288 45196 28328
rect 45236 28288 45237 28328
rect 45195 28279 45237 28288
rect 40972 28194 41012 28279
rect 43948 27749 43988 28279
rect 44908 28194 44948 28279
rect 45292 27749 45332 29800
rect 45579 29840 45621 29849
rect 45579 29800 45580 29840
rect 45620 29800 45621 29840
rect 45579 29791 45621 29800
rect 46731 29840 46773 29849
rect 46731 29800 46732 29840
rect 46772 29800 46773 29840
rect 46731 29791 46773 29800
rect 46924 29840 46964 30388
rect 47308 30379 47348 30388
rect 48472 30260 48840 30269
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48472 30211 48840 30220
rect 49228 30092 49268 30640
rect 63592 30260 63960 30269
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63592 30211 63960 30220
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 93832 30260 94200 30269
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 93832 30211 94200 30220
rect 49324 30092 49364 30101
rect 49228 30052 49324 30092
rect 49324 30043 49364 30052
rect 46924 29791 46964 29800
rect 47308 29840 47348 29849
rect 45772 29672 45812 29681
rect 45483 29168 45525 29177
rect 45483 29128 45484 29168
rect 45524 29128 45525 29168
rect 45483 29119 45525 29128
rect 45484 29034 45524 29119
rect 45579 28328 45621 28337
rect 45579 28288 45580 28328
rect 45620 28288 45621 28328
rect 45579 28279 45621 28288
rect 45772 28328 45812 29632
rect 46923 29168 46965 29177
rect 46923 29128 46924 29168
rect 46964 29128 46965 29168
rect 46923 29119 46965 29128
rect 46924 28580 46964 29119
rect 46924 28531 46964 28540
rect 47308 28337 47348 29800
rect 48171 29840 48213 29849
rect 48171 29800 48172 29840
rect 48212 29800 48213 29840
rect 48171 29791 48213 29800
rect 48172 29706 48212 29791
rect 49712 29504 50080 29513
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 49712 29455 50080 29464
rect 64832 29504 65200 29513
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 64832 29455 65200 29464
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 95072 29504 95440 29513
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95072 29455 95440 29464
rect 48472 28748 48840 28757
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48472 28699 48840 28708
rect 63592 28748 63960 28757
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63592 28699 63960 28708
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 93832 28748 94200 28757
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 93832 28699 94200 28708
rect 45772 28279 45812 28288
rect 47307 28328 47349 28337
rect 47307 28288 47308 28328
rect 47348 28288 47349 28328
rect 47307 28279 47349 28288
rect 40875 27740 40917 27749
rect 40875 27700 40876 27740
rect 40916 27700 40917 27740
rect 40875 27691 40917 27700
rect 43947 27740 43989 27749
rect 43947 27700 43948 27740
rect 43988 27700 43989 27740
rect 43947 27691 43989 27700
rect 45291 27740 45333 27749
rect 45291 27700 45292 27740
rect 45332 27700 45333 27740
rect 45291 27691 45333 27700
rect 40876 27656 40916 27691
rect 40876 27605 40916 27616
rect 42700 26900 42740 26909
rect 42740 26860 42932 26900
rect 42700 26851 42740 26860
rect 40684 26767 40724 26776
rect 41547 26816 41589 26825
rect 41547 26776 41548 26816
rect 41588 26776 41589 26816
rect 41547 26767 41589 26776
rect 42027 26816 42069 26825
rect 42027 26776 42028 26816
rect 42068 26776 42069 26816
rect 42027 26767 42069 26776
rect 42892 26816 42932 26860
rect 42892 26767 42932 26776
rect 41451 26732 41493 26741
rect 41451 26692 41452 26732
rect 41492 26692 41493 26732
rect 41451 26683 41493 26692
rect 40491 26648 40533 26657
rect 40491 26608 40492 26648
rect 40532 26608 40533 26648
rect 40491 26599 40533 26608
rect 41452 26312 41492 26683
rect 41548 26682 41588 26767
rect 41452 26263 41492 26272
rect 35596 26095 35636 26104
rect 36555 26144 36597 26153
rect 36555 26104 36556 26144
rect 36596 26104 36597 26144
rect 36555 26095 36597 26104
rect 34252 26060 34292 26069
rect 34252 25892 34292 26020
rect 34444 25892 34484 25901
rect 34252 25852 34444 25892
rect 33868 24583 33908 24592
rect 34060 24632 34100 24643
rect 31467 24548 31509 24557
rect 31467 24508 31468 24548
rect 31508 24508 31509 24548
rect 31467 24499 31509 24508
rect 31468 24414 31508 24499
rect 31275 24380 31317 24389
rect 31275 24340 31276 24380
rect 31316 24340 31317 24380
rect 31275 24331 31317 24340
rect 31276 24246 31316 24331
rect 30220 23743 30260 23752
rect 30603 23792 30645 23801
rect 30603 23752 30604 23792
rect 30644 23752 30645 23792
rect 30603 23743 30645 23752
rect 31468 23792 31508 23801
rect 30604 23658 30644 23743
rect 29068 21608 29108 21617
rect 28971 21524 29013 21533
rect 29068 21524 29108 21568
rect 31179 21608 31221 21617
rect 31179 21568 31180 21608
rect 31220 21568 31221 21608
rect 31179 21559 31221 21568
rect 28971 21484 28972 21524
rect 29012 21484 29108 21524
rect 28971 21475 29013 21484
rect 31180 21474 31220 21559
rect 28779 21440 28821 21449
rect 28779 21400 28780 21440
rect 28820 21400 28821 21440
rect 28779 21391 28821 21400
rect 31468 21440 31508 23752
rect 31468 21391 31508 21400
rect 28396 21356 28436 21365
rect 28300 21316 28396 21356
rect 28300 20861 28340 21316
rect 28396 21307 28436 21316
rect 27051 20852 27093 20861
rect 27051 20812 27052 20852
rect 27092 20812 27093 20852
rect 27051 20803 27093 20812
rect 28299 20852 28341 20861
rect 28299 20812 28300 20852
rect 28340 20812 28341 20852
rect 28299 20803 28341 20812
rect 27052 20718 27092 20803
rect 28300 20600 28340 20803
rect 28780 20609 28820 21391
rect 28108 20560 28340 20600
rect 28779 20600 28821 20609
rect 28779 20560 28780 20600
rect 28820 20560 28821 20600
rect 27916 20096 27956 20105
rect 27243 18500 27285 18509
rect 27243 18460 27244 18500
rect 27284 18460 27285 18500
rect 27243 18451 27285 18460
rect 27244 18366 27284 18451
rect 27628 18425 27668 18456
rect 27916 18425 27956 20056
rect 28108 20096 28148 20560
rect 28779 20551 28821 20560
rect 29163 20264 29205 20273
rect 29163 20224 29164 20264
rect 29204 20224 29205 20264
rect 29163 20215 29205 20224
rect 28395 20180 28437 20189
rect 28395 20140 28396 20180
rect 28436 20140 28437 20180
rect 28395 20131 28437 20140
rect 28108 20047 28148 20056
rect 28300 20096 28340 20107
rect 28300 20021 28340 20056
rect 28396 20046 28436 20131
rect 28492 20096 28532 20105
rect 28299 20012 28341 20021
rect 28299 19972 28300 20012
rect 28340 19972 28341 20012
rect 28299 19963 28341 19972
rect 28012 19844 28052 19853
rect 28012 19265 28052 19804
rect 28011 19256 28053 19265
rect 28011 19216 28012 19256
rect 28052 19216 28053 19256
rect 28011 19207 28053 19216
rect 28300 18584 28340 18593
rect 28108 18544 28300 18584
rect 27627 18416 27669 18425
rect 27627 18376 27628 18416
rect 27668 18376 27669 18416
rect 27627 18367 27669 18376
rect 27915 18416 27957 18425
rect 27915 18376 27916 18416
rect 27956 18376 27957 18416
rect 27915 18367 27957 18376
rect 27051 18332 27093 18341
rect 27051 18292 27052 18332
rect 27092 18292 27093 18332
rect 27051 18283 27093 18292
rect 27628 18332 27668 18367
rect 27052 18198 27092 18283
rect 27628 17753 27668 18292
rect 28108 17996 28148 18544
rect 28300 18535 28340 18544
rect 28492 18509 28532 20056
rect 28875 19256 28917 19265
rect 28875 19216 28876 19256
rect 28916 19216 28917 19256
rect 28875 19207 28917 19216
rect 29164 19256 29204 20215
rect 32044 20180 32084 24583
rect 34060 24557 34100 24592
rect 34059 24548 34101 24557
rect 34059 24508 34060 24548
rect 34100 24508 34101 24548
rect 34059 24499 34101 24508
rect 34347 24548 34389 24557
rect 34347 24508 34348 24548
rect 34388 24508 34389 24548
rect 34347 24499 34389 24508
rect 33963 24380 34005 24389
rect 33963 24340 33964 24380
rect 34004 24340 34005 24380
rect 33963 24331 34005 24340
rect 33964 24246 34004 24331
rect 33352 24212 33720 24221
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33352 24163 33720 24172
rect 32811 23792 32853 23801
rect 32811 23752 32812 23792
rect 32852 23752 32853 23792
rect 32811 23743 32853 23752
rect 32620 23624 32660 23633
rect 32620 23129 32660 23584
rect 32619 23120 32661 23129
rect 32619 23080 32620 23120
rect 32660 23080 32661 23120
rect 32619 23071 32661 23080
rect 32812 21785 32852 23743
rect 34348 23288 34388 24499
rect 34444 23792 34484 25852
rect 34592 24968 34960 24977
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34592 24919 34960 24928
rect 36556 24641 36596 26095
rect 41643 26060 41685 26069
rect 41643 26020 41644 26060
rect 41684 26020 41685 26060
rect 41643 26011 41685 26020
rect 41644 25926 41684 26011
rect 35115 24632 35157 24641
rect 35115 24592 35116 24632
rect 35156 24592 35157 24632
rect 35115 24583 35157 24592
rect 36555 24632 36597 24641
rect 36555 24592 36556 24632
rect 36596 24592 36597 24632
rect 36555 24583 36597 24592
rect 35116 24498 35156 24583
rect 34924 24380 34964 24389
rect 35211 24380 35253 24389
rect 34964 24340 35156 24380
rect 34924 24331 34964 24340
rect 34828 23792 34868 23801
rect 34444 23752 34828 23792
rect 34828 23743 34868 23752
rect 34923 23792 34965 23801
rect 34923 23752 34924 23792
rect 34964 23752 34965 23792
rect 34923 23743 34965 23752
rect 35020 23792 35060 23801
rect 34924 23658 34964 23743
rect 34592 23456 34960 23465
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34592 23407 34960 23416
rect 34444 23288 34484 23297
rect 34348 23248 34444 23288
rect 34444 23239 34484 23248
rect 33771 23120 33813 23129
rect 33771 23080 33772 23120
rect 33812 23080 33813 23120
rect 33771 23071 33813 23080
rect 33772 22986 33812 23071
rect 34443 22868 34485 22877
rect 34443 22828 34444 22868
rect 34484 22828 34485 22868
rect 34443 22819 34485 22828
rect 34444 22734 34484 22819
rect 33352 22700 33720 22709
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33352 22651 33720 22660
rect 35020 22457 35060 23752
rect 33483 22448 33525 22457
rect 33483 22408 33484 22448
rect 33524 22408 33525 22448
rect 33483 22399 33525 22408
rect 34251 22448 34293 22457
rect 34251 22408 34252 22448
rect 34292 22408 34293 22448
rect 34251 22399 34293 22408
rect 35019 22448 35061 22457
rect 35019 22408 35020 22448
rect 35060 22408 35061 22448
rect 35019 22399 35061 22408
rect 33484 22364 33524 22399
rect 33484 22313 33524 22324
rect 34252 22314 34292 22399
rect 34924 22280 34964 22289
rect 35116 22280 35156 24340
rect 35211 24340 35212 24380
rect 35252 24340 35253 24380
rect 35211 24331 35253 24340
rect 35212 23792 35252 24331
rect 35212 23743 35252 23752
rect 35499 23792 35541 23801
rect 39916 23792 39956 23801
rect 35499 23752 35500 23792
rect 35540 23752 35541 23792
rect 35499 23743 35541 23752
rect 39244 23752 39916 23792
rect 35500 23658 35540 23743
rect 35692 23624 35732 23633
rect 35692 23213 35732 23584
rect 39244 23288 39284 23752
rect 39916 23743 39956 23752
rect 42028 23792 42068 26767
rect 42891 26648 42933 26657
rect 43564 26648 43604 26657
rect 42891 26608 42892 26648
rect 42932 26608 42933 26648
rect 42891 26599 42933 26608
rect 43372 26608 43564 26648
rect 42028 23743 42068 23752
rect 42892 23792 42932 26599
rect 43372 26069 43412 26608
rect 43564 26599 43604 26608
rect 43948 26312 43988 27691
rect 43948 26263 43988 26272
rect 44427 26144 44469 26153
rect 44427 26104 44428 26144
rect 44468 26104 44469 26144
rect 44427 26095 44469 26104
rect 43371 26060 43413 26069
rect 43371 26020 43372 26060
rect 43412 26020 43413 26060
rect 43371 26011 43413 26020
rect 43372 24632 43412 26011
rect 44428 26010 44468 26095
rect 45580 25304 45620 28279
rect 49712 27992 50080 28001
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 49712 27943 50080 27952
rect 64832 27992 65200 28001
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 64832 27943 65200 27952
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 95072 27992 95440 28001
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95072 27943 95440 27952
rect 48472 27236 48840 27245
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48472 27187 48840 27196
rect 63592 27236 63960 27245
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63592 27187 63960 27196
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 93832 27236 94200 27245
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 93832 27187 94200 27196
rect 49712 26480 50080 26489
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 49712 26431 50080 26440
rect 64832 26480 65200 26489
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 64832 26431 65200 26440
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 95072 26480 95440 26489
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95072 26431 95440 26440
rect 46155 26144 46197 26153
rect 46155 26104 46156 26144
rect 46196 26104 46197 26144
rect 46155 26095 46197 26104
rect 47020 26144 47060 26153
rect 47060 26104 47636 26144
rect 47020 26095 47060 26104
rect 45580 25229 45620 25264
rect 45196 25220 45236 25229
rect 45100 24800 45140 24809
rect 45196 24800 45236 25180
rect 45579 25220 45621 25229
rect 45579 25180 45580 25220
rect 45620 25180 45621 25220
rect 45579 25171 45621 25180
rect 45140 24760 45236 24800
rect 45100 24751 45140 24760
rect 43372 24583 43412 24592
rect 43564 24632 43604 24643
rect 43564 24557 43604 24592
rect 46156 24632 46196 26095
rect 46156 24583 46196 24592
rect 46348 25892 46388 25901
rect 46348 24557 46388 25852
rect 47596 25556 47636 26104
rect 48472 25724 48840 25733
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48472 25675 48840 25684
rect 63592 25724 63960 25733
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63592 25675 63960 25684
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 93832 25724 94200 25733
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 93832 25675 94200 25684
rect 47596 25507 47636 25516
rect 46443 25304 46485 25313
rect 46443 25264 46444 25304
rect 46484 25264 46485 25304
rect 46443 25255 46485 25264
rect 47787 25304 47829 25313
rect 47787 25264 47788 25304
rect 47828 25264 47829 25304
rect 47787 25255 47829 25264
rect 46444 25170 46484 25255
rect 46923 25220 46965 25229
rect 46923 25180 46924 25220
rect 46964 25180 46965 25220
rect 46923 25171 46965 25180
rect 46540 24632 46580 24641
rect 43563 24548 43605 24557
rect 43563 24508 43564 24548
rect 43604 24508 43605 24548
rect 43563 24499 43605 24508
rect 44907 24548 44949 24557
rect 44907 24508 44908 24548
rect 44948 24508 44949 24548
rect 44907 24499 44949 24508
rect 46347 24548 46389 24557
rect 46347 24508 46348 24548
rect 46388 24508 46389 24548
rect 46347 24499 46389 24508
rect 42892 23743 42932 23752
rect 43468 24380 43508 24389
rect 43468 23792 43508 24340
rect 44908 23960 44948 24499
rect 45964 24380 46004 24389
rect 44908 23920 45044 23960
rect 43852 23801 43892 23886
rect 43468 23743 43508 23752
rect 43851 23792 43893 23801
rect 43851 23752 43852 23792
rect 43892 23752 43893 23792
rect 43851 23743 43893 23752
rect 43276 23708 43316 23717
rect 43316 23668 43412 23708
rect 43276 23659 43316 23668
rect 39244 23239 39284 23248
rect 40588 23624 40628 23633
rect 35691 23204 35733 23213
rect 35691 23164 35692 23204
rect 35732 23164 35733 23204
rect 35691 23155 35733 23164
rect 36843 23204 36885 23213
rect 36843 23164 36844 23204
rect 36884 23164 36885 23204
rect 36843 23155 36885 23164
rect 40299 23204 40341 23213
rect 40299 23164 40300 23204
rect 40340 23164 40341 23204
rect 40299 23155 40341 23164
rect 36844 23070 36884 23155
rect 37228 23120 37268 23129
rect 35211 22868 35253 22877
rect 35211 22828 35212 22868
rect 35252 22828 35253 22868
rect 35211 22819 35253 22828
rect 34924 22121 34964 22240
rect 35020 22240 35156 22280
rect 35212 22280 35252 22819
rect 33292 22112 33332 22121
rect 32811 21776 32853 21785
rect 32811 21736 32812 21776
rect 32852 21736 32853 21776
rect 32811 21727 32853 21736
rect 32427 21692 32469 21701
rect 32427 21652 32428 21692
rect 32468 21652 32469 21692
rect 32427 21643 32469 21652
rect 32139 21608 32181 21617
rect 32139 21568 32140 21608
rect 32180 21568 32181 21608
rect 32139 21559 32181 21568
rect 32140 21474 32180 21559
rect 32428 21558 32468 21643
rect 32812 21608 32852 21727
rect 33292 21701 33332 22072
rect 34923 22112 34965 22121
rect 34923 22072 34924 22112
rect 34964 22072 34965 22112
rect 34923 22063 34965 22072
rect 34592 21944 34960 21953
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34592 21895 34960 21904
rect 34828 21776 34868 21787
rect 34828 21701 34868 21736
rect 33291 21692 33333 21701
rect 33291 21652 33292 21692
rect 33332 21652 33333 21692
rect 33291 21643 33333 21652
rect 34827 21692 34869 21701
rect 34827 21652 34828 21692
rect 34868 21652 34869 21692
rect 34827 21643 34869 21652
rect 35020 21617 35060 22240
rect 35212 22231 35252 22240
rect 35115 22112 35157 22121
rect 35115 22072 35116 22112
rect 35156 22072 35157 22112
rect 35115 22063 35157 22072
rect 35404 22112 35444 22121
rect 35444 22072 36308 22112
rect 35404 22063 35444 22072
rect 35116 21978 35156 22063
rect 36268 21692 36308 22072
rect 37228 21785 37268 23080
rect 38092 23120 38132 23129
rect 36651 21776 36693 21785
rect 36651 21736 36652 21776
rect 36692 21736 36693 21776
rect 36651 21727 36693 21736
rect 37227 21776 37269 21785
rect 37227 21736 37228 21776
rect 37268 21736 37269 21776
rect 37227 21727 37269 21736
rect 36268 21643 36308 21652
rect 32812 21559 32852 21568
rect 33676 21608 33716 21617
rect 35019 21608 35061 21617
rect 33716 21568 33812 21608
rect 33676 21559 33716 21568
rect 32427 21440 32469 21449
rect 32427 21400 32428 21440
rect 32468 21400 32469 21440
rect 32427 21391 32469 21400
rect 32044 20131 32084 20140
rect 31179 20096 31221 20105
rect 31179 20056 31180 20096
rect 31220 20056 31221 20096
rect 31179 20047 31221 20056
rect 32428 20096 32468 21391
rect 33352 21188 33720 21197
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33352 21139 33720 21148
rect 32428 20047 32468 20056
rect 31180 19962 31220 20047
rect 31467 19844 31509 19853
rect 31467 19804 31468 19844
rect 31508 19804 31509 19844
rect 31467 19795 31509 19804
rect 31660 19844 31700 19853
rect 29164 19207 29204 19216
rect 31468 19256 31508 19795
rect 28876 19122 28916 19207
rect 29355 19172 29397 19181
rect 29355 19132 29356 19172
rect 29396 19132 29397 19172
rect 29355 19123 29397 19132
rect 31083 19172 31125 19181
rect 31083 19132 31084 19172
rect 31124 19132 31125 19172
rect 31083 19123 31125 19132
rect 29356 19038 29396 19123
rect 31084 19038 31124 19123
rect 28491 18500 28533 18509
rect 28491 18460 28492 18500
rect 28532 18460 28533 18500
rect 28491 18451 28533 18460
rect 28492 18005 28532 18451
rect 28108 17947 28148 17956
rect 28491 17996 28533 18005
rect 28491 17956 28492 17996
rect 28532 17956 28533 17996
rect 28491 17947 28533 17956
rect 28971 17996 29013 18005
rect 28971 17956 28972 17996
rect 29012 17956 29013 17996
rect 28971 17947 29013 17956
rect 29163 17996 29205 18005
rect 29163 17956 29164 17996
rect 29204 17956 29205 17996
rect 29163 17947 29205 17956
rect 28972 17862 29012 17947
rect 27627 17744 27669 17753
rect 26667 17704 26668 17744
rect 26708 17704 26709 17744
rect 26667 17695 26709 17704
rect 26764 17704 26956 17744
rect 26996 17704 27476 17744
rect 26571 17660 26613 17669
rect 26571 17620 26572 17660
rect 26612 17620 26613 17660
rect 26571 17611 26613 17620
rect 26188 17107 26228 17116
rect 26572 17072 26612 17611
rect 26572 17023 26612 17032
rect 25227 16232 25269 16241
rect 25227 16192 25228 16232
rect 25268 16192 25269 16232
rect 25227 16183 25269 16192
rect 25707 16232 25749 16241
rect 25707 16192 25708 16232
rect 25748 16192 25749 16232
rect 25707 16183 25749 16192
rect 25323 15644 25365 15653
rect 25323 15604 25324 15644
rect 25364 15604 25365 15644
rect 25323 15595 25365 15604
rect 25324 15510 25364 15595
rect 25708 15569 25748 16183
rect 25707 15560 25749 15569
rect 25707 15520 25708 15560
rect 25748 15520 25749 15560
rect 25707 15511 25749 15520
rect 26572 15560 26612 15569
rect 26764 15560 26804 17704
rect 26956 17695 26996 17704
rect 27436 17072 27476 17704
rect 27627 17704 27628 17744
rect 27668 17704 27669 17744
rect 27627 17695 27669 17704
rect 28300 17744 28340 17753
rect 28340 17704 28628 17744
rect 28300 17695 28340 17704
rect 28588 17240 28628 17704
rect 29164 17576 29204 17947
rect 29259 17744 29301 17753
rect 29259 17704 29260 17744
rect 29300 17704 29301 17744
rect 29259 17695 29301 17704
rect 29260 17610 29300 17695
rect 29164 17527 29204 17536
rect 29452 17576 29492 17585
rect 28588 17191 28628 17200
rect 27436 17023 27476 17032
rect 27723 17072 27765 17081
rect 27723 17032 27724 17072
rect 27764 17032 27765 17072
rect 27723 17023 27765 17032
rect 27724 15728 27764 17023
rect 29452 16241 29492 17536
rect 29451 16232 29493 16241
rect 29451 16192 29452 16232
rect 29492 16192 29493 16232
rect 29451 16183 29493 16192
rect 31083 16232 31125 16241
rect 31083 16192 31084 16232
rect 31124 16192 31125 16232
rect 31083 16183 31125 16192
rect 31468 16232 31508 19216
rect 31468 16183 31508 16192
rect 31084 16098 31124 16183
rect 27724 15679 27764 15688
rect 26612 15520 26804 15560
rect 26859 15560 26901 15569
rect 26859 15520 26860 15560
rect 26900 15520 26901 15560
rect 26572 15511 26612 15520
rect 26859 15511 26901 15520
rect 25708 15426 25748 15511
rect 26860 14048 26900 15511
rect 31660 15140 31700 19804
rect 33099 19844 33141 19853
rect 33099 19804 33100 19844
rect 33140 19804 33141 19844
rect 33099 19795 33141 19804
rect 33100 19710 33140 19795
rect 33352 19676 33720 19685
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33352 19627 33720 19636
rect 33772 19517 33812 21568
rect 35019 21568 35020 21608
rect 35060 21568 35061 21608
rect 35019 21559 35061 21568
rect 36652 21608 36692 21727
rect 38092 21617 38132 23080
rect 40300 23070 40340 23155
rect 40492 23120 40532 23129
rect 40588 23120 40628 23584
rect 40876 23624 40916 23633
rect 43372 23624 43412 23668
rect 43948 23624 43988 23633
rect 43372 23584 43948 23624
rect 40532 23080 40628 23120
rect 40780 23120 40820 23129
rect 40876 23120 40916 23584
rect 43948 23575 43988 23584
rect 41067 23204 41109 23213
rect 41067 23164 41068 23204
rect 41108 23164 41109 23204
rect 41067 23155 41109 23164
rect 40820 23080 40916 23120
rect 40492 23071 40532 23080
rect 40780 23071 40820 23080
rect 41068 22280 41108 23155
rect 41068 22231 41108 22240
rect 45004 22280 45044 23920
rect 45675 23876 45717 23885
rect 45675 23836 45676 23876
rect 45716 23836 45717 23876
rect 45675 23827 45717 23836
rect 45484 23792 45524 23801
rect 45388 23752 45484 23792
rect 45388 22280 45428 23752
rect 45484 23743 45524 23752
rect 45579 23792 45621 23801
rect 45579 23752 45580 23792
rect 45620 23752 45621 23792
rect 45579 23743 45621 23752
rect 45676 23792 45716 23827
rect 45580 23658 45620 23743
rect 45676 23741 45716 23752
rect 45964 22289 46004 24340
rect 46348 24044 46388 24053
rect 46540 24044 46580 24592
rect 46924 24632 46964 25171
rect 47788 24641 47828 25255
rect 49712 24968 50080 24977
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 49712 24919 50080 24928
rect 64832 24968 65200 24977
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 64832 24919 65200 24928
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 95072 24968 95440 24977
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95072 24919 95440 24928
rect 46924 24583 46964 24592
rect 47787 24632 47829 24641
rect 47787 24592 47788 24632
rect 47828 24592 47829 24632
rect 47787 24583 47829 24592
rect 49611 24632 49653 24641
rect 49611 24592 49612 24632
rect 49652 24592 49653 24632
rect 49611 24583 49653 24592
rect 47788 24498 47828 24583
rect 48940 24380 48980 24389
rect 48472 24212 48840 24221
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48472 24163 48840 24172
rect 46388 24004 46580 24044
rect 46348 23995 46388 24004
rect 48940 23960 48980 24340
rect 48364 23920 48980 23960
rect 46155 23876 46197 23885
rect 46155 23836 46156 23876
rect 46196 23836 46197 23876
rect 46155 23827 46197 23836
rect 47691 23876 47733 23885
rect 47691 23836 47692 23876
rect 47732 23836 47733 23876
rect 47691 23827 47733 23836
rect 46156 23742 46196 23827
rect 47692 23742 47732 23827
rect 48364 23792 48404 23920
rect 48364 23743 48404 23752
rect 48472 22700 48840 22709
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48472 22651 48840 22660
rect 49612 22532 49652 24583
rect 63592 24212 63960 24221
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63592 24163 63960 24172
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 93832 24212 94200 24221
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 93832 24163 94200 24172
rect 49712 23456 50080 23465
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 49712 23407 50080 23416
rect 64832 23456 65200 23465
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 64832 23407 65200 23416
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 95072 23456 95440 23465
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95072 23407 95440 23416
rect 63592 22700 63960 22709
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63592 22651 63960 22660
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 93832 22700 94200 22709
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 93832 22651 94200 22660
rect 49612 22483 49652 22492
rect 45004 22231 45044 22240
rect 45100 22240 45428 22280
rect 45963 22280 46005 22289
rect 45963 22240 45964 22280
rect 46004 22240 46005 22280
rect 40396 22112 40436 22121
rect 44908 22112 44948 22121
rect 45100 22112 45140 22240
rect 45963 22231 46005 22240
rect 49323 22280 49365 22289
rect 49323 22240 49324 22280
rect 49364 22240 49365 22280
rect 49323 22231 49365 22240
rect 50284 22280 50324 22289
rect 40436 22072 40532 22112
rect 40396 22063 40436 22072
rect 36652 21559 36692 21568
rect 37515 21608 37557 21617
rect 37515 21568 37516 21608
rect 37556 21568 37557 21608
rect 37515 21559 37557 21568
rect 38091 21608 38133 21617
rect 38091 21568 38092 21608
rect 38132 21568 38133 21608
rect 38091 21559 38133 21568
rect 38956 21608 38996 21617
rect 34592 20432 34960 20441
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34592 20383 34960 20392
rect 33771 19508 33813 19517
rect 33771 19468 33772 19508
rect 33812 19468 33813 19508
rect 33771 19459 33813 19468
rect 32332 19256 32372 19265
rect 32332 19097 32372 19216
rect 33772 19097 33812 19459
rect 35020 19256 35060 21559
rect 37516 21474 37556 21559
rect 38668 21524 38708 21533
rect 38956 21524 38996 21568
rect 38708 21484 38996 21524
rect 38668 21475 38708 21484
rect 39628 21356 39668 21365
rect 39628 20777 39668 21316
rect 38955 20768 38997 20777
rect 38955 20728 38956 20768
rect 38996 20728 38997 20768
rect 38955 20719 38997 20728
rect 39627 20768 39669 20777
rect 39724 20768 39764 20777
rect 39627 20728 39628 20768
rect 39668 20728 39724 20768
rect 39627 20719 39669 20728
rect 39724 20719 39764 20728
rect 39819 20768 39861 20777
rect 39819 20728 39820 20768
rect 39860 20728 39861 20768
rect 39819 20719 39861 20728
rect 39916 20768 39956 20779
rect 38667 20096 38709 20105
rect 38667 20056 38668 20096
rect 38708 20056 38709 20096
rect 38667 20047 38709 20056
rect 38956 20096 38996 20719
rect 39051 20684 39093 20693
rect 39051 20644 39052 20684
rect 39092 20644 39093 20684
rect 39051 20635 39093 20644
rect 39052 20105 39092 20635
rect 39628 20634 39668 20719
rect 39820 20634 39860 20719
rect 39916 20693 39956 20728
rect 40395 20768 40437 20777
rect 40395 20728 40396 20768
rect 40436 20728 40437 20768
rect 40395 20719 40437 20728
rect 40492 20768 40532 22072
rect 44948 22072 45140 22112
rect 45196 22112 45236 22121
rect 44908 22063 44948 22072
rect 44811 21776 44853 21785
rect 44811 21736 44812 21776
rect 44852 21736 44853 21776
rect 44811 21727 44853 21736
rect 41835 21608 41877 21617
rect 41835 21568 41836 21608
rect 41876 21568 41877 21608
rect 41835 21559 41877 21568
rect 43083 21608 43125 21617
rect 43083 21568 43084 21608
rect 43124 21568 43125 21608
rect 43083 21559 43125 21568
rect 44043 21608 44085 21617
rect 44043 21568 44044 21608
rect 44084 21568 44085 21608
rect 44043 21559 44085 21568
rect 44428 21608 44468 21617
rect 44812 21608 44852 21727
rect 44468 21568 44756 21608
rect 44428 21559 44468 21568
rect 40492 20719 40532 20728
rect 39915 20684 39957 20693
rect 39915 20644 39916 20684
rect 39956 20644 39957 20684
rect 39915 20635 39957 20644
rect 40396 20634 40436 20719
rect 40684 20600 40724 20609
rect 40724 20560 40820 20600
rect 40684 20551 40724 20560
rect 39148 20180 39188 20189
rect 39188 20140 40148 20180
rect 39148 20131 39188 20140
rect 38956 20047 38996 20056
rect 39051 20096 39093 20105
rect 39051 20056 39052 20096
rect 39092 20056 39093 20096
rect 39051 20047 39093 20056
rect 40108 20096 40148 20140
rect 40108 20047 40148 20056
rect 40780 20096 40820 20560
rect 40780 20047 40820 20056
rect 38668 19962 38708 20047
rect 39436 19844 39476 19853
rect 35403 19508 35445 19517
rect 35403 19468 35404 19508
rect 35444 19468 35445 19508
rect 35403 19459 35445 19468
rect 35404 19374 35444 19459
rect 35020 19207 35060 19216
rect 35884 19256 35924 19265
rect 32331 19088 32373 19097
rect 32331 19048 32332 19088
rect 32372 19048 32373 19088
rect 32331 19039 32373 19048
rect 33484 19088 33524 19097
rect 32332 16232 32372 19039
rect 33484 18929 33524 19048
rect 33771 19088 33813 19097
rect 33771 19048 33772 19088
rect 33812 19048 33813 19088
rect 33771 19039 33813 19048
rect 35884 18929 35924 19216
rect 33483 18920 33525 18929
rect 33483 18880 33484 18920
rect 33524 18880 33525 18920
rect 33483 18871 33525 18880
rect 34059 18920 34101 18929
rect 34059 18880 34060 18920
rect 34100 18880 34101 18920
rect 34059 18871 34101 18880
rect 34592 18920 34960 18929
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34592 18871 34960 18880
rect 35883 18920 35925 18929
rect 35883 18880 35884 18920
rect 35924 18880 35925 18920
rect 35883 18871 35925 18880
rect 37515 18920 37557 18929
rect 37515 18880 37516 18920
rect 37556 18880 37557 18920
rect 37515 18871 37557 18880
rect 38187 18920 38229 18929
rect 38187 18880 38188 18920
rect 38228 18880 38229 18920
rect 38187 18871 38229 18880
rect 34060 18584 34100 18871
rect 34060 18535 34100 18544
rect 33388 18332 33428 18341
rect 33100 18292 33388 18332
rect 32715 17072 32757 17081
rect 32715 17032 32716 17072
rect 32756 17032 32757 17072
rect 32715 17023 32757 17032
rect 33100 17072 33140 18292
rect 33388 18283 33428 18292
rect 37036 18332 37076 18341
rect 33352 18164 33720 18173
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33352 18115 33720 18124
rect 37036 17753 37076 18292
rect 37035 17744 37077 17753
rect 37035 17704 37036 17744
rect 37076 17704 37077 17744
rect 37035 17695 37077 17704
rect 36651 17660 36693 17669
rect 36651 17620 36652 17660
rect 36692 17620 36693 17660
rect 36651 17611 36693 17620
rect 34592 17408 34960 17417
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34592 17359 34960 17368
rect 33196 17156 33236 17165
rect 33236 17116 33812 17156
rect 33196 17107 33236 17116
rect 33100 17023 33140 17032
rect 33772 17072 33812 17116
rect 33772 17023 33812 17032
rect 35404 17072 35444 17081
rect 32716 16938 32756 17023
rect 34444 16820 34484 16829
rect 34156 16780 34444 16820
rect 33352 16652 33720 16661
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33352 16603 33720 16612
rect 32332 16183 32372 16192
rect 34060 16232 34100 16241
rect 33484 16064 33524 16073
rect 33524 16024 33908 16064
rect 33484 16015 33524 16024
rect 33484 15688 33812 15728
rect 33484 15560 33524 15688
rect 33484 15511 33524 15520
rect 33579 15560 33621 15569
rect 33579 15520 33580 15560
rect 33620 15520 33621 15560
rect 33579 15511 33621 15520
rect 33676 15560 33716 15571
rect 33580 15426 33620 15511
rect 33676 15485 33716 15520
rect 33675 15476 33717 15485
rect 33675 15436 33676 15476
rect 33716 15436 33717 15476
rect 33675 15427 33717 15436
rect 31564 15100 31700 15140
rect 33352 15140 33720 15149
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 26860 13999 26900 14008
rect 27724 14048 27764 14057
rect 26092 13208 26132 13217
rect 24171 13040 24213 13049
rect 24171 13000 24172 13040
rect 24212 13000 24213 13040
rect 24171 12991 24213 13000
rect 24172 12906 24212 12991
rect 26092 12629 26132 13168
rect 26764 13040 26804 13049
rect 26764 12629 26804 13000
rect 26091 12620 26133 12629
rect 26091 12580 26092 12620
rect 26132 12580 26133 12620
rect 26091 12571 26133 12580
rect 26763 12620 26805 12629
rect 26763 12580 26764 12620
rect 26804 12580 26805 12620
rect 26763 12571 26805 12580
rect 23973 12536 24013 12544
rect 23884 12535 24013 12536
rect 23884 12496 23973 12535
rect 23973 12461 24013 12495
rect 24075 12536 24117 12545
rect 24172 12536 24212 12545
rect 24075 12496 24076 12536
rect 24116 12496 24172 12536
rect 24075 12487 24117 12496
rect 24172 12487 24212 12496
rect 24076 12402 24116 12487
rect 23595 12368 23637 12377
rect 23595 12328 23596 12368
rect 23636 12328 23637 12368
rect 23595 12319 23637 12328
rect 23979 12368 24021 12377
rect 23979 12328 23980 12368
rect 24020 12328 24021 12368
rect 23979 12319 24021 12328
rect 23980 12234 24020 12319
rect 27724 12293 27764 14008
rect 28299 12620 28341 12629
rect 28299 12580 28300 12620
rect 28340 12580 28341 12620
rect 28299 12571 28341 12580
rect 28300 12486 28340 12571
rect 28684 12536 28724 12545
rect 27723 12284 27765 12293
rect 27723 12244 27724 12284
rect 27764 12244 27765 12284
rect 27723 12235 27765 12244
rect 23691 11780 23733 11789
rect 23691 11740 23692 11780
rect 23732 11740 23733 11780
rect 23691 11731 23733 11740
rect 22635 11360 22677 11369
rect 22635 11320 22636 11360
rect 22676 11320 22677 11360
rect 22635 11311 22677 11320
rect 23404 10445 23444 11656
rect 23692 11646 23732 11731
rect 24171 11696 24213 11705
rect 24171 11656 24172 11696
rect 24212 11656 24213 11696
rect 24171 11647 24213 11656
rect 24172 11562 24212 11647
rect 24844 11528 24884 11537
rect 24460 11488 24844 11528
rect 24460 11108 24500 11488
rect 24844 11479 24884 11488
rect 28684 11369 28724 12496
rect 29548 12536 29588 12545
rect 29548 11705 29588 12496
rect 29931 12536 29973 12545
rect 29931 12496 29932 12536
rect 29972 12496 29973 12536
rect 29931 12487 29973 12496
rect 30699 12536 30741 12545
rect 30699 12496 30700 12536
rect 30740 12496 30741 12536
rect 30699 12487 30741 12496
rect 31180 12536 31220 12545
rect 29932 11864 29972 12487
rect 30700 12452 30740 12487
rect 30892 12452 30932 12461
rect 30700 12401 30740 12412
rect 30796 12412 30892 12452
rect 30027 11948 30069 11957
rect 30027 11908 30028 11948
rect 30068 11908 30069 11948
rect 30027 11899 30069 11908
rect 30315 11948 30357 11957
rect 30315 11908 30316 11948
rect 30356 11908 30357 11948
rect 30315 11899 30357 11908
rect 29932 11815 29972 11824
rect 29547 11696 29589 11705
rect 29547 11656 29548 11696
rect 29588 11656 29589 11696
rect 29547 11647 29589 11656
rect 29932 11696 29972 11705
rect 30028 11696 30068 11899
rect 30316 11814 30356 11899
rect 29972 11656 30068 11696
rect 29932 11647 29972 11656
rect 30124 11528 30164 11537
rect 24843 11360 24885 11369
rect 24843 11320 24844 11360
rect 24884 11320 24885 11360
rect 24843 11311 24885 11320
rect 28683 11360 28725 11369
rect 28683 11320 28684 11360
rect 28724 11320 28725 11360
rect 28683 11311 28725 11320
rect 24460 11059 24500 11068
rect 24844 11024 24884 11311
rect 30124 11201 30164 11488
rect 30123 11192 30165 11201
rect 30123 11152 30124 11192
rect 30164 11152 30165 11192
rect 30123 11143 30165 11152
rect 23403 10436 23445 10445
rect 23403 10396 23404 10436
rect 23444 10396 23445 10436
rect 23403 10387 23445 10396
rect 22060 10135 22100 10144
rect 21867 9512 21909 9521
rect 21867 9472 21868 9512
rect 21908 9472 21909 9512
rect 21867 9463 21909 9472
rect 21868 9378 21908 9463
rect 22540 9260 22580 9269
rect 21964 9220 22540 9260
rect 21964 8084 22004 9220
rect 22540 9211 22580 9220
rect 23499 8672 23541 8681
rect 23499 8632 23500 8672
rect 23540 8632 23541 8672
rect 23499 8623 23541 8632
rect 24459 8672 24501 8681
rect 24459 8632 24460 8672
rect 24500 8632 24501 8672
rect 24459 8623 24501 8632
rect 23500 8538 23540 8623
rect 24460 8538 24500 8623
rect 21964 8035 22004 8044
rect 23980 8504 24020 8513
rect 23980 8009 24020 8464
rect 22347 8000 22389 8009
rect 22347 7960 22348 8000
rect 22388 7960 22389 8000
rect 22347 7951 22389 7960
rect 23211 8000 23253 8009
rect 23211 7960 23212 8000
rect 23252 7960 23253 8000
rect 23211 7951 23253 7960
rect 23979 8000 24021 8009
rect 23979 7960 23980 8000
rect 24020 7960 24021 8000
rect 23979 7951 24021 7960
rect 24267 8000 24309 8009
rect 24267 7960 24268 8000
rect 24308 7960 24309 8000
rect 24267 7951 24309 7960
rect 22348 7866 22388 7951
rect 23212 7866 23252 7951
rect 23403 7916 23445 7925
rect 23403 7876 23404 7916
rect 23444 7876 23445 7916
rect 23403 7867 23445 7876
rect 23404 7757 23444 7867
rect 23403 7748 23445 7757
rect 23403 7708 23404 7748
rect 23444 7708 23445 7748
rect 23403 7699 23445 7708
rect 23404 7160 23444 7699
rect 23404 7111 23444 7120
rect 24268 7160 24308 7951
rect 24363 7916 24405 7925
rect 24363 7876 24364 7916
rect 24404 7876 24405 7916
rect 24363 7867 24405 7876
rect 24364 7782 24404 7867
rect 24844 7757 24884 10984
rect 25708 11024 25748 11033
rect 25708 8681 25748 10984
rect 26860 10772 26900 10781
rect 26860 10193 26900 10732
rect 27820 10312 28436 10352
rect 26859 10184 26901 10193
rect 26859 10144 26860 10184
rect 26900 10144 26901 10184
rect 26859 10135 26901 10144
rect 27820 10184 27860 10312
rect 27820 10135 27860 10144
rect 28011 10184 28053 10193
rect 28011 10144 28012 10184
rect 28052 10144 28053 10184
rect 28011 10135 28053 10144
rect 28203 10184 28245 10193
rect 28203 10144 28204 10184
rect 28244 10144 28245 10184
rect 28203 10135 28245 10144
rect 28396 10184 28436 10312
rect 27916 10016 27956 10025
rect 27916 8849 27956 9976
rect 27915 8840 27957 8849
rect 27915 8800 27916 8840
rect 27956 8800 27957 8840
rect 27915 8791 27957 8800
rect 25707 8672 25749 8681
rect 25707 8632 25708 8672
rect 25748 8632 25749 8672
rect 25707 8623 25749 8632
rect 25900 8672 25940 8681
rect 25324 8084 25364 8093
rect 24843 7748 24885 7757
rect 24843 7708 24844 7748
rect 24884 7708 24885 7748
rect 24843 7699 24885 7708
rect 23019 7076 23061 7085
rect 23019 7036 23020 7076
rect 23060 7036 23061 7076
rect 23019 7027 23061 7036
rect 23020 6942 23060 7027
rect 20620 5599 20660 5608
rect 21676 6280 21812 6320
rect 21676 3809 21716 6280
rect 24268 4145 24308 7120
rect 21771 4136 21813 4145
rect 21771 4096 21772 4136
rect 21812 4096 21813 4136
rect 21771 4087 21813 4096
rect 22923 4136 22965 4145
rect 22923 4096 22924 4136
rect 22964 4096 22965 4136
rect 22923 4087 22965 4096
rect 24172 4136 24212 4145
rect 21675 3800 21717 3809
rect 21675 3760 21676 3800
rect 21716 3760 21717 3800
rect 21675 3751 21717 3760
rect 19796 3424 19988 3464
rect 20619 3464 20661 3473
rect 20619 3424 20620 3464
rect 20660 3424 20661 3464
rect 19756 3415 19796 3424
rect 20619 3415 20661 3424
rect 20620 3330 20660 3415
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 18124 2876 18164 2885
rect 18164 2836 18740 2876
rect 18124 2827 18164 2836
rect 18028 2668 18164 2708
rect 18124 2624 18164 2668
rect 18220 2624 18260 2633
rect 17740 2611 18059 2624
rect 17740 2584 18019 2611
rect 17644 2575 17684 2584
rect 12268 2540 12308 2549
rect 652 2456 692 2465
rect 652 2297 692 2416
rect 651 2288 693 2297
rect 651 2248 652 2288
rect 692 2248 693 2288
rect 651 2239 693 2248
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 12268 2129 12308 2500
rect 12267 2120 12309 2129
rect 12267 2080 12268 2120
rect 12308 2080 12309 2120
rect 12267 2071 12309 2080
rect 13323 2120 13365 2129
rect 13323 2080 13324 2120
rect 13364 2080 13365 2120
rect 13323 2071 13365 2080
rect 13324 1986 13364 2071
rect 13516 1868 13556 1877
rect 13612 1868 13652 2575
rect 18124 2584 18220 2624
rect 18220 2575 18260 2584
rect 18700 2624 18740 2836
rect 18987 2792 19029 2801
rect 18987 2752 18988 2792
rect 19028 2752 19029 2792
rect 18987 2743 19029 2752
rect 18700 2575 18740 2584
rect 18988 2624 19028 2743
rect 19180 2633 19220 2635
rect 21676 2633 21716 3751
rect 21772 3632 21812 4087
rect 22924 4002 22964 4087
rect 23596 4052 23636 4061
rect 23788 4052 23828 4061
rect 23636 4012 23788 4052
rect 23596 4003 23636 4012
rect 23788 4003 23828 4012
rect 24172 3809 24212 4096
rect 24267 4136 24309 4145
rect 24267 4096 24268 4136
rect 24308 4096 24309 4136
rect 24267 4087 24309 4096
rect 25035 4136 25077 4145
rect 25035 4096 25036 4136
rect 25076 4096 25077 4136
rect 25035 4087 25077 4096
rect 25036 4002 25076 4087
rect 24171 3800 24213 3809
rect 24171 3760 24172 3800
rect 24212 3760 24213 3800
rect 24171 3751 24213 3760
rect 21772 3583 21812 3592
rect 22155 3464 22197 3473
rect 22155 3424 22156 3464
rect 22196 3424 22197 3464
rect 22155 3415 22197 3424
rect 18988 2575 19028 2584
rect 19179 2624 19221 2633
rect 19179 2584 19180 2624
rect 19220 2584 19221 2624
rect 19179 2575 19221 2584
rect 21291 2624 21333 2633
rect 21291 2584 21292 2624
rect 21332 2584 21333 2624
rect 21291 2575 21333 2584
rect 21675 2624 21717 2633
rect 21675 2584 21676 2624
rect 21716 2584 21717 2624
rect 21675 2575 21717 2584
rect 22156 2624 22196 3415
rect 23308 2708 23348 2717
rect 23348 2668 23828 2708
rect 23308 2659 23348 2668
rect 22156 2575 22196 2584
rect 23788 2624 23828 2668
rect 24172 2633 24212 3751
rect 25324 2717 25364 8044
rect 25420 8000 25460 8011
rect 25420 7925 25460 7960
rect 25804 8000 25844 8009
rect 25419 7916 25461 7925
rect 25419 7876 25420 7916
rect 25460 7876 25461 7916
rect 25419 7867 25461 7876
rect 25804 7748 25844 7960
rect 25900 7925 25940 8632
rect 26092 8672 26132 8681
rect 25995 8588 26037 8597
rect 25995 8548 25996 8588
rect 26036 8548 26037 8588
rect 25995 8539 26037 8548
rect 25996 8454 26036 8539
rect 25899 7916 25941 7925
rect 25899 7876 25900 7916
rect 25940 7876 25941 7916
rect 25899 7867 25941 7876
rect 26092 7748 26132 8632
rect 27244 8672 27284 8683
rect 27244 8597 27284 8632
rect 27339 8672 27381 8681
rect 27339 8632 27340 8672
rect 27380 8632 27381 8672
rect 27339 8623 27381 8632
rect 27819 8672 27861 8681
rect 27819 8632 27820 8672
rect 27860 8632 27861 8672
rect 27819 8623 27861 8632
rect 28012 8672 28052 10135
rect 28204 10050 28244 10135
rect 28299 10100 28341 10109
rect 28299 10060 28300 10100
rect 28340 10060 28341 10100
rect 28299 10051 28341 10060
rect 28300 9966 28340 10051
rect 28012 8623 28052 8632
rect 28300 8672 28340 8681
rect 28396 8672 28436 10144
rect 29739 10100 29781 10109
rect 29739 10060 29740 10100
rect 29780 10060 29781 10100
rect 29739 10051 29781 10060
rect 29643 8840 29685 8849
rect 29643 8800 29644 8840
rect 29684 8800 29685 8840
rect 29643 8791 29685 8800
rect 28340 8632 28436 8672
rect 29164 8672 29204 8681
rect 27243 8588 27285 8597
rect 27243 8548 27244 8588
rect 27284 8548 27285 8588
rect 27243 8539 27285 8548
rect 27340 8538 27380 8623
rect 27820 8588 27860 8623
rect 27820 8537 27860 8548
rect 25804 7708 26132 7748
rect 26956 8504 26996 8513
rect 25420 7412 25460 7421
rect 25804 7412 25844 7708
rect 25460 7372 25844 7412
rect 25420 7363 25460 7372
rect 26860 4976 26900 4985
rect 26860 4397 26900 4936
rect 26187 4388 26229 4397
rect 26187 4348 26188 4388
rect 26228 4348 26229 4388
rect 26187 4339 26229 4348
rect 26859 4388 26901 4397
rect 26859 4348 26860 4388
rect 26900 4348 26901 4388
rect 26859 4339 26901 4348
rect 26188 4254 26228 4339
rect 25899 4136 25941 4145
rect 25899 4096 25900 4136
rect 25940 4096 25941 4136
rect 25899 4087 25941 4096
rect 25323 2708 25365 2717
rect 25323 2668 25324 2708
rect 25364 2668 25365 2708
rect 25323 2659 25365 2668
rect 23788 2575 23828 2584
rect 24171 2624 24213 2633
rect 24171 2584 24172 2624
rect 24212 2584 24213 2624
rect 24171 2575 24213 2584
rect 25035 2624 25077 2633
rect 25035 2584 25036 2624
rect 25076 2584 25077 2624
rect 25035 2575 25077 2584
rect 25900 2624 25940 4087
rect 26956 3389 26996 8464
rect 28300 8177 28340 8632
rect 28492 8504 28532 8513
rect 27627 8168 27669 8177
rect 27627 8128 27628 8168
rect 27668 8128 27669 8168
rect 27627 8119 27669 8128
rect 28299 8168 28341 8177
rect 28299 8128 28300 8168
rect 28340 8128 28341 8168
rect 28299 8119 28341 8128
rect 27628 8034 27668 8119
rect 28492 7085 28532 8464
rect 29164 8261 29204 8632
rect 29547 8672 29589 8681
rect 29547 8632 29548 8672
rect 29588 8632 29589 8672
rect 29547 8623 29589 8632
rect 29644 8672 29684 8791
rect 29644 8623 29684 8632
rect 29740 8672 29780 10051
rect 29835 10016 29877 10025
rect 29835 9976 29836 10016
rect 29876 9976 29877 10016
rect 29835 9967 29877 9976
rect 29740 8623 29780 8632
rect 29836 8672 29876 9967
rect 29836 8623 29876 8632
rect 29548 8538 29588 8623
rect 29163 8252 29205 8261
rect 29163 8212 29164 8252
rect 29204 8212 29205 8252
rect 29163 8203 29205 8212
rect 30027 8084 30069 8093
rect 30027 8044 30028 8084
rect 30068 8044 30069 8084
rect 30027 8035 30069 8044
rect 28780 8000 28820 8009
rect 28491 7076 28533 7085
rect 28491 7036 28492 7076
rect 28532 7036 28533 7076
rect 28491 7027 28533 7036
rect 28780 6413 28820 7960
rect 29644 8000 29684 8009
rect 29644 7757 29684 7960
rect 30028 7950 30068 8035
rect 29643 7748 29685 7757
rect 29643 7708 29644 7748
rect 29684 7708 29685 7748
rect 29643 7699 29685 7708
rect 28779 6404 28821 6413
rect 28779 6364 28780 6404
rect 28820 6364 28821 6404
rect 28779 6355 28821 6364
rect 28971 6320 29013 6329
rect 28971 6280 28972 6320
rect 29012 6280 29013 6320
rect 28971 6271 29013 6280
rect 27532 4976 27572 4985
rect 27724 4976 27764 4985
rect 27572 4936 27724 4976
rect 27532 4927 27572 4936
rect 27724 4927 27764 4936
rect 28107 4976 28149 4985
rect 28107 4936 28108 4976
rect 28148 4936 28149 4976
rect 28107 4927 28149 4936
rect 28587 4976 28629 4985
rect 28587 4936 28588 4976
rect 28628 4936 28629 4976
rect 28587 4927 28629 4936
rect 28972 4976 29012 6271
rect 28108 4842 28148 4927
rect 26955 3380 26997 3389
rect 26955 3340 26956 3380
rect 26996 3340 26997 3380
rect 26955 3331 26997 3340
rect 27052 2708 27092 2717
rect 27092 2668 27380 2708
rect 27052 2659 27092 2668
rect 25900 2575 25940 2584
rect 27340 2624 27380 2668
rect 28588 2633 28628 4927
rect 27340 2575 27380 2584
rect 28587 2624 28629 2633
rect 28587 2584 28588 2624
rect 28628 2584 28629 2624
rect 28972 2624 29012 4936
rect 30220 5648 30260 5657
rect 30124 4892 30164 4901
rect 30220 4892 30260 5608
rect 30164 4852 30260 4892
rect 30124 4843 30164 4852
rect 30796 4313 30836 12412
rect 30892 12403 30932 12412
rect 31180 11276 31220 12496
rect 31276 12536 31316 12547
rect 31276 12461 31316 12496
rect 31275 12452 31317 12461
rect 31275 12412 31276 12452
rect 31316 12412 31317 12452
rect 31275 12403 31317 12412
rect 31467 11696 31509 11705
rect 31467 11656 31468 11696
rect 31508 11656 31509 11696
rect 31467 11647 31509 11656
rect 31468 11562 31508 11647
rect 31180 11236 31316 11276
rect 31179 11108 31221 11117
rect 31179 11068 31180 11108
rect 31220 11068 31221 11108
rect 31179 11059 31221 11068
rect 31180 11024 31220 11059
rect 31180 10973 31220 10984
rect 31276 10989 31316 11236
rect 31371 11192 31413 11201
rect 31371 11152 31372 11192
rect 31412 11152 31413 11192
rect 31371 11143 31413 11152
rect 31372 11024 31412 11143
rect 31564 11033 31604 15100
rect 33352 15091 33720 15100
rect 33676 14720 33716 14729
rect 33772 14720 33812 15688
rect 33868 15560 33908 16024
rect 34060 15569 34100 16192
rect 34156 16232 34196 16780
rect 34444 16771 34484 16780
rect 35404 16409 35444 17032
rect 36076 17072 36116 17081
rect 36268 17072 36308 17081
rect 36116 17032 36268 17072
rect 36076 17023 36116 17032
rect 36268 17023 36308 17032
rect 36652 17072 36692 17611
rect 34347 16400 34389 16409
rect 34347 16360 34348 16400
rect 34388 16360 34389 16400
rect 34347 16351 34389 16360
rect 35403 16400 35445 16409
rect 35403 16360 35404 16400
rect 35444 16360 35445 16400
rect 35403 16351 35445 16360
rect 34348 16316 34388 16351
rect 34348 16265 34388 16276
rect 34156 16183 34196 16192
rect 34592 15896 34960 15905
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34592 15847 34960 15856
rect 33868 15511 33908 15520
rect 34059 15560 34101 15569
rect 34059 15520 34060 15560
rect 34100 15520 34101 15560
rect 34059 15511 34101 15520
rect 34539 15476 34581 15485
rect 34539 15436 34540 15476
rect 34580 15436 34581 15476
rect 34539 15427 34581 15436
rect 34059 15392 34101 15401
rect 34059 15352 34060 15392
rect 34100 15352 34101 15392
rect 34059 15343 34101 15352
rect 33716 14680 33812 14720
rect 34060 14720 34100 15343
rect 34540 15342 34580 15427
rect 36652 15140 36692 17032
rect 37516 17072 37556 18871
rect 38188 18584 38228 18871
rect 39436 18668 39476 19804
rect 41452 19844 41492 19853
rect 41452 18677 41492 19804
rect 39436 18619 39476 18628
rect 41451 18668 41493 18677
rect 41451 18628 41452 18668
rect 41492 18628 41493 18668
rect 41451 18619 41493 18628
rect 38188 18535 38228 18544
rect 39052 18584 39092 18593
rect 39052 17753 39092 18544
rect 41836 18584 41876 21559
rect 43084 21474 43124 21559
rect 44044 21474 44084 21559
rect 43755 21440 43797 21449
rect 43755 21400 43756 21440
rect 43796 21400 43797 21440
rect 43755 21391 43797 21400
rect 43756 21306 43796 21391
rect 44427 20600 44469 20609
rect 44427 20560 44428 20600
rect 44468 20560 44469 20600
rect 44427 20551 44469 20560
rect 44428 20466 44468 20551
rect 44716 19928 44756 21568
rect 44812 21559 44852 21568
rect 45004 20189 45044 22072
rect 45196 20777 45236 22072
rect 45964 21617 46004 22231
rect 49324 22146 49364 22231
rect 49712 21944 50080 21953
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 49712 21895 50080 21904
rect 46443 21776 46485 21785
rect 46443 21736 46444 21776
rect 46484 21736 46485 21776
rect 46443 21727 46485 21736
rect 45676 21608 45716 21617
rect 45580 21568 45676 21608
rect 45580 21449 45620 21568
rect 45676 21559 45716 21568
rect 45963 21608 46005 21617
rect 45963 21568 45964 21608
rect 46004 21568 46005 21608
rect 45963 21559 46005 21568
rect 45579 21440 45621 21449
rect 45579 21400 45580 21440
rect 45620 21400 45621 21440
rect 45579 21391 45621 21400
rect 45195 20768 45237 20777
rect 45195 20728 45196 20768
rect 45236 20728 45237 20768
rect 45195 20719 45237 20728
rect 45580 20768 45620 21391
rect 45580 20719 45620 20728
rect 46444 20768 46484 21727
rect 46828 21356 46868 21365
rect 45003 20180 45045 20189
rect 45003 20140 45004 20180
rect 45044 20140 45045 20180
rect 45003 20131 45045 20140
rect 46059 20180 46101 20189
rect 46059 20140 46060 20180
rect 46100 20140 46101 20180
rect 46059 20131 46101 20140
rect 45004 20012 45044 20131
rect 46060 20046 46100 20131
rect 45004 19963 45044 19972
rect 44812 19928 44852 19937
rect 44716 19888 44812 19928
rect 44812 19879 44852 19888
rect 43563 19844 43605 19853
rect 43563 19804 43564 19844
rect 43604 19804 43605 19844
rect 43563 19795 43605 19804
rect 43083 18668 43125 18677
rect 43083 18628 43084 18668
rect 43124 18628 43125 18668
rect 43083 18619 43125 18628
rect 41836 18535 41876 18544
rect 42700 18584 42740 18593
rect 40684 18332 40724 18341
rect 37899 17744 37941 17753
rect 37899 17704 37900 17744
rect 37940 17704 37941 17744
rect 37899 17695 37941 17704
rect 39051 17744 39093 17753
rect 39051 17704 39052 17744
rect 39092 17704 39093 17744
rect 39051 17695 39093 17704
rect 37900 17610 37940 17695
rect 37516 17023 37556 17032
rect 38572 17576 38612 17585
rect 38572 15485 38612 17536
rect 40396 17072 40436 17083
rect 40396 16997 40436 17032
rect 40684 17072 40724 18292
rect 42700 17753 42740 18544
rect 43084 18534 43124 18619
rect 43564 17753 43604 19795
rect 46444 18509 46484 20728
rect 46732 21316 46828 21356
rect 46732 20096 46772 21316
rect 46828 21307 46868 21316
rect 48472 21188 48840 21197
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48472 21139 48840 21148
rect 46827 20768 46869 20777
rect 46827 20728 46828 20768
rect 46868 20728 46869 20768
rect 46827 20719 46869 20728
rect 46828 20634 46868 20719
rect 49712 20432 50080 20441
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 49712 20383 50080 20392
rect 50284 20105 50324 22240
rect 64832 21944 65200 21953
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 64832 21895 65200 21904
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 95072 21944 95440 21953
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95072 21895 95440 21904
rect 63592 21188 63960 21197
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63592 21139 63960 21148
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 93832 21188 94200 21197
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 93832 21139 94200 21148
rect 52684 20852 52724 20861
rect 52492 20600 52532 20609
rect 52108 20560 52492 20600
rect 52108 20180 52148 20560
rect 52492 20551 52532 20560
rect 52108 20131 52148 20140
rect 50283 20096 50325 20105
rect 46732 20047 46772 20056
rect 50188 20056 50284 20096
rect 50324 20056 50325 20096
rect 48472 19676 48840 19685
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48472 19627 48840 19636
rect 49712 18920 50080 18929
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 49712 18871 50080 18880
rect 48747 18584 48789 18593
rect 48747 18544 48748 18584
rect 48788 18544 48789 18584
rect 48747 18535 48789 18544
rect 49132 18584 49172 18595
rect 46443 18500 46485 18509
rect 46443 18460 46444 18500
rect 46484 18460 46485 18500
rect 46443 18451 46485 18460
rect 42219 17744 42261 17753
rect 42219 17704 42220 17744
rect 42260 17704 42261 17744
rect 42219 17695 42261 17704
rect 42699 17744 42741 17753
rect 42699 17704 42700 17744
rect 42740 17704 42741 17744
rect 42699 17695 42741 17704
rect 43563 17744 43605 17753
rect 43563 17704 43564 17744
rect 43604 17704 43605 17744
rect 43563 17695 43605 17704
rect 45099 17744 45141 17753
rect 45099 17704 45100 17744
rect 45140 17704 45141 17744
rect 45099 17695 45141 17704
rect 40684 17023 40724 17032
rect 40876 17156 40916 17165
rect 38667 16988 38709 16997
rect 38667 16948 38668 16988
rect 38708 16948 38709 16988
rect 38667 16939 38709 16948
rect 40395 16988 40437 16997
rect 40395 16948 40396 16988
rect 40436 16948 40437 16988
rect 40395 16939 40437 16948
rect 38668 16854 38708 16939
rect 39340 15728 39380 15737
rect 39380 15688 39764 15728
rect 39340 15679 39380 15688
rect 38668 15560 38708 15569
rect 38571 15476 38613 15485
rect 38571 15436 38572 15476
rect 38612 15436 38613 15476
rect 38571 15427 38613 15436
rect 38668 15140 38708 15520
rect 39532 15560 39572 15571
rect 39532 15485 39572 15520
rect 39627 15560 39669 15569
rect 39627 15520 39628 15560
rect 39668 15520 39669 15560
rect 39627 15511 39669 15520
rect 39724 15560 39764 15688
rect 39724 15511 39764 15520
rect 40683 15560 40725 15569
rect 40683 15520 40684 15560
rect 40724 15520 40725 15560
rect 40683 15511 40725 15520
rect 40780 15560 40820 15569
rect 40876 15560 40916 17116
rect 41452 16232 41492 16241
rect 40972 16192 41452 16232
rect 40972 15728 41012 16192
rect 41452 16183 41492 16192
rect 42124 16064 42164 16073
rect 40972 15679 41012 15688
rect 41740 16024 42124 16064
rect 41740 15644 41780 16024
rect 42124 16015 42164 16024
rect 41740 15595 41780 15604
rect 40820 15520 40916 15560
rect 42124 15560 42164 15569
rect 42220 15560 42260 17695
rect 42700 17610 42740 17695
rect 43564 17610 43604 17695
rect 45100 17072 45140 17695
rect 45100 17023 45140 17032
rect 46059 17072 46101 17081
rect 46059 17032 46060 17072
rect 46100 17032 46101 17072
rect 46059 17023 46101 17032
rect 45964 16232 46004 16241
rect 46060 16232 46100 17023
rect 46444 16400 46484 18451
rect 48748 18450 48788 18535
rect 49132 18509 49172 18544
rect 49323 18584 49365 18593
rect 49323 18544 49324 18584
rect 49364 18544 49365 18584
rect 49323 18535 49365 18544
rect 49996 18584 50036 18593
rect 50188 18584 50228 20056
rect 50283 20047 50325 20056
rect 52492 20096 52532 20105
rect 52492 19265 52532 20056
rect 52491 19256 52533 19265
rect 52491 19216 52492 19256
rect 52532 19216 52533 19256
rect 52491 19207 52533 19216
rect 52492 19013 52532 19207
rect 52491 19004 52533 19013
rect 52491 18964 52492 19004
rect 52532 18964 52533 19004
rect 52491 18955 52533 18964
rect 52684 18929 52724 20812
rect 64832 20432 65200 20441
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 64832 20383 65200 20392
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 95072 20432 95440 20441
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95072 20383 95440 20392
rect 53355 20096 53397 20105
rect 53355 20056 53356 20096
rect 53396 20056 53397 20096
rect 53355 20047 53397 20056
rect 56907 20096 56949 20105
rect 56907 20056 56908 20096
rect 56948 20056 56949 20096
rect 56907 20047 56949 20056
rect 57484 20096 57524 20105
rect 53356 19962 53396 20047
rect 54508 19844 54548 19853
rect 54220 19804 54508 19844
rect 54220 19256 54260 19804
rect 54508 19795 54548 19804
rect 56812 19844 56852 19853
rect 56812 19349 56852 19804
rect 55275 19340 55317 19349
rect 56811 19340 56853 19349
rect 55275 19300 55276 19340
rect 55316 19300 55412 19340
rect 55275 19291 55317 19300
rect 54220 19207 54260 19216
rect 55276 19206 55316 19291
rect 53548 19088 53588 19097
rect 53548 18929 53588 19048
rect 50283 18920 50325 18929
rect 50283 18880 50284 18920
rect 50324 18880 50325 18920
rect 50283 18871 50325 18880
rect 52395 18920 52437 18929
rect 52395 18880 52396 18920
rect 52436 18880 52437 18920
rect 52395 18871 52437 18880
rect 52683 18920 52725 18929
rect 52683 18880 52684 18920
rect 52724 18880 52725 18920
rect 52683 18871 52725 18880
rect 53547 18920 53589 18929
rect 53547 18880 53548 18920
rect 53588 18880 53589 18920
rect 53547 18871 53589 18880
rect 55179 18920 55221 18929
rect 55179 18880 55180 18920
rect 55220 18880 55221 18920
rect 55179 18871 55221 18880
rect 50036 18544 50228 18584
rect 49996 18535 50036 18544
rect 49131 18500 49173 18509
rect 49131 18460 49132 18500
rect 49172 18460 49173 18500
rect 49131 18451 49173 18460
rect 48472 18164 48840 18173
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48472 18115 48840 18124
rect 49324 17996 49364 18535
rect 50284 18509 50324 18871
rect 51340 18584 51380 18593
rect 50283 18500 50325 18509
rect 50283 18460 50284 18500
rect 50324 18460 50325 18500
rect 50283 18451 50325 18460
rect 51148 18500 51188 18509
rect 51340 18500 51380 18544
rect 51188 18460 51380 18500
rect 51148 18451 51188 18460
rect 49324 17947 49364 17956
rect 47787 17912 47829 17921
rect 47787 17872 47788 17912
rect 47828 17872 47829 17912
rect 47787 17863 47829 17872
rect 48843 17912 48885 17921
rect 48843 17872 48844 17912
rect 48884 17872 48885 17912
rect 48843 17863 48885 17872
rect 47788 17156 47828 17863
rect 48844 17778 48884 17863
rect 49036 17828 49076 17839
rect 49036 17753 49076 17788
rect 49515 17828 49557 17837
rect 49515 17788 49516 17828
rect 49556 17788 49557 17828
rect 49515 17779 49557 17788
rect 49035 17744 49077 17753
rect 49035 17704 49036 17744
rect 49076 17704 49077 17744
rect 49035 17695 49077 17704
rect 49516 17694 49556 17779
rect 49707 17744 49749 17753
rect 49707 17704 49708 17744
rect 49748 17704 49749 17744
rect 49707 17695 49749 17704
rect 49708 17610 49748 17695
rect 49712 17408 50080 17417
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 49712 17359 50080 17368
rect 50187 17324 50229 17333
rect 50187 17284 50188 17324
rect 50228 17284 50229 17324
rect 50187 17275 50229 17284
rect 50188 17240 50228 17275
rect 50188 17189 50228 17200
rect 47788 17107 47828 17116
rect 48171 17072 48213 17081
rect 48171 17032 48172 17072
rect 48212 17032 48213 17072
rect 48171 17023 48213 17032
rect 49036 17072 49076 17081
rect 48172 16938 48212 17023
rect 48472 16652 48840 16661
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48472 16603 48840 16612
rect 46540 16400 46580 16409
rect 46444 16360 46540 16400
rect 46540 16351 46580 16360
rect 46004 16192 46100 16232
rect 45964 16183 46004 16192
rect 46348 16064 46388 16073
rect 42164 15520 42260 15560
rect 42988 15560 43028 15569
rect 40780 15511 40820 15520
rect 38763 15476 38805 15485
rect 38763 15436 38764 15476
rect 38804 15436 38805 15476
rect 38763 15427 38805 15436
rect 39531 15476 39573 15485
rect 39531 15436 39532 15476
rect 39572 15436 39573 15476
rect 39531 15427 39573 15436
rect 36652 15100 36788 15140
rect 36748 14729 36788 15100
rect 38284 15100 38708 15140
rect 37804 14804 37844 14813
rect 38284 14804 38324 15100
rect 37844 14764 38324 14804
rect 37804 14755 37844 14764
rect 34540 14720 34580 14729
rect 33676 14561 33716 14680
rect 34060 14671 34100 14680
rect 34156 14680 34540 14720
rect 34156 14636 34196 14680
rect 34540 14671 34580 14680
rect 35787 14720 35829 14729
rect 35787 14680 35788 14720
rect 35828 14680 35829 14720
rect 35787 14671 35829 14680
rect 36652 14720 36692 14729
rect 34156 14587 34196 14596
rect 35212 14636 35252 14645
rect 35404 14636 35444 14645
rect 35252 14596 35404 14636
rect 35212 14587 35252 14596
rect 35404 14587 35444 14596
rect 35788 14586 35828 14671
rect 33675 14552 33717 14561
rect 33675 14512 33676 14552
rect 33716 14512 33717 14552
rect 33675 14503 33717 14512
rect 34592 14384 34960 14393
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34592 14335 34960 14344
rect 33352 13628 33720 13637
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33352 13579 33720 13588
rect 34592 12872 34960 12881
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34592 12823 34960 12832
rect 31660 12704 31700 12713
rect 31660 11957 31700 12664
rect 31755 12536 31797 12545
rect 31755 12496 31756 12536
rect 31796 12496 31797 12536
rect 31755 12487 31797 12496
rect 35883 12536 35925 12545
rect 35883 12496 35884 12536
rect 35924 12496 35925 12536
rect 35883 12487 35925 12496
rect 31756 12402 31796 12487
rect 32235 12452 32277 12461
rect 32235 12412 32236 12452
rect 32276 12412 32277 12452
rect 32235 12403 32277 12412
rect 31948 12284 31988 12293
rect 31659 11948 31701 11957
rect 31659 11908 31660 11948
rect 31700 11908 31701 11948
rect 31659 11899 31701 11908
rect 31948 11117 31988 12244
rect 32043 11192 32085 11201
rect 32043 11152 32044 11192
rect 32084 11152 32085 11192
rect 32043 11143 32085 11152
rect 32236 11192 32276 12403
rect 35884 12402 35924 12487
rect 36652 12293 36692 14680
rect 36747 14720 36789 14729
rect 36747 14680 36748 14720
rect 36788 14680 36789 14720
rect 36747 14671 36789 14680
rect 38284 14720 38324 14764
rect 38284 14671 38324 14680
rect 38668 14720 38708 14729
rect 38764 14720 38804 15427
rect 39628 15426 39668 15511
rect 40684 15426 40724 15511
rect 42124 15140 42164 15520
rect 42124 15100 42260 15140
rect 38708 14680 38804 14720
rect 38668 14671 38708 14680
rect 36748 13217 36788 14671
rect 38764 14552 38804 14561
rect 38764 14057 38804 14512
rect 38763 14048 38805 14057
rect 38763 14008 38764 14048
rect 38804 14008 38805 14048
rect 38763 13999 38805 14008
rect 39147 14048 39189 14057
rect 39147 14008 39148 14048
rect 39188 14008 39189 14048
rect 39147 13999 39189 14008
rect 39148 13914 39188 13999
rect 38476 13796 38516 13805
rect 36747 13208 36789 13217
rect 36747 13168 36748 13208
rect 36788 13168 36789 13208
rect 36747 13159 36789 13168
rect 36939 13208 36981 13217
rect 36939 13168 36940 13208
rect 36980 13168 36981 13208
rect 36939 13159 36981 13168
rect 38476 13208 38516 13756
rect 38476 13159 38516 13168
rect 38859 13208 38901 13217
rect 38859 13168 38860 13208
rect 38900 13168 38901 13208
rect 38859 13159 38901 13168
rect 39723 13208 39765 13217
rect 39723 13168 39724 13208
rect 39764 13168 39765 13208
rect 39723 13159 39765 13168
rect 41163 13208 41205 13217
rect 41163 13168 41164 13208
rect 41204 13168 41205 13208
rect 41163 13159 41205 13168
rect 41644 13208 41684 13217
rect 35211 12284 35253 12293
rect 35211 12244 35212 12284
rect 35252 12244 35253 12284
rect 35211 12235 35253 12244
rect 36651 12284 36693 12293
rect 36651 12244 36652 12284
rect 36692 12244 36693 12284
rect 36651 12235 36693 12244
rect 33352 12116 33720 12125
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33352 12067 33720 12076
rect 35212 11705 35252 12235
rect 32332 11696 32372 11705
rect 32332 11369 32372 11656
rect 35211 11696 35253 11705
rect 35211 11656 35212 11696
rect 35252 11656 35253 11696
rect 35211 11647 35253 11656
rect 32715 11612 32757 11621
rect 32715 11572 32716 11612
rect 32756 11572 32757 11612
rect 32715 11563 32757 11572
rect 33099 11612 33141 11621
rect 33099 11572 33100 11612
rect 33140 11572 33141 11612
rect 33099 11563 33141 11572
rect 32716 11478 32756 11563
rect 32331 11360 32373 11369
rect 32331 11320 32332 11360
rect 32372 11320 32373 11360
rect 32331 11311 32373 11320
rect 32236 11143 32276 11152
rect 33100 11192 33140 11563
rect 34592 11360 34960 11369
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34592 11311 34960 11320
rect 33100 11143 33140 11152
rect 31947 11108 31989 11117
rect 31947 11068 31948 11108
rect 31988 11068 31989 11108
rect 31947 11059 31989 11068
rect 31372 10975 31412 10984
rect 31563 11024 31605 11033
rect 31563 10984 31564 11024
rect 31604 10984 31605 11024
rect 31563 10975 31605 10984
rect 31948 11024 31988 11059
rect 31948 10974 31988 10984
rect 32044 11024 32084 11143
rect 33772 11024 33812 11033
rect 32044 10975 32084 10984
rect 33004 10984 33772 11024
rect 30891 10772 30933 10781
rect 30891 10732 30892 10772
rect 30932 10732 30933 10772
rect 30891 10723 30933 10732
rect 30892 10638 30932 10723
rect 31276 10025 31316 10949
rect 31275 10016 31317 10025
rect 31275 9976 31276 10016
rect 31316 9976 31317 10016
rect 31275 9967 31317 9976
rect 33004 9680 33044 10984
rect 33772 10975 33812 10984
rect 35884 10772 35924 10781
rect 33352 10604 33720 10613
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33352 10555 33720 10564
rect 34592 9848 34960 9857
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34592 9799 34960 9808
rect 33004 9631 33044 9640
rect 33100 9724 33524 9764
rect 33100 9512 33140 9724
rect 33484 9680 33524 9724
rect 33484 9631 33524 9640
rect 33196 9521 33236 9606
rect 33100 9463 33140 9472
rect 33195 9512 33237 9521
rect 33195 9472 33196 9512
rect 33236 9472 33237 9512
rect 33195 9463 33237 9472
rect 33292 9512 33332 9521
rect 33292 9260 33332 9472
rect 33100 9220 33332 9260
rect 34156 9512 34196 9521
rect 32332 8672 32372 8681
rect 31660 8504 31700 8513
rect 31660 8093 31700 8464
rect 32332 8177 32372 8632
rect 33100 8336 33140 9220
rect 33352 9092 33720 9101
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33352 9043 33720 9052
rect 34156 8849 34196 9472
rect 34443 9512 34485 9521
rect 34443 9472 34444 9512
rect 34484 9472 34485 9512
rect 34443 9463 34485 9472
rect 33291 8840 33333 8849
rect 33291 8800 33292 8840
rect 33332 8800 33333 8840
rect 33291 8791 33333 8800
rect 34155 8840 34197 8849
rect 34155 8800 34156 8840
rect 34196 8800 34197 8840
rect 34155 8791 34197 8800
rect 33292 8706 33332 8791
rect 34444 8756 34484 9463
rect 34444 8707 34484 8716
rect 35692 9260 35732 9269
rect 33196 8672 33236 8683
rect 33196 8597 33236 8632
rect 33387 8672 33429 8681
rect 33387 8632 33388 8672
rect 33428 8632 33429 8672
rect 33387 8623 33429 8632
rect 33868 8672 33908 8683
rect 33195 8588 33237 8597
rect 33195 8548 33196 8588
rect 33236 8548 33237 8588
rect 33195 8539 33237 8548
rect 33388 8538 33428 8623
rect 33868 8597 33908 8632
rect 34155 8672 34197 8681
rect 34348 8672 34388 8700
rect 34155 8632 34156 8672
rect 34196 8632 34348 8672
rect 34155 8623 34197 8632
rect 33867 8588 33909 8597
rect 33867 8548 33868 8588
rect 33908 8548 33909 8588
rect 33867 8539 33909 8548
rect 34156 8538 34196 8623
rect 33676 8504 33716 8513
rect 33484 8464 33676 8504
rect 33100 8296 33428 8336
rect 32331 8168 32373 8177
rect 32331 8128 32332 8168
rect 32372 8128 32373 8168
rect 32331 8119 32373 8128
rect 33099 8168 33141 8177
rect 33099 8128 33100 8168
rect 33140 8128 33141 8168
rect 33099 8119 33141 8128
rect 31659 8084 31701 8093
rect 31659 8044 31660 8084
rect 31700 8044 31701 8084
rect 31659 8035 31701 8044
rect 33100 8034 33140 8119
rect 33196 7412 33236 8296
rect 33388 8000 33428 8296
rect 33388 7951 33428 7960
rect 33484 8000 33524 8464
rect 33676 8455 33716 8464
rect 33963 8252 34005 8261
rect 33963 8212 33964 8252
rect 34004 8212 34005 8252
rect 33963 8203 34005 8212
rect 33964 8168 34004 8203
rect 33964 8117 34004 8128
rect 33484 7951 33524 7960
rect 33771 8000 33813 8009
rect 33771 7960 33772 8000
rect 33812 7960 33813 8000
rect 33771 7951 33813 7960
rect 34059 8000 34101 8009
rect 34059 7960 34060 8000
rect 34100 7960 34101 8000
rect 34059 7951 34101 7960
rect 33352 7580 33720 7589
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33352 7531 33720 7540
rect 33292 7412 33332 7421
rect 33772 7412 33812 7951
rect 34060 7866 34100 7951
rect 33196 7372 33292 7412
rect 33292 7363 33332 7372
rect 33388 7372 33812 7412
rect 34252 7412 34292 8632
rect 34348 8623 34388 8632
rect 34539 8672 34581 8681
rect 34539 8632 34540 8672
rect 34580 8632 34581 8672
rect 34539 8623 34581 8632
rect 34540 8538 34580 8623
rect 34592 8336 34960 8345
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34592 8287 34960 8296
rect 35692 8009 35732 9220
rect 35884 8681 35924 10732
rect 36940 10184 36980 13159
rect 38860 13074 38900 13159
rect 39724 13074 39764 13159
rect 40875 13040 40917 13049
rect 40875 13000 40876 13040
rect 40916 13000 40917 13040
rect 40875 12991 40917 13000
rect 40876 12906 40916 12991
rect 38187 12536 38229 12545
rect 38187 12496 38188 12536
rect 38228 12496 38229 12536
rect 38187 12487 38229 12496
rect 37035 12284 37077 12293
rect 37035 12244 37036 12284
rect 37076 12244 37077 12284
rect 37035 12235 37077 12244
rect 37036 11024 37076 12235
rect 38188 11705 38228 12487
rect 41164 12461 41204 13159
rect 41644 13049 41684 13168
rect 41643 13040 41685 13049
rect 41643 13000 41644 13040
rect 41684 13000 41685 13040
rect 41643 12991 41685 13000
rect 41163 12452 41205 12461
rect 41163 12412 41164 12452
rect 41204 12412 41205 12452
rect 41163 12403 41205 12412
rect 41164 12318 41204 12403
rect 41451 12284 41493 12293
rect 41451 12244 41452 12284
rect 41492 12244 41493 12284
rect 41451 12235 41493 12244
rect 41355 11864 41397 11873
rect 41355 11824 41356 11864
rect 41396 11824 41397 11864
rect 41355 11815 41397 11824
rect 38187 11696 38229 11705
rect 38187 11656 38188 11696
rect 38228 11656 38229 11696
rect 38187 11647 38229 11656
rect 41356 11696 41396 11815
rect 41356 11647 41396 11656
rect 37899 11192 37941 11201
rect 37899 11152 37900 11192
rect 37940 11152 37941 11192
rect 37899 11143 37941 11152
rect 37900 11024 37940 11143
rect 37076 10984 37172 11024
rect 37036 10975 37076 10984
rect 37036 10184 37076 10193
rect 36940 10144 37036 10184
rect 37036 10135 37076 10144
rect 37132 9521 37172 10984
rect 37900 10268 37940 10984
rect 37804 10228 37900 10268
rect 36364 9512 36404 9521
rect 36364 9353 36404 9472
rect 37131 9512 37173 9521
rect 37131 9472 37132 9512
rect 37172 9472 37173 9512
rect 37131 9463 37173 9472
rect 36363 9344 36405 9353
rect 36363 9304 36364 9344
rect 36404 9304 36405 9344
rect 36363 9295 36405 9304
rect 37131 9344 37173 9353
rect 37131 9304 37132 9344
rect 37172 9304 37173 9344
rect 37131 9295 37173 9304
rect 37132 9210 37172 9295
rect 35883 8672 35925 8681
rect 35883 8632 35884 8672
rect 35924 8632 35925 8672
rect 35883 8623 35925 8632
rect 34444 8000 34484 8009
rect 33196 7160 33236 7169
rect 33196 6656 33236 7120
rect 33388 7160 33428 7372
rect 34252 7363 34292 7372
rect 34348 7960 34444 8000
rect 33388 7111 33428 7120
rect 33580 7160 33620 7169
rect 33484 6656 33524 6665
rect 33196 6616 33484 6656
rect 33484 6607 33524 6616
rect 32331 6404 32373 6413
rect 32331 6364 32332 6404
rect 32372 6364 32373 6404
rect 32331 6355 32373 6364
rect 31468 5648 31508 5657
rect 30892 5564 30932 5573
rect 31084 5564 31124 5573
rect 30932 5524 31084 5564
rect 30892 5515 30932 5524
rect 31084 5515 31124 5524
rect 31468 4985 31508 5608
rect 32332 5648 32372 6355
rect 33580 6320 33620 7120
rect 34348 6908 34388 7960
rect 34444 7951 34484 7960
rect 35691 8000 35733 8009
rect 35691 7960 35692 8000
rect 35732 7960 35733 8000
rect 35691 7951 35733 7960
rect 35307 7580 35349 7589
rect 35307 7540 35308 7580
rect 35348 7540 35349 7580
rect 35307 7531 35349 7540
rect 34156 6868 34388 6908
rect 34156 6488 34196 6868
rect 34592 6824 34960 6833
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34592 6775 34960 6784
rect 33964 6448 34156 6488
rect 33580 6280 33812 6320
rect 33352 6068 33720 6077
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33352 6019 33720 6028
rect 33483 5900 33525 5909
rect 33483 5860 33484 5900
rect 33524 5860 33525 5900
rect 33483 5851 33525 5860
rect 33484 5766 33524 5851
rect 31467 4976 31509 4985
rect 31467 4936 31468 4976
rect 31508 4936 31509 4976
rect 31467 4927 31509 4936
rect 30795 4304 30837 4313
rect 30795 4264 30796 4304
rect 30836 4264 30837 4304
rect 30795 4255 30837 4264
rect 30988 4136 31028 4145
rect 30604 4096 30988 4136
rect 30604 2876 30644 4096
rect 30988 4087 31028 4096
rect 31083 3968 31125 3977
rect 31083 3928 31084 3968
rect 31124 3928 31125 3968
rect 31083 3919 31125 3928
rect 31084 3464 31124 3919
rect 31084 3415 31124 3424
rect 31468 3464 31508 4927
rect 31659 3968 31701 3977
rect 31659 3928 31660 3968
rect 31700 3928 31701 3968
rect 31659 3919 31701 3928
rect 31660 3834 31700 3919
rect 31468 3415 31508 3424
rect 32332 3464 32372 5608
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 32332 3415 32372 3424
rect 33580 3464 33620 3473
rect 33772 3464 33812 6280
rect 33964 5909 34004 6448
rect 34156 6439 34196 6448
rect 34347 6488 34389 6497
rect 34347 6448 34348 6488
rect 34388 6448 34389 6488
rect 34347 6439 34389 6448
rect 35308 6488 35348 7531
rect 35308 6439 35348 6448
rect 34348 6354 34388 6439
rect 37804 6320 37844 10228
rect 37900 10219 37940 10228
rect 38188 10184 38228 11647
rect 40684 11528 40724 11537
rect 39147 11192 39189 11201
rect 39147 11152 39148 11192
rect 39188 11152 39189 11192
rect 39147 11143 39189 11152
rect 38283 11108 38325 11117
rect 38283 11068 38284 11108
rect 38324 11068 38325 11108
rect 38283 11059 38325 11068
rect 38284 11024 38324 11059
rect 38284 10973 38324 10984
rect 38379 11024 38421 11033
rect 38379 10984 38380 11024
rect 38420 10984 38421 11024
rect 38379 10975 38421 10984
rect 39051 11024 39093 11033
rect 39051 10984 39052 11024
rect 39092 10984 39093 11024
rect 39051 10975 39093 10984
rect 38188 10135 38228 10144
rect 38283 9512 38325 9521
rect 38283 9472 38284 9512
rect 38324 9472 38325 9512
rect 38283 9463 38325 9472
rect 38284 9378 38324 9463
rect 38380 8672 38420 10975
rect 39052 10193 39092 10975
rect 39051 10184 39093 10193
rect 39051 10144 39052 10184
rect 39092 10144 39093 10184
rect 39051 10135 39093 10144
rect 39052 10050 39092 10135
rect 39148 9512 39188 11143
rect 40684 11117 40724 11488
rect 40683 11108 40725 11117
rect 40683 11068 40684 11108
rect 40724 11068 40725 11108
rect 40683 11059 40725 11068
rect 41164 11024 41204 11033
rect 39531 10772 39573 10781
rect 39531 10732 39532 10772
rect 39572 10732 39573 10772
rect 39531 10723 39573 10732
rect 40491 10772 40533 10781
rect 40491 10732 40492 10772
rect 40532 10732 40533 10772
rect 40491 10723 40533 10732
rect 39532 9596 39572 10723
rect 40492 10638 40532 10723
rect 41164 10100 41204 10984
rect 41452 10184 41492 12235
rect 41644 12116 41684 12991
rect 41740 12536 41780 12545
rect 41780 12496 41876 12536
rect 41740 12487 41780 12496
rect 41644 12076 41780 12116
rect 41643 11696 41685 11705
rect 41643 11656 41644 11696
rect 41684 11656 41685 11696
rect 41643 11647 41685 11656
rect 41644 11562 41684 11647
rect 41452 10135 41492 10144
rect 41740 10184 41780 12076
rect 41836 11192 41876 12496
rect 41931 12452 41973 12461
rect 41931 12412 41932 12452
rect 41972 12412 41973 12452
rect 41931 12403 41973 12412
rect 41932 11948 41972 12403
rect 41932 11899 41972 11908
rect 41932 11192 41972 11201
rect 41836 11152 41932 11192
rect 41932 11143 41972 11152
rect 41740 10135 41780 10144
rect 41260 10100 41300 10109
rect 41164 10060 41260 10100
rect 41260 10051 41300 10060
rect 39532 9547 39572 9556
rect 39148 9463 39188 9472
rect 42220 8672 42260 15100
rect 42316 13040 42356 13049
rect 42356 13000 42836 13040
rect 42316 12991 42356 13000
rect 42699 12620 42741 12629
rect 42699 12580 42700 12620
rect 42740 12580 42741 12620
rect 42699 12571 42741 12580
rect 42604 12536 42644 12545
rect 42604 12293 42644 12496
rect 42700 12486 42740 12571
rect 42796 12536 42836 13000
rect 42796 12487 42836 12496
rect 42988 12461 43028 15520
rect 44140 15308 44180 15317
rect 44140 15140 44180 15268
rect 46348 15140 46388 16024
rect 44044 15100 44180 15140
rect 46252 15100 46388 15140
rect 48472 15140 48840 15149
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 43564 14132 43604 14141
rect 43180 14092 43564 14132
rect 43083 12620 43125 12629
rect 43083 12580 43084 12620
rect 43124 12580 43125 12620
rect 43083 12571 43125 12580
rect 42987 12452 43029 12461
rect 42987 12412 42988 12452
rect 43028 12412 43029 12452
rect 42987 12403 43029 12412
rect 42411 12284 42453 12293
rect 42411 12244 42412 12284
rect 42452 12244 42453 12284
rect 42411 12235 42453 12244
rect 42603 12284 42645 12293
rect 42603 12244 42604 12284
rect 42644 12244 42645 12284
rect 42603 12235 42645 12244
rect 42412 12150 42452 12235
rect 42891 11864 42933 11873
rect 42891 11824 42892 11864
rect 42932 11824 42933 11864
rect 42891 11815 42933 11824
rect 42892 11730 42932 11815
rect 42604 11696 42644 11705
rect 42604 11537 42644 11656
rect 43084 11696 43124 12571
rect 43084 11647 43124 11656
rect 43180 11696 43220 14092
rect 43564 14083 43604 14092
rect 43756 14048 43796 14059
rect 43756 13973 43796 14008
rect 44044 14048 44084 15100
rect 44044 13999 44084 14008
rect 45387 14048 45429 14057
rect 45387 14008 45388 14048
rect 45428 14008 45429 14048
rect 45387 13999 45429 14008
rect 46252 14048 46292 15100
rect 48472 15091 48840 15100
rect 49036 14057 49076 17032
rect 49712 15896 50080 15905
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 49712 15847 50080 15856
rect 50284 15140 50324 18451
rect 52012 18332 52052 18341
rect 52012 17921 52052 18292
rect 51339 17912 51381 17921
rect 51339 17872 51340 17912
rect 51380 17872 51381 17912
rect 51339 17863 51381 17872
rect 52011 17912 52053 17921
rect 52011 17872 52012 17912
rect 52052 17872 52053 17912
rect 52011 17863 52053 17872
rect 52299 17912 52341 17921
rect 52299 17872 52300 17912
rect 52340 17872 52341 17912
rect 52299 17863 52341 17872
rect 51147 17744 51189 17753
rect 50380 17711 50420 17720
rect 51147 17704 51148 17744
rect 51188 17704 51189 17744
rect 51147 17695 51189 17704
rect 51340 17744 51380 17863
rect 51340 17695 51380 17704
rect 50380 17417 50420 17671
rect 51148 17610 51188 17695
rect 51243 17660 51285 17669
rect 51243 17620 51244 17660
rect 51284 17620 51285 17660
rect 51243 17611 51285 17620
rect 51244 17526 51284 17611
rect 52300 17576 52340 17863
rect 52396 17744 52436 18871
rect 55180 18584 55220 18871
rect 55180 18535 55220 18544
rect 55372 18584 55412 19300
rect 56811 19300 56812 19340
rect 56852 19300 56853 19340
rect 56811 19291 56853 19300
rect 56043 19256 56085 19265
rect 56043 19216 56044 19256
rect 56084 19216 56085 19256
rect 56043 19207 56085 19216
rect 56908 19256 56948 20047
rect 57484 19517 57524 20056
rect 63592 19676 63960 19685
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63592 19627 63960 19636
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 93832 19676 94200 19685
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 93832 19627 94200 19636
rect 57483 19508 57525 19517
rect 57483 19468 57484 19508
rect 57524 19468 57525 19508
rect 57483 19459 57525 19468
rect 58059 19508 58101 19517
rect 58059 19468 58060 19508
rect 58100 19468 58101 19508
rect 58059 19459 58101 19468
rect 58060 19374 58100 19459
rect 56908 19207 56948 19216
rect 57003 19256 57045 19265
rect 57003 19216 57004 19256
rect 57044 19216 57045 19256
rect 57003 19207 57045 19216
rect 55660 19172 55700 19181
rect 55468 19088 55508 19097
rect 55660 19088 55700 19132
rect 56044 19122 56084 19207
rect 55508 19048 55700 19088
rect 55468 19039 55508 19048
rect 55372 18535 55412 18544
rect 55276 18332 55316 18341
rect 52396 17695 52436 17704
rect 55180 17744 55220 17753
rect 55276 17744 55316 18292
rect 55220 17704 55316 17744
rect 55468 17744 55508 17755
rect 55180 17695 55220 17704
rect 55468 17669 55508 17704
rect 55467 17660 55509 17669
rect 55467 17620 55468 17660
rect 55508 17620 55509 17660
rect 55467 17611 55509 17620
rect 52300 17527 52340 17536
rect 52588 17576 52628 17585
rect 50379 17408 50421 17417
rect 50379 17368 50380 17408
rect 50420 17368 50421 17408
rect 50379 17359 50421 17368
rect 52588 17156 52628 17536
rect 55660 17576 55700 17585
rect 55700 17536 56660 17576
rect 55660 17527 55700 17536
rect 52780 17156 52820 17165
rect 52588 17116 52780 17156
rect 52780 17107 52820 17116
rect 56620 17156 56660 17536
rect 56620 17107 56660 17116
rect 53163 17072 53205 17081
rect 53163 17032 53164 17072
rect 53204 17032 53205 17072
rect 53163 17023 53205 17032
rect 54028 17072 54068 17081
rect 50188 15100 50324 15140
rect 49712 14384 50080 14393
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 49712 14335 50080 14344
rect 46252 13999 46292 14008
rect 46636 14048 46676 14057
rect 47308 14048 47348 14057
rect 46676 14008 47308 14048
rect 46636 13999 46676 14008
rect 47308 13999 47348 14008
rect 47980 14048 48020 14057
rect 43755 13964 43797 13973
rect 43755 13924 43756 13964
rect 43796 13924 43797 13964
rect 43755 13915 43797 13924
rect 44235 13964 44277 13973
rect 44235 13924 44236 13964
rect 44276 13924 44277 13964
rect 44235 13915 44277 13924
rect 44236 13830 44276 13915
rect 45388 13914 45428 13999
rect 47980 13889 48020 14008
rect 49035 14048 49077 14057
rect 49035 14008 49036 14048
rect 49076 14008 49077 14048
rect 49035 13999 49077 14008
rect 49323 14048 49365 14057
rect 49323 14008 49324 14048
rect 49364 14008 49365 14048
rect 49323 13999 49365 14008
rect 50188 14048 50228 15100
rect 51531 14888 51573 14897
rect 51531 14848 51532 14888
rect 51572 14848 51573 14888
rect 51531 14839 51573 14848
rect 51532 14754 51572 14839
rect 51244 14720 51284 14729
rect 50571 14132 50613 14141
rect 50571 14092 50572 14132
rect 50612 14092 50613 14132
rect 50571 14083 50613 14092
rect 50188 13999 50228 14008
rect 49324 13914 49364 13999
rect 50572 13998 50612 14083
rect 51244 14057 51284 14680
rect 52203 14720 52245 14729
rect 52203 14680 52204 14720
rect 52244 14680 52245 14720
rect 52203 14671 52245 14680
rect 52204 14586 52244 14671
rect 52972 14552 53012 14561
rect 52972 14141 53012 14512
rect 52971 14132 53013 14141
rect 52971 14092 52972 14132
rect 53012 14092 53013 14132
rect 52971 14083 53013 14092
rect 51243 14048 51285 14057
rect 51243 14008 51244 14048
rect 51284 14008 51285 14048
rect 51243 13999 51285 14008
rect 47979 13880 48021 13889
rect 47979 13840 47980 13880
rect 48020 13840 48021 13880
rect 47979 13831 48021 13840
rect 49611 13880 49653 13889
rect 49611 13840 49612 13880
rect 49652 13840 49653 13880
rect 49611 13831 49653 13840
rect 48172 13796 48212 13805
rect 48212 13756 48404 13796
rect 48172 13747 48212 13756
rect 48364 13208 48404 13756
rect 48472 13628 48840 13637
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48472 13579 48840 13588
rect 49612 13460 49652 13831
rect 49612 13411 49652 13420
rect 48652 13208 48692 13217
rect 49804 13208 49844 13217
rect 48364 13168 48652 13208
rect 48652 13159 48692 13168
rect 49420 13168 49804 13208
rect 49324 13040 49364 13049
rect 49324 12536 49364 13000
rect 49420 12620 49460 13168
rect 49804 13159 49844 13168
rect 49900 13208 49940 13217
rect 49940 13168 50516 13208
rect 49900 13159 49940 13168
rect 49712 12872 50080 12881
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 49712 12823 50080 12832
rect 50476 12704 50516 13168
rect 50476 12655 50516 12664
rect 49420 12571 49460 12580
rect 49036 12496 49324 12536
rect 48472 12116 48840 12125
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48472 12067 48840 12076
rect 43180 11647 43220 11656
rect 47307 11696 47349 11705
rect 47307 11656 47308 11696
rect 47348 11656 47349 11696
rect 47307 11647 47349 11656
rect 48843 11696 48885 11705
rect 48843 11656 48844 11696
rect 48884 11656 48885 11696
rect 48843 11647 48885 11656
rect 49036 11696 49076 12496
rect 49324 12487 49364 12496
rect 49516 12536 49556 12545
rect 49516 11948 49556 12496
rect 50571 12536 50613 12545
rect 50956 12536 50996 12545
rect 50571 12496 50572 12536
rect 50612 12496 50613 12536
rect 50571 12487 50613 12496
rect 50668 12496 50956 12536
rect 50572 12402 50612 12487
rect 49516 11899 49556 11908
rect 49324 11696 49364 11705
rect 50188 11696 50228 11705
rect 49036 11647 49076 11656
rect 49228 11656 49324 11696
rect 49364 11656 50188 11696
rect 47308 11562 47348 11647
rect 48844 11612 48884 11647
rect 48844 11561 48884 11572
rect 42603 11528 42645 11537
rect 42603 11488 42604 11528
rect 42644 11488 42645 11528
rect 42603 11479 42645 11488
rect 43083 11528 43125 11537
rect 43083 11488 43084 11528
rect 43124 11488 43125 11528
rect 43083 11479 43125 11488
rect 46636 11528 46676 11537
rect 43084 11024 43124 11479
rect 43947 11192 43989 11201
rect 43947 11152 43948 11192
rect 43988 11152 43989 11192
rect 43947 11143 43989 11152
rect 42508 8672 42548 8681
rect 42220 8632 42508 8672
rect 43084 8672 43124 10984
rect 43948 11024 43988 11143
rect 46636 11117 46676 11488
rect 44331 11108 44373 11117
rect 44331 11068 44332 11108
rect 44372 11068 44373 11108
rect 44331 11059 44373 11068
rect 46635 11108 46677 11117
rect 46635 11068 46636 11108
rect 46676 11068 46677 11108
rect 46635 11059 46677 11068
rect 43948 10975 43988 10984
rect 44332 10974 44372 11059
rect 48472 10604 48840 10613
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48472 10555 48840 10564
rect 49228 10436 49268 11656
rect 49324 11647 49364 11656
rect 50188 11647 50228 11656
rect 49712 11360 50080 11369
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 49712 11311 50080 11320
rect 50668 10856 50708 12496
rect 50956 12487 50996 12496
rect 53164 12536 53204 17023
rect 54028 14897 54068 17032
rect 57004 17072 57044 19207
rect 64832 18920 65200 18929
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 64832 18871 65200 18880
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 95072 18920 95440 18929
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95072 18871 95440 18880
rect 63592 18164 63960 18173
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63592 18115 63960 18124
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 93832 18164 94200 18173
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 93832 18115 94200 18124
rect 64832 17408 65200 17417
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 64832 17359 65200 17368
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 95072 17408 95440 17417
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95072 17359 95440 17368
rect 57004 17023 57044 17032
rect 57868 17072 57908 17081
rect 55179 16820 55221 16829
rect 55179 16780 55180 16820
rect 55220 16780 55221 16820
rect 55179 16771 55221 16780
rect 56043 16820 56085 16829
rect 56043 16780 56044 16820
rect 56084 16780 56085 16820
rect 56043 16771 56085 16780
rect 55180 16686 55220 16771
rect 56044 16232 56084 16771
rect 56044 16183 56084 16192
rect 55372 16064 55412 16073
rect 54027 14888 54069 14897
rect 54027 14848 54028 14888
rect 54068 14848 54069 14888
rect 54027 14839 54069 14848
rect 53644 14720 53684 14729
rect 53644 14225 53684 14680
rect 53835 14720 53877 14729
rect 53835 14680 53836 14720
rect 53876 14680 53877 14720
rect 53835 14671 53877 14680
rect 53643 14216 53685 14225
rect 53643 14176 53644 14216
rect 53684 14176 53685 14216
rect 53643 14167 53685 14176
rect 53836 14057 53876 14671
rect 54028 14309 54068 14839
rect 55372 14720 55412 16024
rect 55468 14888 55508 14897
rect 55508 14848 56084 14888
rect 55468 14839 55508 14848
rect 54027 14300 54069 14309
rect 54027 14260 54028 14300
rect 54068 14260 54069 14300
rect 54027 14251 54069 14260
rect 54795 14300 54837 14309
rect 54795 14260 54796 14300
rect 54836 14260 54837 14300
rect 54795 14251 54837 14260
rect 53835 14048 53877 14057
rect 53835 14008 53836 14048
rect 53876 14008 53877 14048
rect 53835 13999 53877 14008
rect 53644 13040 53684 13049
rect 53644 12545 53684 13000
rect 53164 11033 53204 12496
rect 53643 12536 53685 12545
rect 53643 12496 53644 12536
rect 53684 12496 53685 12536
rect 53643 12487 53685 12496
rect 53836 11948 53876 13999
rect 54796 13208 54836 14251
rect 55179 14216 55221 14225
rect 55179 14176 55180 14216
rect 55220 14176 55221 14216
rect 55179 14167 55221 14176
rect 55180 14082 55220 14167
rect 55372 14048 55412 14680
rect 55563 14720 55605 14729
rect 55563 14680 55564 14720
rect 55604 14680 55605 14720
rect 55563 14671 55605 14680
rect 56044 14720 56084 14848
rect 56523 14804 56565 14813
rect 56523 14764 56524 14804
rect 56564 14764 56565 14804
rect 56523 14755 56565 14764
rect 56044 14671 56084 14680
rect 56139 14720 56181 14729
rect 56139 14680 56140 14720
rect 56180 14680 56181 14720
rect 56139 14671 56181 14680
rect 55564 14586 55604 14671
rect 56140 14586 56180 14671
rect 56524 14670 56564 14755
rect 57196 14720 57236 14729
rect 56331 14552 56373 14561
rect 56331 14512 56332 14552
rect 56372 14512 56373 14552
rect 56331 14503 56373 14512
rect 56715 14552 56757 14561
rect 56715 14512 56716 14552
rect 56756 14512 56757 14552
rect 56715 14503 56757 14512
rect 56332 14418 56372 14503
rect 55659 14132 55701 14141
rect 55659 14092 55660 14132
rect 55700 14092 55701 14132
rect 55659 14083 55701 14092
rect 55372 13999 55412 14008
rect 55660 14048 55700 14083
rect 55660 13997 55700 14008
rect 56716 14048 56756 14503
rect 57196 14141 57236 14680
rect 56811 14132 56853 14141
rect 56811 14092 56812 14132
rect 56852 14092 56853 14132
rect 56811 14083 56853 14092
rect 57195 14132 57237 14141
rect 57195 14092 57196 14132
rect 57236 14092 57237 14132
rect 57195 14083 57237 14092
rect 57868 14132 57908 17032
rect 59020 16820 59060 16829
rect 59020 14729 59060 16780
rect 63592 16652 63960 16661
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63592 16603 63960 16612
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 93832 16652 94200 16661
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 93832 16603 94200 16612
rect 64832 15896 65200 15905
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 64832 15847 65200 15856
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 95072 15896 95440 15905
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95072 15847 95440 15856
rect 63592 15140 63960 15149
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63592 15091 63960 15100
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 93832 15140 94200 15149
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 93832 15091 94200 15100
rect 59019 14720 59061 14729
rect 59019 14680 59020 14720
rect 59060 14680 59061 14720
rect 59019 14671 59061 14680
rect 59403 14720 59445 14729
rect 59403 14680 59404 14720
rect 59444 14680 59445 14720
rect 59403 14671 59445 14680
rect 59788 14720 59828 14729
rect 59307 14636 59349 14645
rect 59307 14596 59308 14636
rect 59348 14596 59349 14636
rect 59307 14587 59349 14596
rect 59308 14502 59348 14587
rect 59404 14586 59444 14671
rect 59788 14225 59828 14680
rect 64832 14384 65200 14393
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 64832 14335 65200 14344
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 95072 14384 95440 14393
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95072 14335 95440 14344
rect 59787 14216 59829 14225
rect 59787 14176 59788 14216
rect 59828 14176 59829 14216
rect 59787 14167 59829 14176
rect 61419 14216 61461 14225
rect 61419 14176 61420 14216
rect 61460 14176 61461 14216
rect 61419 14167 61461 14176
rect 56716 13999 56756 14008
rect 56619 13880 56661 13889
rect 56619 13840 56620 13880
rect 56660 13840 56661 13880
rect 56619 13831 56661 13840
rect 56044 13796 56084 13805
rect 55660 13208 55700 13217
rect 54796 13159 54836 13168
rect 55564 13168 55660 13208
rect 54124 12536 54164 12545
rect 54124 12377 54164 12496
rect 54412 12536 54452 12545
rect 54796 12536 54836 12545
rect 54452 12496 54740 12536
rect 54412 12487 54452 12496
rect 54123 12368 54165 12377
rect 54123 12328 54124 12368
rect 54164 12328 54165 12368
rect 54123 12319 54165 12328
rect 53836 11899 53876 11908
rect 53548 11696 53588 11705
rect 53452 11656 53548 11696
rect 52587 11024 52629 11033
rect 52587 10984 52588 11024
rect 52628 10984 52629 11024
rect 52587 10975 52629 10984
rect 53163 11024 53205 11033
rect 53163 10984 53164 11024
rect 53204 10984 53205 11024
rect 53163 10975 53205 10984
rect 49228 10387 49268 10396
rect 50476 10816 50708 10856
rect 51724 10940 51764 10949
rect 47212 10184 47252 10195
rect 47212 10109 47252 10144
rect 48076 10184 48116 10193
rect 46828 10100 46868 10109
rect 47211 10100 47253 10109
rect 46868 10060 47060 10100
rect 46828 10051 46868 10060
rect 47020 9680 47060 10060
rect 47211 10060 47212 10100
rect 47252 10060 47253 10100
rect 47211 10051 47253 10060
rect 48076 9689 48116 10144
rect 48459 10100 48501 10109
rect 48459 10060 48460 10100
rect 48500 10060 48501 10100
rect 48459 10051 48501 10060
rect 47020 9631 47060 9640
rect 48075 9680 48117 9689
rect 48075 9640 48076 9680
rect 48116 9640 48117 9680
rect 48075 9631 48117 9640
rect 46348 9512 46388 9521
rect 47212 9512 47252 9521
rect 47884 9512 47924 9521
rect 48076 9512 48116 9521
rect 48460 9512 48500 10051
rect 49712 9848 50080 9857
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 49712 9799 50080 9808
rect 49323 9680 49365 9689
rect 49323 9640 49324 9680
rect 49364 9640 49365 9680
rect 49323 9631 49365 9640
rect 50476 9680 50516 10816
rect 51724 10109 51764 10900
rect 52588 10890 52628 10975
rect 53452 10193 53492 11656
rect 53548 11647 53588 11656
rect 54700 10436 54740 12496
rect 54796 12377 54836 12496
rect 54795 12368 54837 12377
rect 54795 12328 54796 12368
rect 54836 12328 54837 12368
rect 55564 12368 55604 13168
rect 55660 13159 55700 13168
rect 56044 13208 56084 13756
rect 56044 13159 56084 13168
rect 56620 13208 56660 13831
rect 55660 12536 55700 12545
rect 56620 12536 56660 13168
rect 55700 12496 56660 12536
rect 55660 12487 55700 12496
rect 56812 12452 56852 14083
rect 57868 14057 57908 14092
rect 61420 14082 61460 14167
rect 57003 14048 57045 14057
rect 57003 14008 57004 14048
rect 57044 14008 57045 14048
rect 57003 13999 57045 14008
rect 57867 14048 57909 14057
rect 57867 14008 57868 14048
rect 57908 14008 57909 14048
rect 57867 13999 57909 14008
rect 59020 14048 59060 14057
rect 59404 14048 59444 14057
rect 60267 14048 60309 14057
rect 59060 14008 59252 14048
rect 59020 13999 59060 14008
rect 57004 13914 57044 13999
rect 57868 13968 57908 13999
rect 57291 13880 57333 13889
rect 57291 13840 57292 13880
rect 57332 13840 57333 13880
rect 57291 13831 57333 13840
rect 57292 13746 57332 13831
rect 56812 12403 56852 12412
rect 55659 12368 55701 12377
rect 55564 12328 55660 12368
rect 55700 12328 55701 12368
rect 54795 12319 54837 12328
rect 55659 12319 55701 12328
rect 55180 10436 55220 10445
rect 54700 10396 55180 10436
rect 55180 10387 55220 10396
rect 55467 10352 55509 10361
rect 55467 10312 55468 10352
rect 55508 10312 55509 10352
rect 55467 10303 55509 10312
rect 53451 10184 53493 10193
rect 53451 10144 53452 10184
rect 53492 10144 53493 10184
rect 53451 10135 53493 10144
rect 55371 10184 55413 10193
rect 55371 10144 55372 10184
rect 55412 10144 55413 10184
rect 55371 10135 55413 10144
rect 51723 10100 51765 10109
rect 51723 10060 51724 10100
rect 51764 10060 51765 10100
rect 51723 10051 51765 10060
rect 52395 10100 52437 10109
rect 52395 10060 52396 10100
rect 52436 10060 52437 10100
rect 52395 10051 52437 10060
rect 50476 9631 50516 9640
rect 46388 9472 46484 9512
rect 46348 9463 46388 9472
rect 44523 8756 44565 8765
rect 44523 8716 44524 8756
rect 44564 8716 44565 8756
rect 44523 8707 44565 8716
rect 45675 8756 45717 8765
rect 45675 8716 45676 8756
rect 45716 8716 45717 8756
rect 45675 8707 45717 8716
rect 43372 8672 43412 8681
rect 43084 8632 43372 8672
rect 38380 8623 38420 8632
rect 42508 8623 42548 8632
rect 40971 8588 41013 8597
rect 40971 8548 40972 8588
rect 41012 8548 41013 8588
rect 40971 8539 41013 8548
rect 42123 8588 42165 8597
rect 42123 8548 42124 8588
rect 42164 8548 42165 8588
rect 42123 8539 42165 8548
rect 37996 8504 38036 8513
rect 37996 7589 38036 8464
rect 37995 7580 38037 7589
rect 37995 7540 37996 7580
rect 38036 7540 38037 7580
rect 37995 7531 38037 7540
rect 39915 7580 39957 7589
rect 39915 7540 39916 7580
rect 39956 7540 39957 7580
rect 39915 7531 39957 7540
rect 38859 7244 38901 7253
rect 38859 7204 38860 7244
rect 38900 7204 38901 7244
rect 38859 7195 38901 7204
rect 39531 7244 39573 7253
rect 39531 7204 39532 7244
rect 39572 7204 39573 7244
rect 39531 7195 39573 7204
rect 39723 7244 39765 7253
rect 39723 7204 39724 7244
rect 39764 7204 39765 7244
rect 39723 7195 39765 7204
rect 38860 7110 38900 7195
rect 38668 6992 38708 7001
rect 37900 6952 38668 6992
rect 37900 6572 37940 6952
rect 38668 6943 38708 6952
rect 39532 6581 39572 7195
rect 39724 7110 39764 7195
rect 37900 6523 37940 6532
rect 39531 6572 39573 6581
rect 39531 6532 39532 6572
rect 39572 6532 39573 6572
rect 39531 6523 39573 6532
rect 38284 6488 38324 6497
rect 38284 6320 38324 6448
rect 39147 6488 39189 6497
rect 39147 6448 39148 6488
rect 39188 6448 39189 6488
rect 39147 6439 39189 6448
rect 39148 6354 39188 6439
rect 37804 6280 38324 6320
rect 33963 5900 34005 5909
rect 33963 5860 33964 5900
rect 34004 5860 34005 5900
rect 33963 5851 34005 5860
rect 37420 5732 37460 5743
rect 37420 5657 37460 5692
rect 35979 5648 36021 5657
rect 35979 5608 35980 5648
rect 36020 5608 36021 5648
rect 35979 5599 36021 5608
rect 36555 5648 36597 5657
rect 36555 5608 36556 5648
rect 36596 5608 36597 5648
rect 36555 5599 36597 5608
rect 37227 5648 37269 5657
rect 37227 5608 37228 5648
rect 37268 5608 37269 5648
rect 37227 5599 37269 5608
rect 37419 5648 37461 5657
rect 37419 5608 37420 5648
rect 37460 5608 37461 5648
rect 37419 5599 37461 5608
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 35980 4892 36020 5599
rect 36556 5514 36596 5599
rect 37228 5514 37268 5599
rect 37612 5480 37652 5489
rect 37612 5069 37652 5440
rect 37611 5060 37653 5069
rect 37611 5020 37612 5060
rect 37652 5020 37653 5060
rect 37611 5011 37653 5020
rect 37132 4976 37172 4987
rect 37132 4901 37172 4936
rect 37996 4976 38036 6280
rect 39339 5648 39381 5657
rect 39339 5608 39340 5648
rect 39380 5608 39381 5648
rect 39339 5599 39381 5608
rect 39532 5648 39572 6523
rect 39532 5599 39572 5608
rect 39340 5514 39380 5599
rect 39435 5564 39477 5573
rect 39435 5524 39436 5564
rect 39476 5524 39477 5564
rect 39435 5515 39477 5524
rect 39436 5430 39476 5515
rect 38379 5060 38421 5069
rect 38379 5020 38380 5060
rect 38420 5020 38421 5060
rect 38379 5011 38421 5020
rect 35980 4843 36020 4852
rect 37131 4892 37173 4901
rect 37131 4852 37132 4892
rect 37172 4852 37173 4892
rect 37131 4843 37173 4852
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 33620 3424 33812 3464
rect 33580 3415 33620 3424
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 30604 2827 30644 2836
rect 37996 2717 38036 4936
rect 38380 4926 38420 5011
rect 39916 4976 39956 7531
rect 40396 7160 40436 7169
rect 40300 6656 40340 6665
rect 40396 6656 40436 7120
rect 40340 6616 40436 6656
rect 40684 6656 40724 6665
rect 40300 6607 40340 6616
rect 39916 4927 39956 4936
rect 39435 4892 39477 4901
rect 39435 4852 39436 4892
rect 39476 4852 39477 4892
rect 39435 4843 39477 4852
rect 40203 4892 40245 4901
rect 40203 4852 40204 4892
rect 40244 4852 40245 4892
rect 40203 4843 40245 4852
rect 39436 4758 39476 4843
rect 40204 4724 40244 4843
rect 39435 4136 39477 4145
rect 39435 4096 39436 4136
rect 39476 4096 39477 4136
rect 39435 4087 39477 4096
rect 40107 4136 40149 4145
rect 40107 4096 40108 4136
rect 40148 4096 40149 4136
rect 40107 4087 40149 4096
rect 39436 3380 39476 4087
rect 40108 3632 40148 4087
rect 40108 3583 40148 3592
rect 39436 3331 39476 3340
rect 38091 3212 38133 3221
rect 38091 3172 38092 3212
rect 38132 3172 38133 3212
rect 38091 3163 38133 3172
rect 39243 3212 39285 3221
rect 39243 3172 39244 3212
rect 39284 3172 39285 3212
rect 39243 3163 39285 3172
rect 37995 2708 38037 2717
rect 37995 2668 37996 2708
rect 38036 2668 38037 2708
rect 37995 2659 38037 2668
rect 29452 2624 29492 2633
rect 28972 2584 29452 2624
rect 28587 2575 28629 2584
rect 29452 2575 29492 2584
rect 38092 2624 38132 3163
rect 39244 3078 39284 3163
rect 38475 2708 38517 2717
rect 38475 2668 38476 2708
rect 38516 2668 38517 2708
rect 38475 2659 38517 2668
rect 38092 2575 38132 2584
rect 38476 2624 38516 2659
rect 40204 2633 40244 4684
rect 40684 4145 40724 6616
rect 40972 6656 41012 8539
rect 42124 8454 42164 8539
rect 40972 6607 41012 6616
rect 40779 6572 40821 6581
rect 40779 6532 40780 6572
rect 40820 6532 40821 6572
rect 40779 6523 40821 6532
rect 40780 6488 40820 6523
rect 43372 6497 43412 8632
rect 44524 8622 44564 8707
rect 45676 8672 45716 8707
rect 45676 8621 45716 8632
rect 46444 8588 46484 9472
rect 47252 9472 47540 9512
rect 47212 9463 47252 9472
rect 47115 8756 47157 8765
rect 47115 8716 47116 8756
rect 47156 8716 47157 8756
rect 47115 8707 47157 8716
rect 46732 8672 46772 8681
rect 46636 8588 46676 8597
rect 46444 8548 46636 8588
rect 46636 8539 46676 8548
rect 46348 8504 46388 8513
rect 46388 8464 46580 8504
rect 46348 8455 46388 8464
rect 46540 8000 46580 8464
rect 46732 8093 46772 8632
rect 47116 8672 47156 8707
rect 47116 8621 47156 8632
rect 47500 8168 47540 9472
rect 47924 9472 48076 9512
rect 47884 9463 47924 9472
rect 48076 9463 48116 9472
rect 48364 9472 48460 9512
rect 47500 8119 47540 8128
rect 46731 8084 46773 8093
rect 46731 8044 46732 8084
rect 46772 8044 46773 8084
rect 46731 8035 46773 8044
rect 46540 7951 46580 7960
rect 46635 8000 46677 8009
rect 46635 7960 46636 8000
rect 46676 7960 46677 8000
rect 46635 7951 46677 7960
rect 46732 8000 46772 8035
rect 47116 8000 47156 8009
rect 46636 7866 46676 7951
rect 46732 7949 46772 7960
rect 46924 7960 47116 8000
rect 46924 6656 46964 7960
rect 47116 7951 47156 7960
rect 47211 8000 47253 8009
rect 47211 7960 47212 8000
rect 47252 7960 47253 8000
rect 47211 7951 47253 7960
rect 47212 7866 47252 7951
rect 46924 6607 46964 6616
rect 40780 6437 40820 6448
rect 43371 6488 43413 6497
rect 43371 6448 43372 6488
rect 43412 6448 43413 6488
rect 43371 6439 43413 6448
rect 46347 6488 46389 6497
rect 46347 6448 46348 6488
rect 46388 6448 46389 6488
rect 46347 6439 46389 6448
rect 46444 6488 46484 6497
rect 44619 6236 44661 6245
rect 44619 6196 44620 6236
rect 44660 6196 44661 6236
rect 44619 6187 44661 6196
rect 44620 5900 44660 6187
rect 44620 5851 44660 5860
rect 46348 5900 46388 6439
rect 46444 6329 46484 6448
rect 46731 6488 46773 6497
rect 46731 6448 46732 6488
rect 46772 6448 46773 6488
rect 46731 6439 46773 6448
rect 46732 6354 46772 6439
rect 46443 6320 46485 6329
rect 46443 6280 46444 6320
rect 46484 6280 46485 6320
rect 46443 6271 46485 6280
rect 46348 5851 46388 5860
rect 42604 5648 42644 5657
rect 43468 5648 43508 5657
rect 42644 5608 42740 5648
rect 42604 5599 42644 5608
rect 41067 5564 41109 5573
rect 42220 5564 42260 5573
rect 41067 5524 41068 5564
rect 41108 5524 41109 5564
rect 41067 5515 41109 5524
rect 41740 5524 42220 5564
rect 41068 4976 41108 5515
rect 41548 5144 41588 5172
rect 41740 5144 41780 5524
rect 42220 5515 42260 5524
rect 41588 5104 41780 5144
rect 41548 5095 41588 5104
rect 41068 4927 41108 4936
rect 41356 4976 41396 4985
rect 41164 4388 41204 4397
rect 41356 4388 41396 4936
rect 41204 4348 41396 4388
rect 41164 4339 41204 4348
rect 40683 4136 40725 4145
rect 40683 4096 40684 4136
rect 40724 4096 40725 4136
rect 40683 4087 40725 4096
rect 41067 4136 41109 4145
rect 41067 4096 41068 4136
rect 41108 4096 41109 4136
rect 41067 4087 41109 4096
rect 41259 4136 41301 4145
rect 41259 4096 41260 4136
rect 41300 4096 41301 4136
rect 41259 4087 41301 4096
rect 41643 4136 41685 4145
rect 41643 4096 41644 4136
rect 41684 4096 41685 4136
rect 41643 4087 41685 4096
rect 41068 4002 41108 4087
rect 41260 4002 41300 4087
rect 41644 3632 41684 4087
rect 41684 3592 41876 3632
rect 41644 3583 41684 3592
rect 40780 3464 40820 3473
rect 40972 3464 41012 3473
rect 40492 3424 40780 3464
rect 40492 2876 40532 3424
rect 40780 3415 40820 3424
rect 40876 3424 40972 3464
rect 40492 2827 40532 2836
rect 40684 2876 40724 2885
rect 40876 2876 40916 3424
rect 40972 3415 41012 3424
rect 41836 3380 41876 3592
rect 41836 3331 41876 3340
rect 42027 3212 42069 3221
rect 42027 3172 42028 3212
rect 42068 3172 42069 3212
rect 42027 3163 42069 3172
rect 42028 3078 42068 3163
rect 40724 2836 40916 2876
rect 40684 2827 40724 2836
rect 42700 2717 42740 5608
rect 43083 3212 43125 3221
rect 43083 3172 43084 3212
rect 43124 3172 43125 3212
rect 43083 3163 43125 3172
rect 42699 2708 42741 2717
rect 42699 2668 42700 2708
rect 42740 2668 42741 2708
rect 42699 2659 42741 2668
rect 18019 2562 18059 2571
rect 19180 2540 19220 2575
rect 19180 2491 19220 2500
rect 20907 2540 20949 2549
rect 20907 2500 20908 2540
rect 20948 2500 20949 2540
rect 20907 2491 20949 2500
rect 20908 2406 20948 2491
rect 21292 2490 21332 2575
rect 24460 2540 24500 2549
rect 24652 2540 24692 2549
rect 24500 2500 24652 2540
rect 24460 2491 24500 2500
rect 24652 2491 24692 2500
rect 25036 2490 25076 2575
rect 28012 2540 28052 2549
rect 28204 2540 28244 2549
rect 28052 2500 28204 2540
rect 28012 2491 28052 2500
rect 28204 2491 28244 2500
rect 28588 2490 28628 2575
rect 38476 2573 38516 2584
rect 39339 2624 39381 2633
rect 39339 2584 39340 2624
rect 39380 2584 39381 2624
rect 39339 2575 39381 2584
rect 40203 2624 40245 2633
rect 40203 2584 40204 2624
rect 40244 2584 40245 2624
rect 40203 2575 40245 2584
rect 41835 2624 41877 2633
rect 41835 2584 41836 2624
rect 41876 2584 41877 2624
rect 41835 2575 41877 2584
rect 42700 2624 42740 2659
rect 39340 2490 39380 2575
rect 41836 2490 41876 2575
rect 42700 2574 42740 2584
rect 43084 2624 43124 3163
rect 43468 2633 43508 5608
rect 47499 5648 47541 5657
rect 47499 5608 47500 5648
rect 47540 5608 47541 5648
rect 47499 5599 47541 5608
rect 48364 5648 48404 9472
rect 48460 9463 48500 9472
rect 49324 9512 49364 9631
rect 48472 9092 48840 9101
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48472 9043 48840 9052
rect 48555 8084 48597 8093
rect 48555 8044 48556 8084
rect 48596 8044 48597 8084
rect 48555 8035 48597 8044
rect 48556 7950 48596 8035
rect 49228 8000 49268 8009
rect 48472 7580 48840 7589
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48472 7531 48840 7540
rect 49228 7421 49268 7960
rect 49324 7505 49364 9472
rect 49712 8336 50080 8345
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 49712 8287 50080 8296
rect 49323 7496 49365 7505
rect 49323 7456 49324 7496
rect 49364 7456 49365 7496
rect 49323 7447 49365 7456
rect 51531 7496 51573 7505
rect 51531 7456 51532 7496
rect 51572 7456 51573 7496
rect 51531 7447 51573 7456
rect 49227 7412 49269 7421
rect 49227 7372 49228 7412
rect 49268 7372 49269 7412
rect 49227 7363 49269 7372
rect 49324 7412 49364 7447
rect 49324 7362 49364 7372
rect 50379 7412 50421 7421
rect 50379 7372 50380 7412
rect 50420 7372 50421 7412
rect 50379 7363 50421 7372
rect 50380 7278 50420 7363
rect 49803 7160 49845 7169
rect 49803 7120 49804 7160
rect 49844 7120 49845 7160
rect 49803 7111 49845 7120
rect 51532 7160 51572 7447
rect 52396 7160 52436 10051
rect 53452 9512 53492 10135
rect 55372 10050 55412 10135
rect 55468 10025 55508 10303
rect 54891 10016 54933 10025
rect 54891 9976 54892 10016
rect 54932 9976 54933 10016
rect 54891 9967 54933 9976
rect 55467 10016 55509 10025
rect 55467 9976 55468 10016
rect 55508 9976 55509 10016
rect 55467 9967 55509 9976
rect 53452 9463 53492 9472
rect 54507 9512 54549 9521
rect 54507 9472 54508 9512
rect 54548 9472 54549 9512
rect 54507 9463 54549 9472
rect 53260 9260 53300 9269
rect 53260 7169 53300 9220
rect 54123 9260 54165 9269
rect 54123 9220 54124 9260
rect 54164 9220 54165 9260
rect 54123 9211 54165 9220
rect 54124 8672 54164 9211
rect 54124 8623 54164 8632
rect 54508 8672 54548 9463
rect 54892 9428 54932 9967
rect 55468 9882 55508 9967
rect 55660 9521 55700 12319
rect 59212 11192 59252 14008
rect 59444 14008 60020 14048
rect 59404 13999 59444 14008
rect 59212 11143 59252 11152
rect 58732 11024 58772 11033
rect 58540 10436 58580 10445
rect 58732 10436 58772 10984
rect 59020 11024 59060 11033
rect 58580 10396 58772 10436
rect 58924 10436 58964 10445
rect 59020 10436 59060 10984
rect 59596 11024 59636 11033
rect 59980 11024 60020 14008
rect 60267 14008 60268 14048
rect 60308 14008 60309 14048
rect 60267 13999 60309 14008
rect 60843 14048 60885 14057
rect 60843 14008 60844 14048
rect 60884 14008 60885 14048
rect 60843 13999 60885 14008
rect 60268 13914 60308 13999
rect 59636 10984 59828 11024
rect 59596 10975 59636 10984
rect 58964 10396 59060 10436
rect 59788 10436 59828 10984
rect 58540 10387 58580 10396
rect 58924 10387 58964 10396
rect 59788 10387 59828 10396
rect 59884 10984 59980 11024
rect 55851 10352 55893 10361
rect 55851 10312 55852 10352
rect 55892 10312 55893 10352
rect 55851 10303 55893 10312
rect 58827 10352 58869 10361
rect 58827 10312 58828 10352
rect 58868 10312 58869 10352
rect 58827 10303 58869 10312
rect 55852 10218 55892 10303
rect 56427 10184 56469 10193
rect 56427 10144 56428 10184
rect 56468 10144 56469 10184
rect 56427 10135 56469 10144
rect 56524 10184 56564 10193
rect 58443 10184 58485 10193
rect 56564 10144 56660 10184
rect 56524 10135 56564 10144
rect 55276 9512 55316 9521
rect 55659 9512 55701 9521
rect 55316 9472 55604 9512
rect 55276 9463 55316 9472
rect 54892 9379 54932 9388
rect 54699 9260 54741 9269
rect 54699 9220 54700 9260
rect 54740 9220 54741 9260
rect 54699 9211 54741 9220
rect 54700 9126 54740 9211
rect 55371 8756 55413 8765
rect 55371 8716 55372 8756
rect 55412 8716 55413 8756
rect 55371 8707 55413 8716
rect 54508 8623 54548 8632
rect 55372 8672 55412 8707
rect 51532 7111 51572 7120
rect 52300 7120 52396 7160
rect 48940 7076 48980 7085
rect 48472 6068 48840 6077
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48472 6019 48840 6028
rect 48940 5657 48980 7036
rect 49804 7026 49844 7111
rect 49712 6824 50080 6833
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 49712 6775 50080 6784
rect 47500 5514 47540 5599
rect 45772 3464 45812 3473
rect 45772 2885 45812 3424
rect 46443 3464 46485 3473
rect 46443 3424 46444 3464
rect 46484 3424 46485 3464
rect 46443 3415 46485 3424
rect 46635 3464 46677 3473
rect 46635 3424 46636 3464
rect 46676 3424 46677 3464
rect 46635 3415 46677 3424
rect 46444 3330 46484 3415
rect 46636 3380 46676 3415
rect 46636 3329 46676 3340
rect 46828 3212 46868 3221
rect 47595 3212 47637 3221
rect 46868 3172 47444 3212
rect 46828 3163 46868 3172
rect 45003 2876 45045 2885
rect 45003 2836 45004 2876
rect 45044 2836 45045 2876
rect 45003 2827 45045 2836
rect 45771 2876 45813 2885
rect 45771 2836 45772 2876
rect 45812 2836 45813 2876
rect 45771 2827 45813 2836
rect 45004 2742 45044 2827
rect 43084 2575 43124 2584
rect 43467 2624 43509 2633
rect 43467 2584 43468 2624
rect 43508 2584 43509 2624
rect 43467 2575 43509 2584
rect 46155 2624 46197 2633
rect 46155 2584 46156 2624
rect 46196 2584 46197 2624
rect 46155 2575 46197 2584
rect 47019 2624 47061 2633
rect 47019 2584 47020 2624
rect 47060 2584 47061 2624
rect 47019 2575 47061 2584
rect 47404 2624 47444 3172
rect 47595 3172 47596 3212
rect 47636 3172 47637 3212
rect 47595 3163 47637 3172
rect 47404 2575 47444 2584
rect 47596 2624 47636 3163
rect 48364 2633 48404 5608
rect 48939 5648 48981 5657
rect 48939 5608 48940 5648
rect 48980 5608 48981 5648
rect 48939 5599 48981 5608
rect 48747 5564 48789 5573
rect 48747 5524 48748 5564
rect 48788 5524 48789 5564
rect 48747 5515 48789 5524
rect 48748 5430 48788 5515
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 48747 3632 48789 3641
rect 48747 3592 48748 3632
rect 48788 3592 48789 3632
rect 48747 3583 48789 3592
rect 48748 3380 48788 3583
rect 48748 3331 48788 3340
rect 48556 3221 48596 3306
rect 48555 3212 48597 3221
rect 48555 3172 48556 3212
rect 48596 3172 48597 3212
rect 48555 3163 48597 3172
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 47596 2575 47636 2584
rect 47979 2624 48021 2633
rect 47979 2584 47980 2624
rect 48020 2584 48021 2624
rect 47979 2575 48021 2584
rect 48363 2624 48405 2633
rect 48363 2584 48364 2624
rect 48404 2584 48405 2624
rect 48363 2575 48405 2584
rect 48844 2624 48884 2633
rect 48940 2624 48980 5599
rect 49035 5564 49077 5573
rect 49035 5524 49036 5564
rect 49076 5524 49077 5564
rect 49035 5515 49077 5524
rect 49036 4052 49076 5515
rect 52107 5480 52149 5489
rect 52107 5440 52108 5480
rect 52148 5440 52149 5480
rect 52107 5431 52149 5440
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 52108 5153 52148 5431
rect 49323 5144 49365 5153
rect 49323 5104 49324 5144
rect 49364 5104 49365 5144
rect 49323 5095 49365 5104
rect 50091 5144 50133 5153
rect 50091 5104 50092 5144
rect 50132 5104 50133 5144
rect 50091 5095 50133 5104
rect 52107 5144 52149 5153
rect 52107 5104 52108 5144
rect 52148 5104 52149 5144
rect 52107 5095 52149 5104
rect 49228 4136 49268 4145
rect 49132 4052 49172 4061
rect 49036 4012 49132 4052
rect 49132 4003 49172 4012
rect 49228 3548 49268 4096
rect 49228 3499 49268 3508
rect 49131 3464 49173 3473
rect 49131 3424 49132 3464
rect 49172 3424 49173 3464
rect 49131 3415 49173 3424
rect 49324 3464 49364 5095
rect 50092 5010 50132 5095
rect 50379 5060 50421 5069
rect 50379 5020 50380 5060
rect 50420 5020 50421 5060
rect 50379 5011 50421 5020
rect 50188 4976 50228 4985
rect 49611 4136 49653 4145
rect 49611 4096 49612 4136
rect 49652 4096 49653 4136
rect 49611 4087 49653 4096
rect 49612 4002 49652 4087
rect 50188 3884 50228 4936
rect 50380 4926 50420 5011
rect 51916 4976 51956 4985
rect 51916 4388 51956 4936
rect 51916 4339 51956 4348
rect 52108 4220 52148 5095
rect 52108 4171 52148 4180
rect 52300 4976 52340 7120
rect 52396 7111 52436 7120
rect 53259 7160 53301 7169
rect 53259 7120 53260 7160
rect 53300 7120 53301 7160
rect 53259 7111 53301 7120
rect 52780 7076 52820 7085
rect 52780 5069 52820 7036
rect 54028 5648 54068 5657
rect 54068 5608 54356 5648
rect 54028 5599 54068 5608
rect 53355 5480 53397 5489
rect 53355 5440 53356 5480
rect 53396 5440 53397 5480
rect 53355 5431 53397 5440
rect 53356 5346 53396 5431
rect 52779 5060 52821 5069
rect 52779 5020 52780 5060
rect 52820 5020 52821 5060
rect 52779 5011 52821 5020
rect 50475 4136 50517 4145
rect 50475 4096 50476 4136
rect 50516 4096 50517 4136
rect 50475 4087 50517 4096
rect 50188 3844 50419 3884
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 50379 3641 50419 3844
rect 49515 3632 49557 3641
rect 49515 3592 49516 3632
rect 49556 3592 49557 3632
rect 49515 3583 49557 3592
rect 50378 3632 50420 3641
rect 50378 3592 50379 3632
rect 50419 3592 50420 3632
rect 50378 3583 50420 3592
rect 49516 3498 49556 3583
rect 50379 3485 50419 3583
rect 50476 3548 50516 4087
rect 50476 3499 50516 3508
rect 50188 3464 50228 3473
rect 49324 3415 49364 3424
rect 49996 3424 50188 3464
rect 50379 3436 50419 3445
rect 50572 3464 50612 3473
rect 49132 3330 49172 3415
rect 49996 2876 50036 3424
rect 50188 3415 50228 3424
rect 49996 2827 50036 2836
rect 50572 2717 50612 3424
rect 52012 2792 52052 2801
rect 52052 2752 52244 2792
rect 52012 2743 52052 2752
rect 50571 2708 50613 2717
rect 50571 2668 50572 2708
rect 50612 2668 50613 2708
rect 50571 2659 50613 2668
rect 51819 2708 51861 2717
rect 51819 2668 51820 2708
rect 51860 2668 51861 2708
rect 51819 2659 51861 2668
rect 48884 2584 48980 2624
rect 48844 2575 48884 2584
rect 46156 2490 46196 2575
rect 47020 2490 47060 2575
rect 47980 2490 48020 2575
rect 51820 2574 51860 2659
rect 52204 2624 52244 2752
rect 52300 2624 52340 4936
rect 53163 4976 53205 4985
rect 53163 4936 53164 4976
rect 53204 4936 53205 4976
rect 53163 4927 53205 4936
rect 53451 4976 53493 4985
rect 53451 4936 53452 4976
rect 53492 4936 53493 4976
rect 53451 4927 53493 4936
rect 53164 4842 53204 4927
rect 53356 3212 53396 3221
rect 53356 2717 53396 3172
rect 53355 2708 53397 2717
rect 53355 2668 53356 2708
rect 53396 2668 53397 2708
rect 53355 2659 53397 2668
rect 52588 2624 52628 2633
rect 52300 2584 52588 2624
rect 52204 2575 52244 2584
rect 52588 2575 52628 2584
rect 53452 2624 53492 4927
rect 54316 4892 54356 5608
rect 55372 4985 55412 8632
rect 55564 8168 55604 9472
rect 55659 9472 55660 9512
rect 55700 9472 55701 9512
rect 55659 9463 55701 9472
rect 55660 9378 55700 9463
rect 56428 8849 56468 10135
rect 56524 9512 56564 9521
rect 55755 8840 55797 8849
rect 55755 8800 55756 8840
rect 55796 8800 55797 8840
rect 55755 8791 55797 8800
rect 56427 8840 56469 8849
rect 56427 8800 56428 8840
rect 56468 8800 56469 8840
rect 56427 8791 56469 8800
rect 55564 8119 55604 8128
rect 55756 7916 55796 8791
rect 56524 8765 56564 9472
rect 56523 8756 56565 8765
rect 56523 8716 56524 8756
rect 56564 8716 56565 8756
rect 56523 8707 56565 8716
rect 56524 8504 56564 8513
rect 56620 8504 56660 10144
rect 58443 10144 58444 10184
rect 58484 10144 58485 10184
rect 58443 10135 58485 10144
rect 58635 10184 58677 10193
rect 58635 10144 58636 10184
rect 58676 10144 58677 10184
rect 58635 10135 58677 10144
rect 58828 10184 58868 10303
rect 58828 10135 58868 10144
rect 59019 10184 59061 10193
rect 59019 10144 59020 10184
rect 59060 10144 59061 10184
rect 59019 10135 59061 10144
rect 58444 10050 58484 10135
rect 58636 10050 58676 10135
rect 59020 10050 59060 10135
rect 59211 10100 59253 10109
rect 59211 10060 59212 10100
rect 59252 10060 59253 10100
rect 59211 10051 59253 10060
rect 59212 9428 59252 10051
rect 59404 9680 59444 9689
rect 59444 9640 59636 9680
rect 59404 9631 59444 9640
rect 59596 9596 59636 9640
rect 59596 9547 59636 9556
rect 59884 9521 59924 10984
rect 59980 10975 60020 10984
rect 60844 11024 60884 13999
rect 63592 13628 63960 13637
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63592 13579 63960 13588
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 93832 13628 94200 13637
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 93832 13579 94200 13588
rect 64832 12872 65200 12881
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 64832 12823 65200 12832
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 95072 12872 95440 12881
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95072 12823 95440 12832
rect 63592 12116 63960 12125
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63592 12067 63960 12076
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 93832 12116 94200 12125
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 93832 12067 94200 12076
rect 61804 11696 61844 11705
rect 61844 11656 62036 11696
rect 61804 11647 61844 11656
rect 60844 10975 60884 10984
rect 61132 11528 61172 11537
rect 61132 10277 61172 11488
rect 61996 11192 62036 11656
rect 64832 11360 65200 11369
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 64832 11311 65200 11320
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 95072 11360 95440 11369
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95072 11311 95440 11320
rect 61996 11143 62036 11152
rect 63592 10604 63960 10613
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63592 10555 63960 10564
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 93832 10604 94200 10613
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 93832 10555 94200 10564
rect 59979 10268 60021 10277
rect 59979 10228 59980 10268
rect 60020 10228 60021 10268
rect 59979 10219 60021 10228
rect 61131 10268 61173 10277
rect 61131 10228 61132 10268
rect 61172 10228 61173 10268
rect 61131 10219 61173 10228
rect 59980 10134 60020 10219
rect 61419 10184 61461 10193
rect 61419 10144 61420 10184
rect 61460 10144 61461 10184
rect 61419 10135 61461 10144
rect 61995 10184 62037 10193
rect 61995 10144 61996 10184
rect 62036 10144 62037 10184
rect 61995 10135 62037 10144
rect 60747 10100 60789 10109
rect 60747 10060 60748 10100
rect 60788 10060 60789 10100
rect 60747 10051 60789 10060
rect 60748 9966 60788 10051
rect 61420 10050 61460 10135
rect 61996 9680 62036 10135
rect 64832 9848 65200 9857
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 64832 9799 65200 9808
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 95072 9848 95440 9857
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95072 9799 95440 9808
rect 61996 9631 62036 9640
rect 59883 9512 59925 9521
rect 59980 9512 60020 9521
rect 59883 9472 59884 9512
rect 59924 9472 59980 9512
rect 59883 9463 59925 9472
rect 59980 9463 60020 9472
rect 60844 9512 60884 9521
rect 59212 9379 59252 9388
rect 59884 9378 59924 9463
rect 57676 9260 57716 9269
rect 57484 9220 57676 9260
rect 56811 8840 56853 8849
rect 56811 8800 56812 8840
rect 56852 8800 56853 8840
rect 56811 8791 56853 8800
rect 56715 8756 56757 8765
rect 56715 8716 56716 8756
rect 56756 8716 56757 8756
rect 56715 8707 56757 8716
rect 56564 8464 56660 8504
rect 56524 8455 56564 8464
rect 55756 7867 55796 7876
rect 56716 7412 56756 8707
rect 56812 8706 56852 8791
rect 57484 8672 57524 9220
rect 57676 9211 57716 9220
rect 60844 8765 60884 9472
rect 63592 9092 63960 9101
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63592 9043 63960 9052
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 93832 9092 94200 9101
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 93832 9043 94200 9052
rect 60843 8756 60885 8765
rect 60843 8716 60844 8756
rect 60884 8716 60885 8756
rect 60843 8707 60885 8716
rect 57484 8623 57524 8632
rect 64832 8336 65200 8345
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 64832 8287 65200 8296
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 95072 8336 95440 8345
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95072 8287 95440 8296
rect 63592 7580 63960 7589
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63592 7531 63960 7540
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 93832 7580 94200 7589
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 93832 7531 94200 7540
rect 56716 7363 56756 7372
rect 56427 7160 56469 7169
rect 56427 7120 56428 7160
rect 56468 7120 56469 7160
rect 56427 7111 56469 7120
rect 56428 7026 56468 7111
rect 64832 6824 65200 6833
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 64832 6775 65200 6784
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 95072 6824 95440 6833
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95072 6775 95440 6784
rect 63592 6068 63960 6077
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63592 6019 63960 6028
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 93832 6068 94200 6077
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 93832 6019 94200 6028
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 95072 5312 95440 5321
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95072 5263 95440 5272
rect 55371 4976 55413 4985
rect 55371 4936 55372 4976
rect 55412 4936 55413 4976
rect 55371 4927 55413 4936
rect 54316 4843 54356 4852
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 93832 4556 94200 4565
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 93832 4507 94200 4516
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 95072 3800 95440 3809
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95072 3751 95440 3760
rect 54028 3464 54068 3473
rect 54028 2885 54068 3424
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 93832 3044 94200 3053
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 93832 2995 94200 3004
rect 54027 2876 54069 2885
rect 54027 2836 54028 2876
rect 54068 2836 54069 2876
rect 54027 2827 54069 2836
rect 54603 2876 54645 2885
rect 54603 2836 54604 2876
rect 54644 2836 54645 2876
rect 54603 2827 54645 2836
rect 54604 2742 54644 2827
rect 53452 2575 53492 2584
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 95072 2288 95440 2297
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95072 2239 95440 2248
rect 13556 1828 13652 1868
rect 13516 1819 13556 1828
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 93832 1532 94200 1541
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 93832 1483 94200 1492
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
rect 95072 776 95440 785
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95072 727 95440 736
<< via2 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 20620 37528 20660 37568
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 76 36688 116 36728
rect 5836 36604 5876 36644
rect 4684 36520 4724 36560
rect 5644 36520 5684 36560
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 6604 36520 6644 36560
rect 7372 36520 7412 36560
rect 5068 35848 5108 35888
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 5068 35176 5108 35216
rect 4300 34336 4340 34376
rect 4972 34336 5012 34376
rect 5836 35176 5876 35216
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 9100 35848 9140 35888
rect 8716 35764 8756 35804
rect 7372 35260 7412 35300
rect 8428 35260 8468 35300
rect 7468 35176 7508 35216
rect 7948 35176 7988 35216
rect 8044 35092 8084 35132
rect 8236 34168 8276 34208
rect 8812 34168 8852 34208
rect 4108 32740 4148 32780
rect 5932 32740 5972 32780
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 2860 30640 2900 30680
rect 7468 32824 7508 32864
rect 6508 32656 6548 32696
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 18316 37276 18356 37316
rect 10348 36856 10388 36896
rect 11788 36856 11828 36896
rect 9772 35848 9812 35888
rect 9964 35848 10004 35888
rect 19276 37276 19316 37316
rect 18796 36688 18836 36728
rect 18700 36520 18740 36560
rect 19180 36520 19220 36560
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 19852 36688 19892 36728
rect 20044 35932 20084 35972
rect 9292 35764 9332 35804
rect 10348 35680 10388 35720
rect 9292 35092 9332 35132
rect 9676 35092 9716 35132
rect 9676 33664 9716 33704
rect 19468 35848 19508 35888
rect 11980 35680 12020 35720
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 16876 34420 16916 34460
rect 17740 34420 17780 34460
rect 14476 34252 14516 34292
rect 11116 33664 11156 33704
rect 10060 33496 10100 33536
rect 10732 33496 10772 33536
rect 11404 33496 11444 33536
rect 6988 32152 7028 32192
rect 9676 32824 9716 32864
rect 15436 34252 15476 34292
rect 14956 33076 14996 33116
rect 12076 32824 12116 32864
rect 9196 31480 9236 31520
rect 4876 31144 4916 31184
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 3916 30640 3956 30680
rect 3244 30556 3284 30596
rect 3628 30556 3668 30596
rect 3820 30556 3860 30596
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 3724 29884 3764 29924
rect 8236 30556 8276 30596
rect 4108 29968 4148 30008
rect 5068 29968 5108 30008
rect 5452 29968 5492 30008
rect 4588 29884 4628 29924
rect 4972 29884 5012 29924
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 4972 27868 5012 27908
rect 4396 27784 4436 27824
rect 4684 27784 4724 27824
rect 4300 27700 4340 27740
rect 3820 27616 3860 27656
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 3436 26860 3476 26900
rect 4588 27616 4628 27656
rect 5932 29128 5972 29168
rect 7852 29128 7892 29168
rect 15724 34168 15764 34208
rect 16204 34168 16244 34208
rect 15916 33076 15956 33116
rect 20332 34168 20372 34208
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 15628 32908 15668 32948
rect 15628 32740 15668 32780
rect 10060 32152 10100 32192
rect 11212 31900 11252 31940
rect 10156 29800 10196 29840
rect 5740 27784 5780 27824
rect 5452 27700 5492 27740
rect 8236 29044 8276 29084
rect 5068 27448 5108 27488
rect 5260 27364 5300 27404
rect 7084 27364 7124 27404
rect 4204 26860 4244 26900
rect 2476 26608 2516 26648
rect 2380 26440 2420 26480
rect 3628 26608 3668 26648
rect 3244 26440 3284 26480
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 2860 26104 2900 26144
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 4876 26440 4916 26480
rect 5740 26440 5780 26480
rect 6796 26440 6836 26480
rect 6124 25516 6164 25556
rect 3724 25264 3764 25304
rect 5068 25264 5108 25304
rect 5836 25264 5876 25304
rect 7468 26104 7508 26144
rect 8332 25516 8372 25556
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 1228 23080 1268 23120
rect 2092 23080 2132 23120
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 4492 22996 4532 23036
rect 2764 22828 2804 22868
rect 2956 22828 2996 22868
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 2668 22324 2708 22364
rect 3244 22324 3284 22364
rect 2380 22240 2420 22280
rect 3724 22324 3764 22364
rect 652 21568 692 21608
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 652 20728 692 20768
rect 76 20056 116 20096
rect 652 19888 692 19928
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 4108 22660 4148 22700
rect 4204 22324 4244 22364
rect 11020 29128 11060 29168
rect 9772 27616 9812 27656
rect 10156 27616 10196 27656
rect 9580 26776 9620 26816
rect 10156 26776 10196 26816
rect 11788 31900 11828 31940
rect 12076 31480 12116 31520
rect 11884 29128 11924 29168
rect 9484 26440 9524 26480
rect 11884 26440 11924 26480
rect 11692 26188 11732 26228
rect 11788 25264 11828 25304
rect 14380 30388 14420 30428
rect 15436 30640 15476 30680
rect 15244 30388 15284 30428
rect 17068 32908 17108 32948
rect 16108 32152 16148 32192
rect 17164 32152 17204 32192
rect 17068 31900 17108 31940
rect 17740 31900 17780 31940
rect 17164 31564 17204 31604
rect 16204 30640 16244 30680
rect 16396 30220 16436 30260
rect 15052 29128 15092 29168
rect 15244 29044 15284 29084
rect 12268 26188 12308 26228
rect 12076 25264 12116 25304
rect 14092 24676 14132 24716
rect 13804 24592 13844 24632
rect 15244 24592 15284 24632
rect 9100 24424 9140 24464
rect 12172 24424 12212 24464
rect 14860 24424 14900 24464
rect 5452 22996 5492 23036
rect 5068 22240 5108 22280
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 8428 21568 8468 21608
rect 9964 22240 10004 22280
rect 9484 21568 9524 21608
rect 10444 21568 10484 21608
rect 11020 21568 11060 21608
rect 11788 21568 11828 21608
rect 12268 21568 12308 21608
rect 13036 21568 13076 21608
rect 5836 20980 5876 21020
rect 8044 20980 8084 21020
rect 4780 20140 4820 20180
rect 5164 20140 5204 20180
rect 2668 19468 2708 19508
rect 3724 19468 3764 19508
rect 652 19048 692 19088
rect 2284 19048 2324 19088
rect 3148 19300 3188 19340
rect 2764 19216 2804 19256
rect 652 18208 692 18248
rect 652 17368 692 17408
rect 2188 17200 2228 17240
rect 652 16528 692 16568
rect 556 15688 596 15728
rect 652 14848 692 14888
rect 3436 19216 3476 19256
rect 2956 19048 2996 19088
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 3436 17704 3476 17744
rect 3052 17200 3092 17240
rect 4588 19972 4628 20012
rect 4876 19972 4916 20012
rect 4684 19384 4724 19424
rect 5260 19300 5300 19340
rect 4396 19048 4436 19088
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 5548 19300 5588 19340
rect 5356 19216 5396 19256
rect 7372 19216 7412 19256
rect 7756 19048 7796 19088
rect 11404 20728 11444 20768
rect 12172 20728 12212 20768
rect 14764 22240 14804 22280
rect 15820 29128 15860 29168
rect 17068 30640 17108 30680
rect 17260 30640 17300 30680
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 20524 32824 20564 32864
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 18124 31564 18164 31604
rect 18316 31564 18356 31604
rect 17932 30724 17972 30764
rect 18220 30640 18260 30680
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 20140 30724 20180 30764
rect 17260 30220 17300 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 20524 29968 20564 30008
rect 18700 29884 18740 29924
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 16684 29128 16724 29168
rect 19276 29128 19316 29168
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 23980 36520 24020 36560
rect 22156 35932 22196 35972
rect 21292 35848 21332 35888
rect 21484 35848 21524 35888
rect 23212 35848 23252 35888
rect 22348 35260 22388 35300
rect 23020 34168 23060 34208
rect 20812 34000 20852 34040
rect 22348 34000 22388 34040
rect 22156 32824 22196 32864
rect 24940 36688 24980 36728
rect 24940 36520 24980 36560
rect 25804 36520 25844 36560
rect 24748 35848 24788 35888
rect 35596 37360 35636 37400
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 30220 36520 30260 36560
rect 31180 36520 31220 36560
rect 31372 36520 31412 36560
rect 32140 36520 32180 36560
rect 24844 35260 24884 35300
rect 24556 34000 24596 34040
rect 24268 33664 24308 33704
rect 25228 35848 25268 35888
rect 33100 36520 33140 36560
rect 25324 35260 25364 35300
rect 26188 35260 26228 35300
rect 25036 33664 25076 33704
rect 23980 32824 24020 32864
rect 25036 32824 25076 32864
rect 30316 34924 30356 34964
rect 31468 35092 31508 35132
rect 31276 34924 31316 34964
rect 30700 34336 30740 34376
rect 32236 35092 32276 35132
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 36460 36688 36500 36728
rect 35404 36184 35444 36224
rect 36076 36184 36116 36224
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 33196 35176 33236 35216
rect 33292 35092 33332 35132
rect 33772 35092 33812 35132
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 25996 32908 26036 32948
rect 22540 30808 22580 30848
rect 21196 29968 21236 30008
rect 20812 29884 20852 29924
rect 24364 31144 24404 31184
rect 25708 31144 25748 31184
rect 23884 30808 23924 30848
rect 25324 30724 25364 30764
rect 25612 30724 25652 30764
rect 25228 30640 25268 30680
rect 23212 30052 23252 30092
rect 24268 30052 24308 30092
rect 25324 30052 25364 30092
rect 22636 29800 22676 29840
rect 25804 30640 25844 30680
rect 26860 32824 26900 32864
rect 28588 32824 28628 32864
rect 27628 32656 27668 32696
rect 28012 32656 28052 32696
rect 26956 30724 26996 30764
rect 26092 30556 26132 30596
rect 26764 30556 26804 30596
rect 27052 29800 27092 29840
rect 27724 29800 27764 29840
rect 28972 29800 29012 29840
rect 32428 34336 32468 34376
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 36940 37360 36980 37400
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 37804 36688 37844 36728
rect 38572 36688 38612 36728
rect 36940 36604 36980 36644
rect 37708 36604 37748 36644
rect 37516 36520 37556 36560
rect 36652 36184 36692 36224
rect 36268 35932 36308 35972
rect 36652 35932 36691 35972
rect 36691 35932 36692 35972
rect 36844 35932 36884 35972
rect 35788 35176 35828 35216
rect 33868 34336 33908 34376
rect 35404 34336 35444 34376
rect 36268 34336 36308 34376
rect 37324 34336 37364 34376
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 34252 32236 34292 32276
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 33772 31480 33812 31520
rect 34252 31480 34292 31520
rect 32428 31312 32468 31352
rect 33100 31312 33140 31352
rect 31564 30640 31604 30680
rect 32812 30724 32852 30764
rect 33772 30640 33812 30680
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 22636 29212 22676 29252
rect 21388 29128 21428 29168
rect 22060 29128 22100 29168
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 19084 26104 19124 26144
rect 20620 28288 20660 28328
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 16876 25516 16916 25556
rect 17836 25516 17876 25556
rect 15916 24424 15956 24464
rect 15916 23752 15956 23792
rect 15436 23668 15476 23708
rect 16012 22492 16052 22532
rect 14764 21988 14804 22028
rect 15340 21988 15380 22028
rect 15724 21568 15764 21608
rect 13996 21400 14036 21440
rect 15244 21400 15284 21440
rect 9484 19132 9524 19172
rect 8620 17788 8660 17828
rect 4204 17704 4244 17744
rect 9772 19048 9812 19088
rect 10732 19048 10772 19088
rect 16396 24592 16436 24632
rect 17068 24424 17108 24464
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 23116 29128 23156 29168
rect 22636 29044 22676 29084
rect 24268 28960 24308 29000
rect 22156 28288 22196 28328
rect 23980 28120 24020 28160
rect 21100 25264 21140 25304
rect 21772 25264 21812 25304
rect 23596 26104 23636 26144
rect 22732 25432 22772 25472
rect 20908 24676 20948 24716
rect 17068 23752 17108 23792
rect 17644 23752 17684 23792
rect 18316 23752 18356 23792
rect 19084 23752 19124 23792
rect 20332 23836 20372 23876
rect 16204 23668 16244 23708
rect 16204 22492 16244 22532
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 20044 21988 20084 22028
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 17644 21568 17684 21608
rect 19948 21316 19988 21356
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 9868 17788 9908 17828
rect 10828 17788 10868 17828
rect 3244 16948 3284 16988
rect 4012 16948 4052 16988
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 4012 14512 4052 14552
rect 2956 14092 2996 14132
rect 3820 14092 3860 14132
rect 652 14008 692 14048
rect 2764 14008 2804 14048
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 4492 14512 4532 14552
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 3340 14008 3380 14048
rect 4204 14008 4244 14048
rect 5836 14008 5876 14048
rect 4396 13924 4436 13964
rect 5740 13924 5780 13964
rect 4012 13840 4052 13880
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 652 13168 692 13208
rect 5548 13840 5588 13880
rect 7276 14512 7316 14552
rect 7180 14092 7220 14132
rect 14860 17872 14900 17912
rect 11980 17620 12020 17660
rect 12844 17620 12884 17660
rect 8908 14680 8948 14720
rect 9100 14680 9140 14720
rect 8812 14512 8852 14552
rect 8044 14092 8084 14132
rect 8428 14092 8468 14132
rect 9196 14092 9236 14132
rect 6892 13924 6932 13964
rect 7084 13924 7124 13964
rect 6412 13840 6452 13880
rect 9004 13840 9044 13880
rect 5260 13168 5300 13208
rect 5836 13168 5876 13208
rect 8044 13168 8084 13208
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 652 12328 692 12368
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 652 11488 692 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 652 10648 692 10688
rect 844 10648 884 10688
rect 652 9808 692 9848
rect 652 8968 692 9008
rect 556 8128 596 8168
rect 652 7288 692 7328
rect 652 6448 692 6488
rect 652 5608 692 5648
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 2284 10312 2324 10352
rect 3148 10312 3188 10352
rect 3340 10228 3380 10268
rect 4108 10228 4148 10268
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 2764 5608 2804 5648
rect 2476 4936 2516 4976
rect 3532 8632 3572 8672
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 6124 9472 6164 9512
rect 6796 9472 6836 9512
rect 4204 8632 4244 8672
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 4492 7960 4532 8000
rect 6604 8632 6644 8672
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 4588 6616 4628 6656
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 5932 7960 5972 8000
rect 5644 6616 5684 6656
rect 2956 5608 2996 5648
rect 4492 5608 4532 5648
rect 4780 5608 4820 5648
rect 5164 5608 5204 5648
rect 5068 5440 5108 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 2860 4852 2900 4892
rect 3340 4852 3380 4892
rect 652 4768 692 4808
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 4300 4852 4340 4892
rect 844 4180 884 4220
rect 5548 5440 5588 5480
rect 5356 5020 5396 5060
rect 5164 4936 5204 4976
rect 9292 14008 9332 14048
rect 9580 14008 9620 14048
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 20332 21316 20372 21356
rect 20812 23836 20852 23876
rect 21100 24592 21140 24632
rect 21484 24592 21524 24632
rect 21004 24340 21044 24380
rect 21964 24340 22004 24380
rect 21004 23836 21044 23876
rect 21964 20560 22004 20600
rect 26476 28120 26516 28160
rect 27148 28372 27188 28412
rect 28780 28372 28820 28412
rect 28876 28288 28916 28328
rect 26188 27700 26228 27740
rect 26764 27700 26804 27740
rect 26572 26524 26612 26564
rect 26092 26104 26132 26144
rect 24556 25432 24596 25472
rect 22924 24676 22964 24716
rect 27148 25852 27188 25892
rect 26092 24676 26132 24716
rect 26764 24676 26804 24716
rect 23596 24592 23636 24632
rect 25228 24592 25268 24632
rect 25900 24592 25940 24632
rect 24748 24508 24788 24548
rect 28876 26776 28916 26816
rect 28684 26692 28724 26732
rect 28876 26524 28916 26564
rect 27724 25852 27764 25892
rect 31564 29128 31604 29168
rect 29068 28288 29108 28328
rect 29164 26776 29204 26816
rect 30604 26608 30644 26648
rect 29644 25264 29684 25304
rect 26956 24592 26996 24632
rect 27436 24592 27476 24632
rect 25708 22156 25748 22196
rect 25804 21568 25844 21608
rect 26476 22156 26516 22196
rect 26860 21568 26900 21608
rect 27052 21568 27092 21608
rect 22252 20056 22292 20096
rect 22732 20056 22772 20096
rect 20332 19972 20372 20012
rect 21388 19972 21428 20012
rect 25228 19972 25268 20012
rect 26668 19972 26708 20012
rect 20428 19804 20468 19844
rect 20812 19804 20852 19844
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 15820 17872 15860 17912
rect 16012 17620 16052 17660
rect 16780 17620 16820 17660
rect 17548 17620 17588 17660
rect 14956 16360 14996 16400
rect 15820 16360 15860 16400
rect 14956 16192 14996 16232
rect 15244 16192 15284 16232
rect 10636 14680 10676 14720
rect 14572 15688 14612 15728
rect 15628 15688 15668 15728
rect 16972 15520 17012 15560
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 20140 16360 20180 16400
rect 18028 16276 18068 16316
rect 18508 16276 18548 16316
rect 19468 16276 19508 16316
rect 20044 16276 20084 16316
rect 15820 15436 15860 15476
rect 17548 15352 17588 15392
rect 11308 14176 11348 14216
rect 11884 14176 11924 14216
rect 10252 13840 10292 13880
rect 12076 14008 12116 14048
rect 12268 14008 12308 14048
rect 12748 14008 12788 14048
rect 9484 12496 9524 12536
rect 10252 12496 10292 12536
rect 19276 16192 19316 16232
rect 18796 15940 18836 15980
rect 18700 15604 18740 15644
rect 17836 15436 17876 15476
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 18796 15520 18836 15560
rect 18508 15352 18548 15392
rect 18700 15352 18740 15392
rect 17644 15268 17684 15308
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 18124 14512 18164 14552
rect 17548 13924 17588 13964
rect 17260 13168 17300 13208
rect 18508 13924 18548 13964
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 18700 12412 18740 12452
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 9196 9640 9236 9680
rect 12748 10228 12788 10268
rect 10732 10060 10772 10100
rect 12652 10060 12692 10100
rect 9868 9640 9908 9680
rect 16492 10984 16532 11024
rect 13132 10228 13172 10268
rect 7564 7960 7604 8000
rect 9580 7960 9620 8000
rect 11212 7960 11252 8000
rect 11020 7372 11060 7412
rect 7180 6364 7220 6404
rect 10156 6364 10196 6404
rect 7372 6280 7412 6320
rect 6988 5020 7028 5060
rect 6892 4936 6932 4976
rect 8236 4936 8276 4976
rect 7372 4852 7412 4892
rect 9772 6196 9812 6236
rect 10348 6280 10388 6320
rect 11500 7372 11540 7412
rect 12172 7120 12212 7160
rect 12172 6364 12212 6404
rect 14188 10144 14228 10184
rect 16492 10144 16532 10184
rect 13324 10060 13364 10100
rect 17548 10984 17588 11024
rect 19948 15352 19988 15392
rect 20332 15940 20372 15980
rect 20140 15016 20180 15056
rect 20428 15016 20468 15056
rect 20236 14680 20276 14720
rect 20140 14512 20180 14552
rect 21292 16360 21332 16400
rect 26860 18376 26900 18416
rect 26188 18292 26228 18332
rect 25708 17704 25748 17744
rect 25228 17620 25268 17660
rect 22444 15520 22484 15560
rect 22636 15520 22676 15560
rect 22924 15520 22964 15560
rect 21292 14680 21332 14720
rect 20812 14428 20852 14468
rect 21292 14428 21332 14468
rect 21676 14428 21716 14468
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 18988 13168 19028 13208
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 18988 12580 19028 12620
rect 21292 12580 21332 12620
rect 19372 12496 19412 12536
rect 21676 12496 21716 12536
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 21100 11320 21140 11360
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 18124 10228 18164 10268
rect 16684 10060 16724 10100
rect 17068 10060 17108 10100
rect 14764 7960 14804 8000
rect 15820 7960 15860 8000
rect 13516 7120 13556 7160
rect 12172 5692 12212 5732
rect 13036 5692 13076 5732
rect 12940 4180 12980 4220
rect 652 3928 692 3968
rect 11788 3928 11828 3968
rect 12748 3928 12788 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 12172 3424 12212 3464
rect 12652 3424 12692 3464
rect 844 3340 884 3380
rect 652 3172 692 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 844 2668 884 2708
rect 13132 3424 13172 3464
rect 17644 6196 17684 6236
rect 16780 5692 16820 5732
rect 17068 5692 17108 5732
rect 14188 4096 14228 4136
rect 16300 4096 16340 4136
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 19084 8800 19124 8840
rect 20332 8800 20372 8840
rect 21004 10144 21044 10184
rect 21772 12244 21812 12284
rect 21676 10984 21716 11024
rect 21484 10144 21524 10184
rect 21580 9472 21620 9512
rect 20620 8632 20660 8672
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 18700 7960 18740 8000
rect 18124 7624 18164 7664
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 18124 6196 18164 6236
rect 17932 5608 17972 5648
rect 16972 4180 17012 4220
rect 17644 4096 17684 4136
rect 17548 3963 17588 3968
rect 17548 3928 17588 3963
rect 17644 3844 17684 3884
rect 17548 3760 17588 3800
rect 17548 3424 17588 3464
rect 16300 2836 16340 2876
rect 16876 2836 16916 2876
rect 13612 2584 13652 2624
rect 17548 2752 17588 2792
rect 15532 2584 15572 2624
rect 17452 2584 17492 2624
rect 17836 3928 17876 3968
rect 18028 4012 18068 4052
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 19948 7624 19988 7664
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 18700 5692 18740 5732
rect 19660 5608 19700 5648
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 17932 3760 17972 3800
rect 19372 3928 19412 3968
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 21964 10396 22004 10436
rect 21868 10144 21908 10184
rect 22540 15016 22580 15056
rect 23692 14512 23732 14552
rect 23020 12580 23060 12620
rect 22732 12496 22772 12536
rect 23020 12412 23060 12452
rect 23692 13000 23732 13040
rect 23308 12496 23348 12536
rect 23884 12664 23924 12704
rect 23788 12580 23828 12620
rect 26092 17620 26132 17660
rect 28204 21484 28244 21524
rect 30604 25264 30644 25304
rect 30220 24340 30260 24380
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 32524 26776 32564 26816
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 37228 32152 37268 32192
rect 38956 36520 38996 36560
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 37708 32236 37748 32276
rect 36268 32068 36308 32108
rect 36940 32068 36980 32108
rect 37612 32068 37652 32108
rect 37324 31900 37364 31940
rect 37996 32152 38036 32192
rect 36172 31396 36212 31436
rect 34636 30808 34676 30848
rect 35116 30808 35156 30848
rect 35980 30808 36020 30848
rect 35500 30724 35540 30764
rect 35788 30724 35828 30764
rect 34156 30640 34196 30680
rect 35116 30640 35156 30680
rect 35596 30640 35636 30680
rect 37420 31312 37460 31352
rect 37612 30808 37652 30848
rect 37132 30724 37172 30764
rect 34060 30220 34100 30260
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 33196 26776 33236 26816
rect 32908 26524 32948 26564
rect 33580 26440 33620 26480
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 31564 24592 31604 24632
rect 32044 24592 32084 24632
rect 35308 26776 35348 26816
rect 34444 26608 34484 26648
rect 34924 26608 34964 26648
rect 35116 26608 35156 26648
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 36460 30640 36500 30680
rect 38284 32152 38324 32192
rect 38476 31396 38516 31436
rect 38860 32236 38900 32276
rect 38764 31900 38804 31940
rect 38572 31312 38612 31352
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 45676 33412 45716 33452
rect 46828 33412 46868 33452
rect 42508 32992 42548 33032
rect 43372 32992 43412 33032
rect 39916 32236 39956 32276
rect 43564 32908 43604 32948
rect 44332 32908 44372 32948
rect 39724 32152 39764 32192
rect 40396 32152 40436 32192
rect 42892 31564 42932 31604
rect 41836 30724 41876 30764
rect 38380 30640 38420 30680
rect 39916 30220 39956 30260
rect 38092 29800 38132 29840
rect 39628 29800 39668 29840
rect 40204 27700 40244 27740
rect 39628 27616 39668 27656
rect 40300 27616 40340 27656
rect 40684 30220 40724 30260
rect 41452 30220 41492 30260
rect 39628 26776 39668 26816
rect 38476 26692 38516 26732
rect 40300 26692 40340 26732
rect 36460 26608 36500 26648
rect 44524 31480 44564 31520
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 45196 31564 45236 31604
rect 44332 30640 44372 30680
rect 43756 29800 43796 29840
rect 44524 29800 44564 29840
rect 40876 29548 40916 29588
rect 42892 29548 42932 29588
rect 40972 28288 41012 28328
rect 43948 28288 43988 28328
rect 45772 31564 45812 31604
rect 45676 31480 45716 31520
rect 46444 31480 46484 31520
rect 45484 30724 45524 30764
rect 45388 30640 45428 30680
rect 46540 30640 46580 30680
rect 46636 30556 46676 30596
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 47500 30556 47540 30596
rect 48556 30556 48596 30596
rect 44908 28288 44948 28328
rect 45196 28288 45236 28328
rect 45580 29800 45620 29840
rect 46732 29800 46772 29840
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 45484 29128 45524 29168
rect 45580 28288 45620 28328
rect 46924 29128 46964 29168
rect 48172 29800 48212 29840
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 47308 28288 47348 28328
rect 40876 27700 40916 27740
rect 43948 27700 43988 27740
rect 45292 27700 45332 27740
rect 41548 26776 41588 26816
rect 42028 26776 42068 26816
rect 41452 26692 41492 26732
rect 40492 26608 40532 26648
rect 36556 26104 36596 26144
rect 31468 24508 31508 24548
rect 31276 24340 31316 24380
rect 30604 23752 30644 23792
rect 31180 21568 31220 21608
rect 28972 21484 29012 21524
rect 28780 21400 28820 21440
rect 27052 20812 27092 20852
rect 28300 20812 28340 20852
rect 28780 20560 28820 20600
rect 27244 18460 27284 18500
rect 29164 20224 29204 20264
rect 28396 20140 28436 20180
rect 28300 19972 28340 20012
rect 28012 19216 28052 19256
rect 27628 18376 27668 18416
rect 27916 18376 27956 18416
rect 27052 18292 27092 18332
rect 28876 19216 28916 19256
rect 34060 24508 34100 24548
rect 34348 24508 34388 24548
rect 33964 24340 34004 24380
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 32812 23752 32852 23792
rect 32620 23080 32660 23120
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 41644 26020 41684 26060
rect 35116 24592 35156 24632
rect 36556 24592 36596 24632
rect 34924 23752 34964 23792
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 33772 23080 33812 23120
rect 34444 22828 34484 22868
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 33484 22408 33524 22448
rect 34252 22408 34292 22448
rect 35020 22408 35060 22448
rect 35212 24340 35252 24380
rect 35500 23752 35540 23792
rect 42892 26608 42932 26648
rect 44428 26104 44468 26144
rect 43372 26020 43412 26060
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 46156 26104 46196 26144
rect 45580 25180 45620 25220
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 46444 25264 46484 25304
rect 47788 25264 47828 25304
rect 46924 25180 46964 25220
rect 43564 24508 43604 24548
rect 44908 24508 44948 24548
rect 46348 24508 46388 24548
rect 43852 23752 43892 23792
rect 35692 23164 35732 23204
rect 36844 23164 36884 23204
rect 40300 23164 40340 23204
rect 35212 22828 35252 22868
rect 32812 21736 32852 21776
rect 32428 21652 32468 21692
rect 32140 21568 32180 21608
rect 34924 22072 34964 22112
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 33292 21652 33332 21692
rect 34828 21652 34868 21692
rect 35116 22072 35156 22112
rect 36652 21736 36692 21776
rect 37228 21736 37268 21776
rect 32428 21400 32468 21440
rect 31180 20056 31220 20096
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 31468 19804 31508 19844
rect 29356 19132 29396 19172
rect 31084 19132 31124 19172
rect 28492 18460 28532 18500
rect 28492 17956 28532 17996
rect 28972 17956 29012 17996
rect 29164 17956 29204 17996
rect 26668 17704 26708 17744
rect 26572 17620 26612 17660
rect 25228 16192 25268 16232
rect 25708 16192 25748 16232
rect 25324 15604 25364 15644
rect 25708 15520 25748 15560
rect 27628 17704 27668 17744
rect 29260 17704 29300 17744
rect 27724 17032 27764 17072
rect 29452 16192 29492 16232
rect 31084 16192 31124 16232
rect 26860 15520 26900 15560
rect 33100 19804 33140 19844
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 35020 21568 35060 21608
rect 41068 23164 41108 23204
rect 45676 23836 45716 23876
rect 45580 23752 45620 23792
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 47788 24592 47828 24632
rect 49612 24592 49652 24632
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 46156 23836 46196 23876
rect 47692 23836 47732 23876
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 45964 22240 46004 22280
rect 49324 22240 49364 22280
rect 37516 21568 37556 21608
rect 38092 21568 38132 21608
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 33772 19468 33812 19508
rect 38956 20728 38996 20768
rect 39628 20728 39668 20768
rect 39820 20728 39860 20768
rect 38668 20056 38708 20096
rect 39052 20644 39092 20684
rect 40396 20728 40436 20768
rect 44812 21736 44852 21776
rect 41836 21568 41876 21608
rect 43084 21568 43124 21608
rect 44044 21568 44084 21608
rect 39916 20644 39956 20684
rect 39052 20056 39092 20096
rect 35404 19468 35444 19508
rect 32332 19048 32372 19088
rect 33772 19048 33812 19088
rect 33484 18880 33524 18920
rect 34060 18880 34100 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 35884 18880 35924 18920
rect 37516 18880 37556 18920
rect 38188 18880 38228 18920
rect 32716 17032 32756 17072
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 37036 17704 37076 17744
rect 36652 17620 36692 17660
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 33580 15520 33620 15560
rect 33676 15436 33716 15476
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 24172 13000 24212 13040
rect 26092 12580 26132 12620
rect 26764 12580 26804 12620
rect 24076 12496 24116 12536
rect 23596 12328 23636 12368
rect 23980 12328 24020 12368
rect 28300 12580 28340 12620
rect 27724 12244 27764 12284
rect 23692 11740 23732 11780
rect 22636 11320 22676 11360
rect 24172 11656 24212 11696
rect 29932 12496 29972 12536
rect 30700 12496 30740 12536
rect 30028 11908 30068 11948
rect 30316 11908 30356 11948
rect 29548 11656 29588 11696
rect 24844 11320 24884 11360
rect 28684 11320 28724 11360
rect 30124 11152 30164 11192
rect 23404 10396 23444 10436
rect 21868 9472 21908 9512
rect 23500 8632 23540 8672
rect 24460 8632 24500 8672
rect 22348 7960 22388 8000
rect 23212 7960 23252 8000
rect 23980 7960 24020 8000
rect 24268 7960 24308 8000
rect 23404 7876 23444 7916
rect 23404 7708 23444 7748
rect 24364 7876 24404 7916
rect 26860 10144 26900 10184
rect 28012 10144 28052 10184
rect 28204 10144 28244 10184
rect 27916 8800 27956 8840
rect 25708 8632 25748 8672
rect 24844 7708 24884 7748
rect 23020 7036 23060 7076
rect 21772 4096 21812 4136
rect 22924 4096 22964 4136
rect 21676 3760 21716 3800
rect 20620 3424 20660 3464
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 652 2248 692 2288
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 12268 2080 12308 2120
rect 13324 2080 13364 2120
rect 18988 2752 19028 2792
rect 24268 4096 24308 4136
rect 25036 4096 25076 4136
rect 24172 3760 24212 3800
rect 22156 3424 22196 3464
rect 19180 2584 19220 2624
rect 21292 2584 21332 2624
rect 21676 2584 21716 2624
rect 25420 7876 25460 7916
rect 25996 8548 26036 8588
rect 25900 7876 25940 7916
rect 27340 8632 27380 8672
rect 27820 8632 27860 8672
rect 28300 10060 28340 10100
rect 29740 10060 29780 10100
rect 29644 8800 29684 8840
rect 27244 8548 27284 8588
rect 26188 4348 26228 4388
rect 26860 4348 26900 4388
rect 25900 4096 25940 4136
rect 25324 2668 25364 2708
rect 24172 2584 24212 2624
rect 25036 2584 25076 2624
rect 27628 8128 27668 8168
rect 28300 8128 28340 8168
rect 29548 8632 29588 8672
rect 29836 9976 29876 10016
rect 29164 8212 29204 8252
rect 30028 8044 30068 8084
rect 28492 7036 28532 7076
rect 29644 7708 29684 7748
rect 28780 6364 28820 6404
rect 28972 6280 29012 6320
rect 28108 4936 28148 4976
rect 28588 4936 28628 4976
rect 26956 3340 26996 3380
rect 28588 2584 28628 2624
rect 31276 12412 31316 12452
rect 31468 11656 31508 11696
rect 31180 11068 31220 11108
rect 31372 11152 31412 11192
rect 34348 16360 34388 16400
rect 35404 16360 35444 16400
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 34060 15520 34100 15560
rect 34540 15436 34580 15476
rect 34060 15352 34100 15392
rect 41452 18628 41492 18668
rect 43756 21400 43796 21440
rect 44428 20560 44468 20600
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 46444 21736 46484 21776
rect 45964 21568 46004 21608
rect 45580 21400 45620 21440
rect 45196 20728 45236 20768
rect 45004 20140 45044 20180
rect 46060 20140 46100 20180
rect 43564 19804 43604 19844
rect 43084 18628 43124 18668
rect 37900 17704 37940 17744
rect 39052 17704 39092 17744
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 46828 20728 46868 20768
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 50284 20056 50324 20096
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 48748 18544 48788 18584
rect 46444 18460 46484 18500
rect 42220 17704 42260 17744
rect 42700 17704 42740 17744
rect 43564 17704 43604 17744
rect 45100 17704 45140 17744
rect 38668 16948 38708 16988
rect 40396 16948 40436 16988
rect 38572 15436 38612 15476
rect 39628 15520 39668 15560
rect 40684 15520 40724 15560
rect 46060 17032 46100 17072
rect 49324 18544 49364 18584
rect 52492 19216 52532 19256
rect 52492 18964 52532 19004
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 53356 20056 53396 20096
rect 56908 20056 56948 20096
rect 55276 19300 55316 19340
rect 50284 18880 50324 18920
rect 52396 18880 52436 18920
rect 52684 18880 52724 18920
rect 53548 18880 53588 18920
rect 55180 18880 55220 18920
rect 49132 18460 49172 18500
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 50284 18460 50324 18500
rect 47788 17872 47828 17912
rect 48844 17872 48884 17912
rect 49516 17788 49556 17828
rect 49036 17704 49076 17744
rect 49708 17704 49748 17744
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 50188 17284 50228 17324
rect 48172 17032 48212 17072
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 38764 15436 38804 15476
rect 39532 15436 39572 15476
rect 35788 14680 35828 14720
rect 33676 14512 33716 14552
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 31756 12496 31796 12536
rect 35884 12496 35924 12536
rect 32236 12412 32276 12452
rect 31660 11908 31700 11948
rect 32044 11152 32084 11192
rect 36748 14680 36788 14720
rect 38764 14008 38804 14048
rect 39148 14008 39188 14048
rect 36748 13168 36788 13208
rect 36940 13168 36980 13208
rect 38860 13168 38900 13208
rect 39724 13168 39764 13208
rect 41164 13168 41204 13208
rect 35212 12244 35252 12284
rect 36652 12244 36692 12284
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 35212 11656 35252 11696
rect 32716 11572 32756 11612
rect 33100 11572 33140 11612
rect 32332 11320 32372 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 31948 11068 31988 11108
rect 31564 10984 31604 11024
rect 30892 10732 30932 10772
rect 31276 9976 31316 10016
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 33196 9472 33236 9512
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 34444 9472 34484 9512
rect 33292 8800 33332 8840
rect 34156 8800 34196 8840
rect 33388 8632 33428 8672
rect 33196 8548 33236 8588
rect 34156 8632 34196 8672
rect 33868 8548 33908 8588
rect 32332 8128 32372 8168
rect 33100 8128 33140 8168
rect 31660 8044 31700 8084
rect 33964 8212 34004 8252
rect 33772 7960 33812 8000
rect 34060 7960 34100 8000
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 34540 8632 34580 8672
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 40876 13000 40916 13040
rect 38188 12496 38228 12536
rect 37036 12244 37076 12284
rect 41644 13000 41684 13040
rect 41164 12412 41204 12452
rect 41452 12244 41492 12284
rect 41356 11824 41396 11864
rect 38188 11656 38228 11696
rect 37900 11152 37940 11192
rect 37132 9472 37172 9512
rect 36364 9304 36404 9344
rect 37132 9304 37172 9344
rect 35884 8632 35924 8672
rect 32332 6364 32372 6404
rect 35692 7960 35732 8000
rect 35308 7540 35348 7580
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 33484 5860 33524 5900
rect 31468 4936 31508 4976
rect 30796 4264 30836 4304
rect 31084 3928 31124 3968
rect 31660 3928 31700 3968
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 34348 6448 34388 6488
rect 39148 11152 39188 11192
rect 38284 11068 38324 11108
rect 38380 10984 38420 11024
rect 39052 10984 39092 11024
rect 38284 9472 38324 9512
rect 39052 10144 39092 10184
rect 40684 11068 40724 11108
rect 39532 10732 39572 10772
rect 40492 10732 40532 10772
rect 41644 11656 41684 11696
rect 41932 12412 41972 12452
rect 42700 12580 42740 12620
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 43084 12580 43124 12620
rect 42988 12412 43028 12452
rect 42412 12244 42452 12284
rect 42604 12244 42644 12284
rect 42892 11824 42932 11864
rect 45388 14008 45428 14048
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 51340 17872 51380 17912
rect 52012 17872 52052 17912
rect 52300 17872 52340 17912
rect 51148 17704 51188 17744
rect 51244 17620 51284 17660
rect 56812 19300 56852 19340
rect 56044 19216 56084 19256
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 57484 19468 57524 19508
rect 58060 19468 58100 19508
rect 57004 19216 57044 19256
rect 55468 17620 55508 17660
rect 50380 17368 50420 17408
rect 53164 17032 53204 17072
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 43756 13924 43796 13964
rect 44236 13924 44276 13964
rect 49036 14008 49076 14048
rect 49324 14008 49364 14048
rect 51532 14848 51572 14888
rect 50572 14092 50612 14132
rect 52204 14680 52244 14720
rect 52972 14092 53012 14132
rect 51244 14008 51284 14048
rect 47980 13840 48020 13880
rect 49612 13840 49652 13880
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 47308 11656 47348 11696
rect 48844 11656 48884 11696
rect 50572 12496 50612 12536
rect 42604 11488 42644 11528
rect 43084 11488 43124 11528
rect 43948 11152 43988 11192
rect 44332 11068 44372 11108
rect 46636 11068 46676 11108
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 55180 16780 55220 16820
rect 56044 16780 56084 16820
rect 54028 14848 54068 14888
rect 53836 14680 53876 14720
rect 53644 14176 53684 14216
rect 54028 14260 54068 14300
rect 54796 14260 54836 14300
rect 53836 14008 53876 14048
rect 53644 12496 53684 12536
rect 55180 14176 55220 14216
rect 55564 14680 55604 14720
rect 56524 14764 56564 14804
rect 56140 14680 56180 14720
rect 56332 14512 56372 14552
rect 56716 14512 56756 14552
rect 55660 14092 55700 14132
rect 56812 14092 56852 14132
rect 57196 14092 57236 14132
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 59020 14680 59060 14720
rect 59404 14680 59444 14720
rect 59308 14596 59348 14636
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 59788 14176 59828 14216
rect 61420 14176 61460 14216
rect 56620 13840 56660 13880
rect 54124 12328 54164 12368
rect 52588 10984 52628 11024
rect 53164 10984 53204 11024
rect 47212 10060 47252 10100
rect 48460 10060 48500 10100
rect 48076 9640 48116 9680
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 49324 9640 49364 9680
rect 54796 12328 54836 12368
rect 57004 14008 57044 14048
rect 57868 14008 57908 14048
rect 57292 13840 57332 13880
rect 55660 12328 55700 12368
rect 55468 10312 55508 10352
rect 53452 10144 53492 10184
rect 55372 10144 55412 10184
rect 51724 10060 51764 10100
rect 52396 10060 52436 10100
rect 44524 8716 44564 8756
rect 45676 8716 45716 8756
rect 40972 8548 41012 8588
rect 42124 8548 42164 8588
rect 37996 7540 38036 7580
rect 39916 7540 39956 7580
rect 38860 7204 38900 7244
rect 39532 7204 39572 7244
rect 39724 7204 39764 7244
rect 39532 6532 39572 6572
rect 39148 6448 39188 6488
rect 33964 5860 34004 5900
rect 35980 5608 36020 5648
rect 36556 5608 36596 5648
rect 37228 5608 37268 5648
rect 37420 5608 37460 5648
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 37612 5020 37652 5060
rect 39340 5608 39380 5648
rect 39436 5524 39476 5564
rect 38380 5020 38420 5060
rect 37132 4852 37172 4892
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 39436 4852 39476 4892
rect 40204 4852 40244 4892
rect 39436 4096 39476 4136
rect 40108 4096 40148 4136
rect 38092 3172 38132 3212
rect 39244 3172 39284 3212
rect 37996 2668 38036 2708
rect 38476 2668 38516 2708
rect 40780 6532 40820 6572
rect 47116 8716 47156 8756
rect 46732 8044 46772 8084
rect 46636 7960 46676 8000
rect 47212 7960 47252 8000
rect 43372 6448 43412 6488
rect 46348 6448 46388 6488
rect 44620 6196 44660 6236
rect 46732 6448 46772 6488
rect 46444 6280 46484 6320
rect 41068 5524 41108 5564
rect 40684 4096 40724 4136
rect 41068 4096 41108 4136
rect 41260 4096 41300 4136
rect 41644 4096 41684 4136
rect 42028 3172 42068 3212
rect 43084 3172 43124 3212
rect 42700 2668 42740 2708
rect 20908 2500 20948 2540
rect 39340 2584 39380 2624
rect 40204 2584 40244 2624
rect 41836 2584 41876 2624
rect 47500 5608 47540 5648
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 48556 8044 48596 8084
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 49324 7456 49364 7496
rect 51532 7456 51572 7496
rect 49228 7372 49268 7412
rect 50380 7372 50420 7412
rect 49804 7120 49844 7160
rect 54892 9976 54932 10016
rect 55468 9976 55508 10016
rect 54508 9472 54548 9512
rect 54124 9220 54164 9260
rect 60268 14008 60308 14048
rect 60844 14008 60884 14048
rect 55852 10312 55892 10352
rect 58828 10312 58868 10352
rect 56428 10144 56468 10184
rect 54700 9220 54740 9260
rect 55372 8716 55412 8756
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 46444 3424 46484 3464
rect 46636 3424 46676 3464
rect 45004 2836 45044 2876
rect 45772 2836 45812 2876
rect 43468 2584 43508 2624
rect 46156 2584 46196 2624
rect 47020 2584 47060 2624
rect 47596 3172 47636 3212
rect 48940 5608 48980 5648
rect 48748 5524 48788 5564
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 48748 3592 48788 3632
rect 48556 3172 48596 3212
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 47980 2584 48020 2624
rect 48364 2584 48404 2624
rect 49036 5524 49076 5564
rect 52108 5440 52148 5480
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 49324 5104 49364 5144
rect 50092 5104 50132 5144
rect 52108 5104 52148 5144
rect 49132 3424 49172 3464
rect 50380 5020 50420 5060
rect 49612 4096 49652 4136
rect 53260 7120 53300 7160
rect 53356 5440 53396 5480
rect 52780 5020 52820 5060
rect 50476 4096 50516 4136
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 49516 3592 49556 3632
rect 50379 3592 50419 3632
rect 50572 2668 50612 2708
rect 51820 2668 51860 2708
rect 53164 4936 53204 4976
rect 53452 4936 53492 4976
rect 53356 2668 53396 2708
rect 55660 9472 55700 9512
rect 55756 8800 55796 8840
rect 56428 8800 56468 8840
rect 56524 8716 56564 8756
rect 58444 10144 58484 10184
rect 58636 10144 58676 10184
rect 59020 10144 59060 10184
rect 59212 10060 59252 10100
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 59980 10228 60020 10268
rect 61132 10228 61172 10268
rect 61420 10144 61460 10184
rect 61996 10144 62036 10184
rect 60748 10060 60788 10100
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 59884 9472 59924 9512
rect 56812 8800 56852 8840
rect 56716 8716 56756 8756
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 60844 8716 60884 8756
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 56428 7120 56468 7160
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 55372 4936 55412 4976
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 54028 2836 54068 2876
rect 54604 2836 54644 2876
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal3 >>
rect 4343 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 4729 38576
rect 19463 38536 19472 38576
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19840 38536 19849 38576
rect 34583 38536 34592 38576
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34960 38536 34969 38576
rect 49703 38536 49712 38576
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 50080 38536 50089 38576
rect 64823 38536 64832 38576
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 65200 38536 65209 38576
rect 79943 38536 79952 38576
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 80320 38536 80329 38576
rect 95063 38536 95072 38576
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95440 38536 95449 38576
rect 3103 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 3489 37820
rect 18223 37780 18232 37820
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18600 37780 18609 37820
rect 33343 37780 33352 37820
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33720 37780 33729 37820
rect 48463 37780 48472 37820
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48840 37780 48849 37820
rect 63583 37780 63592 37820
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63960 37780 63969 37820
rect 78703 37780 78712 37820
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 79080 37780 79089 37820
rect 93823 37780 93832 37820
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 94200 37780 94209 37820
rect 0 37568 80 37588
rect 0 37528 20620 37568
rect 20660 37528 20669 37568
rect 0 37508 80 37528
rect 35587 37360 35596 37400
rect 35636 37360 36940 37400
rect 36980 37360 36989 37400
rect 18307 37276 18316 37316
rect 18356 37276 19276 37316
rect 19316 37276 19325 37316
rect 4343 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 4729 37064
rect 19463 37024 19472 37064
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19840 37024 19849 37064
rect 34583 37024 34592 37064
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34960 37024 34969 37064
rect 49703 37024 49712 37064
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 50080 37024 50089 37064
rect 64823 37024 64832 37064
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 65200 37024 65209 37064
rect 79943 37024 79952 37064
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 80320 37024 80329 37064
rect 95063 37024 95072 37064
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95440 37024 95449 37064
rect 10339 36856 10348 36896
rect 10388 36856 11788 36896
rect 11828 36856 11837 36896
rect 0 36728 80 36748
rect 0 36688 76 36728
rect 116 36688 125 36728
rect 18787 36688 18796 36728
rect 18836 36688 19852 36728
rect 19892 36688 19901 36728
rect 23980 36688 24940 36728
rect 24980 36688 24989 36728
rect 36451 36688 36460 36728
rect 36500 36688 37804 36728
rect 37844 36688 38572 36728
rect 38612 36688 38621 36728
rect 0 36668 80 36688
rect 5827 36604 5836 36644
rect 5876 36604 6320 36644
rect 6280 36560 6320 36604
rect 23980 36560 24020 36688
rect 36931 36604 36940 36644
rect 36980 36604 37708 36644
rect 37748 36604 37757 36644
rect 4675 36520 4684 36560
rect 4724 36520 5644 36560
rect 5684 36520 5693 36560
rect 6280 36520 6604 36560
rect 6644 36520 7372 36560
rect 7412 36520 7421 36560
rect 18691 36520 18700 36560
rect 18740 36520 19180 36560
rect 19220 36520 23980 36560
rect 24020 36520 24029 36560
rect 24931 36520 24940 36560
rect 24980 36520 25804 36560
rect 25844 36520 25853 36560
rect 30211 36520 30220 36560
rect 30260 36520 31180 36560
rect 31220 36520 31229 36560
rect 31363 36520 31372 36560
rect 31412 36520 32140 36560
rect 32180 36520 33100 36560
rect 33140 36520 33149 36560
rect 37507 36520 37516 36560
rect 37556 36520 38956 36560
rect 38996 36520 39005 36560
rect 3103 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 3489 36308
rect 18223 36268 18232 36308
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18600 36268 18609 36308
rect 33343 36268 33352 36308
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33720 36268 33729 36308
rect 48463 36268 48472 36308
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48840 36268 48849 36308
rect 63583 36268 63592 36308
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63960 36268 63969 36308
rect 78703 36268 78712 36308
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 79080 36268 79089 36308
rect 93823 36268 93832 36308
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 94200 36268 94209 36308
rect 35395 36184 35404 36224
rect 35444 36184 36076 36224
rect 36116 36184 36652 36224
rect 36692 36184 36701 36224
rect 20035 35932 20044 35972
rect 20084 35932 22156 35972
rect 22196 35932 22205 35972
rect 36259 35932 36268 35972
rect 36308 35932 36652 35972
rect 36692 35932 36844 35972
rect 36884 35932 36893 35972
rect 0 35828 80 35908
rect 5059 35848 5068 35888
rect 5108 35848 9100 35888
rect 9140 35848 9772 35888
rect 9812 35848 9964 35888
rect 10004 35848 10013 35888
rect 19459 35848 19468 35888
rect 19508 35848 21292 35888
rect 21332 35848 21341 35888
rect 21475 35848 21484 35888
rect 21524 35848 23212 35888
rect 23252 35848 24748 35888
rect 24788 35848 25228 35888
rect 25268 35848 25277 35888
rect 8707 35764 8716 35804
rect 8756 35764 9292 35804
rect 9332 35764 9341 35804
rect 10339 35680 10348 35720
rect 10388 35680 11980 35720
rect 12020 35680 12029 35720
rect 4343 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 4729 35552
rect 19463 35512 19472 35552
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19840 35512 19849 35552
rect 34583 35512 34592 35552
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34960 35512 34969 35552
rect 49703 35512 49712 35552
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 50080 35512 50089 35552
rect 64823 35512 64832 35552
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 65200 35512 65209 35552
rect 79943 35512 79952 35552
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 80320 35512 80329 35552
rect 95063 35512 95072 35552
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95440 35512 95449 35552
rect 7363 35260 7372 35300
rect 7412 35260 8428 35300
rect 8468 35260 8477 35300
rect 22339 35260 22348 35300
rect 22388 35260 24844 35300
rect 24884 35260 25324 35300
rect 25364 35260 26188 35300
rect 26228 35260 26237 35300
rect 5059 35176 5068 35216
rect 5108 35176 5836 35216
rect 5876 35176 7468 35216
rect 7508 35176 7948 35216
rect 7988 35176 7997 35216
rect 33187 35176 33196 35216
rect 33236 35176 35788 35216
rect 35828 35176 35837 35216
rect 8035 35092 8044 35132
rect 8084 35092 9292 35132
rect 9332 35092 9676 35132
rect 9716 35092 9725 35132
rect 31459 35092 31468 35132
rect 31508 35092 32236 35132
rect 32276 35092 33292 35132
rect 33332 35092 33772 35132
rect 33812 35092 33821 35132
rect 0 34988 80 35068
rect 30307 34924 30316 34964
rect 30356 34924 31276 34964
rect 31316 34924 31325 34964
rect 3103 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 3489 34796
rect 18223 34756 18232 34796
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18600 34756 18609 34796
rect 33343 34756 33352 34796
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33720 34756 33729 34796
rect 48463 34756 48472 34796
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48840 34756 48849 34796
rect 63583 34756 63592 34796
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63960 34756 63969 34796
rect 78703 34756 78712 34796
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 79080 34756 79089 34796
rect 93823 34756 93832 34796
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 94200 34756 94209 34796
rect 16867 34420 16876 34460
rect 16916 34420 17740 34460
rect 17780 34420 17789 34460
rect 4291 34336 4300 34376
rect 4340 34336 4972 34376
rect 5012 34336 5021 34376
rect 30691 34336 30700 34376
rect 30740 34336 32428 34376
rect 32468 34336 32477 34376
rect 33859 34336 33868 34376
rect 33908 34336 35404 34376
rect 35444 34336 35453 34376
rect 36259 34336 36268 34376
rect 36308 34336 37324 34376
rect 37364 34336 37373 34376
rect 14467 34252 14476 34292
rect 14516 34252 15436 34292
rect 15476 34252 15485 34292
rect 0 34148 80 34228
rect 8227 34168 8236 34208
rect 8276 34168 8812 34208
rect 8852 34168 8861 34208
rect 15715 34168 15724 34208
rect 15764 34168 16204 34208
rect 16244 34168 20332 34208
rect 20372 34168 23020 34208
rect 23060 34168 23069 34208
rect 4343 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 4729 34040
rect 19463 34000 19472 34040
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19840 34000 19849 34040
rect 20803 34000 20812 34040
rect 20852 34000 22348 34040
rect 22388 34000 24556 34040
rect 24596 34000 24605 34040
rect 34583 34000 34592 34040
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34960 34000 34969 34040
rect 49703 34000 49712 34040
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 50080 34000 50089 34040
rect 64823 34000 64832 34040
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 65200 34000 65209 34040
rect 79943 34000 79952 34040
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 80320 34000 80329 34040
rect 95063 34000 95072 34040
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95440 34000 95449 34040
rect 9667 33664 9676 33704
rect 9716 33664 11116 33704
rect 11156 33664 11165 33704
rect 24259 33664 24268 33704
rect 24308 33664 25036 33704
rect 25076 33664 25085 33704
rect 10051 33496 10060 33536
rect 10100 33496 10732 33536
rect 10772 33496 11404 33536
rect 11444 33496 11453 33536
rect 45667 33412 45676 33452
rect 45716 33412 46828 33452
rect 46868 33412 46877 33452
rect 0 33308 80 33388
rect 3103 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 3489 33284
rect 18223 33244 18232 33284
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18600 33244 18609 33284
rect 33343 33244 33352 33284
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33720 33244 33729 33284
rect 48463 33244 48472 33284
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48840 33244 48849 33284
rect 63583 33244 63592 33284
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63960 33244 63969 33284
rect 78703 33244 78712 33284
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 79080 33244 79089 33284
rect 93823 33244 93832 33284
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 94200 33244 94209 33284
rect 14947 33076 14956 33116
rect 14996 33076 15916 33116
rect 15956 33076 15965 33116
rect 42499 32992 42508 33032
rect 42548 32992 43372 33032
rect 43412 32992 43421 33032
rect 15619 32908 15628 32948
rect 15668 32908 17068 32948
rect 17108 32908 17117 32948
rect 23980 32908 25996 32948
rect 26036 32908 26045 32948
rect 43555 32908 43564 32948
rect 43604 32908 44332 32948
rect 44372 32908 44381 32948
rect 23980 32864 24020 32908
rect 4108 32824 5972 32864
rect 7459 32824 7468 32864
rect 7508 32824 9676 32864
rect 9716 32824 9725 32864
rect 12067 32824 12076 32864
rect 12116 32824 15668 32864
rect 20515 32824 20524 32864
rect 20564 32824 22156 32864
rect 22196 32824 23980 32864
rect 24020 32824 24029 32864
rect 25027 32824 25036 32864
rect 25076 32824 26860 32864
rect 26900 32824 28588 32864
rect 28628 32824 28637 32864
rect 4108 32780 4148 32824
rect 5932 32780 5972 32824
rect 15628 32780 15668 32824
rect 4068 32740 4108 32780
rect 4148 32740 4157 32780
rect 5892 32740 5932 32780
rect 5972 32740 5981 32780
rect 15588 32740 15628 32780
rect 15668 32740 15677 32780
rect 5932 32696 5972 32740
rect 5932 32656 6508 32696
rect 6548 32656 6557 32696
rect 27619 32656 27628 32696
rect 27668 32656 28012 32696
rect 28052 32656 28061 32696
rect 0 32468 80 32548
rect 4343 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 4729 32528
rect 19463 32488 19472 32528
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19840 32488 19849 32528
rect 34583 32488 34592 32528
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34960 32488 34969 32528
rect 49703 32488 49712 32528
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 50080 32488 50089 32528
rect 64823 32488 64832 32528
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 65200 32488 65209 32528
rect 79943 32488 79952 32528
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 80320 32488 80329 32528
rect 95063 32488 95072 32528
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95440 32488 95449 32528
rect 34243 32236 34252 32276
rect 34292 32236 37708 32276
rect 37748 32236 37757 32276
rect 38851 32236 38860 32276
rect 38900 32236 39916 32276
rect 39956 32236 39965 32276
rect 6979 32152 6988 32192
rect 7028 32152 10060 32192
rect 10100 32152 10109 32192
rect 16099 32152 16108 32192
rect 16148 32152 17164 32192
rect 17204 32152 17213 32192
rect 37219 32152 37228 32192
rect 37268 32152 37996 32192
rect 38036 32152 38284 32192
rect 38324 32152 38333 32192
rect 39715 32152 39724 32192
rect 39764 32152 40396 32192
rect 40436 32152 40445 32192
rect 36259 32068 36268 32108
rect 36308 32068 36940 32108
rect 36980 32068 37612 32108
rect 37652 32068 37661 32108
rect 11203 31900 11212 31940
rect 11252 31900 11788 31940
rect 11828 31900 11837 31940
rect 17059 31900 17068 31940
rect 17108 31900 17740 31940
rect 17780 31900 17789 31940
rect 37315 31900 37324 31940
rect 37364 31900 38764 31940
rect 38804 31900 38813 31940
rect 3103 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 3489 31772
rect 18223 31732 18232 31772
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18600 31732 18609 31772
rect 33343 31732 33352 31772
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33720 31732 33729 31772
rect 48463 31732 48472 31772
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48840 31732 48849 31772
rect 63583 31732 63592 31772
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63960 31732 63969 31772
rect 78703 31732 78712 31772
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 79080 31732 79089 31772
rect 93823 31732 93832 31772
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 94200 31732 94209 31772
rect 0 31628 80 31708
rect 17155 31564 17164 31604
rect 17204 31564 18124 31604
rect 18164 31564 18316 31604
rect 18356 31564 18365 31604
rect 42883 31564 42892 31604
rect 42932 31564 45196 31604
rect 45236 31564 45772 31604
rect 45812 31564 45821 31604
rect 9187 31480 9196 31520
rect 9236 31480 12076 31520
rect 12116 31480 12125 31520
rect 33763 31480 33772 31520
rect 33812 31480 34252 31520
rect 34292 31480 34301 31520
rect 44515 31480 44524 31520
rect 44564 31480 45676 31520
rect 45716 31480 46444 31520
rect 46484 31480 46493 31520
rect 9196 31184 9236 31480
rect 36163 31396 36172 31436
rect 36212 31396 38476 31436
rect 38516 31396 38525 31436
rect 32419 31312 32428 31352
rect 32468 31312 33100 31352
rect 33140 31312 33149 31352
rect 37411 31312 37420 31352
rect 37460 31312 38572 31352
rect 38612 31312 38621 31352
rect 4867 31144 4876 31184
rect 4916 31144 9236 31184
rect 24355 31144 24364 31184
rect 24404 31144 25708 31184
rect 25748 31144 25757 31184
rect 4343 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 4729 31016
rect 19463 30976 19472 31016
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19840 30976 19849 31016
rect 34583 30976 34592 31016
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34960 30976 34969 31016
rect 49703 30976 49712 31016
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 50080 30976 50089 31016
rect 64823 30976 64832 31016
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 65200 30976 65209 31016
rect 79943 30976 79952 31016
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 80320 30976 80329 31016
rect 95063 30976 95072 31016
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95440 30976 95449 31016
rect 0 30788 80 30868
rect 22531 30808 22540 30848
rect 22580 30808 23884 30848
rect 23924 30808 23933 30848
rect 34627 30808 34636 30848
rect 34676 30808 35116 30848
rect 35156 30808 35165 30848
rect 35971 30808 35980 30848
rect 36020 30808 37612 30848
rect 37652 30808 37661 30848
rect 17923 30724 17932 30764
rect 17972 30724 20140 30764
rect 20180 30724 20189 30764
rect 25315 30724 25324 30764
rect 25364 30724 25612 30764
rect 25652 30724 26956 30764
rect 26996 30724 27005 30764
rect 32803 30724 32812 30764
rect 32852 30724 35500 30764
rect 35540 30724 35549 30764
rect 35779 30724 35788 30764
rect 35828 30724 37132 30764
rect 37172 30724 37181 30764
rect 41827 30724 41836 30764
rect 41876 30724 45484 30764
rect 45524 30724 45533 30764
rect 2851 30640 2860 30680
rect 2900 30640 3916 30680
rect 3956 30640 3965 30680
rect 15427 30640 15436 30680
rect 15476 30640 16204 30680
rect 16244 30640 17068 30680
rect 17108 30640 17117 30680
rect 17251 30640 17260 30680
rect 17300 30640 18220 30680
rect 18260 30640 18269 30680
rect 25219 30640 25228 30680
rect 25268 30640 25804 30680
rect 25844 30640 25853 30680
rect 31555 30640 31564 30680
rect 31604 30640 33772 30680
rect 33812 30640 34156 30680
rect 34196 30640 34205 30680
rect 35107 30640 35116 30680
rect 35156 30640 35596 30680
rect 35636 30640 36460 30680
rect 36500 30640 36509 30680
rect 38371 30640 38380 30680
rect 38420 30640 44332 30680
rect 44372 30640 44381 30680
rect 45379 30640 45388 30680
rect 45428 30640 46540 30680
rect 46580 30640 46589 30680
rect 3235 30556 3244 30596
rect 3284 30556 3628 30596
rect 3668 30556 3820 30596
rect 3860 30556 8236 30596
rect 8276 30556 8285 30596
rect 14371 30388 14380 30428
rect 14420 30388 15244 30428
rect 15284 30388 15293 30428
rect 17260 30260 17300 30640
rect 26083 30556 26092 30596
rect 26132 30556 26764 30596
rect 26804 30556 26813 30596
rect 46627 30556 46636 30596
rect 46676 30556 47500 30596
rect 47540 30556 48556 30596
rect 48596 30556 48605 30596
rect 3103 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 3489 30260
rect 16387 30220 16396 30260
rect 16436 30220 17260 30260
rect 17300 30220 17309 30260
rect 18223 30220 18232 30260
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18600 30220 18609 30260
rect 33343 30220 33352 30260
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33720 30220 33729 30260
rect 34051 30220 34060 30260
rect 34100 30220 39916 30260
rect 39956 30220 40684 30260
rect 40724 30220 41452 30260
rect 41492 30220 41501 30260
rect 48463 30220 48472 30260
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48840 30220 48849 30260
rect 63583 30220 63592 30260
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63960 30220 63969 30260
rect 78703 30220 78712 30260
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 79080 30220 79089 30260
rect 93823 30220 93832 30260
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 94200 30220 94209 30260
rect 23203 30052 23212 30092
rect 23252 30052 24268 30092
rect 24308 30052 25324 30092
rect 25364 30052 25373 30092
rect 0 29948 80 30028
rect 4099 29968 4108 30008
rect 4148 29968 5068 30008
rect 5108 29968 5452 30008
rect 5492 29968 5501 30008
rect 20515 29968 20524 30008
rect 20564 29968 21196 30008
rect 21236 29968 21245 30008
rect 3715 29884 3724 29924
rect 3764 29884 4588 29924
rect 4628 29884 4972 29924
rect 5012 29884 5021 29924
rect 18691 29884 18700 29924
rect 18740 29884 20812 29924
rect 20852 29884 20861 29924
rect 10147 29800 10156 29840
rect 10196 29800 22636 29840
rect 22676 29800 22685 29840
rect 27043 29800 27052 29840
rect 27092 29800 27724 29840
rect 27764 29800 28972 29840
rect 29012 29800 29021 29840
rect 38083 29800 38092 29840
rect 38132 29800 39628 29840
rect 39668 29800 39677 29840
rect 43747 29800 43756 29840
rect 43796 29800 44524 29840
rect 44564 29800 45580 29840
rect 45620 29800 46732 29840
rect 46772 29800 48172 29840
rect 48212 29800 48221 29840
rect 40867 29548 40876 29588
rect 40916 29548 42892 29588
rect 42932 29548 42941 29588
rect 4343 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 4729 29504
rect 19463 29464 19472 29504
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19840 29464 19849 29504
rect 34583 29464 34592 29504
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34960 29464 34969 29504
rect 49703 29464 49712 29504
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 50080 29464 50089 29504
rect 64823 29464 64832 29504
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 65200 29464 65209 29504
rect 79943 29464 79952 29504
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 80320 29464 80329 29504
rect 95063 29464 95072 29504
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95440 29464 95449 29504
rect 22627 29212 22636 29252
rect 22676 29212 22685 29252
rect 0 29108 80 29188
rect 22636 29168 22676 29212
rect 5923 29128 5932 29168
rect 5972 29128 7852 29168
rect 7892 29128 7901 29168
rect 11011 29128 11020 29168
rect 11060 29128 11884 29168
rect 11924 29128 11933 29168
rect 15043 29128 15052 29168
rect 15092 29128 15820 29168
rect 15860 29128 15869 29168
rect 16675 29128 16684 29168
rect 16724 29128 19276 29168
rect 19316 29128 21388 29168
rect 21428 29128 22060 29168
rect 22100 29128 22109 29168
rect 22636 29128 23116 29168
rect 23156 29128 31564 29168
rect 31604 29128 31613 29168
rect 45475 29128 45484 29168
rect 45524 29128 46924 29168
rect 46964 29128 46973 29168
rect 8227 29044 8236 29084
rect 8276 29044 15244 29084
rect 15284 29044 15293 29084
rect 22627 29044 22636 29084
rect 22676 29044 24308 29084
rect 24268 29000 24308 29044
rect 24259 28960 24268 29000
rect 24308 28960 24317 29000
rect 3103 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 3489 28748
rect 18223 28708 18232 28748
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18600 28708 18609 28748
rect 33343 28708 33352 28748
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33720 28708 33729 28748
rect 48463 28708 48472 28748
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48840 28708 48849 28748
rect 63583 28708 63592 28748
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63960 28708 63969 28748
rect 78703 28708 78712 28748
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 79080 28708 79089 28748
rect 93823 28708 93832 28748
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 94200 28708 94209 28748
rect 27139 28372 27148 28412
rect 27188 28372 28780 28412
rect 28820 28372 28829 28412
rect 0 28268 80 28348
rect 20611 28288 20620 28328
rect 20660 28288 22156 28328
rect 22196 28288 22205 28328
rect 28867 28288 28876 28328
rect 28916 28288 29068 28328
rect 29108 28288 29117 28328
rect 40963 28288 40972 28328
rect 41012 28288 43948 28328
rect 43988 28288 43997 28328
rect 44899 28288 44908 28328
rect 44948 28288 45196 28328
rect 45236 28288 45580 28328
rect 45620 28288 47308 28328
rect 47348 28288 47357 28328
rect 23971 28120 23980 28160
rect 24020 28120 26476 28160
rect 26516 28120 26525 28160
rect 4343 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 4729 27992
rect 19463 27952 19472 27992
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19840 27952 19849 27992
rect 34583 27952 34592 27992
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34960 27952 34969 27992
rect 49703 27952 49712 27992
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 50080 27952 50089 27992
rect 64823 27952 64832 27992
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 65200 27952 65209 27992
rect 79943 27952 79952 27992
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 80320 27952 80329 27992
rect 95063 27952 95072 27992
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95440 27952 95449 27992
rect 4396 27868 4972 27908
rect 5012 27868 5021 27908
rect 4396 27824 4436 27868
rect 4387 27784 4396 27824
rect 4436 27784 4445 27824
rect 4675 27784 4684 27824
rect 4724 27784 5740 27824
rect 5780 27784 5789 27824
rect 4291 27700 4300 27740
rect 4340 27700 5452 27740
rect 5492 27700 5501 27740
rect 26179 27700 26188 27740
rect 26228 27700 26764 27740
rect 26804 27700 26813 27740
rect 40195 27700 40204 27740
rect 40244 27700 40876 27740
rect 40916 27700 40925 27740
rect 43939 27700 43948 27740
rect 43988 27700 45292 27740
rect 45332 27700 45341 27740
rect 3811 27616 3820 27656
rect 3860 27616 4588 27656
rect 4628 27616 5108 27656
rect 9763 27616 9772 27656
rect 9812 27616 10156 27656
rect 10196 27616 10205 27656
rect 39619 27616 39628 27656
rect 39668 27616 40300 27656
rect 40340 27616 40349 27656
rect 0 27428 80 27508
rect 5068 27488 5108 27616
rect 5059 27448 5068 27488
rect 5108 27448 5117 27488
rect 5251 27364 5260 27404
rect 5300 27364 7084 27404
rect 7124 27364 7133 27404
rect 3103 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 3489 27236
rect 18223 27196 18232 27236
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18600 27196 18609 27236
rect 33343 27196 33352 27236
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33720 27196 33729 27236
rect 48463 27196 48472 27236
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48840 27196 48849 27236
rect 63583 27196 63592 27236
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63960 27196 63969 27236
rect 78703 27196 78712 27236
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 79080 27196 79089 27236
rect 93823 27196 93832 27236
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 94200 27196 94209 27236
rect 3427 26860 3436 26900
rect 3476 26860 4204 26900
rect 4244 26860 4253 26900
rect 9571 26776 9580 26816
rect 9620 26776 10156 26816
rect 10196 26776 10205 26816
rect 28867 26776 28876 26816
rect 28916 26776 29164 26816
rect 29204 26776 29213 26816
rect 32515 26776 32524 26816
rect 32564 26776 33196 26816
rect 33236 26776 33245 26816
rect 35299 26776 35308 26816
rect 35348 26776 39628 26816
rect 39668 26776 41548 26816
rect 41588 26776 42028 26816
rect 42068 26776 42077 26816
rect 28675 26692 28684 26732
rect 28724 26692 38476 26732
rect 38516 26692 38525 26732
rect 40291 26692 40300 26732
rect 40340 26692 41452 26732
rect 41492 26692 41501 26732
rect 0 26588 80 26668
rect 2467 26608 2476 26648
rect 2516 26608 3628 26648
rect 3668 26608 3677 26648
rect 30595 26608 30604 26648
rect 30644 26608 34444 26648
rect 34484 26608 34493 26648
rect 34915 26608 34924 26648
rect 34964 26608 34973 26648
rect 35107 26608 35116 26648
rect 35156 26608 36460 26648
rect 36500 26608 36509 26648
rect 40483 26608 40492 26648
rect 40532 26608 42892 26648
rect 42932 26608 42941 26648
rect 34924 26564 34964 26608
rect 26563 26524 26572 26564
rect 26612 26524 28876 26564
rect 28916 26524 32908 26564
rect 32948 26524 32957 26564
rect 33580 26524 34964 26564
rect 33580 26480 33620 26524
rect 2371 26440 2380 26480
rect 2420 26440 3244 26480
rect 3284 26440 3293 26480
rect 4343 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 4729 26480
rect 4867 26440 4876 26480
rect 4916 26440 5740 26480
rect 5780 26440 5789 26480
rect 6787 26440 6796 26480
rect 6836 26440 9484 26480
rect 9524 26440 11884 26480
rect 11924 26440 11933 26480
rect 19463 26440 19472 26480
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19840 26440 19849 26480
rect 33571 26440 33580 26480
rect 33620 26440 33629 26480
rect 34583 26440 34592 26480
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34960 26440 34969 26480
rect 49703 26440 49712 26480
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 50080 26440 50089 26480
rect 64823 26440 64832 26480
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 65200 26440 65209 26480
rect 79943 26440 79952 26480
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 80320 26440 80329 26480
rect 95063 26440 95072 26480
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95440 26440 95449 26480
rect 11683 26188 11692 26228
rect 11732 26188 12268 26228
rect 12308 26188 12317 26228
rect 2851 26104 2860 26144
rect 2900 26104 7468 26144
rect 7508 26104 7517 26144
rect 19075 26104 19084 26144
rect 19124 26104 23596 26144
rect 23636 26104 26092 26144
rect 26132 26104 26141 26144
rect 36547 26104 36556 26144
rect 36596 26104 44428 26144
rect 44468 26104 46156 26144
rect 46196 26104 46205 26144
rect 41635 26020 41644 26060
rect 41684 26020 43372 26060
rect 43412 26020 43421 26060
rect 27139 25852 27148 25892
rect 27188 25852 27724 25892
rect 27764 25852 27773 25892
rect 0 25748 80 25828
rect 3103 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 3489 25724
rect 18223 25684 18232 25724
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18600 25684 18609 25724
rect 33343 25684 33352 25724
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33720 25684 33729 25724
rect 48463 25684 48472 25724
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48840 25684 48849 25724
rect 63583 25684 63592 25724
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63960 25684 63969 25724
rect 78703 25684 78712 25724
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 79080 25684 79089 25724
rect 93823 25684 93832 25724
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 94200 25684 94209 25724
rect 6115 25516 6124 25556
rect 6164 25516 8332 25556
rect 8372 25516 8381 25556
rect 16867 25516 16876 25556
rect 16916 25516 17836 25556
rect 17876 25516 17885 25556
rect 22723 25432 22732 25472
rect 22772 25432 24556 25472
rect 24596 25432 24605 25472
rect 3715 25264 3724 25304
rect 3764 25264 5068 25304
rect 5108 25264 5836 25304
rect 5876 25264 5885 25304
rect 11779 25264 11788 25304
rect 11828 25264 12076 25304
rect 12116 25264 12125 25304
rect 21091 25264 21100 25304
rect 21140 25264 21772 25304
rect 21812 25264 21821 25304
rect 29635 25264 29644 25304
rect 29684 25264 30604 25304
rect 30644 25264 30653 25304
rect 46435 25264 46444 25304
rect 46484 25264 47788 25304
rect 47828 25264 47837 25304
rect 45571 25180 45580 25220
rect 45620 25180 46924 25220
rect 46964 25180 46973 25220
rect 0 24908 80 24988
rect 4343 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 4729 24968
rect 19463 24928 19472 24968
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19840 24928 19849 24968
rect 34583 24928 34592 24968
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34960 24928 34969 24968
rect 49703 24928 49712 24968
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 50080 24928 50089 24968
rect 64823 24928 64832 24968
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 65200 24928 65209 24968
rect 79943 24928 79952 24968
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 80320 24928 80329 24968
rect 95063 24928 95072 24968
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95440 24928 95449 24968
rect 14083 24676 14092 24716
rect 14132 24676 16436 24716
rect 20899 24676 20908 24716
rect 20948 24676 22924 24716
rect 22964 24676 22973 24716
rect 26083 24676 26092 24716
rect 26132 24676 26764 24716
rect 26804 24676 26813 24716
rect 16396 24632 16436 24676
rect 13795 24592 13804 24632
rect 13844 24592 15244 24632
rect 15284 24592 15293 24632
rect 16387 24592 16396 24632
rect 16436 24592 16445 24632
rect 21091 24592 21100 24632
rect 21140 24592 21484 24632
rect 21524 24592 21533 24632
rect 23587 24592 23596 24632
rect 23636 24592 23960 24632
rect 25219 24592 25228 24632
rect 25268 24592 25900 24632
rect 25940 24592 26956 24632
rect 26996 24592 27436 24632
rect 27476 24592 27485 24632
rect 31555 24592 31564 24632
rect 31604 24592 32044 24632
rect 32084 24592 35116 24632
rect 35156 24592 36556 24632
rect 36596 24592 36605 24632
rect 47779 24592 47788 24632
rect 47828 24592 49612 24632
rect 49652 24592 49661 24632
rect 23920 24548 23960 24592
rect 23920 24508 24748 24548
rect 24788 24508 24797 24548
rect 31459 24508 31468 24548
rect 31508 24508 34060 24548
rect 34100 24508 34348 24548
rect 34388 24508 34397 24548
rect 43555 24508 43564 24548
rect 43604 24508 44908 24548
rect 44948 24508 46348 24548
rect 46388 24508 46397 24548
rect 9091 24424 9100 24464
rect 9140 24424 12172 24464
rect 12212 24424 14860 24464
rect 14900 24424 14909 24464
rect 15907 24424 15916 24464
rect 15956 24424 17068 24464
rect 17108 24424 17117 24464
rect 20995 24340 21004 24380
rect 21044 24340 21964 24380
rect 22004 24340 22013 24380
rect 30211 24340 30220 24380
rect 30260 24340 31276 24380
rect 31316 24340 31325 24380
rect 33955 24340 33964 24380
rect 34004 24340 35212 24380
rect 35252 24340 35261 24380
rect 3103 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 3489 24212
rect 18223 24172 18232 24212
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18600 24172 18609 24212
rect 33343 24172 33352 24212
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33720 24172 33729 24212
rect 48463 24172 48472 24212
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48840 24172 48849 24212
rect 63583 24172 63592 24212
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63960 24172 63969 24212
rect 78703 24172 78712 24212
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 79080 24172 79089 24212
rect 93823 24172 93832 24212
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 94200 24172 94209 24212
rect 0 24068 80 24148
rect 20323 23836 20332 23876
rect 20372 23836 20812 23876
rect 20852 23836 21004 23876
rect 21044 23836 21053 23876
rect 45667 23836 45676 23876
rect 45716 23836 46156 23876
rect 46196 23836 47692 23876
rect 47732 23836 47741 23876
rect 15907 23752 15916 23792
rect 15956 23752 17068 23792
rect 17108 23752 17117 23792
rect 17635 23752 17644 23792
rect 17684 23752 18316 23792
rect 18356 23752 19084 23792
rect 19124 23752 19133 23792
rect 30595 23752 30604 23792
rect 30644 23752 32812 23792
rect 32852 23752 32861 23792
rect 34915 23752 34924 23792
rect 34964 23752 35500 23792
rect 35540 23752 35549 23792
rect 43843 23752 43852 23792
rect 43892 23752 45580 23792
rect 45620 23752 45629 23792
rect 15427 23668 15436 23708
rect 15476 23668 16204 23708
rect 16244 23668 16253 23708
rect 4343 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 4729 23456
rect 19463 23416 19472 23456
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19840 23416 19849 23456
rect 34583 23416 34592 23456
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34960 23416 34969 23456
rect 49703 23416 49712 23456
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 50080 23416 50089 23456
rect 64823 23416 64832 23456
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 65200 23416 65209 23456
rect 79943 23416 79952 23456
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 80320 23416 80329 23456
rect 95063 23416 95072 23456
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95440 23416 95449 23456
rect 0 23228 80 23308
rect 35683 23164 35692 23204
rect 35732 23164 36844 23204
rect 36884 23164 36893 23204
rect 40291 23164 40300 23204
rect 40340 23164 41068 23204
rect 41108 23164 41117 23204
rect 1219 23080 1228 23120
rect 1268 23080 2092 23120
rect 2132 23080 2141 23120
rect 32611 23080 32620 23120
rect 32660 23080 33772 23120
rect 33812 23080 33821 23120
rect 4483 22996 4492 23036
rect 4532 22996 5452 23036
rect 5492 22996 5501 23036
rect 2755 22828 2764 22868
rect 2804 22828 2956 22868
rect 2996 22828 4148 22868
rect 34435 22828 34444 22868
rect 34484 22828 35212 22868
rect 35252 22828 35261 22868
rect 4108 22700 4148 22828
rect 3103 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 3489 22700
rect 4099 22660 4108 22700
rect 4148 22660 4157 22700
rect 18223 22660 18232 22700
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18600 22660 18609 22700
rect 33343 22660 33352 22700
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33720 22660 33729 22700
rect 48463 22660 48472 22700
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48840 22660 48849 22700
rect 63583 22660 63592 22700
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63960 22660 63969 22700
rect 78703 22660 78712 22700
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 79080 22660 79089 22700
rect 93823 22660 93832 22700
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 94200 22660 94209 22700
rect 16003 22492 16012 22532
rect 16052 22492 16204 22532
rect 16244 22492 16253 22532
rect 0 22388 80 22468
rect 33475 22408 33484 22448
rect 33524 22408 34252 22448
rect 34292 22408 35020 22448
rect 35060 22408 35069 22448
rect 2659 22324 2668 22364
rect 2708 22324 3244 22364
rect 3284 22324 3724 22364
rect 3764 22324 4204 22364
rect 4244 22324 4253 22364
rect 2371 22240 2380 22280
rect 2420 22240 5068 22280
rect 5108 22240 5117 22280
rect 9955 22240 9964 22280
rect 10004 22240 14764 22280
rect 14804 22240 14813 22280
rect 25699 22156 25708 22196
rect 25748 22156 26476 22196
rect 26516 22156 26525 22196
rect 35020 22112 35060 22408
rect 45955 22240 45964 22280
rect 46004 22240 49324 22280
rect 49364 22240 49373 22280
rect 34915 22072 34924 22112
rect 34964 22072 34973 22112
rect 35020 22072 35116 22112
rect 35156 22072 35165 22112
rect 34924 22028 34964 22072
rect 35011 22028 35069 22029
rect 14755 21988 14764 22028
rect 14804 21988 15340 22028
rect 15380 21988 20044 22028
rect 20084 21988 20093 22028
rect 34924 21988 35020 22028
rect 35060 21988 35069 22028
rect 35011 21987 35069 21988
rect 4343 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 4729 21944
rect 19463 21904 19472 21944
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19840 21904 19849 21944
rect 34583 21904 34592 21944
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34960 21904 34969 21944
rect 49703 21904 49712 21944
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 50080 21904 50089 21944
rect 64823 21904 64832 21944
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 65200 21904 65209 21944
rect 79943 21904 79952 21944
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 80320 21904 80329 21944
rect 95063 21904 95072 21944
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95440 21904 95449 21944
rect 32803 21736 32812 21776
rect 32852 21736 36652 21776
rect 36692 21736 37228 21776
rect 37268 21736 37277 21776
rect 44803 21736 44812 21776
rect 44852 21736 46444 21776
rect 46484 21736 46493 21776
rect 35011 21692 35069 21693
rect 32419 21652 32428 21692
rect 32468 21652 33292 21692
rect 33332 21652 33341 21692
rect 34819 21652 34828 21692
rect 34868 21652 35020 21692
rect 35060 21652 35069 21692
rect 35011 21651 35069 21652
rect 0 21608 80 21628
rect 0 21568 652 21608
rect 692 21568 701 21608
rect 8419 21568 8428 21608
rect 8468 21568 9484 21608
rect 9524 21568 9533 21608
rect 10435 21568 10444 21608
rect 10484 21568 11020 21608
rect 11060 21568 11788 21608
rect 11828 21568 11837 21608
rect 12259 21568 12268 21608
rect 12308 21568 13036 21608
rect 13076 21568 13085 21608
rect 15715 21568 15724 21608
rect 15764 21568 17644 21608
rect 17684 21568 17693 21608
rect 25795 21568 25804 21608
rect 25844 21568 26860 21608
rect 26900 21568 26909 21608
rect 27043 21568 27052 21608
rect 27092 21568 31180 21608
rect 31220 21568 31229 21608
rect 32131 21568 32140 21608
rect 32180 21568 35020 21608
rect 35060 21568 35069 21608
rect 37507 21568 37516 21608
rect 37556 21568 38092 21608
rect 38132 21568 41836 21608
rect 41876 21568 43084 21608
rect 43124 21568 43133 21608
rect 44035 21568 44044 21608
rect 44084 21568 45964 21608
rect 46004 21568 46013 21608
rect 0 21548 80 21568
rect 28195 21484 28204 21524
rect 28244 21484 28972 21524
rect 29012 21484 29021 21524
rect 13987 21400 13996 21440
rect 14036 21400 15244 21440
rect 15284 21400 15293 21440
rect 28771 21400 28780 21440
rect 28820 21400 32428 21440
rect 32468 21400 32477 21440
rect 43747 21400 43756 21440
rect 43796 21400 45580 21440
rect 45620 21400 45629 21440
rect 19939 21316 19948 21356
rect 19988 21316 20332 21356
rect 20372 21316 20381 21356
rect 3103 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 3489 21188
rect 18223 21148 18232 21188
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18600 21148 18609 21188
rect 33343 21148 33352 21188
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33720 21148 33729 21188
rect 48463 21148 48472 21188
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48840 21148 48849 21188
rect 63583 21148 63592 21188
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63960 21148 63969 21188
rect 78703 21148 78712 21188
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 79080 21148 79089 21188
rect 93823 21148 93832 21188
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 94200 21148 94209 21188
rect 5827 20980 5836 21020
rect 5876 20980 8044 21020
rect 8084 20980 8093 21020
rect 27043 20812 27052 20852
rect 27092 20812 28300 20852
rect 28340 20812 28349 20852
rect 0 20768 80 20788
rect 0 20728 652 20768
rect 692 20728 701 20768
rect 11395 20728 11404 20768
rect 11444 20728 12172 20768
rect 12212 20728 12221 20768
rect 38947 20728 38956 20768
rect 38996 20728 39628 20768
rect 39668 20728 39677 20768
rect 39811 20728 39820 20768
rect 39860 20728 40396 20768
rect 40436 20728 40445 20768
rect 45187 20728 45196 20768
rect 45236 20728 46828 20768
rect 46868 20728 46877 20768
rect 0 20708 80 20728
rect 39043 20644 39052 20684
rect 39092 20644 39916 20684
rect 39956 20644 41600 20684
rect 41560 20600 41600 20644
rect 21955 20560 21964 20600
rect 22004 20560 28780 20600
rect 28820 20560 28829 20600
rect 41560 20560 44428 20600
rect 44468 20560 44477 20600
rect 4343 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 4729 20432
rect 19463 20392 19472 20432
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19840 20392 19849 20432
rect 34583 20392 34592 20432
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34960 20392 34969 20432
rect 49703 20392 49712 20432
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 50080 20392 50089 20432
rect 64823 20392 64832 20432
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 65200 20392 65209 20432
rect 79943 20392 79952 20432
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 80320 20392 80329 20432
rect 95063 20392 95072 20432
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95440 20392 95449 20432
rect 28960 20224 29164 20264
rect 29204 20224 29213 20264
rect 28960 20180 29000 20224
rect 4771 20140 4780 20180
rect 4820 20140 5164 20180
rect 5204 20140 5213 20180
rect 6280 20140 23960 20180
rect 28387 20140 28396 20180
rect 28436 20140 29000 20180
rect 44995 20140 45004 20180
rect 45044 20140 46060 20180
rect 46100 20140 46109 20180
rect 6280 20096 6320 20140
rect 23920 20096 23960 20140
rect 67 20056 76 20096
rect 116 20056 6320 20096
rect 22243 20056 22252 20096
rect 22292 20056 22732 20096
rect 22772 20056 22781 20096
rect 23920 20056 31180 20096
rect 31220 20056 31229 20096
rect 38659 20056 38668 20096
rect 38708 20056 39052 20096
rect 39092 20056 39101 20096
rect 50275 20056 50284 20096
rect 50324 20056 53356 20096
rect 53396 20056 56908 20096
rect 56948 20056 56957 20096
rect 4579 19972 4588 20012
rect 4628 19972 4876 20012
rect 4916 19972 4925 20012
rect 20323 19972 20332 20012
rect 20372 19972 21388 20012
rect 21428 19972 25228 20012
rect 25268 19972 25277 20012
rect 26659 19972 26668 20012
rect 26708 19972 28300 20012
rect 28340 19972 28349 20012
rect 0 19928 80 19948
rect 0 19888 652 19928
rect 692 19888 701 19928
rect 0 19868 80 19888
rect 20419 19804 20428 19844
rect 20468 19804 20812 19844
rect 20852 19804 20861 19844
rect 31459 19804 31468 19844
rect 31508 19804 33100 19844
rect 33140 19804 43564 19844
rect 43604 19804 43613 19844
rect 3103 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 3489 19676
rect 18223 19636 18232 19676
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18600 19636 18609 19676
rect 33343 19636 33352 19676
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33720 19636 33729 19676
rect 48463 19636 48472 19676
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48840 19636 48849 19676
rect 63583 19636 63592 19676
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63960 19636 63969 19676
rect 78703 19636 78712 19676
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 79080 19636 79089 19676
rect 93823 19636 93832 19676
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 94200 19636 94209 19676
rect 2659 19468 2668 19508
rect 2708 19468 3724 19508
rect 3764 19468 3773 19508
rect 33763 19468 33772 19508
rect 33812 19468 35404 19508
rect 35444 19468 35453 19508
rect 57475 19468 57484 19508
rect 57524 19468 58060 19508
rect 58100 19468 58109 19508
rect 4675 19384 4684 19424
rect 4724 19384 4764 19424
rect 4684 19340 4724 19384
rect 3139 19300 3148 19340
rect 3188 19300 5260 19340
rect 5300 19300 5548 19340
rect 5588 19300 5597 19340
rect 55267 19300 55276 19340
rect 55316 19300 56812 19340
rect 56852 19300 56861 19340
rect 2755 19216 2764 19256
rect 2804 19216 3436 19256
rect 3476 19216 3485 19256
rect 5347 19216 5356 19256
rect 5396 19216 7372 19256
rect 7412 19216 7421 19256
rect 28003 19216 28012 19256
rect 28052 19216 28876 19256
rect 28916 19216 28925 19256
rect 52483 19216 52492 19256
rect 52532 19216 56044 19256
rect 56084 19216 57004 19256
rect 57044 19216 57053 19256
rect 3436 19172 3476 19216
rect 3436 19132 9484 19172
rect 9524 19132 9533 19172
rect 29347 19132 29356 19172
rect 29396 19132 31084 19172
rect 31124 19132 31133 19172
rect 0 19088 80 19108
rect 0 19048 652 19088
rect 692 19048 701 19088
rect 2275 19048 2284 19088
rect 2324 19048 2956 19088
rect 2996 19048 3005 19088
rect 4387 19048 4396 19088
rect 4436 19048 7756 19088
rect 7796 19048 7805 19088
rect 9763 19048 9772 19088
rect 9812 19048 10732 19088
rect 10772 19048 10781 19088
rect 32323 19048 32332 19088
rect 32372 19048 33772 19088
rect 33812 19048 33821 19088
rect 0 19028 80 19048
rect 52300 18964 52492 19004
rect 52532 18964 52541 19004
rect 52300 18920 52340 18964
rect 4343 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 4729 18920
rect 19463 18880 19472 18920
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19840 18880 19849 18920
rect 33475 18880 33484 18920
rect 33524 18880 34060 18920
rect 34100 18880 34109 18920
rect 34583 18880 34592 18920
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34960 18880 34969 18920
rect 35875 18880 35884 18920
rect 35924 18880 37516 18920
rect 37556 18880 38188 18920
rect 38228 18880 38237 18920
rect 49703 18880 49712 18920
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 50080 18880 50089 18920
rect 50275 18880 50284 18920
rect 50324 18880 52340 18920
rect 52387 18880 52396 18920
rect 52436 18880 52684 18920
rect 52724 18880 53548 18920
rect 53588 18880 55180 18920
rect 55220 18880 55229 18920
rect 64823 18880 64832 18920
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 65200 18880 65209 18920
rect 79943 18880 79952 18920
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 80320 18880 80329 18920
rect 95063 18880 95072 18920
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95440 18880 95449 18920
rect 41443 18628 41452 18668
rect 41492 18628 43084 18668
rect 43124 18628 43133 18668
rect 48739 18544 48748 18584
rect 48788 18544 49324 18584
rect 49364 18544 49373 18584
rect 27235 18460 27244 18500
rect 27284 18460 28492 18500
rect 28532 18460 28541 18500
rect 46435 18460 46444 18500
rect 46484 18460 49132 18500
rect 49172 18460 50284 18500
rect 50324 18460 50333 18500
rect 26851 18376 26860 18416
rect 26900 18376 27628 18416
rect 27668 18376 27916 18416
rect 27956 18376 27965 18416
rect 26179 18292 26188 18332
rect 26228 18292 27052 18332
rect 27092 18292 27101 18332
rect 0 18248 80 18268
rect 0 18208 652 18248
rect 692 18208 701 18248
rect 0 18188 80 18208
rect 3103 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 3489 18164
rect 18223 18124 18232 18164
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18600 18124 18609 18164
rect 33343 18124 33352 18164
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33720 18124 33729 18164
rect 48463 18124 48472 18164
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48840 18124 48849 18164
rect 63583 18124 63592 18164
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63960 18124 63969 18164
rect 78703 18124 78712 18164
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 79080 18124 79089 18164
rect 93823 18124 93832 18164
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 94200 18124 94209 18164
rect 28483 17956 28492 17996
rect 28532 17956 28972 17996
rect 29012 17956 29164 17996
rect 29204 17956 29213 17996
rect 14851 17872 14860 17912
rect 14900 17872 15820 17912
rect 15860 17872 15869 17912
rect 47779 17872 47788 17912
rect 47828 17872 48844 17912
rect 48884 17872 48893 17912
rect 50380 17872 51340 17912
rect 51380 17872 52012 17912
rect 52052 17872 52300 17912
rect 52340 17872 52349 17912
rect 50380 17828 50420 17872
rect 8611 17788 8620 17828
rect 8660 17788 9868 17828
rect 9908 17788 10828 17828
rect 10868 17788 10877 17828
rect 49507 17788 49516 17828
rect 49556 17788 50420 17828
rect 3427 17704 3436 17744
rect 3476 17704 4204 17744
rect 4244 17704 4253 17744
rect 25699 17704 25708 17744
rect 25748 17704 26668 17744
rect 26708 17704 26717 17744
rect 27619 17704 27628 17744
rect 27668 17704 29260 17744
rect 29300 17704 29309 17744
rect 37027 17704 37036 17744
rect 37076 17704 37900 17744
rect 37940 17704 37949 17744
rect 39043 17704 39052 17744
rect 39092 17704 42220 17744
rect 42260 17704 42700 17744
rect 42740 17704 42749 17744
rect 43555 17704 43564 17744
rect 43604 17704 45100 17744
rect 45140 17704 45149 17744
rect 49027 17704 49036 17744
rect 49076 17704 49708 17744
rect 49748 17704 51148 17744
rect 51188 17704 51197 17744
rect 39052 17660 39092 17704
rect 11971 17620 11980 17660
rect 12020 17620 12844 17660
rect 12884 17620 12893 17660
rect 16003 17620 16012 17660
rect 16052 17620 16780 17660
rect 16820 17620 17548 17660
rect 17588 17620 17597 17660
rect 25219 17620 25228 17660
rect 25268 17620 26092 17660
rect 26132 17620 26572 17660
rect 26612 17620 26621 17660
rect 36643 17620 36652 17660
rect 36692 17620 39092 17660
rect 51235 17620 51244 17660
rect 51284 17620 55468 17660
rect 55508 17620 55517 17660
rect 0 17408 80 17428
rect 0 17368 652 17408
rect 692 17368 701 17408
rect 4343 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 4729 17408
rect 19463 17368 19472 17408
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19840 17368 19849 17408
rect 34583 17368 34592 17408
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34960 17368 34969 17408
rect 49703 17368 49712 17408
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 50080 17368 50089 17408
rect 50188 17368 50380 17408
rect 50420 17368 50429 17408
rect 64823 17368 64832 17408
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 65200 17368 65209 17408
rect 79943 17368 79952 17408
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 80320 17368 80329 17408
rect 95063 17368 95072 17408
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95440 17368 95449 17408
rect 0 17348 80 17368
rect 50188 17324 50228 17368
rect 50179 17284 50188 17324
rect 50228 17284 50237 17324
rect 2179 17200 2188 17240
rect 2228 17200 3052 17240
rect 3092 17200 3101 17240
rect 27715 17032 27724 17072
rect 27764 17032 32716 17072
rect 32756 17032 32765 17072
rect 46051 17032 46060 17072
rect 46100 17032 48172 17072
rect 48212 17032 53164 17072
rect 53204 17032 53213 17072
rect 3235 16948 3244 16988
rect 3284 16948 4012 16988
rect 4052 16948 4061 16988
rect 38659 16948 38668 16988
rect 38708 16948 40396 16988
rect 40436 16948 40445 16988
rect 55171 16780 55180 16820
rect 55220 16780 56044 16820
rect 56084 16780 56093 16820
rect 3103 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 3489 16652
rect 18223 16612 18232 16652
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18600 16612 18609 16652
rect 33343 16612 33352 16652
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33720 16612 33729 16652
rect 48463 16612 48472 16652
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48840 16612 48849 16652
rect 63583 16612 63592 16652
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63960 16612 63969 16652
rect 78703 16612 78712 16652
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 79080 16612 79089 16652
rect 93823 16612 93832 16652
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 94200 16612 94209 16652
rect 0 16568 80 16588
rect 0 16528 652 16568
rect 692 16528 701 16568
rect 0 16508 80 16528
rect 14947 16360 14956 16400
rect 14996 16360 15820 16400
rect 15860 16360 15869 16400
rect 20131 16360 20140 16400
rect 20180 16360 21292 16400
rect 21332 16360 21341 16400
rect 34339 16360 34348 16400
rect 34388 16360 35404 16400
rect 35444 16360 35453 16400
rect 18019 16276 18028 16316
rect 18068 16276 18508 16316
rect 18548 16276 19468 16316
rect 19508 16276 20044 16316
rect 20084 16276 20093 16316
rect 14947 16192 14956 16232
rect 14996 16192 15244 16232
rect 15284 16192 19276 16232
rect 19316 16192 25228 16232
rect 25268 16192 25708 16232
rect 25748 16192 25757 16232
rect 29443 16192 29452 16232
rect 29492 16192 31084 16232
rect 31124 16192 31133 16232
rect 18787 15940 18796 15980
rect 18836 15940 20332 15980
rect 20372 15940 20381 15980
rect 4343 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 4729 15896
rect 19463 15856 19472 15896
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19840 15856 19849 15896
rect 34583 15856 34592 15896
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34960 15856 34969 15896
rect 49703 15856 49712 15896
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 50080 15856 50089 15896
rect 64823 15856 64832 15896
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 65200 15856 65209 15896
rect 79943 15856 79952 15896
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 80320 15856 80329 15896
rect 95063 15856 95072 15896
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95440 15856 95449 15896
rect 0 15728 80 15748
rect 0 15688 556 15728
rect 596 15688 605 15728
rect 14563 15688 14572 15728
rect 14612 15688 15628 15728
rect 15668 15688 15677 15728
rect 0 15668 80 15688
rect 18691 15604 18700 15644
rect 18740 15604 25324 15644
rect 25364 15604 25373 15644
rect 16963 15520 16972 15560
rect 17012 15520 18796 15560
rect 18836 15520 18845 15560
rect 22435 15520 22444 15560
rect 22484 15520 22636 15560
rect 22676 15520 22924 15560
rect 22964 15520 22973 15560
rect 25699 15520 25708 15560
rect 25748 15520 26860 15560
rect 26900 15520 26909 15560
rect 33571 15520 33580 15560
rect 33620 15520 34060 15560
rect 34100 15520 34109 15560
rect 39619 15520 39628 15560
rect 39668 15520 40684 15560
rect 40724 15520 40733 15560
rect 15811 15436 15820 15476
rect 15860 15436 17836 15476
rect 17876 15436 17885 15476
rect 33667 15436 33676 15476
rect 33716 15436 34540 15476
rect 34580 15436 34589 15476
rect 38563 15436 38572 15476
rect 38612 15436 38764 15476
rect 38804 15436 39532 15476
rect 39572 15436 39581 15476
rect 34060 15392 34100 15436
rect 17539 15352 17548 15392
rect 17588 15352 18508 15392
rect 18548 15352 18557 15392
rect 18691 15352 18700 15392
rect 18740 15352 19948 15392
rect 19988 15352 19997 15392
rect 34051 15352 34060 15392
rect 34100 15352 34140 15392
rect 18700 15308 18740 15352
rect 17635 15268 17644 15308
rect 17684 15268 18740 15308
rect 3103 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 3489 15140
rect 18223 15100 18232 15140
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18600 15100 18609 15140
rect 33343 15100 33352 15140
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33720 15100 33729 15140
rect 48463 15100 48472 15140
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48840 15100 48849 15140
rect 63583 15100 63592 15140
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63960 15100 63969 15140
rect 78703 15100 78712 15140
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 79080 15100 79089 15140
rect 93823 15100 93832 15140
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 94200 15100 94209 15140
rect 20131 15016 20140 15056
rect 20180 15016 20428 15056
rect 20468 15016 22540 15056
rect 22580 15016 22589 15056
rect 0 14888 80 14908
rect 0 14848 652 14888
rect 692 14848 701 14888
rect 51523 14848 51532 14888
rect 51572 14848 54028 14888
rect 54068 14848 54077 14888
rect 0 14828 80 14848
rect 55564 14764 56524 14804
rect 56564 14764 56573 14804
rect 55564 14720 55604 14764
rect 8899 14680 8908 14720
rect 8948 14680 9100 14720
rect 9140 14680 10636 14720
rect 10676 14680 10685 14720
rect 20227 14680 20236 14720
rect 20276 14680 21292 14720
rect 21332 14680 21341 14720
rect 35779 14680 35788 14720
rect 35828 14680 36748 14720
rect 36788 14680 36797 14720
rect 52195 14680 52204 14720
rect 52244 14680 53836 14720
rect 53876 14680 53885 14720
rect 55555 14680 55564 14720
rect 55604 14680 55613 14720
rect 56131 14680 56140 14720
rect 56180 14680 56189 14720
rect 59011 14680 59020 14720
rect 59060 14680 59404 14720
rect 59444 14680 59453 14720
rect 56140 14636 56180 14680
rect 56140 14596 59308 14636
rect 59348 14596 59357 14636
rect 4003 14512 4012 14552
rect 4052 14512 4492 14552
rect 4532 14512 7276 14552
rect 7316 14512 8812 14552
rect 8852 14512 8861 14552
rect 18115 14512 18124 14552
rect 18164 14512 20140 14552
rect 20180 14512 20189 14552
rect 23683 14512 23692 14552
rect 23732 14512 33676 14552
rect 33716 14512 33725 14552
rect 56323 14512 56332 14552
rect 56372 14512 56716 14552
rect 56756 14512 56765 14552
rect 20803 14428 20812 14468
rect 20852 14428 21292 14468
rect 21332 14428 21676 14468
rect 21716 14428 21725 14468
rect 4343 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 4729 14384
rect 19463 14344 19472 14384
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19840 14344 19849 14384
rect 34583 14344 34592 14384
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34960 14344 34969 14384
rect 49703 14344 49712 14384
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 50080 14344 50089 14384
rect 64823 14344 64832 14384
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 65200 14344 65209 14384
rect 79943 14344 79952 14384
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 80320 14344 80329 14384
rect 95063 14344 95072 14384
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95440 14344 95449 14384
rect 54019 14260 54028 14300
rect 54068 14260 54796 14300
rect 54836 14260 54845 14300
rect 11299 14176 11308 14216
rect 11348 14176 11884 14216
rect 11924 14176 11933 14216
rect 53635 14176 53644 14216
rect 53684 14176 55180 14216
rect 55220 14176 55229 14216
rect 59779 14176 59788 14216
rect 59828 14176 61420 14216
rect 61460 14176 61469 14216
rect 2947 14092 2956 14132
rect 2996 14092 3820 14132
rect 3860 14092 3869 14132
rect 7171 14092 7180 14132
rect 7220 14092 8044 14132
rect 8084 14092 8093 14132
rect 8419 14092 8428 14132
rect 8468 14092 9196 14132
rect 9236 14092 9245 14132
rect 50563 14092 50572 14132
rect 50612 14092 52972 14132
rect 53012 14092 53021 14132
rect 55651 14092 55660 14132
rect 55700 14092 56812 14132
rect 56852 14092 57196 14132
rect 57236 14092 57245 14132
rect 0 14048 80 14068
rect 0 14008 652 14048
rect 692 14008 701 14048
rect 2755 14008 2764 14048
rect 2804 14008 3340 14048
rect 3380 14008 3389 14048
rect 4195 14008 4204 14048
rect 4244 14008 5836 14048
rect 5876 14008 5885 14048
rect 9283 14008 9292 14048
rect 9332 14008 9580 14048
rect 9620 14008 12076 14048
rect 12116 14008 12125 14048
rect 12259 14008 12268 14048
rect 12308 14008 12748 14048
rect 12788 14008 12797 14048
rect 38755 14008 38764 14048
rect 38804 14008 39148 14048
rect 39188 14008 39197 14048
rect 45379 14008 45388 14048
rect 45428 14008 49036 14048
rect 49076 14008 49324 14048
rect 49364 14008 51244 14048
rect 51284 14008 51293 14048
rect 53827 14008 53836 14048
rect 53876 14008 57004 14048
rect 57044 14008 57053 14048
rect 57859 14008 57868 14048
rect 57908 14008 60268 14048
rect 60308 14008 60844 14048
rect 60884 14008 60893 14048
rect 0 13988 80 14008
rect 3340 13964 3380 14008
rect 3340 13924 4396 13964
rect 4436 13924 4445 13964
rect 5731 13924 5740 13964
rect 5780 13924 6892 13964
rect 6932 13924 7084 13964
rect 7124 13924 7133 13964
rect 17539 13924 17548 13964
rect 17588 13924 18508 13964
rect 18548 13924 18557 13964
rect 43747 13924 43756 13964
rect 43796 13924 44236 13964
rect 44276 13924 44285 13964
rect 4003 13840 4012 13880
rect 4052 13840 5548 13880
rect 5588 13840 5597 13880
rect 6403 13840 6412 13880
rect 6452 13840 9004 13880
rect 9044 13840 10252 13880
rect 10292 13840 10301 13880
rect 47971 13840 47980 13880
rect 48020 13840 49612 13880
rect 49652 13840 49661 13880
rect 56611 13840 56620 13880
rect 56660 13840 57292 13880
rect 57332 13840 57341 13880
rect 3103 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 3489 13628
rect 18223 13588 18232 13628
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18600 13588 18609 13628
rect 33343 13588 33352 13628
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33720 13588 33729 13628
rect 48463 13588 48472 13628
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48840 13588 48849 13628
rect 63583 13588 63592 13628
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63960 13588 63969 13628
rect 78703 13588 78712 13628
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 79080 13588 79089 13628
rect 93823 13588 93832 13628
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 94200 13588 94209 13628
rect 0 13208 80 13228
rect 0 13168 652 13208
rect 692 13168 701 13208
rect 5251 13168 5260 13208
rect 5300 13168 5836 13208
rect 5876 13168 8044 13208
rect 8084 13168 8093 13208
rect 17251 13168 17260 13208
rect 17300 13168 18988 13208
rect 19028 13168 19037 13208
rect 36739 13168 36748 13208
rect 36788 13168 36940 13208
rect 36980 13168 38860 13208
rect 38900 13168 38909 13208
rect 39715 13168 39724 13208
rect 39764 13168 41164 13208
rect 41204 13168 41213 13208
rect 0 13148 80 13168
rect 23683 13000 23692 13040
rect 23732 13000 24172 13040
rect 24212 13000 24221 13040
rect 40867 13000 40876 13040
rect 40916 13000 41644 13040
rect 41684 13000 41693 13040
rect 4343 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 4729 12872
rect 19463 12832 19472 12872
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19840 12832 19849 12872
rect 34583 12832 34592 12872
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34960 12832 34969 12872
rect 49703 12832 49712 12872
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 50080 12832 50089 12872
rect 64823 12832 64832 12872
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 65200 12832 65209 12872
rect 79943 12832 79952 12872
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 80320 12832 80329 12872
rect 95063 12832 95072 12872
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95440 12832 95449 12872
rect 23692 12664 23884 12704
rect 23924 12664 23933 12704
rect 23692 12620 23732 12664
rect 18979 12580 18988 12620
rect 19028 12580 21292 12620
rect 21332 12580 21341 12620
rect 23011 12580 23020 12620
rect 23060 12580 23732 12620
rect 23779 12580 23788 12620
rect 23828 12580 26092 12620
rect 26132 12580 26141 12620
rect 26755 12580 26764 12620
rect 26804 12580 28300 12620
rect 28340 12580 28349 12620
rect 42691 12580 42700 12620
rect 42740 12580 43084 12620
rect 43124 12580 43133 12620
rect 9475 12496 9484 12536
rect 9524 12496 10252 12536
rect 10292 12496 19372 12536
rect 19412 12496 21676 12536
rect 21716 12496 21725 12536
rect 22723 12496 22732 12536
rect 22772 12496 23308 12536
rect 23348 12496 24076 12536
rect 24116 12496 24125 12536
rect 29923 12496 29932 12536
rect 29972 12496 30700 12536
rect 30740 12496 31756 12536
rect 31796 12496 31805 12536
rect 35875 12496 35884 12536
rect 35924 12496 38188 12536
rect 38228 12496 38237 12536
rect 50563 12496 50572 12536
rect 50612 12496 53644 12536
rect 53684 12496 53693 12536
rect 18691 12412 18700 12452
rect 18740 12412 23020 12452
rect 23060 12412 23069 12452
rect 31267 12412 31276 12452
rect 31316 12412 32236 12452
rect 32276 12412 32285 12452
rect 41155 12412 41164 12452
rect 41204 12412 41932 12452
rect 41972 12412 42988 12452
rect 43028 12412 43037 12452
rect 0 12368 80 12388
rect 0 12328 652 12368
rect 692 12328 701 12368
rect 23587 12328 23596 12368
rect 23636 12328 23980 12368
rect 24020 12328 24029 12368
rect 54115 12328 54124 12368
rect 54164 12328 54796 12368
rect 54836 12328 55660 12368
rect 55700 12328 55709 12368
rect 0 12308 80 12328
rect 21763 12244 21772 12284
rect 21812 12244 27724 12284
rect 27764 12244 27773 12284
rect 35203 12244 35212 12284
rect 35252 12244 36652 12284
rect 36692 12244 37036 12284
rect 37076 12244 37085 12284
rect 41443 12244 41452 12284
rect 41492 12244 42412 12284
rect 42452 12244 42604 12284
rect 42644 12244 42653 12284
rect 3103 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 3489 12116
rect 18223 12076 18232 12116
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18600 12076 18609 12116
rect 33343 12076 33352 12116
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33720 12076 33729 12116
rect 48463 12076 48472 12116
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48840 12076 48849 12116
rect 63583 12076 63592 12116
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63960 12076 63969 12116
rect 78703 12076 78712 12116
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 79080 12076 79089 12116
rect 93823 12076 93832 12116
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 94200 12076 94209 12116
rect 30019 11908 30028 11948
rect 30068 11908 30316 11948
rect 30356 11908 31660 11948
rect 31700 11908 31709 11948
rect 41347 11824 41356 11864
rect 41396 11824 42892 11864
rect 42932 11824 42941 11864
rect 23683 11740 23692 11780
rect 23732 11740 23960 11780
rect 23920 11696 23960 11740
rect 23920 11656 24172 11696
rect 24212 11656 24221 11696
rect 29539 11656 29548 11696
rect 29588 11656 31468 11696
rect 31508 11656 35212 11696
rect 35252 11656 35261 11696
rect 38179 11656 38188 11696
rect 38228 11656 41644 11696
rect 41684 11656 41693 11696
rect 47299 11656 47308 11696
rect 47348 11656 48844 11696
rect 48884 11656 48893 11696
rect 32707 11572 32716 11612
rect 32756 11572 33100 11612
rect 33140 11572 33149 11612
rect 0 11528 80 11548
rect 0 11488 652 11528
rect 692 11488 701 11528
rect 42595 11488 42604 11528
rect 42644 11488 43084 11528
rect 43124 11488 43133 11528
rect 0 11468 80 11488
rect 4343 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 4729 11360
rect 19463 11320 19472 11360
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19840 11320 19849 11360
rect 21091 11320 21100 11360
rect 21140 11320 22636 11360
rect 22676 11320 22685 11360
rect 24835 11320 24844 11360
rect 24884 11320 28684 11360
rect 28724 11320 32332 11360
rect 32372 11320 32381 11360
rect 34583 11320 34592 11360
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34960 11320 34969 11360
rect 49703 11320 49712 11360
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 50080 11320 50089 11360
rect 64823 11320 64832 11360
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 65200 11320 65209 11360
rect 79943 11320 79952 11360
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 80320 11320 80329 11360
rect 95063 11320 95072 11360
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95440 11320 95449 11360
rect 30115 11152 30124 11192
rect 30164 11152 31372 11192
rect 31412 11152 32044 11192
rect 32084 11152 32093 11192
rect 37891 11152 37900 11192
rect 37940 11152 39148 11192
rect 39188 11152 43948 11192
rect 43988 11152 43997 11192
rect 31171 11068 31180 11108
rect 31220 11068 31948 11108
rect 31988 11068 31997 11108
rect 38275 11068 38284 11108
rect 38324 11068 40684 11108
rect 40724 11068 40733 11108
rect 44323 11068 44332 11108
rect 44372 11068 46636 11108
rect 46676 11068 46685 11108
rect 16483 10984 16492 11024
rect 16532 10984 17548 11024
rect 17588 10984 17597 11024
rect 21667 10984 21676 11024
rect 21716 10984 31564 11024
rect 31604 10984 38380 11024
rect 38420 10984 39052 11024
rect 39092 10984 39101 11024
rect 52579 10984 52588 11024
rect 52628 10984 53164 11024
rect 53204 10984 53213 11024
rect 23920 10732 30892 10772
rect 30932 10732 30941 10772
rect 39523 10732 39532 10772
rect 39572 10732 40492 10772
rect 40532 10732 40541 10772
rect 0 10688 80 10708
rect 23920 10688 23960 10732
rect 0 10648 652 10688
rect 692 10648 701 10688
rect 835 10648 844 10688
rect 884 10648 23960 10688
rect 0 10628 80 10648
rect 3103 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 3489 10604
rect 18223 10564 18232 10604
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18600 10564 18609 10604
rect 33343 10564 33352 10604
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33720 10564 33729 10604
rect 48463 10564 48472 10604
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48840 10564 48849 10604
rect 63583 10564 63592 10604
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63960 10564 63969 10604
rect 78703 10564 78712 10604
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 79080 10564 79089 10604
rect 93823 10564 93832 10604
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 94200 10564 94209 10604
rect 21955 10396 21964 10436
rect 22004 10396 23404 10436
rect 23444 10396 23453 10436
rect 2275 10312 2284 10352
rect 2324 10312 3148 10352
rect 3188 10312 3197 10352
rect 55459 10312 55468 10352
rect 55508 10312 55852 10352
rect 55892 10312 58828 10352
rect 58868 10312 58877 10352
rect 3331 10228 3340 10268
rect 3380 10228 4108 10268
rect 4148 10228 4157 10268
rect 12739 10228 12748 10268
rect 12788 10228 13132 10268
rect 13172 10228 18124 10268
rect 18164 10228 18173 10268
rect 59971 10228 59980 10268
rect 60020 10228 61132 10268
rect 61172 10228 61181 10268
rect 59980 10184 60020 10228
rect 14179 10144 14188 10184
rect 14228 10144 16492 10184
rect 16532 10144 16541 10184
rect 20995 10144 21004 10184
rect 21044 10144 21484 10184
rect 21524 10144 21868 10184
rect 21908 10144 21917 10184
rect 26851 10144 26860 10184
rect 26900 10144 28012 10184
rect 28052 10144 28204 10184
rect 28244 10144 28253 10184
rect 39043 10144 39052 10184
rect 39092 10144 53452 10184
rect 53492 10144 53501 10184
rect 55363 10144 55372 10184
rect 55412 10144 56428 10184
rect 56468 10144 58444 10184
rect 58484 10144 58493 10184
rect 58627 10144 58636 10184
rect 58676 10144 58685 10184
rect 59011 10144 59020 10184
rect 59060 10144 60020 10184
rect 61411 10144 61420 10184
rect 61460 10144 61996 10184
rect 62036 10144 62045 10184
rect 58636 10100 58676 10144
rect 10723 10060 10732 10100
rect 10772 10060 12652 10100
rect 12692 10060 13324 10100
rect 13364 10060 16684 10100
rect 16724 10060 17068 10100
rect 17108 10060 17117 10100
rect 28291 10060 28300 10100
rect 28340 10060 29740 10100
rect 29780 10060 29789 10100
rect 47203 10060 47212 10100
rect 47252 10060 48460 10100
rect 48500 10060 51724 10100
rect 51764 10060 52396 10100
rect 52436 10060 52445 10100
rect 58636 10060 59212 10100
rect 59252 10060 60748 10100
rect 60788 10060 60797 10100
rect 29827 9976 29836 10016
rect 29876 9976 31276 10016
rect 31316 9976 31325 10016
rect 54883 9976 54892 10016
rect 54932 9976 55468 10016
rect 55508 9976 55517 10016
rect 0 9848 80 9868
rect 0 9808 652 9848
rect 692 9808 701 9848
rect 4343 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 4729 9848
rect 19463 9808 19472 9848
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19840 9808 19849 9848
rect 34583 9808 34592 9848
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34960 9808 34969 9848
rect 49703 9808 49712 9848
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 50080 9808 50089 9848
rect 64823 9808 64832 9848
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 65200 9808 65209 9848
rect 79943 9808 79952 9848
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 80320 9808 80329 9848
rect 95063 9808 95072 9848
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95440 9808 95449 9848
rect 0 9788 80 9808
rect 9187 9640 9196 9680
rect 9236 9640 9868 9680
rect 9908 9640 9917 9680
rect 48067 9640 48076 9680
rect 48116 9640 49324 9680
rect 49364 9640 49373 9680
rect 6115 9472 6124 9512
rect 6164 9472 6796 9512
rect 6836 9472 6845 9512
rect 21571 9472 21580 9512
rect 21620 9472 21868 9512
rect 21908 9472 21917 9512
rect 33187 9472 33196 9512
rect 33236 9472 34444 9512
rect 34484 9472 34493 9512
rect 37123 9472 37132 9512
rect 37172 9472 38284 9512
rect 38324 9472 38333 9512
rect 54499 9472 54508 9512
rect 54548 9472 55660 9512
rect 55700 9472 59884 9512
rect 59924 9472 59933 9512
rect 36355 9304 36364 9344
rect 36404 9304 37132 9344
rect 37172 9304 37181 9344
rect 54115 9220 54124 9260
rect 54164 9220 54700 9260
rect 54740 9220 54749 9260
rect 3103 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3489 9092
rect 18223 9052 18232 9092
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18600 9052 18609 9092
rect 33343 9052 33352 9092
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33720 9052 33729 9092
rect 48463 9052 48472 9092
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48840 9052 48849 9092
rect 63583 9052 63592 9092
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63960 9052 63969 9092
rect 78703 9052 78712 9092
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 79080 9052 79089 9092
rect 93823 9052 93832 9092
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 94200 9052 94209 9092
rect 0 9008 80 9028
rect 0 8968 652 9008
rect 692 8968 701 9008
rect 0 8948 80 8968
rect 19075 8800 19084 8840
rect 19124 8800 20332 8840
rect 20372 8800 20381 8840
rect 27907 8800 27916 8840
rect 27956 8800 29644 8840
rect 29684 8800 29693 8840
rect 33283 8800 33292 8840
rect 33332 8800 34156 8840
rect 34196 8800 34205 8840
rect 55747 8800 55756 8840
rect 55796 8800 56428 8840
rect 56468 8800 56812 8840
rect 56852 8800 56861 8840
rect 44515 8716 44524 8756
rect 44564 8716 45676 8756
rect 45716 8716 47116 8756
rect 47156 8716 47165 8756
rect 55363 8716 55372 8756
rect 55412 8716 56524 8756
rect 56564 8716 56716 8756
rect 56756 8716 60844 8756
rect 60884 8716 60893 8756
rect 3523 8632 3532 8672
rect 3572 8632 4204 8672
rect 4244 8632 6604 8672
rect 6644 8632 6653 8672
rect 20611 8632 20620 8672
rect 20660 8632 23500 8672
rect 23540 8632 23549 8672
rect 24451 8632 24460 8672
rect 24500 8632 25708 8672
rect 25748 8632 25757 8672
rect 27331 8632 27340 8672
rect 27380 8632 27820 8672
rect 27860 8632 27869 8672
rect 29539 8632 29548 8672
rect 29588 8632 29597 8672
rect 33379 8632 33388 8672
rect 33428 8632 34156 8672
rect 34196 8632 34205 8672
rect 34531 8632 34540 8672
rect 34580 8632 35884 8672
rect 35924 8632 35933 8672
rect 29548 8588 29588 8632
rect 34540 8588 34580 8632
rect 25987 8548 25996 8588
rect 26036 8548 27244 8588
rect 27284 8548 29588 8588
rect 33187 8548 33196 8588
rect 33236 8548 33868 8588
rect 33908 8548 34580 8588
rect 40963 8548 40972 8588
rect 41012 8548 42124 8588
rect 42164 8548 42173 8588
rect 4343 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4729 8336
rect 19463 8296 19472 8336
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19840 8296 19849 8336
rect 34583 8296 34592 8336
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34960 8296 34969 8336
rect 49703 8296 49712 8336
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 50080 8296 50089 8336
rect 64823 8296 64832 8336
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 65200 8296 65209 8336
rect 79943 8296 79952 8336
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 80320 8296 80329 8336
rect 95063 8296 95072 8336
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95440 8296 95449 8336
rect 29155 8212 29164 8252
rect 29204 8212 33964 8252
rect 34004 8212 34013 8252
rect 0 8168 80 8188
rect 0 8128 556 8168
rect 596 8128 605 8168
rect 27619 8128 27628 8168
rect 27668 8128 28300 8168
rect 28340 8128 28349 8168
rect 32323 8128 32332 8168
rect 32372 8128 33100 8168
rect 33140 8128 33149 8168
rect 0 8108 80 8128
rect 30019 8044 30028 8084
rect 30068 8044 31660 8084
rect 31700 8044 31709 8084
rect 46723 8044 46732 8084
rect 46772 8044 48556 8084
rect 48596 8044 48605 8084
rect 4483 7960 4492 8000
rect 4532 7960 5932 8000
rect 5972 7960 5981 8000
rect 7555 7960 7564 8000
rect 7604 7960 9580 8000
rect 9620 7960 11212 8000
rect 11252 7960 11261 8000
rect 14755 7960 14764 8000
rect 14804 7960 15820 8000
rect 15860 7960 15869 8000
rect 18691 7960 18700 8000
rect 18740 7960 22348 8000
rect 22388 7960 22397 8000
rect 23203 7960 23212 8000
rect 23252 7960 23980 8000
rect 24020 7960 24268 8000
rect 24308 7960 24317 8000
rect 33763 7960 33772 8000
rect 33812 7960 34060 8000
rect 34100 7960 35692 8000
rect 35732 7960 35741 8000
rect 46627 7960 46636 8000
rect 46676 7960 47212 8000
rect 47252 7960 47261 8000
rect 22348 7916 22388 7960
rect 22348 7876 23404 7916
rect 23444 7876 23453 7916
rect 24355 7876 24364 7916
rect 24404 7876 25420 7916
rect 25460 7876 25900 7916
rect 25940 7876 25949 7916
rect 23395 7708 23404 7748
rect 23444 7708 24844 7748
rect 24884 7708 29644 7748
rect 29684 7708 29693 7748
rect 18115 7624 18124 7664
rect 18164 7624 19948 7664
rect 19988 7624 19997 7664
rect 3103 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3489 7580
rect 18223 7540 18232 7580
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18600 7540 18609 7580
rect 33343 7540 33352 7580
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33720 7540 33729 7580
rect 35299 7540 35308 7580
rect 35348 7540 37996 7580
rect 38036 7540 39916 7580
rect 39956 7540 39965 7580
rect 48463 7540 48472 7580
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48840 7540 48849 7580
rect 63583 7540 63592 7580
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63960 7540 63969 7580
rect 78703 7540 78712 7580
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 79080 7540 79089 7580
rect 93823 7540 93832 7580
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 94200 7540 94209 7580
rect 49315 7456 49324 7496
rect 49364 7456 51532 7496
rect 51572 7456 51581 7496
rect 11011 7372 11020 7412
rect 11060 7372 11500 7412
rect 11540 7372 11549 7412
rect 49219 7372 49228 7412
rect 49268 7372 50380 7412
rect 50420 7372 50429 7412
rect 0 7328 80 7348
rect 0 7288 652 7328
rect 692 7288 701 7328
rect 0 7268 80 7288
rect 38851 7204 38860 7244
rect 38900 7204 39532 7244
rect 39572 7204 39724 7244
rect 39764 7204 39773 7244
rect 12163 7120 12172 7160
rect 12212 7120 13516 7160
rect 13556 7120 13565 7160
rect 49795 7120 49804 7160
rect 49844 7120 53260 7160
rect 53300 7120 56428 7160
rect 56468 7120 56477 7160
rect 23011 7036 23020 7076
rect 23060 7036 28492 7076
rect 28532 7036 28541 7076
rect 4343 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4729 6824
rect 19463 6784 19472 6824
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19840 6784 19849 6824
rect 34583 6784 34592 6824
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34960 6784 34969 6824
rect 49703 6784 49712 6824
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 50080 6784 50089 6824
rect 64823 6784 64832 6824
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 65200 6784 65209 6824
rect 79943 6784 79952 6824
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 80320 6784 80329 6824
rect 95063 6784 95072 6824
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95440 6784 95449 6824
rect 4579 6616 4588 6656
rect 4628 6616 5644 6656
rect 5684 6616 5693 6656
rect 39523 6532 39532 6572
rect 39572 6532 40780 6572
rect 40820 6532 40829 6572
rect 0 6488 80 6508
rect 0 6448 652 6488
rect 692 6448 701 6488
rect 32740 6448 34348 6488
rect 34388 6448 34397 6488
rect 39139 6448 39148 6488
rect 39188 6448 43372 6488
rect 43412 6448 43421 6488
rect 46339 6448 46348 6488
rect 46388 6448 46732 6488
rect 46772 6448 46781 6488
rect 0 6428 80 6448
rect 32740 6404 32780 6448
rect 7171 6364 7180 6404
rect 7220 6364 10156 6404
rect 10196 6364 12172 6404
rect 12212 6364 12221 6404
rect 28771 6364 28780 6404
rect 28820 6364 32332 6404
rect 32372 6364 32780 6404
rect 7372 6320 7412 6364
rect 28972 6320 29012 6364
rect 7363 6280 7372 6320
rect 7412 6280 7421 6320
rect 10308 6280 10348 6320
rect 10388 6280 10397 6320
rect 28963 6280 28972 6320
rect 29012 6280 29021 6320
rect 46404 6280 46444 6320
rect 46484 6280 46493 6320
rect 10348 6236 10388 6280
rect 46444 6236 46484 6280
rect 9763 6196 9772 6236
rect 9812 6196 10388 6236
rect 17635 6196 17644 6236
rect 17684 6196 18124 6236
rect 18164 6196 18173 6236
rect 44611 6196 44620 6236
rect 44660 6196 46484 6236
rect 3103 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3489 6068
rect 18223 6028 18232 6068
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18600 6028 18609 6068
rect 33343 6028 33352 6068
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33720 6028 33729 6068
rect 48463 6028 48472 6068
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48840 6028 48849 6068
rect 63583 6028 63592 6068
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63960 6028 63969 6068
rect 78703 6028 78712 6068
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 79080 6028 79089 6068
rect 93823 6028 93832 6068
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 94200 6028 94209 6068
rect 33475 5860 33484 5900
rect 33524 5860 33964 5900
rect 34004 5860 34013 5900
rect 12163 5692 12172 5732
rect 12212 5692 13036 5732
rect 13076 5692 13085 5732
rect 16771 5692 16780 5732
rect 16820 5692 17068 5732
rect 17108 5692 18700 5732
rect 18740 5692 18749 5732
rect 0 5648 80 5668
rect 0 5608 652 5648
rect 692 5608 701 5648
rect 2755 5608 2764 5648
rect 2804 5608 2956 5648
rect 2996 5608 4492 5648
rect 4532 5608 4541 5648
rect 4771 5608 4780 5648
rect 4820 5608 5164 5648
rect 5204 5608 5213 5648
rect 17923 5608 17932 5648
rect 17972 5608 19660 5648
rect 19700 5608 19709 5648
rect 35971 5608 35980 5648
rect 36020 5608 36556 5648
rect 36596 5608 36605 5648
rect 37219 5608 37228 5648
rect 37268 5608 37420 5648
rect 37460 5608 39340 5648
rect 39380 5608 39389 5648
rect 47491 5608 47500 5648
rect 47540 5608 48940 5648
rect 48980 5608 48989 5648
rect 0 5588 80 5608
rect 39427 5524 39436 5564
rect 39476 5524 41068 5564
rect 41108 5524 41117 5564
rect 48739 5524 48748 5564
rect 48788 5524 49036 5564
rect 49076 5524 49085 5564
rect 5059 5440 5068 5480
rect 5108 5440 5548 5480
rect 5588 5440 5597 5480
rect 52099 5440 52108 5480
rect 52148 5440 53356 5480
rect 53396 5440 53405 5480
rect 4343 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4729 5312
rect 19463 5272 19472 5312
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19840 5272 19849 5312
rect 34583 5272 34592 5312
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34960 5272 34969 5312
rect 49703 5272 49712 5312
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 50080 5272 50089 5312
rect 64823 5272 64832 5312
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 65200 5272 65209 5312
rect 79943 5272 79952 5312
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 80320 5272 80329 5312
rect 95063 5272 95072 5312
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95440 5272 95449 5312
rect 49315 5104 49324 5144
rect 49364 5104 50092 5144
rect 50132 5104 52108 5144
rect 52148 5104 52157 5144
rect 5347 5020 5356 5060
rect 5396 5020 6988 5060
rect 7028 5020 7037 5060
rect 37603 5020 37612 5060
rect 37652 5020 38380 5060
rect 38420 5020 38429 5060
rect 50371 5020 50380 5060
rect 50420 5020 52780 5060
rect 52820 5020 52829 5060
rect 2467 4936 2476 4976
rect 2516 4936 5164 4976
rect 5204 4936 6892 4976
rect 6932 4936 8236 4976
rect 8276 4936 8285 4976
rect 28099 4936 28108 4976
rect 28148 4936 28588 4976
rect 28628 4936 31468 4976
rect 31508 4936 31517 4976
rect 53155 4936 53164 4976
rect 53204 4936 53452 4976
rect 53492 4936 55372 4976
rect 55412 4936 55421 4976
rect 2851 4852 2860 4892
rect 2900 4852 3340 4892
rect 3380 4852 4300 4892
rect 4340 4852 7372 4892
rect 7412 4852 7421 4892
rect 37123 4852 37132 4892
rect 37172 4852 39436 4892
rect 39476 4852 40204 4892
rect 40244 4852 40253 4892
rect 0 4808 80 4828
rect 0 4768 652 4808
rect 692 4768 701 4808
rect 0 4748 80 4768
rect 3103 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3489 4556
rect 18223 4516 18232 4556
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18600 4516 18609 4556
rect 33343 4516 33352 4556
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33720 4516 33729 4556
rect 48463 4516 48472 4556
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48840 4516 48849 4556
rect 63583 4516 63592 4556
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63960 4516 63969 4556
rect 78703 4516 78712 4556
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 79080 4516 79089 4556
rect 93823 4516 93832 4556
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 94200 4516 94209 4556
rect 26179 4348 26188 4388
rect 26228 4348 26860 4388
rect 26900 4348 26909 4388
rect 6280 4264 30796 4304
rect 30836 4264 30845 4304
rect 6280 4220 6320 4264
rect 835 4180 844 4220
rect 884 4180 6320 4220
rect 12931 4180 12940 4220
rect 12980 4180 16972 4220
rect 17012 4180 17684 4220
rect 17644 4136 17684 4180
rect 14179 4096 14188 4136
rect 14228 4096 16300 4136
rect 16340 4096 16349 4136
rect 17635 4096 17644 4136
rect 17684 4096 17693 4136
rect 21763 4096 21772 4136
rect 21812 4096 22924 4136
rect 22964 4096 22973 4136
rect 24259 4096 24268 4136
rect 24308 4096 25036 4136
rect 25076 4096 25900 4136
rect 25940 4096 25949 4136
rect 39427 4096 39436 4136
rect 39476 4096 40108 4136
rect 40148 4096 40684 4136
rect 40724 4096 41068 4136
rect 41108 4096 41117 4136
rect 41251 4096 41260 4136
rect 41300 4096 41644 4136
rect 41684 4096 41693 4136
rect 49603 4096 49612 4136
rect 49652 4096 50476 4136
rect 50516 4096 50525 4136
rect 17548 4012 18028 4052
rect 18068 4012 18077 4052
rect 0 3968 80 3988
rect 17548 3968 17588 4012
rect 0 3928 652 3968
rect 692 3928 701 3968
rect 11779 3928 11788 3968
rect 11828 3928 12748 3968
rect 12788 3928 12797 3968
rect 17539 3928 17548 3968
rect 17588 3928 17684 3968
rect 17827 3928 17836 3968
rect 17876 3928 19372 3968
rect 19412 3928 19421 3968
rect 31075 3928 31084 3968
rect 31124 3928 31660 3968
rect 31700 3928 31709 3968
rect 0 3908 80 3928
rect 17644 3884 17684 3928
rect 17635 3844 17644 3884
rect 17684 3844 17693 3884
rect 4343 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4729 3800
rect 17539 3760 17548 3800
rect 17588 3760 17932 3800
rect 17972 3760 17981 3800
rect 19463 3760 19472 3800
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19840 3760 19849 3800
rect 21667 3760 21676 3800
rect 21716 3760 24172 3800
rect 24212 3760 24221 3800
rect 34583 3760 34592 3800
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34960 3760 34969 3800
rect 49703 3760 49712 3800
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 50080 3760 50089 3800
rect 64823 3760 64832 3800
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 65200 3760 65209 3800
rect 79943 3760 79952 3800
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 80320 3760 80329 3800
rect 95063 3760 95072 3800
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95440 3760 95449 3800
rect 48739 3592 48748 3632
rect 48788 3592 49516 3632
rect 49556 3592 50379 3632
rect 50419 3592 50428 3632
rect 12163 3424 12172 3464
rect 12212 3424 12652 3464
rect 12692 3424 13132 3464
rect 13172 3424 13181 3464
rect 17539 3424 17548 3464
rect 17588 3424 20620 3464
rect 20660 3424 22156 3464
rect 22196 3424 22205 3464
rect 46435 3424 46444 3464
rect 46484 3424 46636 3464
rect 46676 3424 49132 3464
rect 49172 3424 49181 3464
rect 835 3340 844 3380
rect 884 3340 26956 3380
rect 26996 3340 27005 3380
rect 643 3172 652 3212
rect 692 3172 701 3212
rect 38083 3172 38092 3212
rect 38132 3172 39244 3212
rect 39284 3172 39293 3212
rect 42019 3172 42028 3212
rect 42068 3172 43084 3212
rect 43124 3172 43133 3212
rect 47587 3172 47596 3212
rect 47636 3172 48556 3212
rect 48596 3172 48605 3212
rect 0 3128 80 3148
rect 652 3128 692 3172
rect 0 3088 692 3128
rect 0 3068 80 3088
rect 3103 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3489 3044
rect 18223 3004 18232 3044
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18600 3004 18609 3044
rect 33343 3004 33352 3044
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33720 3004 33729 3044
rect 48463 3004 48472 3044
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48840 3004 48849 3044
rect 63583 3004 63592 3044
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63960 3004 63969 3044
rect 78703 3004 78712 3044
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 79080 3004 79089 3044
rect 93823 3004 93832 3044
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 94200 3004 94209 3044
rect 16291 2836 16300 2876
rect 16340 2836 16876 2876
rect 16916 2836 16925 2876
rect 44995 2836 45004 2876
rect 45044 2836 45772 2876
rect 45812 2836 45821 2876
rect 54019 2836 54028 2876
rect 54068 2836 54604 2876
rect 54644 2836 54653 2876
rect 17539 2752 17548 2792
rect 17588 2752 18988 2792
rect 19028 2752 19037 2792
rect 835 2668 844 2708
rect 884 2668 25324 2708
rect 25364 2668 25373 2708
rect 37987 2668 37996 2708
rect 38036 2668 38476 2708
rect 38516 2668 42700 2708
rect 42740 2668 42749 2708
rect 50563 2668 50572 2708
rect 50612 2668 51820 2708
rect 51860 2668 53356 2708
rect 53396 2668 53405 2708
rect 13603 2584 13612 2624
rect 13652 2584 15532 2624
rect 15572 2584 17452 2624
rect 17492 2584 17501 2624
rect 19171 2584 19180 2624
rect 19220 2584 20180 2624
rect 21283 2584 21292 2624
rect 21332 2584 21676 2624
rect 21716 2584 21725 2624
rect 24163 2584 24172 2624
rect 24212 2584 25036 2624
rect 25076 2584 28588 2624
rect 28628 2584 28637 2624
rect 39331 2584 39340 2624
rect 39380 2584 40204 2624
rect 40244 2584 41836 2624
rect 41876 2584 43468 2624
rect 43508 2584 46156 2624
rect 46196 2584 46205 2624
rect 47011 2584 47020 2624
rect 47060 2584 47980 2624
rect 48020 2584 48364 2624
rect 48404 2584 48413 2624
rect 20140 2540 20180 2584
rect 20140 2500 20908 2540
rect 20948 2500 20957 2540
rect 0 2288 80 2308
rect 0 2248 652 2288
rect 692 2248 701 2288
rect 4343 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4729 2288
rect 19463 2248 19472 2288
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19840 2248 19849 2288
rect 34583 2248 34592 2288
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34960 2248 34969 2288
rect 49703 2248 49712 2288
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 50080 2248 50089 2288
rect 64823 2248 64832 2288
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 65200 2248 65209 2288
rect 79943 2248 79952 2288
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 80320 2248 80329 2288
rect 95063 2248 95072 2288
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95440 2248 95449 2288
rect 0 2228 80 2248
rect 12259 2080 12268 2120
rect 12308 2080 13324 2120
rect 13364 2080 13373 2120
rect 3103 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3489 1532
rect 18223 1492 18232 1532
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18600 1492 18609 1532
rect 33343 1492 33352 1532
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33720 1492 33729 1532
rect 48463 1492 48472 1532
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48840 1492 48849 1532
rect 63583 1492 63592 1532
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63960 1492 63969 1532
rect 78703 1492 78712 1532
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 79080 1492 79089 1532
rect 93823 1492 93832 1532
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 94200 1492 94209 1532
rect 4343 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4729 776
rect 19463 736 19472 776
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19840 736 19849 776
rect 34583 736 34592 776
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34960 736 34969 776
rect 49703 736 49712 776
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 50080 736 50089 776
rect 64823 736 64832 776
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 65200 736 65209 776
rect 79943 736 79952 776
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 80320 736 80329 776
rect 95063 736 95072 776
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95440 736 95449 776
<< via3 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 35020 21988 35060 22028
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 35020 21652 35060 21692
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal4 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 19472 38576 19840 38585
rect 19512 38536 19554 38576
rect 19594 38536 19636 38576
rect 19676 38536 19718 38576
rect 19758 38536 19800 38576
rect 19472 38527 19840 38536
rect 34592 38576 34960 38585
rect 34632 38536 34674 38576
rect 34714 38536 34756 38576
rect 34796 38536 34838 38576
rect 34878 38536 34920 38576
rect 34592 38527 34960 38536
rect 49712 38576 50080 38585
rect 49752 38536 49794 38576
rect 49834 38536 49876 38576
rect 49916 38536 49958 38576
rect 49998 38536 50040 38576
rect 49712 38527 50080 38536
rect 64832 38576 65200 38585
rect 64872 38536 64914 38576
rect 64954 38536 64996 38576
rect 65036 38536 65078 38576
rect 65118 38536 65160 38576
rect 64832 38527 65200 38536
rect 79952 38576 80320 38585
rect 79992 38536 80034 38576
rect 80074 38536 80116 38576
rect 80156 38536 80198 38576
rect 80238 38536 80280 38576
rect 79952 38527 80320 38536
rect 95072 38576 95440 38585
rect 95112 38536 95154 38576
rect 95194 38536 95236 38576
rect 95276 38536 95318 38576
rect 95358 38536 95400 38576
rect 95072 38527 95440 38536
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 18232 37820 18600 37829
rect 18272 37780 18314 37820
rect 18354 37780 18396 37820
rect 18436 37780 18478 37820
rect 18518 37780 18560 37820
rect 18232 37771 18600 37780
rect 33352 37820 33720 37829
rect 33392 37780 33434 37820
rect 33474 37780 33516 37820
rect 33556 37780 33598 37820
rect 33638 37780 33680 37820
rect 33352 37771 33720 37780
rect 48472 37820 48840 37829
rect 48512 37780 48554 37820
rect 48594 37780 48636 37820
rect 48676 37780 48718 37820
rect 48758 37780 48800 37820
rect 48472 37771 48840 37780
rect 63592 37820 63960 37829
rect 63632 37780 63674 37820
rect 63714 37780 63756 37820
rect 63796 37780 63838 37820
rect 63878 37780 63920 37820
rect 63592 37771 63960 37780
rect 78712 37820 79080 37829
rect 78752 37780 78794 37820
rect 78834 37780 78876 37820
rect 78916 37780 78958 37820
rect 78998 37780 79040 37820
rect 78712 37771 79080 37780
rect 93832 37820 94200 37829
rect 93872 37780 93914 37820
rect 93954 37780 93996 37820
rect 94036 37780 94078 37820
rect 94118 37780 94160 37820
rect 93832 37771 94200 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 19472 37064 19840 37073
rect 19512 37024 19554 37064
rect 19594 37024 19636 37064
rect 19676 37024 19718 37064
rect 19758 37024 19800 37064
rect 19472 37015 19840 37024
rect 34592 37064 34960 37073
rect 34632 37024 34674 37064
rect 34714 37024 34756 37064
rect 34796 37024 34838 37064
rect 34878 37024 34920 37064
rect 34592 37015 34960 37024
rect 49712 37064 50080 37073
rect 49752 37024 49794 37064
rect 49834 37024 49876 37064
rect 49916 37024 49958 37064
rect 49998 37024 50040 37064
rect 49712 37015 50080 37024
rect 64832 37064 65200 37073
rect 64872 37024 64914 37064
rect 64954 37024 64996 37064
rect 65036 37024 65078 37064
rect 65118 37024 65160 37064
rect 64832 37015 65200 37024
rect 79952 37064 80320 37073
rect 79992 37024 80034 37064
rect 80074 37024 80116 37064
rect 80156 37024 80198 37064
rect 80238 37024 80280 37064
rect 79952 37015 80320 37024
rect 95072 37064 95440 37073
rect 95112 37024 95154 37064
rect 95194 37024 95236 37064
rect 95276 37024 95318 37064
rect 95358 37024 95400 37064
rect 95072 37015 95440 37024
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 18232 36308 18600 36317
rect 18272 36268 18314 36308
rect 18354 36268 18396 36308
rect 18436 36268 18478 36308
rect 18518 36268 18560 36308
rect 18232 36259 18600 36268
rect 33352 36308 33720 36317
rect 33392 36268 33434 36308
rect 33474 36268 33516 36308
rect 33556 36268 33598 36308
rect 33638 36268 33680 36308
rect 33352 36259 33720 36268
rect 48472 36308 48840 36317
rect 48512 36268 48554 36308
rect 48594 36268 48636 36308
rect 48676 36268 48718 36308
rect 48758 36268 48800 36308
rect 48472 36259 48840 36268
rect 63592 36308 63960 36317
rect 63632 36268 63674 36308
rect 63714 36268 63756 36308
rect 63796 36268 63838 36308
rect 63878 36268 63920 36308
rect 63592 36259 63960 36268
rect 78712 36308 79080 36317
rect 78752 36268 78794 36308
rect 78834 36268 78876 36308
rect 78916 36268 78958 36308
rect 78998 36268 79040 36308
rect 78712 36259 79080 36268
rect 93832 36308 94200 36317
rect 93872 36268 93914 36308
rect 93954 36268 93996 36308
rect 94036 36268 94078 36308
rect 94118 36268 94160 36308
rect 93832 36259 94200 36268
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 19472 35552 19840 35561
rect 19512 35512 19554 35552
rect 19594 35512 19636 35552
rect 19676 35512 19718 35552
rect 19758 35512 19800 35552
rect 19472 35503 19840 35512
rect 34592 35552 34960 35561
rect 34632 35512 34674 35552
rect 34714 35512 34756 35552
rect 34796 35512 34838 35552
rect 34878 35512 34920 35552
rect 34592 35503 34960 35512
rect 49712 35552 50080 35561
rect 49752 35512 49794 35552
rect 49834 35512 49876 35552
rect 49916 35512 49958 35552
rect 49998 35512 50040 35552
rect 49712 35503 50080 35512
rect 64832 35552 65200 35561
rect 64872 35512 64914 35552
rect 64954 35512 64996 35552
rect 65036 35512 65078 35552
rect 65118 35512 65160 35552
rect 64832 35503 65200 35512
rect 79952 35552 80320 35561
rect 79992 35512 80034 35552
rect 80074 35512 80116 35552
rect 80156 35512 80198 35552
rect 80238 35512 80280 35552
rect 79952 35503 80320 35512
rect 95072 35552 95440 35561
rect 95112 35512 95154 35552
rect 95194 35512 95236 35552
rect 95276 35512 95318 35552
rect 95358 35512 95400 35552
rect 95072 35503 95440 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 18232 34796 18600 34805
rect 18272 34756 18314 34796
rect 18354 34756 18396 34796
rect 18436 34756 18478 34796
rect 18518 34756 18560 34796
rect 18232 34747 18600 34756
rect 33352 34796 33720 34805
rect 33392 34756 33434 34796
rect 33474 34756 33516 34796
rect 33556 34756 33598 34796
rect 33638 34756 33680 34796
rect 33352 34747 33720 34756
rect 48472 34796 48840 34805
rect 48512 34756 48554 34796
rect 48594 34756 48636 34796
rect 48676 34756 48718 34796
rect 48758 34756 48800 34796
rect 48472 34747 48840 34756
rect 63592 34796 63960 34805
rect 63632 34756 63674 34796
rect 63714 34756 63756 34796
rect 63796 34756 63838 34796
rect 63878 34756 63920 34796
rect 63592 34747 63960 34756
rect 78712 34796 79080 34805
rect 78752 34756 78794 34796
rect 78834 34756 78876 34796
rect 78916 34756 78958 34796
rect 78998 34756 79040 34796
rect 78712 34747 79080 34756
rect 93832 34796 94200 34805
rect 93872 34756 93914 34796
rect 93954 34756 93996 34796
rect 94036 34756 94078 34796
rect 94118 34756 94160 34796
rect 93832 34747 94200 34756
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 19472 34040 19840 34049
rect 19512 34000 19554 34040
rect 19594 34000 19636 34040
rect 19676 34000 19718 34040
rect 19758 34000 19800 34040
rect 19472 33991 19840 34000
rect 34592 34040 34960 34049
rect 34632 34000 34674 34040
rect 34714 34000 34756 34040
rect 34796 34000 34838 34040
rect 34878 34000 34920 34040
rect 34592 33991 34960 34000
rect 49712 34040 50080 34049
rect 49752 34000 49794 34040
rect 49834 34000 49876 34040
rect 49916 34000 49958 34040
rect 49998 34000 50040 34040
rect 49712 33991 50080 34000
rect 64832 34040 65200 34049
rect 64872 34000 64914 34040
rect 64954 34000 64996 34040
rect 65036 34000 65078 34040
rect 65118 34000 65160 34040
rect 64832 33991 65200 34000
rect 79952 34040 80320 34049
rect 79992 34000 80034 34040
rect 80074 34000 80116 34040
rect 80156 34000 80198 34040
rect 80238 34000 80280 34040
rect 79952 33991 80320 34000
rect 95072 34040 95440 34049
rect 95112 34000 95154 34040
rect 95194 34000 95236 34040
rect 95276 34000 95318 34040
rect 95358 34000 95400 34040
rect 95072 33991 95440 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 18232 33284 18600 33293
rect 18272 33244 18314 33284
rect 18354 33244 18396 33284
rect 18436 33244 18478 33284
rect 18518 33244 18560 33284
rect 18232 33235 18600 33244
rect 33352 33284 33720 33293
rect 33392 33244 33434 33284
rect 33474 33244 33516 33284
rect 33556 33244 33598 33284
rect 33638 33244 33680 33284
rect 33352 33235 33720 33244
rect 48472 33284 48840 33293
rect 48512 33244 48554 33284
rect 48594 33244 48636 33284
rect 48676 33244 48718 33284
rect 48758 33244 48800 33284
rect 48472 33235 48840 33244
rect 63592 33284 63960 33293
rect 63632 33244 63674 33284
rect 63714 33244 63756 33284
rect 63796 33244 63838 33284
rect 63878 33244 63920 33284
rect 63592 33235 63960 33244
rect 78712 33284 79080 33293
rect 78752 33244 78794 33284
rect 78834 33244 78876 33284
rect 78916 33244 78958 33284
rect 78998 33244 79040 33284
rect 78712 33235 79080 33244
rect 93832 33284 94200 33293
rect 93872 33244 93914 33284
rect 93954 33244 93996 33284
rect 94036 33244 94078 33284
rect 94118 33244 94160 33284
rect 93832 33235 94200 33244
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 19472 32528 19840 32537
rect 19512 32488 19554 32528
rect 19594 32488 19636 32528
rect 19676 32488 19718 32528
rect 19758 32488 19800 32528
rect 19472 32479 19840 32488
rect 34592 32528 34960 32537
rect 34632 32488 34674 32528
rect 34714 32488 34756 32528
rect 34796 32488 34838 32528
rect 34878 32488 34920 32528
rect 34592 32479 34960 32488
rect 49712 32528 50080 32537
rect 49752 32488 49794 32528
rect 49834 32488 49876 32528
rect 49916 32488 49958 32528
rect 49998 32488 50040 32528
rect 49712 32479 50080 32488
rect 64832 32528 65200 32537
rect 64872 32488 64914 32528
rect 64954 32488 64996 32528
rect 65036 32488 65078 32528
rect 65118 32488 65160 32528
rect 64832 32479 65200 32488
rect 79952 32528 80320 32537
rect 79992 32488 80034 32528
rect 80074 32488 80116 32528
rect 80156 32488 80198 32528
rect 80238 32488 80280 32528
rect 79952 32479 80320 32488
rect 95072 32528 95440 32537
rect 95112 32488 95154 32528
rect 95194 32488 95236 32528
rect 95276 32488 95318 32528
rect 95358 32488 95400 32528
rect 95072 32479 95440 32488
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 18232 31772 18600 31781
rect 18272 31732 18314 31772
rect 18354 31732 18396 31772
rect 18436 31732 18478 31772
rect 18518 31732 18560 31772
rect 18232 31723 18600 31732
rect 33352 31772 33720 31781
rect 33392 31732 33434 31772
rect 33474 31732 33516 31772
rect 33556 31732 33598 31772
rect 33638 31732 33680 31772
rect 33352 31723 33720 31732
rect 48472 31772 48840 31781
rect 48512 31732 48554 31772
rect 48594 31732 48636 31772
rect 48676 31732 48718 31772
rect 48758 31732 48800 31772
rect 48472 31723 48840 31732
rect 63592 31772 63960 31781
rect 63632 31732 63674 31772
rect 63714 31732 63756 31772
rect 63796 31732 63838 31772
rect 63878 31732 63920 31772
rect 63592 31723 63960 31732
rect 78712 31772 79080 31781
rect 78752 31732 78794 31772
rect 78834 31732 78876 31772
rect 78916 31732 78958 31772
rect 78998 31732 79040 31772
rect 78712 31723 79080 31732
rect 93832 31772 94200 31781
rect 93872 31732 93914 31772
rect 93954 31732 93996 31772
rect 94036 31732 94078 31772
rect 94118 31732 94160 31772
rect 93832 31723 94200 31732
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 19472 31016 19840 31025
rect 19512 30976 19554 31016
rect 19594 30976 19636 31016
rect 19676 30976 19718 31016
rect 19758 30976 19800 31016
rect 19472 30967 19840 30976
rect 34592 31016 34960 31025
rect 34632 30976 34674 31016
rect 34714 30976 34756 31016
rect 34796 30976 34838 31016
rect 34878 30976 34920 31016
rect 34592 30967 34960 30976
rect 49712 31016 50080 31025
rect 49752 30976 49794 31016
rect 49834 30976 49876 31016
rect 49916 30976 49958 31016
rect 49998 30976 50040 31016
rect 49712 30967 50080 30976
rect 64832 31016 65200 31025
rect 64872 30976 64914 31016
rect 64954 30976 64996 31016
rect 65036 30976 65078 31016
rect 65118 30976 65160 31016
rect 64832 30967 65200 30976
rect 79952 31016 80320 31025
rect 79992 30976 80034 31016
rect 80074 30976 80116 31016
rect 80156 30976 80198 31016
rect 80238 30976 80280 31016
rect 79952 30967 80320 30976
rect 95072 31016 95440 31025
rect 95112 30976 95154 31016
rect 95194 30976 95236 31016
rect 95276 30976 95318 31016
rect 95358 30976 95400 31016
rect 95072 30967 95440 30976
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 18232 30260 18600 30269
rect 18272 30220 18314 30260
rect 18354 30220 18396 30260
rect 18436 30220 18478 30260
rect 18518 30220 18560 30260
rect 18232 30211 18600 30220
rect 33352 30260 33720 30269
rect 33392 30220 33434 30260
rect 33474 30220 33516 30260
rect 33556 30220 33598 30260
rect 33638 30220 33680 30260
rect 33352 30211 33720 30220
rect 48472 30260 48840 30269
rect 48512 30220 48554 30260
rect 48594 30220 48636 30260
rect 48676 30220 48718 30260
rect 48758 30220 48800 30260
rect 48472 30211 48840 30220
rect 63592 30260 63960 30269
rect 63632 30220 63674 30260
rect 63714 30220 63756 30260
rect 63796 30220 63838 30260
rect 63878 30220 63920 30260
rect 63592 30211 63960 30220
rect 78712 30260 79080 30269
rect 78752 30220 78794 30260
rect 78834 30220 78876 30260
rect 78916 30220 78958 30260
rect 78998 30220 79040 30260
rect 78712 30211 79080 30220
rect 93832 30260 94200 30269
rect 93872 30220 93914 30260
rect 93954 30220 93996 30260
rect 94036 30220 94078 30260
rect 94118 30220 94160 30260
rect 93832 30211 94200 30220
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 19472 29504 19840 29513
rect 19512 29464 19554 29504
rect 19594 29464 19636 29504
rect 19676 29464 19718 29504
rect 19758 29464 19800 29504
rect 19472 29455 19840 29464
rect 34592 29504 34960 29513
rect 34632 29464 34674 29504
rect 34714 29464 34756 29504
rect 34796 29464 34838 29504
rect 34878 29464 34920 29504
rect 34592 29455 34960 29464
rect 49712 29504 50080 29513
rect 49752 29464 49794 29504
rect 49834 29464 49876 29504
rect 49916 29464 49958 29504
rect 49998 29464 50040 29504
rect 49712 29455 50080 29464
rect 64832 29504 65200 29513
rect 64872 29464 64914 29504
rect 64954 29464 64996 29504
rect 65036 29464 65078 29504
rect 65118 29464 65160 29504
rect 64832 29455 65200 29464
rect 79952 29504 80320 29513
rect 79992 29464 80034 29504
rect 80074 29464 80116 29504
rect 80156 29464 80198 29504
rect 80238 29464 80280 29504
rect 79952 29455 80320 29464
rect 95072 29504 95440 29513
rect 95112 29464 95154 29504
rect 95194 29464 95236 29504
rect 95276 29464 95318 29504
rect 95358 29464 95400 29504
rect 95072 29455 95440 29464
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 18232 28748 18600 28757
rect 18272 28708 18314 28748
rect 18354 28708 18396 28748
rect 18436 28708 18478 28748
rect 18518 28708 18560 28748
rect 18232 28699 18600 28708
rect 33352 28748 33720 28757
rect 33392 28708 33434 28748
rect 33474 28708 33516 28748
rect 33556 28708 33598 28748
rect 33638 28708 33680 28748
rect 33352 28699 33720 28708
rect 48472 28748 48840 28757
rect 48512 28708 48554 28748
rect 48594 28708 48636 28748
rect 48676 28708 48718 28748
rect 48758 28708 48800 28748
rect 48472 28699 48840 28708
rect 63592 28748 63960 28757
rect 63632 28708 63674 28748
rect 63714 28708 63756 28748
rect 63796 28708 63838 28748
rect 63878 28708 63920 28748
rect 63592 28699 63960 28708
rect 78712 28748 79080 28757
rect 78752 28708 78794 28748
rect 78834 28708 78876 28748
rect 78916 28708 78958 28748
rect 78998 28708 79040 28748
rect 78712 28699 79080 28708
rect 93832 28748 94200 28757
rect 93872 28708 93914 28748
rect 93954 28708 93996 28748
rect 94036 28708 94078 28748
rect 94118 28708 94160 28748
rect 93832 28699 94200 28708
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 19472 27992 19840 28001
rect 19512 27952 19554 27992
rect 19594 27952 19636 27992
rect 19676 27952 19718 27992
rect 19758 27952 19800 27992
rect 19472 27943 19840 27952
rect 34592 27992 34960 28001
rect 34632 27952 34674 27992
rect 34714 27952 34756 27992
rect 34796 27952 34838 27992
rect 34878 27952 34920 27992
rect 34592 27943 34960 27952
rect 49712 27992 50080 28001
rect 49752 27952 49794 27992
rect 49834 27952 49876 27992
rect 49916 27952 49958 27992
rect 49998 27952 50040 27992
rect 49712 27943 50080 27952
rect 64832 27992 65200 28001
rect 64872 27952 64914 27992
rect 64954 27952 64996 27992
rect 65036 27952 65078 27992
rect 65118 27952 65160 27992
rect 64832 27943 65200 27952
rect 79952 27992 80320 28001
rect 79992 27952 80034 27992
rect 80074 27952 80116 27992
rect 80156 27952 80198 27992
rect 80238 27952 80280 27992
rect 79952 27943 80320 27952
rect 95072 27992 95440 28001
rect 95112 27952 95154 27992
rect 95194 27952 95236 27992
rect 95276 27952 95318 27992
rect 95358 27952 95400 27992
rect 95072 27943 95440 27952
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 18232 27236 18600 27245
rect 18272 27196 18314 27236
rect 18354 27196 18396 27236
rect 18436 27196 18478 27236
rect 18518 27196 18560 27236
rect 18232 27187 18600 27196
rect 33352 27236 33720 27245
rect 33392 27196 33434 27236
rect 33474 27196 33516 27236
rect 33556 27196 33598 27236
rect 33638 27196 33680 27236
rect 33352 27187 33720 27196
rect 48472 27236 48840 27245
rect 48512 27196 48554 27236
rect 48594 27196 48636 27236
rect 48676 27196 48718 27236
rect 48758 27196 48800 27236
rect 48472 27187 48840 27196
rect 63592 27236 63960 27245
rect 63632 27196 63674 27236
rect 63714 27196 63756 27236
rect 63796 27196 63838 27236
rect 63878 27196 63920 27236
rect 63592 27187 63960 27196
rect 78712 27236 79080 27245
rect 78752 27196 78794 27236
rect 78834 27196 78876 27236
rect 78916 27196 78958 27236
rect 78998 27196 79040 27236
rect 78712 27187 79080 27196
rect 93832 27236 94200 27245
rect 93872 27196 93914 27236
rect 93954 27196 93996 27236
rect 94036 27196 94078 27236
rect 94118 27196 94160 27236
rect 93832 27187 94200 27196
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 19472 26480 19840 26489
rect 19512 26440 19554 26480
rect 19594 26440 19636 26480
rect 19676 26440 19718 26480
rect 19758 26440 19800 26480
rect 19472 26431 19840 26440
rect 34592 26480 34960 26489
rect 34632 26440 34674 26480
rect 34714 26440 34756 26480
rect 34796 26440 34838 26480
rect 34878 26440 34920 26480
rect 34592 26431 34960 26440
rect 49712 26480 50080 26489
rect 49752 26440 49794 26480
rect 49834 26440 49876 26480
rect 49916 26440 49958 26480
rect 49998 26440 50040 26480
rect 49712 26431 50080 26440
rect 64832 26480 65200 26489
rect 64872 26440 64914 26480
rect 64954 26440 64996 26480
rect 65036 26440 65078 26480
rect 65118 26440 65160 26480
rect 64832 26431 65200 26440
rect 79952 26480 80320 26489
rect 79992 26440 80034 26480
rect 80074 26440 80116 26480
rect 80156 26440 80198 26480
rect 80238 26440 80280 26480
rect 79952 26431 80320 26440
rect 95072 26480 95440 26489
rect 95112 26440 95154 26480
rect 95194 26440 95236 26480
rect 95276 26440 95318 26480
rect 95358 26440 95400 26480
rect 95072 26431 95440 26440
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 18232 25724 18600 25733
rect 18272 25684 18314 25724
rect 18354 25684 18396 25724
rect 18436 25684 18478 25724
rect 18518 25684 18560 25724
rect 18232 25675 18600 25684
rect 33352 25724 33720 25733
rect 33392 25684 33434 25724
rect 33474 25684 33516 25724
rect 33556 25684 33598 25724
rect 33638 25684 33680 25724
rect 33352 25675 33720 25684
rect 48472 25724 48840 25733
rect 48512 25684 48554 25724
rect 48594 25684 48636 25724
rect 48676 25684 48718 25724
rect 48758 25684 48800 25724
rect 48472 25675 48840 25684
rect 63592 25724 63960 25733
rect 63632 25684 63674 25724
rect 63714 25684 63756 25724
rect 63796 25684 63838 25724
rect 63878 25684 63920 25724
rect 63592 25675 63960 25684
rect 78712 25724 79080 25733
rect 78752 25684 78794 25724
rect 78834 25684 78876 25724
rect 78916 25684 78958 25724
rect 78998 25684 79040 25724
rect 78712 25675 79080 25684
rect 93832 25724 94200 25733
rect 93872 25684 93914 25724
rect 93954 25684 93996 25724
rect 94036 25684 94078 25724
rect 94118 25684 94160 25724
rect 93832 25675 94200 25684
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 19472 24968 19840 24977
rect 19512 24928 19554 24968
rect 19594 24928 19636 24968
rect 19676 24928 19718 24968
rect 19758 24928 19800 24968
rect 19472 24919 19840 24928
rect 34592 24968 34960 24977
rect 34632 24928 34674 24968
rect 34714 24928 34756 24968
rect 34796 24928 34838 24968
rect 34878 24928 34920 24968
rect 34592 24919 34960 24928
rect 49712 24968 50080 24977
rect 49752 24928 49794 24968
rect 49834 24928 49876 24968
rect 49916 24928 49958 24968
rect 49998 24928 50040 24968
rect 49712 24919 50080 24928
rect 64832 24968 65200 24977
rect 64872 24928 64914 24968
rect 64954 24928 64996 24968
rect 65036 24928 65078 24968
rect 65118 24928 65160 24968
rect 64832 24919 65200 24928
rect 79952 24968 80320 24977
rect 79992 24928 80034 24968
rect 80074 24928 80116 24968
rect 80156 24928 80198 24968
rect 80238 24928 80280 24968
rect 79952 24919 80320 24928
rect 95072 24968 95440 24977
rect 95112 24928 95154 24968
rect 95194 24928 95236 24968
rect 95276 24928 95318 24968
rect 95358 24928 95400 24968
rect 95072 24919 95440 24928
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 18232 24212 18600 24221
rect 18272 24172 18314 24212
rect 18354 24172 18396 24212
rect 18436 24172 18478 24212
rect 18518 24172 18560 24212
rect 18232 24163 18600 24172
rect 33352 24212 33720 24221
rect 33392 24172 33434 24212
rect 33474 24172 33516 24212
rect 33556 24172 33598 24212
rect 33638 24172 33680 24212
rect 33352 24163 33720 24172
rect 48472 24212 48840 24221
rect 48512 24172 48554 24212
rect 48594 24172 48636 24212
rect 48676 24172 48718 24212
rect 48758 24172 48800 24212
rect 48472 24163 48840 24172
rect 63592 24212 63960 24221
rect 63632 24172 63674 24212
rect 63714 24172 63756 24212
rect 63796 24172 63838 24212
rect 63878 24172 63920 24212
rect 63592 24163 63960 24172
rect 78712 24212 79080 24221
rect 78752 24172 78794 24212
rect 78834 24172 78876 24212
rect 78916 24172 78958 24212
rect 78998 24172 79040 24212
rect 78712 24163 79080 24172
rect 93832 24212 94200 24221
rect 93872 24172 93914 24212
rect 93954 24172 93996 24212
rect 94036 24172 94078 24212
rect 94118 24172 94160 24212
rect 93832 24163 94200 24172
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 19472 23456 19840 23465
rect 19512 23416 19554 23456
rect 19594 23416 19636 23456
rect 19676 23416 19718 23456
rect 19758 23416 19800 23456
rect 19472 23407 19840 23416
rect 34592 23456 34960 23465
rect 34632 23416 34674 23456
rect 34714 23416 34756 23456
rect 34796 23416 34838 23456
rect 34878 23416 34920 23456
rect 34592 23407 34960 23416
rect 49712 23456 50080 23465
rect 49752 23416 49794 23456
rect 49834 23416 49876 23456
rect 49916 23416 49958 23456
rect 49998 23416 50040 23456
rect 49712 23407 50080 23416
rect 64832 23456 65200 23465
rect 64872 23416 64914 23456
rect 64954 23416 64996 23456
rect 65036 23416 65078 23456
rect 65118 23416 65160 23456
rect 64832 23407 65200 23416
rect 79952 23456 80320 23465
rect 79992 23416 80034 23456
rect 80074 23416 80116 23456
rect 80156 23416 80198 23456
rect 80238 23416 80280 23456
rect 79952 23407 80320 23416
rect 95072 23456 95440 23465
rect 95112 23416 95154 23456
rect 95194 23416 95236 23456
rect 95276 23416 95318 23456
rect 95358 23416 95400 23456
rect 95072 23407 95440 23416
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 18232 22700 18600 22709
rect 18272 22660 18314 22700
rect 18354 22660 18396 22700
rect 18436 22660 18478 22700
rect 18518 22660 18560 22700
rect 18232 22651 18600 22660
rect 33352 22700 33720 22709
rect 33392 22660 33434 22700
rect 33474 22660 33516 22700
rect 33556 22660 33598 22700
rect 33638 22660 33680 22700
rect 33352 22651 33720 22660
rect 48472 22700 48840 22709
rect 48512 22660 48554 22700
rect 48594 22660 48636 22700
rect 48676 22660 48718 22700
rect 48758 22660 48800 22700
rect 48472 22651 48840 22660
rect 63592 22700 63960 22709
rect 63632 22660 63674 22700
rect 63714 22660 63756 22700
rect 63796 22660 63838 22700
rect 63878 22660 63920 22700
rect 63592 22651 63960 22660
rect 78712 22700 79080 22709
rect 78752 22660 78794 22700
rect 78834 22660 78876 22700
rect 78916 22660 78958 22700
rect 78998 22660 79040 22700
rect 78712 22651 79080 22660
rect 93832 22700 94200 22709
rect 93872 22660 93914 22700
rect 93954 22660 93996 22700
rect 94036 22660 94078 22700
rect 94118 22660 94160 22700
rect 93832 22651 94200 22660
rect 35020 22028 35060 22037
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 19472 21944 19840 21953
rect 19512 21904 19554 21944
rect 19594 21904 19636 21944
rect 19676 21904 19718 21944
rect 19758 21904 19800 21944
rect 19472 21895 19840 21904
rect 34592 21944 34960 21953
rect 34632 21904 34674 21944
rect 34714 21904 34756 21944
rect 34796 21904 34838 21944
rect 34878 21904 34920 21944
rect 34592 21895 34960 21904
rect 35020 21692 35060 21988
rect 49712 21944 50080 21953
rect 49752 21904 49794 21944
rect 49834 21904 49876 21944
rect 49916 21904 49958 21944
rect 49998 21904 50040 21944
rect 49712 21895 50080 21904
rect 64832 21944 65200 21953
rect 64872 21904 64914 21944
rect 64954 21904 64996 21944
rect 65036 21904 65078 21944
rect 65118 21904 65160 21944
rect 64832 21895 65200 21904
rect 79952 21944 80320 21953
rect 79992 21904 80034 21944
rect 80074 21904 80116 21944
rect 80156 21904 80198 21944
rect 80238 21904 80280 21944
rect 79952 21895 80320 21904
rect 95072 21944 95440 21953
rect 95112 21904 95154 21944
rect 95194 21904 95236 21944
rect 95276 21904 95318 21944
rect 95358 21904 95400 21944
rect 95072 21895 95440 21904
rect 35020 21643 35060 21652
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 18232 21188 18600 21197
rect 18272 21148 18314 21188
rect 18354 21148 18396 21188
rect 18436 21148 18478 21188
rect 18518 21148 18560 21188
rect 18232 21139 18600 21148
rect 33352 21188 33720 21197
rect 33392 21148 33434 21188
rect 33474 21148 33516 21188
rect 33556 21148 33598 21188
rect 33638 21148 33680 21188
rect 33352 21139 33720 21148
rect 48472 21188 48840 21197
rect 48512 21148 48554 21188
rect 48594 21148 48636 21188
rect 48676 21148 48718 21188
rect 48758 21148 48800 21188
rect 48472 21139 48840 21148
rect 63592 21188 63960 21197
rect 63632 21148 63674 21188
rect 63714 21148 63756 21188
rect 63796 21148 63838 21188
rect 63878 21148 63920 21188
rect 63592 21139 63960 21148
rect 78712 21188 79080 21197
rect 78752 21148 78794 21188
rect 78834 21148 78876 21188
rect 78916 21148 78958 21188
rect 78998 21148 79040 21188
rect 78712 21139 79080 21148
rect 93832 21188 94200 21197
rect 93872 21148 93914 21188
rect 93954 21148 93996 21188
rect 94036 21148 94078 21188
rect 94118 21148 94160 21188
rect 93832 21139 94200 21148
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 19472 20432 19840 20441
rect 19512 20392 19554 20432
rect 19594 20392 19636 20432
rect 19676 20392 19718 20432
rect 19758 20392 19800 20432
rect 19472 20383 19840 20392
rect 34592 20432 34960 20441
rect 34632 20392 34674 20432
rect 34714 20392 34756 20432
rect 34796 20392 34838 20432
rect 34878 20392 34920 20432
rect 34592 20383 34960 20392
rect 49712 20432 50080 20441
rect 49752 20392 49794 20432
rect 49834 20392 49876 20432
rect 49916 20392 49958 20432
rect 49998 20392 50040 20432
rect 49712 20383 50080 20392
rect 64832 20432 65200 20441
rect 64872 20392 64914 20432
rect 64954 20392 64996 20432
rect 65036 20392 65078 20432
rect 65118 20392 65160 20432
rect 64832 20383 65200 20392
rect 79952 20432 80320 20441
rect 79992 20392 80034 20432
rect 80074 20392 80116 20432
rect 80156 20392 80198 20432
rect 80238 20392 80280 20432
rect 79952 20383 80320 20392
rect 95072 20432 95440 20441
rect 95112 20392 95154 20432
rect 95194 20392 95236 20432
rect 95276 20392 95318 20432
rect 95358 20392 95400 20432
rect 95072 20383 95440 20392
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 18232 19676 18600 19685
rect 18272 19636 18314 19676
rect 18354 19636 18396 19676
rect 18436 19636 18478 19676
rect 18518 19636 18560 19676
rect 18232 19627 18600 19636
rect 33352 19676 33720 19685
rect 33392 19636 33434 19676
rect 33474 19636 33516 19676
rect 33556 19636 33598 19676
rect 33638 19636 33680 19676
rect 33352 19627 33720 19636
rect 48472 19676 48840 19685
rect 48512 19636 48554 19676
rect 48594 19636 48636 19676
rect 48676 19636 48718 19676
rect 48758 19636 48800 19676
rect 48472 19627 48840 19636
rect 63592 19676 63960 19685
rect 63632 19636 63674 19676
rect 63714 19636 63756 19676
rect 63796 19636 63838 19676
rect 63878 19636 63920 19676
rect 63592 19627 63960 19636
rect 78712 19676 79080 19685
rect 78752 19636 78794 19676
rect 78834 19636 78876 19676
rect 78916 19636 78958 19676
rect 78998 19636 79040 19676
rect 78712 19627 79080 19636
rect 93832 19676 94200 19685
rect 93872 19636 93914 19676
rect 93954 19636 93996 19676
rect 94036 19636 94078 19676
rect 94118 19636 94160 19676
rect 93832 19627 94200 19636
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 19472 18920 19840 18929
rect 19512 18880 19554 18920
rect 19594 18880 19636 18920
rect 19676 18880 19718 18920
rect 19758 18880 19800 18920
rect 19472 18871 19840 18880
rect 34592 18920 34960 18929
rect 34632 18880 34674 18920
rect 34714 18880 34756 18920
rect 34796 18880 34838 18920
rect 34878 18880 34920 18920
rect 34592 18871 34960 18880
rect 49712 18920 50080 18929
rect 49752 18880 49794 18920
rect 49834 18880 49876 18920
rect 49916 18880 49958 18920
rect 49998 18880 50040 18920
rect 49712 18871 50080 18880
rect 64832 18920 65200 18929
rect 64872 18880 64914 18920
rect 64954 18880 64996 18920
rect 65036 18880 65078 18920
rect 65118 18880 65160 18920
rect 64832 18871 65200 18880
rect 79952 18920 80320 18929
rect 79992 18880 80034 18920
rect 80074 18880 80116 18920
rect 80156 18880 80198 18920
rect 80238 18880 80280 18920
rect 79952 18871 80320 18880
rect 95072 18920 95440 18929
rect 95112 18880 95154 18920
rect 95194 18880 95236 18920
rect 95276 18880 95318 18920
rect 95358 18880 95400 18920
rect 95072 18871 95440 18880
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 18232 18164 18600 18173
rect 18272 18124 18314 18164
rect 18354 18124 18396 18164
rect 18436 18124 18478 18164
rect 18518 18124 18560 18164
rect 18232 18115 18600 18124
rect 33352 18164 33720 18173
rect 33392 18124 33434 18164
rect 33474 18124 33516 18164
rect 33556 18124 33598 18164
rect 33638 18124 33680 18164
rect 33352 18115 33720 18124
rect 48472 18164 48840 18173
rect 48512 18124 48554 18164
rect 48594 18124 48636 18164
rect 48676 18124 48718 18164
rect 48758 18124 48800 18164
rect 48472 18115 48840 18124
rect 63592 18164 63960 18173
rect 63632 18124 63674 18164
rect 63714 18124 63756 18164
rect 63796 18124 63838 18164
rect 63878 18124 63920 18164
rect 63592 18115 63960 18124
rect 78712 18164 79080 18173
rect 78752 18124 78794 18164
rect 78834 18124 78876 18164
rect 78916 18124 78958 18164
rect 78998 18124 79040 18164
rect 78712 18115 79080 18124
rect 93832 18164 94200 18173
rect 93872 18124 93914 18164
rect 93954 18124 93996 18164
rect 94036 18124 94078 18164
rect 94118 18124 94160 18164
rect 93832 18115 94200 18124
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 19472 17408 19840 17417
rect 19512 17368 19554 17408
rect 19594 17368 19636 17408
rect 19676 17368 19718 17408
rect 19758 17368 19800 17408
rect 19472 17359 19840 17368
rect 34592 17408 34960 17417
rect 34632 17368 34674 17408
rect 34714 17368 34756 17408
rect 34796 17368 34838 17408
rect 34878 17368 34920 17408
rect 34592 17359 34960 17368
rect 49712 17408 50080 17417
rect 49752 17368 49794 17408
rect 49834 17368 49876 17408
rect 49916 17368 49958 17408
rect 49998 17368 50040 17408
rect 49712 17359 50080 17368
rect 64832 17408 65200 17417
rect 64872 17368 64914 17408
rect 64954 17368 64996 17408
rect 65036 17368 65078 17408
rect 65118 17368 65160 17408
rect 64832 17359 65200 17368
rect 79952 17408 80320 17417
rect 79992 17368 80034 17408
rect 80074 17368 80116 17408
rect 80156 17368 80198 17408
rect 80238 17368 80280 17408
rect 79952 17359 80320 17368
rect 95072 17408 95440 17417
rect 95112 17368 95154 17408
rect 95194 17368 95236 17408
rect 95276 17368 95318 17408
rect 95358 17368 95400 17408
rect 95072 17359 95440 17368
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 18232 16652 18600 16661
rect 18272 16612 18314 16652
rect 18354 16612 18396 16652
rect 18436 16612 18478 16652
rect 18518 16612 18560 16652
rect 18232 16603 18600 16612
rect 33352 16652 33720 16661
rect 33392 16612 33434 16652
rect 33474 16612 33516 16652
rect 33556 16612 33598 16652
rect 33638 16612 33680 16652
rect 33352 16603 33720 16612
rect 48472 16652 48840 16661
rect 48512 16612 48554 16652
rect 48594 16612 48636 16652
rect 48676 16612 48718 16652
rect 48758 16612 48800 16652
rect 48472 16603 48840 16612
rect 63592 16652 63960 16661
rect 63632 16612 63674 16652
rect 63714 16612 63756 16652
rect 63796 16612 63838 16652
rect 63878 16612 63920 16652
rect 63592 16603 63960 16612
rect 78712 16652 79080 16661
rect 78752 16612 78794 16652
rect 78834 16612 78876 16652
rect 78916 16612 78958 16652
rect 78998 16612 79040 16652
rect 78712 16603 79080 16612
rect 93832 16652 94200 16661
rect 93872 16612 93914 16652
rect 93954 16612 93996 16652
rect 94036 16612 94078 16652
rect 94118 16612 94160 16652
rect 93832 16603 94200 16612
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 19472 15896 19840 15905
rect 19512 15856 19554 15896
rect 19594 15856 19636 15896
rect 19676 15856 19718 15896
rect 19758 15856 19800 15896
rect 19472 15847 19840 15856
rect 34592 15896 34960 15905
rect 34632 15856 34674 15896
rect 34714 15856 34756 15896
rect 34796 15856 34838 15896
rect 34878 15856 34920 15896
rect 34592 15847 34960 15856
rect 49712 15896 50080 15905
rect 49752 15856 49794 15896
rect 49834 15856 49876 15896
rect 49916 15856 49958 15896
rect 49998 15856 50040 15896
rect 49712 15847 50080 15856
rect 64832 15896 65200 15905
rect 64872 15856 64914 15896
rect 64954 15856 64996 15896
rect 65036 15856 65078 15896
rect 65118 15856 65160 15896
rect 64832 15847 65200 15856
rect 79952 15896 80320 15905
rect 79992 15856 80034 15896
rect 80074 15856 80116 15896
rect 80156 15856 80198 15896
rect 80238 15856 80280 15896
rect 79952 15847 80320 15856
rect 95072 15896 95440 15905
rect 95112 15856 95154 15896
rect 95194 15856 95236 15896
rect 95276 15856 95318 15896
rect 95358 15856 95400 15896
rect 95072 15847 95440 15856
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 18232 15140 18600 15149
rect 18272 15100 18314 15140
rect 18354 15100 18396 15140
rect 18436 15100 18478 15140
rect 18518 15100 18560 15140
rect 18232 15091 18600 15100
rect 33352 15140 33720 15149
rect 33392 15100 33434 15140
rect 33474 15100 33516 15140
rect 33556 15100 33598 15140
rect 33638 15100 33680 15140
rect 33352 15091 33720 15100
rect 48472 15140 48840 15149
rect 48512 15100 48554 15140
rect 48594 15100 48636 15140
rect 48676 15100 48718 15140
rect 48758 15100 48800 15140
rect 48472 15091 48840 15100
rect 63592 15140 63960 15149
rect 63632 15100 63674 15140
rect 63714 15100 63756 15140
rect 63796 15100 63838 15140
rect 63878 15100 63920 15140
rect 63592 15091 63960 15100
rect 78712 15140 79080 15149
rect 78752 15100 78794 15140
rect 78834 15100 78876 15140
rect 78916 15100 78958 15140
rect 78998 15100 79040 15140
rect 78712 15091 79080 15100
rect 93832 15140 94200 15149
rect 93872 15100 93914 15140
rect 93954 15100 93996 15140
rect 94036 15100 94078 15140
rect 94118 15100 94160 15140
rect 93832 15091 94200 15100
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 19472 14384 19840 14393
rect 19512 14344 19554 14384
rect 19594 14344 19636 14384
rect 19676 14344 19718 14384
rect 19758 14344 19800 14384
rect 19472 14335 19840 14344
rect 34592 14384 34960 14393
rect 34632 14344 34674 14384
rect 34714 14344 34756 14384
rect 34796 14344 34838 14384
rect 34878 14344 34920 14384
rect 34592 14335 34960 14344
rect 49712 14384 50080 14393
rect 49752 14344 49794 14384
rect 49834 14344 49876 14384
rect 49916 14344 49958 14384
rect 49998 14344 50040 14384
rect 49712 14335 50080 14344
rect 64832 14384 65200 14393
rect 64872 14344 64914 14384
rect 64954 14344 64996 14384
rect 65036 14344 65078 14384
rect 65118 14344 65160 14384
rect 64832 14335 65200 14344
rect 79952 14384 80320 14393
rect 79992 14344 80034 14384
rect 80074 14344 80116 14384
rect 80156 14344 80198 14384
rect 80238 14344 80280 14384
rect 79952 14335 80320 14344
rect 95072 14384 95440 14393
rect 95112 14344 95154 14384
rect 95194 14344 95236 14384
rect 95276 14344 95318 14384
rect 95358 14344 95400 14384
rect 95072 14335 95440 14344
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 18232 13628 18600 13637
rect 18272 13588 18314 13628
rect 18354 13588 18396 13628
rect 18436 13588 18478 13628
rect 18518 13588 18560 13628
rect 18232 13579 18600 13588
rect 33352 13628 33720 13637
rect 33392 13588 33434 13628
rect 33474 13588 33516 13628
rect 33556 13588 33598 13628
rect 33638 13588 33680 13628
rect 33352 13579 33720 13588
rect 48472 13628 48840 13637
rect 48512 13588 48554 13628
rect 48594 13588 48636 13628
rect 48676 13588 48718 13628
rect 48758 13588 48800 13628
rect 48472 13579 48840 13588
rect 63592 13628 63960 13637
rect 63632 13588 63674 13628
rect 63714 13588 63756 13628
rect 63796 13588 63838 13628
rect 63878 13588 63920 13628
rect 63592 13579 63960 13588
rect 78712 13628 79080 13637
rect 78752 13588 78794 13628
rect 78834 13588 78876 13628
rect 78916 13588 78958 13628
rect 78998 13588 79040 13628
rect 78712 13579 79080 13588
rect 93832 13628 94200 13637
rect 93872 13588 93914 13628
rect 93954 13588 93996 13628
rect 94036 13588 94078 13628
rect 94118 13588 94160 13628
rect 93832 13579 94200 13588
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 19472 12872 19840 12881
rect 19512 12832 19554 12872
rect 19594 12832 19636 12872
rect 19676 12832 19718 12872
rect 19758 12832 19800 12872
rect 19472 12823 19840 12832
rect 34592 12872 34960 12881
rect 34632 12832 34674 12872
rect 34714 12832 34756 12872
rect 34796 12832 34838 12872
rect 34878 12832 34920 12872
rect 34592 12823 34960 12832
rect 49712 12872 50080 12881
rect 49752 12832 49794 12872
rect 49834 12832 49876 12872
rect 49916 12832 49958 12872
rect 49998 12832 50040 12872
rect 49712 12823 50080 12832
rect 64832 12872 65200 12881
rect 64872 12832 64914 12872
rect 64954 12832 64996 12872
rect 65036 12832 65078 12872
rect 65118 12832 65160 12872
rect 64832 12823 65200 12832
rect 79952 12872 80320 12881
rect 79992 12832 80034 12872
rect 80074 12832 80116 12872
rect 80156 12832 80198 12872
rect 80238 12832 80280 12872
rect 79952 12823 80320 12832
rect 95072 12872 95440 12881
rect 95112 12832 95154 12872
rect 95194 12832 95236 12872
rect 95276 12832 95318 12872
rect 95358 12832 95400 12872
rect 95072 12823 95440 12832
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 18232 12116 18600 12125
rect 18272 12076 18314 12116
rect 18354 12076 18396 12116
rect 18436 12076 18478 12116
rect 18518 12076 18560 12116
rect 18232 12067 18600 12076
rect 33352 12116 33720 12125
rect 33392 12076 33434 12116
rect 33474 12076 33516 12116
rect 33556 12076 33598 12116
rect 33638 12076 33680 12116
rect 33352 12067 33720 12076
rect 48472 12116 48840 12125
rect 48512 12076 48554 12116
rect 48594 12076 48636 12116
rect 48676 12076 48718 12116
rect 48758 12076 48800 12116
rect 48472 12067 48840 12076
rect 63592 12116 63960 12125
rect 63632 12076 63674 12116
rect 63714 12076 63756 12116
rect 63796 12076 63838 12116
rect 63878 12076 63920 12116
rect 63592 12067 63960 12076
rect 78712 12116 79080 12125
rect 78752 12076 78794 12116
rect 78834 12076 78876 12116
rect 78916 12076 78958 12116
rect 78998 12076 79040 12116
rect 78712 12067 79080 12076
rect 93832 12116 94200 12125
rect 93872 12076 93914 12116
rect 93954 12076 93996 12116
rect 94036 12076 94078 12116
rect 94118 12076 94160 12116
rect 93832 12067 94200 12076
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 19472 11360 19840 11369
rect 19512 11320 19554 11360
rect 19594 11320 19636 11360
rect 19676 11320 19718 11360
rect 19758 11320 19800 11360
rect 19472 11311 19840 11320
rect 34592 11360 34960 11369
rect 34632 11320 34674 11360
rect 34714 11320 34756 11360
rect 34796 11320 34838 11360
rect 34878 11320 34920 11360
rect 34592 11311 34960 11320
rect 49712 11360 50080 11369
rect 49752 11320 49794 11360
rect 49834 11320 49876 11360
rect 49916 11320 49958 11360
rect 49998 11320 50040 11360
rect 49712 11311 50080 11320
rect 64832 11360 65200 11369
rect 64872 11320 64914 11360
rect 64954 11320 64996 11360
rect 65036 11320 65078 11360
rect 65118 11320 65160 11360
rect 64832 11311 65200 11320
rect 79952 11360 80320 11369
rect 79992 11320 80034 11360
rect 80074 11320 80116 11360
rect 80156 11320 80198 11360
rect 80238 11320 80280 11360
rect 79952 11311 80320 11320
rect 95072 11360 95440 11369
rect 95112 11320 95154 11360
rect 95194 11320 95236 11360
rect 95276 11320 95318 11360
rect 95358 11320 95400 11360
rect 95072 11311 95440 11320
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 18232 10604 18600 10613
rect 18272 10564 18314 10604
rect 18354 10564 18396 10604
rect 18436 10564 18478 10604
rect 18518 10564 18560 10604
rect 18232 10555 18600 10564
rect 33352 10604 33720 10613
rect 33392 10564 33434 10604
rect 33474 10564 33516 10604
rect 33556 10564 33598 10604
rect 33638 10564 33680 10604
rect 33352 10555 33720 10564
rect 48472 10604 48840 10613
rect 48512 10564 48554 10604
rect 48594 10564 48636 10604
rect 48676 10564 48718 10604
rect 48758 10564 48800 10604
rect 48472 10555 48840 10564
rect 63592 10604 63960 10613
rect 63632 10564 63674 10604
rect 63714 10564 63756 10604
rect 63796 10564 63838 10604
rect 63878 10564 63920 10604
rect 63592 10555 63960 10564
rect 78712 10604 79080 10613
rect 78752 10564 78794 10604
rect 78834 10564 78876 10604
rect 78916 10564 78958 10604
rect 78998 10564 79040 10604
rect 78712 10555 79080 10564
rect 93832 10604 94200 10613
rect 93872 10564 93914 10604
rect 93954 10564 93996 10604
rect 94036 10564 94078 10604
rect 94118 10564 94160 10604
rect 93832 10555 94200 10564
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 19472 9848 19840 9857
rect 19512 9808 19554 9848
rect 19594 9808 19636 9848
rect 19676 9808 19718 9848
rect 19758 9808 19800 9848
rect 19472 9799 19840 9808
rect 34592 9848 34960 9857
rect 34632 9808 34674 9848
rect 34714 9808 34756 9848
rect 34796 9808 34838 9848
rect 34878 9808 34920 9848
rect 34592 9799 34960 9808
rect 49712 9848 50080 9857
rect 49752 9808 49794 9848
rect 49834 9808 49876 9848
rect 49916 9808 49958 9848
rect 49998 9808 50040 9848
rect 49712 9799 50080 9808
rect 64832 9848 65200 9857
rect 64872 9808 64914 9848
rect 64954 9808 64996 9848
rect 65036 9808 65078 9848
rect 65118 9808 65160 9848
rect 64832 9799 65200 9808
rect 79952 9848 80320 9857
rect 79992 9808 80034 9848
rect 80074 9808 80116 9848
rect 80156 9808 80198 9848
rect 80238 9808 80280 9848
rect 79952 9799 80320 9808
rect 95072 9848 95440 9857
rect 95112 9808 95154 9848
rect 95194 9808 95236 9848
rect 95276 9808 95318 9848
rect 95358 9808 95400 9848
rect 95072 9799 95440 9808
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 18232 9092 18600 9101
rect 18272 9052 18314 9092
rect 18354 9052 18396 9092
rect 18436 9052 18478 9092
rect 18518 9052 18560 9092
rect 18232 9043 18600 9052
rect 33352 9092 33720 9101
rect 33392 9052 33434 9092
rect 33474 9052 33516 9092
rect 33556 9052 33598 9092
rect 33638 9052 33680 9092
rect 33352 9043 33720 9052
rect 48472 9092 48840 9101
rect 48512 9052 48554 9092
rect 48594 9052 48636 9092
rect 48676 9052 48718 9092
rect 48758 9052 48800 9092
rect 48472 9043 48840 9052
rect 63592 9092 63960 9101
rect 63632 9052 63674 9092
rect 63714 9052 63756 9092
rect 63796 9052 63838 9092
rect 63878 9052 63920 9092
rect 63592 9043 63960 9052
rect 78712 9092 79080 9101
rect 78752 9052 78794 9092
rect 78834 9052 78876 9092
rect 78916 9052 78958 9092
rect 78998 9052 79040 9092
rect 78712 9043 79080 9052
rect 93832 9092 94200 9101
rect 93872 9052 93914 9092
rect 93954 9052 93996 9092
rect 94036 9052 94078 9092
rect 94118 9052 94160 9092
rect 93832 9043 94200 9052
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 19472 8336 19840 8345
rect 19512 8296 19554 8336
rect 19594 8296 19636 8336
rect 19676 8296 19718 8336
rect 19758 8296 19800 8336
rect 19472 8287 19840 8296
rect 34592 8336 34960 8345
rect 34632 8296 34674 8336
rect 34714 8296 34756 8336
rect 34796 8296 34838 8336
rect 34878 8296 34920 8336
rect 34592 8287 34960 8296
rect 49712 8336 50080 8345
rect 49752 8296 49794 8336
rect 49834 8296 49876 8336
rect 49916 8296 49958 8336
rect 49998 8296 50040 8336
rect 49712 8287 50080 8296
rect 64832 8336 65200 8345
rect 64872 8296 64914 8336
rect 64954 8296 64996 8336
rect 65036 8296 65078 8336
rect 65118 8296 65160 8336
rect 64832 8287 65200 8296
rect 79952 8336 80320 8345
rect 79992 8296 80034 8336
rect 80074 8296 80116 8336
rect 80156 8296 80198 8336
rect 80238 8296 80280 8336
rect 79952 8287 80320 8296
rect 95072 8336 95440 8345
rect 95112 8296 95154 8336
rect 95194 8296 95236 8336
rect 95276 8296 95318 8336
rect 95358 8296 95400 8336
rect 95072 8287 95440 8296
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 18232 7580 18600 7589
rect 18272 7540 18314 7580
rect 18354 7540 18396 7580
rect 18436 7540 18478 7580
rect 18518 7540 18560 7580
rect 18232 7531 18600 7540
rect 33352 7580 33720 7589
rect 33392 7540 33434 7580
rect 33474 7540 33516 7580
rect 33556 7540 33598 7580
rect 33638 7540 33680 7580
rect 33352 7531 33720 7540
rect 48472 7580 48840 7589
rect 48512 7540 48554 7580
rect 48594 7540 48636 7580
rect 48676 7540 48718 7580
rect 48758 7540 48800 7580
rect 48472 7531 48840 7540
rect 63592 7580 63960 7589
rect 63632 7540 63674 7580
rect 63714 7540 63756 7580
rect 63796 7540 63838 7580
rect 63878 7540 63920 7580
rect 63592 7531 63960 7540
rect 78712 7580 79080 7589
rect 78752 7540 78794 7580
rect 78834 7540 78876 7580
rect 78916 7540 78958 7580
rect 78998 7540 79040 7580
rect 78712 7531 79080 7540
rect 93832 7580 94200 7589
rect 93872 7540 93914 7580
rect 93954 7540 93996 7580
rect 94036 7540 94078 7580
rect 94118 7540 94160 7580
rect 93832 7531 94200 7540
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 19472 6824 19840 6833
rect 19512 6784 19554 6824
rect 19594 6784 19636 6824
rect 19676 6784 19718 6824
rect 19758 6784 19800 6824
rect 19472 6775 19840 6784
rect 34592 6824 34960 6833
rect 34632 6784 34674 6824
rect 34714 6784 34756 6824
rect 34796 6784 34838 6824
rect 34878 6784 34920 6824
rect 34592 6775 34960 6784
rect 49712 6824 50080 6833
rect 49752 6784 49794 6824
rect 49834 6784 49876 6824
rect 49916 6784 49958 6824
rect 49998 6784 50040 6824
rect 49712 6775 50080 6784
rect 64832 6824 65200 6833
rect 64872 6784 64914 6824
rect 64954 6784 64996 6824
rect 65036 6784 65078 6824
rect 65118 6784 65160 6824
rect 64832 6775 65200 6784
rect 79952 6824 80320 6833
rect 79992 6784 80034 6824
rect 80074 6784 80116 6824
rect 80156 6784 80198 6824
rect 80238 6784 80280 6824
rect 79952 6775 80320 6784
rect 95072 6824 95440 6833
rect 95112 6784 95154 6824
rect 95194 6784 95236 6824
rect 95276 6784 95318 6824
rect 95358 6784 95400 6824
rect 95072 6775 95440 6784
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 18232 6068 18600 6077
rect 18272 6028 18314 6068
rect 18354 6028 18396 6068
rect 18436 6028 18478 6068
rect 18518 6028 18560 6068
rect 18232 6019 18600 6028
rect 33352 6068 33720 6077
rect 33392 6028 33434 6068
rect 33474 6028 33516 6068
rect 33556 6028 33598 6068
rect 33638 6028 33680 6068
rect 33352 6019 33720 6028
rect 48472 6068 48840 6077
rect 48512 6028 48554 6068
rect 48594 6028 48636 6068
rect 48676 6028 48718 6068
rect 48758 6028 48800 6068
rect 48472 6019 48840 6028
rect 63592 6068 63960 6077
rect 63632 6028 63674 6068
rect 63714 6028 63756 6068
rect 63796 6028 63838 6068
rect 63878 6028 63920 6068
rect 63592 6019 63960 6028
rect 78712 6068 79080 6077
rect 78752 6028 78794 6068
rect 78834 6028 78876 6068
rect 78916 6028 78958 6068
rect 78998 6028 79040 6068
rect 78712 6019 79080 6028
rect 93832 6068 94200 6077
rect 93872 6028 93914 6068
rect 93954 6028 93996 6068
rect 94036 6028 94078 6068
rect 94118 6028 94160 6068
rect 93832 6019 94200 6028
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 19472 5312 19840 5321
rect 19512 5272 19554 5312
rect 19594 5272 19636 5312
rect 19676 5272 19718 5312
rect 19758 5272 19800 5312
rect 19472 5263 19840 5272
rect 34592 5312 34960 5321
rect 34632 5272 34674 5312
rect 34714 5272 34756 5312
rect 34796 5272 34838 5312
rect 34878 5272 34920 5312
rect 34592 5263 34960 5272
rect 49712 5312 50080 5321
rect 49752 5272 49794 5312
rect 49834 5272 49876 5312
rect 49916 5272 49958 5312
rect 49998 5272 50040 5312
rect 49712 5263 50080 5272
rect 64832 5312 65200 5321
rect 64872 5272 64914 5312
rect 64954 5272 64996 5312
rect 65036 5272 65078 5312
rect 65118 5272 65160 5312
rect 64832 5263 65200 5272
rect 79952 5312 80320 5321
rect 79992 5272 80034 5312
rect 80074 5272 80116 5312
rect 80156 5272 80198 5312
rect 80238 5272 80280 5312
rect 79952 5263 80320 5272
rect 95072 5312 95440 5321
rect 95112 5272 95154 5312
rect 95194 5272 95236 5312
rect 95276 5272 95318 5312
rect 95358 5272 95400 5312
rect 95072 5263 95440 5272
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 18232 4556 18600 4565
rect 18272 4516 18314 4556
rect 18354 4516 18396 4556
rect 18436 4516 18478 4556
rect 18518 4516 18560 4556
rect 18232 4507 18600 4516
rect 33352 4556 33720 4565
rect 33392 4516 33434 4556
rect 33474 4516 33516 4556
rect 33556 4516 33598 4556
rect 33638 4516 33680 4556
rect 33352 4507 33720 4516
rect 48472 4556 48840 4565
rect 48512 4516 48554 4556
rect 48594 4516 48636 4556
rect 48676 4516 48718 4556
rect 48758 4516 48800 4556
rect 48472 4507 48840 4516
rect 63592 4556 63960 4565
rect 63632 4516 63674 4556
rect 63714 4516 63756 4556
rect 63796 4516 63838 4556
rect 63878 4516 63920 4556
rect 63592 4507 63960 4516
rect 78712 4556 79080 4565
rect 78752 4516 78794 4556
rect 78834 4516 78876 4556
rect 78916 4516 78958 4556
rect 78998 4516 79040 4556
rect 78712 4507 79080 4516
rect 93832 4556 94200 4565
rect 93872 4516 93914 4556
rect 93954 4516 93996 4556
rect 94036 4516 94078 4556
rect 94118 4516 94160 4556
rect 93832 4507 94200 4516
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 19472 3800 19840 3809
rect 19512 3760 19554 3800
rect 19594 3760 19636 3800
rect 19676 3760 19718 3800
rect 19758 3760 19800 3800
rect 19472 3751 19840 3760
rect 34592 3800 34960 3809
rect 34632 3760 34674 3800
rect 34714 3760 34756 3800
rect 34796 3760 34838 3800
rect 34878 3760 34920 3800
rect 34592 3751 34960 3760
rect 49712 3800 50080 3809
rect 49752 3760 49794 3800
rect 49834 3760 49876 3800
rect 49916 3760 49958 3800
rect 49998 3760 50040 3800
rect 49712 3751 50080 3760
rect 64832 3800 65200 3809
rect 64872 3760 64914 3800
rect 64954 3760 64996 3800
rect 65036 3760 65078 3800
rect 65118 3760 65160 3800
rect 64832 3751 65200 3760
rect 79952 3800 80320 3809
rect 79992 3760 80034 3800
rect 80074 3760 80116 3800
rect 80156 3760 80198 3800
rect 80238 3760 80280 3800
rect 79952 3751 80320 3760
rect 95072 3800 95440 3809
rect 95112 3760 95154 3800
rect 95194 3760 95236 3800
rect 95276 3760 95318 3800
rect 95358 3760 95400 3800
rect 95072 3751 95440 3760
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 18232 3044 18600 3053
rect 18272 3004 18314 3044
rect 18354 3004 18396 3044
rect 18436 3004 18478 3044
rect 18518 3004 18560 3044
rect 18232 2995 18600 3004
rect 33352 3044 33720 3053
rect 33392 3004 33434 3044
rect 33474 3004 33516 3044
rect 33556 3004 33598 3044
rect 33638 3004 33680 3044
rect 33352 2995 33720 3004
rect 48472 3044 48840 3053
rect 48512 3004 48554 3044
rect 48594 3004 48636 3044
rect 48676 3004 48718 3044
rect 48758 3004 48800 3044
rect 48472 2995 48840 3004
rect 63592 3044 63960 3053
rect 63632 3004 63674 3044
rect 63714 3004 63756 3044
rect 63796 3004 63838 3044
rect 63878 3004 63920 3044
rect 63592 2995 63960 3004
rect 78712 3044 79080 3053
rect 78752 3004 78794 3044
rect 78834 3004 78876 3044
rect 78916 3004 78958 3044
rect 78998 3004 79040 3044
rect 78712 2995 79080 3004
rect 93832 3044 94200 3053
rect 93872 3004 93914 3044
rect 93954 3004 93996 3044
rect 94036 3004 94078 3044
rect 94118 3004 94160 3044
rect 93832 2995 94200 3004
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 19472 2288 19840 2297
rect 19512 2248 19554 2288
rect 19594 2248 19636 2288
rect 19676 2248 19718 2288
rect 19758 2248 19800 2288
rect 19472 2239 19840 2248
rect 34592 2288 34960 2297
rect 34632 2248 34674 2288
rect 34714 2248 34756 2288
rect 34796 2248 34838 2288
rect 34878 2248 34920 2288
rect 34592 2239 34960 2248
rect 49712 2288 50080 2297
rect 49752 2248 49794 2288
rect 49834 2248 49876 2288
rect 49916 2248 49958 2288
rect 49998 2248 50040 2288
rect 49712 2239 50080 2248
rect 64832 2288 65200 2297
rect 64872 2248 64914 2288
rect 64954 2248 64996 2288
rect 65036 2248 65078 2288
rect 65118 2248 65160 2288
rect 64832 2239 65200 2248
rect 79952 2288 80320 2297
rect 79992 2248 80034 2288
rect 80074 2248 80116 2288
rect 80156 2248 80198 2288
rect 80238 2248 80280 2288
rect 79952 2239 80320 2248
rect 95072 2288 95440 2297
rect 95112 2248 95154 2288
rect 95194 2248 95236 2288
rect 95276 2248 95318 2288
rect 95358 2248 95400 2288
rect 95072 2239 95440 2248
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 18232 1532 18600 1541
rect 18272 1492 18314 1532
rect 18354 1492 18396 1532
rect 18436 1492 18478 1532
rect 18518 1492 18560 1532
rect 18232 1483 18600 1492
rect 33352 1532 33720 1541
rect 33392 1492 33434 1532
rect 33474 1492 33516 1532
rect 33556 1492 33598 1532
rect 33638 1492 33680 1532
rect 33352 1483 33720 1492
rect 48472 1532 48840 1541
rect 48512 1492 48554 1532
rect 48594 1492 48636 1532
rect 48676 1492 48718 1532
rect 48758 1492 48800 1532
rect 48472 1483 48840 1492
rect 63592 1532 63960 1541
rect 63632 1492 63674 1532
rect 63714 1492 63756 1532
rect 63796 1492 63838 1532
rect 63878 1492 63920 1532
rect 63592 1483 63960 1492
rect 78712 1532 79080 1541
rect 78752 1492 78794 1532
rect 78834 1492 78876 1532
rect 78916 1492 78958 1532
rect 78998 1492 79040 1532
rect 78712 1483 79080 1492
rect 93832 1532 94200 1541
rect 93872 1492 93914 1532
rect 93954 1492 93996 1532
rect 94036 1492 94078 1532
rect 94118 1492 94160 1532
rect 93832 1483 94200 1492
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 19472 776 19840 785
rect 19512 736 19554 776
rect 19594 736 19636 776
rect 19676 736 19718 776
rect 19758 736 19800 776
rect 19472 727 19840 736
rect 34592 776 34960 785
rect 34632 736 34674 776
rect 34714 736 34756 776
rect 34796 736 34838 776
rect 34878 736 34920 776
rect 34592 727 34960 736
rect 49712 776 50080 785
rect 49752 736 49794 776
rect 49834 736 49876 776
rect 49916 736 49958 776
rect 49998 736 50040 776
rect 49712 727 50080 736
rect 64832 776 65200 785
rect 64872 736 64914 776
rect 64954 736 64996 776
rect 65036 736 65078 776
rect 65118 736 65160 776
rect 64832 727 65200 736
rect 79952 776 80320 785
rect 79992 736 80034 776
rect 80074 736 80116 776
rect 80156 736 80198 776
rect 80238 736 80280 776
rect 79952 727 80320 736
rect 95072 776 95440 785
rect 95112 736 95154 776
rect 95194 736 95236 776
rect 95276 736 95318 776
rect 95358 736 95400 776
rect 95072 727 95440 736
<< via4 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 19472 38536 19512 38576
rect 19554 38536 19594 38576
rect 19636 38536 19676 38576
rect 19718 38536 19758 38576
rect 19800 38536 19840 38576
rect 34592 38536 34632 38576
rect 34674 38536 34714 38576
rect 34756 38536 34796 38576
rect 34838 38536 34878 38576
rect 34920 38536 34960 38576
rect 49712 38536 49752 38576
rect 49794 38536 49834 38576
rect 49876 38536 49916 38576
rect 49958 38536 49998 38576
rect 50040 38536 50080 38576
rect 64832 38536 64872 38576
rect 64914 38536 64954 38576
rect 64996 38536 65036 38576
rect 65078 38536 65118 38576
rect 65160 38536 65200 38576
rect 79952 38536 79992 38576
rect 80034 38536 80074 38576
rect 80116 38536 80156 38576
rect 80198 38536 80238 38576
rect 80280 38536 80320 38576
rect 95072 38536 95112 38576
rect 95154 38536 95194 38576
rect 95236 38536 95276 38576
rect 95318 38536 95358 38576
rect 95400 38536 95440 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 18232 37780 18272 37820
rect 18314 37780 18354 37820
rect 18396 37780 18436 37820
rect 18478 37780 18518 37820
rect 18560 37780 18600 37820
rect 33352 37780 33392 37820
rect 33434 37780 33474 37820
rect 33516 37780 33556 37820
rect 33598 37780 33638 37820
rect 33680 37780 33720 37820
rect 48472 37780 48512 37820
rect 48554 37780 48594 37820
rect 48636 37780 48676 37820
rect 48718 37780 48758 37820
rect 48800 37780 48840 37820
rect 63592 37780 63632 37820
rect 63674 37780 63714 37820
rect 63756 37780 63796 37820
rect 63838 37780 63878 37820
rect 63920 37780 63960 37820
rect 78712 37780 78752 37820
rect 78794 37780 78834 37820
rect 78876 37780 78916 37820
rect 78958 37780 78998 37820
rect 79040 37780 79080 37820
rect 93832 37780 93872 37820
rect 93914 37780 93954 37820
rect 93996 37780 94036 37820
rect 94078 37780 94118 37820
rect 94160 37780 94200 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 19472 37024 19512 37064
rect 19554 37024 19594 37064
rect 19636 37024 19676 37064
rect 19718 37024 19758 37064
rect 19800 37024 19840 37064
rect 34592 37024 34632 37064
rect 34674 37024 34714 37064
rect 34756 37024 34796 37064
rect 34838 37024 34878 37064
rect 34920 37024 34960 37064
rect 49712 37024 49752 37064
rect 49794 37024 49834 37064
rect 49876 37024 49916 37064
rect 49958 37024 49998 37064
rect 50040 37024 50080 37064
rect 64832 37024 64872 37064
rect 64914 37024 64954 37064
rect 64996 37024 65036 37064
rect 65078 37024 65118 37064
rect 65160 37024 65200 37064
rect 79952 37024 79992 37064
rect 80034 37024 80074 37064
rect 80116 37024 80156 37064
rect 80198 37024 80238 37064
rect 80280 37024 80320 37064
rect 95072 37024 95112 37064
rect 95154 37024 95194 37064
rect 95236 37024 95276 37064
rect 95318 37024 95358 37064
rect 95400 37024 95440 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 18232 36268 18272 36308
rect 18314 36268 18354 36308
rect 18396 36268 18436 36308
rect 18478 36268 18518 36308
rect 18560 36268 18600 36308
rect 33352 36268 33392 36308
rect 33434 36268 33474 36308
rect 33516 36268 33556 36308
rect 33598 36268 33638 36308
rect 33680 36268 33720 36308
rect 48472 36268 48512 36308
rect 48554 36268 48594 36308
rect 48636 36268 48676 36308
rect 48718 36268 48758 36308
rect 48800 36268 48840 36308
rect 63592 36268 63632 36308
rect 63674 36268 63714 36308
rect 63756 36268 63796 36308
rect 63838 36268 63878 36308
rect 63920 36268 63960 36308
rect 78712 36268 78752 36308
rect 78794 36268 78834 36308
rect 78876 36268 78916 36308
rect 78958 36268 78998 36308
rect 79040 36268 79080 36308
rect 93832 36268 93872 36308
rect 93914 36268 93954 36308
rect 93996 36268 94036 36308
rect 94078 36268 94118 36308
rect 94160 36268 94200 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 19472 35512 19512 35552
rect 19554 35512 19594 35552
rect 19636 35512 19676 35552
rect 19718 35512 19758 35552
rect 19800 35512 19840 35552
rect 34592 35512 34632 35552
rect 34674 35512 34714 35552
rect 34756 35512 34796 35552
rect 34838 35512 34878 35552
rect 34920 35512 34960 35552
rect 49712 35512 49752 35552
rect 49794 35512 49834 35552
rect 49876 35512 49916 35552
rect 49958 35512 49998 35552
rect 50040 35512 50080 35552
rect 64832 35512 64872 35552
rect 64914 35512 64954 35552
rect 64996 35512 65036 35552
rect 65078 35512 65118 35552
rect 65160 35512 65200 35552
rect 79952 35512 79992 35552
rect 80034 35512 80074 35552
rect 80116 35512 80156 35552
rect 80198 35512 80238 35552
rect 80280 35512 80320 35552
rect 95072 35512 95112 35552
rect 95154 35512 95194 35552
rect 95236 35512 95276 35552
rect 95318 35512 95358 35552
rect 95400 35512 95440 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 18232 34756 18272 34796
rect 18314 34756 18354 34796
rect 18396 34756 18436 34796
rect 18478 34756 18518 34796
rect 18560 34756 18600 34796
rect 33352 34756 33392 34796
rect 33434 34756 33474 34796
rect 33516 34756 33556 34796
rect 33598 34756 33638 34796
rect 33680 34756 33720 34796
rect 48472 34756 48512 34796
rect 48554 34756 48594 34796
rect 48636 34756 48676 34796
rect 48718 34756 48758 34796
rect 48800 34756 48840 34796
rect 63592 34756 63632 34796
rect 63674 34756 63714 34796
rect 63756 34756 63796 34796
rect 63838 34756 63878 34796
rect 63920 34756 63960 34796
rect 78712 34756 78752 34796
rect 78794 34756 78834 34796
rect 78876 34756 78916 34796
rect 78958 34756 78998 34796
rect 79040 34756 79080 34796
rect 93832 34756 93872 34796
rect 93914 34756 93954 34796
rect 93996 34756 94036 34796
rect 94078 34756 94118 34796
rect 94160 34756 94200 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 19472 34000 19512 34040
rect 19554 34000 19594 34040
rect 19636 34000 19676 34040
rect 19718 34000 19758 34040
rect 19800 34000 19840 34040
rect 34592 34000 34632 34040
rect 34674 34000 34714 34040
rect 34756 34000 34796 34040
rect 34838 34000 34878 34040
rect 34920 34000 34960 34040
rect 49712 34000 49752 34040
rect 49794 34000 49834 34040
rect 49876 34000 49916 34040
rect 49958 34000 49998 34040
rect 50040 34000 50080 34040
rect 64832 34000 64872 34040
rect 64914 34000 64954 34040
rect 64996 34000 65036 34040
rect 65078 34000 65118 34040
rect 65160 34000 65200 34040
rect 79952 34000 79992 34040
rect 80034 34000 80074 34040
rect 80116 34000 80156 34040
rect 80198 34000 80238 34040
rect 80280 34000 80320 34040
rect 95072 34000 95112 34040
rect 95154 34000 95194 34040
rect 95236 34000 95276 34040
rect 95318 34000 95358 34040
rect 95400 34000 95440 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 18232 33244 18272 33284
rect 18314 33244 18354 33284
rect 18396 33244 18436 33284
rect 18478 33244 18518 33284
rect 18560 33244 18600 33284
rect 33352 33244 33392 33284
rect 33434 33244 33474 33284
rect 33516 33244 33556 33284
rect 33598 33244 33638 33284
rect 33680 33244 33720 33284
rect 48472 33244 48512 33284
rect 48554 33244 48594 33284
rect 48636 33244 48676 33284
rect 48718 33244 48758 33284
rect 48800 33244 48840 33284
rect 63592 33244 63632 33284
rect 63674 33244 63714 33284
rect 63756 33244 63796 33284
rect 63838 33244 63878 33284
rect 63920 33244 63960 33284
rect 78712 33244 78752 33284
rect 78794 33244 78834 33284
rect 78876 33244 78916 33284
rect 78958 33244 78998 33284
rect 79040 33244 79080 33284
rect 93832 33244 93872 33284
rect 93914 33244 93954 33284
rect 93996 33244 94036 33284
rect 94078 33244 94118 33284
rect 94160 33244 94200 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 19472 32488 19512 32528
rect 19554 32488 19594 32528
rect 19636 32488 19676 32528
rect 19718 32488 19758 32528
rect 19800 32488 19840 32528
rect 34592 32488 34632 32528
rect 34674 32488 34714 32528
rect 34756 32488 34796 32528
rect 34838 32488 34878 32528
rect 34920 32488 34960 32528
rect 49712 32488 49752 32528
rect 49794 32488 49834 32528
rect 49876 32488 49916 32528
rect 49958 32488 49998 32528
rect 50040 32488 50080 32528
rect 64832 32488 64872 32528
rect 64914 32488 64954 32528
rect 64996 32488 65036 32528
rect 65078 32488 65118 32528
rect 65160 32488 65200 32528
rect 79952 32488 79992 32528
rect 80034 32488 80074 32528
rect 80116 32488 80156 32528
rect 80198 32488 80238 32528
rect 80280 32488 80320 32528
rect 95072 32488 95112 32528
rect 95154 32488 95194 32528
rect 95236 32488 95276 32528
rect 95318 32488 95358 32528
rect 95400 32488 95440 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 18232 31732 18272 31772
rect 18314 31732 18354 31772
rect 18396 31732 18436 31772
rect 18478 31732 18518 31772
rect 18560 31732 18600 31772
rect 33352 31732 33392 31772
rect 33434 31732 33474 31772
rect 33516 31732 33556 31772
rect 33598 31732 33638 31772
rect 33680 31732 33720 31772
rect 48472 31732 48512 31772
rect 48554 31732 48594 31772
rect 48636 31732 48676 31772
rect 48718 31732 48758 31772
rect 48800 31732 48840 31772
rect 63592 31732 63632 31772
rect 63674 31732 63714 31772
rect 63756 31732 63796 31772
rect 63838 31732 63878 31772
rect 63920 31732 63960 31772
rect 78712 31732 78752 31772
rect 78794 31732 78834 31772
rect 78876 31732 78916 31772
rect 78958 31732 78998 31772
rect 79040 31732 79080 31772
rect 93832 31732 93872 31772
rect 93914 31732 93954 31772
rect 93996 31732 94036 31772
rect 94078 31732 94118 31772
rect 94160 31732 94200 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 19472 30976 19512 31016
rect 19554 30976 19594 31016
rect 19636 30976 19676 31016
rect 19718 30976 19758 31016
rect 19800 30976 19840 31016
rect 34592 30976 34632 31016
rect 34674 30976 34714 31016
rect 34756 30976 34796 31016
rect 34838 30976 34878 31016
rect 34920 30976 34960 31016
rect 49712 30976 49752 31016
rect 49794 30976 49834 31016
rect 49876 30976 49916 31016
rect 49958 30976 49998 31016
rect 50040 30976 50080 31016
rect 64832 30976 64872 31016
rect 64914 30976 64954 31016
rect 64996 30976 65036 31016
rect 65078 30976 65118 31016
rect 65160 30976 65200 31016
rect 79952 30976 79992 31016
rect 80034 30976 80074 31016
rect 80116 30976 80156 31016
rect 80198 30976 80238 31016
rect 80280 30976 80320 31016
rect 95072 30976 95112 31016
rect 95154 30976 95194 31016
rect 95236 30976 95276 31016
rect 95318 30976 95358 31016
rect 95400 30976 95440 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 18232 30220 18272 30260
rect 18314 30220 18354 30260
rect 18396 30220 18436 30260
rect 18478 30220 18518 30260
rect 18560 30220 18600 30260
rect 33352 30220 33392 30260
rect 33434 30220 33474 30260
rect 33516 30220 33556 30260
rect 33598 30220 33638 30260
rect 33680 30220 33720 30260
rect 48472 30220 48512 30260
rect 48554 30220 48594 30260
rect 48636 30220 48676 30260
rect 48718 30220 48758 30260
rect 48800 30220 48840 30260
rect 63592 30220 63632 30260
rect 63674 30220 63714 30260
rect 63756 30220 63796 30260
rect 63838 30220 63878 30260
rect 63920 30220 63960 30260
rect 78712 30220 78752 30260
rect 78794 30220 78834 30260
rect 78876 30220 78916 30260
rect 78958 30220 78998 30260
rect 79040 30220 79080 30260
rect 93832 30220 93872 30260
rect 93914 30220 93954 30260
rect 93996 30220 94036 30260
rect 94078 30220 94118 30260
rect 94160 30220 94200 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 19472 29464 19512 29504
rect 19554 29464 19594 29504
rect 19636 29464 19676 29504
rect 19718 29464 19758 29504
rect 19800 29464 19840 29504
rect 34592 29464 34632 29504
rect 34674 29464 34714 29504
rect 34756 29464 34796 29504
rect 34838 29464 34878 29504
rect 34920 29464 34960 29504
rect 49712 29464 49752 29504
rect 49794 29464 49834 29504
rect 49876 29464 49916 29504
rect 49958 29464 49998 29504
rect 50040 29464 50080 29504
rect 64832 29464 64872 29504
rect 64914 29464 64954 29504
rect 64996 29464 65036 29504
rect 65078 29464 65118 29504
rect 65160 29464 65200 29504
rect 79952 29464 79992 29504
rect 80034 29464 80074 29504
rect 80116 29464 80156 29504
rect 80198 29464 80238 29504
rect 80280 29464 80320 29504
rect 95072 29464 95112 29504
rect 95154 29464 95194 29504
rect 95236 29464 95276 29504
rect 95318 29464 95358 29504
rect 95400 29464 95440 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 18232 28708 18272 28748
rect 18314 28708 18354 28748
rect 18396 28708 18436 28748
rect 18478 28708 18518 28748
rect 18560 28708 18600 28748
rect 33352 28708 33392 28748
rect 33434 28708 33474 28748
rect 33516 28708 33556 28748
rect 33598 28708 33638 28748
rect 33680 28708 33720 28748
rect 48472 28708 48512 28748
rect 48554 28708 48594 28748
rect 48636 28708 48676 28748
rect 48718 28708 48758 28748
rect 48800 28708 48840 28748
rect 63592 28708 63632 28748
rect 63674 28708 63714 28748
rect 63756 28708 63796 28748
rect 63838 28708 63878 28748
rect 63920 28708 63960 28748
rect 78712 28708 78752 28748
rect 78794 28708 78834 28748
rect 78876 28708 78916 28748
rect 78958 28708 78998 28748
rect 79040 28708 79080 28748
rect 93832 28708 93872 28748
rect 93914 28708 93954 28748
rect 93996 28708 94036 28748
rect 94078 28708 94118 28748
rect 94160 28708 94200 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 19472 27952 19512 27992
rect 19554 27952 19594 27992
rect 19636 27952 19676 27992
rect 19718 27952 19758 27992
rect 19800 27952 19840 27992
rect 34592 27952 34632 27992
rect 34674 27952 34714 27992
rect 34756 27952 34796 27992
rect 34838 27952 34878 27992
rect 34920 27952 34960 27992
rect 49712 27952 49752 27992
rect 49794 27952 49834 27992
rect 49876 27952 49916 27992
rect 49958 27952 49998 27992
rect 50040 27952 50080 27992
rect 64832 27952 64872 27992
rect 64914 27952 64954 27992
rect 64996 27952 65036 27992
rect 65078 27952 65118 27992
rect 65160 27952 65200 27992
rect 79952 27952 79992 27992
rect 80034 27952 80074 27992
rect 80116 27952 80156 27992
rect 80198 27952 80238 27992
rect 80280 27952 80320 27992
rect 95072 27952 95112 27992
rect 95154 27952 95194 27992
rect 95236 27952 95276 27992
rect 95318 27952 95358 27992
rect 95400 27952 95440 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 18232 27196 18272 27236
rect 18314 27196 18354 27236
rect 18396 27196 18436 27236
rect 18478 27196 18518 27236
rect 18560 27196 18600 27236
rect 33352 27196 33392 27236
rect 33434 27196 33474 27236
rect 33516 27196 33556 27236
rect 33598 27196 33638 27236
rect 33680 27196 33720 27236
rect 48472 27196 48512 27236
rect 48554 27196 48594 27236
rect 48636 27196 48676 27236
rect 48718 27196 48758 27236
rect 48800 27196 48840 27236
rect 63592 27196 63632 27236
rect 63674 27196 63714 27236
rect 63756 27196 63796 27236
rect 63838 27196 63878 27236
rect 63920 27196 63960 27236
rect 78712 27196 78752 27236
rect 78794 27196 78834 27236
rect 78876 27196 78916 27236
rect 78958 27196 78998 27236
rect 79040 27196 79080 27236
rect 93832 27196 93872 27236
rect 93914 27196 93954 27236
rect 93996 27196 94036 27236
rect 94078 27196 94118 27236
rect 94160 27196 94200 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 19472 26440 19512 26480
rect 19554 26440 19594 26480
rect 19636 26440 19676 26480
rect 19718 26440 19758 26480
rect 19800 26440 19840 26480
rect 34592 26440 34632 26480
rect 34674 26440 34714 26480
rect 34756 26440 34796 26480
rect 34838 26440 34878 26480
rect 34920 26440 34960 26480
rect 49712 26440 49752 26480
rect 49794 26440 49834 26480
rect 49876 26440 49916 26480
rect 49958 26440 49998 26480
rect 50040 26440 50080 26480
rect 64832 26440 64872 26480
rect 64914 26440 64954 26480
rect 64996 26440 65036 26480
rect 65078 26440 65118 26480
rect 65160 26440 65200 26480
rect 79952 26440 79992 26480
rect 80034 26440 80074 26480
rect 80116 26440 80156 26480
rect 80198 26440 80238 26480
rect 80280 26440 80320 26480
rect 95072 26440 95112 26480
rect 95154 26440 95194 26480
rect 95236 26440 95276 26480
rect 95318 26440 95358 26480
rect 95400 26440 95440 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 18232 25684 18272 25724
rect 18314 25684 18354 25724
rect 18396 25684 18436 25724
rect 18478 25684 18518 25724
rect 18560 25684 18600 25724
rect 33352 25684 33392 25724
rect 33434 25684 33474 25724
rect 33516 25684 33556 25724
rect 33598 25684 33638 25724
rect 33680 25684 33720 25724
rect 48472 25684 48512 25724
rect 48554 25684 48594 25724
rect 48636 25684 48676 25724
rect 48718 25684 48758 25724
rect 48800 25684 48840 25724
rect 63592 25684 63632 25724
rect 63674 25684 63714 25724
rect 63756 25684 63796 25724
rect 63838 25684 63878 25724
rect 63920 25684 63960 25724
rect 78712 25684 78752 25724
rect 78794 25684 78834 25724
rect 78876 25684 78916 25724
rect 78958 25684 78998 25724
rect 79040 25684 79080 25724
rect 93832 25684 93872 25724
rect 93914 25684 93954 25724
rect 93996 25684 94036 25724
rect 94078 25684 94118 25724
rect 94160 25684 94200 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 19472 24928 19512 24968
rect 19554 24928 19594 24968
rect 19636 24928 19676 24968
rect 19718 24928 19758 24968
rect 19800 24928 19840 24968
rect 34592 24928 34632 24968
rect 34674 24928 34714 24968
rect 34756 24928 34796 24968
rect 34838 24928 34878 24968
rect 34920 24928 34960 24968
rect 49712 24928 49752 24968
rect 49794 24928 49834 24968
rect 49876 24928 49916 24968
rect 49958 24928 49998 24968
rect 50040 24928 50080 24968
rect 64832 24928 64872 24968
rect 64914 24928 64954 24968
rect 64996 24928 65036 24968
rect 65078 24928 65118 24968
rect 65160 24928 65200 24968
rect 79952 24928 79992 24968
rect 80034 24928 80074 24968
rect 80116 24928 80156 24968
rect 80198 24928 80238 24968
rect 80280 24928 80320 24968
rect 95072 24928 95112 24968
rect 95154 24928 95194 24968
rect 95236 24928 95276 24968
rect 95318 24928 95358 24968
rect 95400 24928 95440 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 18232 24172 18272 24212
rect 18314 24172 18354 24212
rect 18396 24172 18436 24212
rect 18478 24172 18518 24212
rect 18560 24172 18600 24212
rect 33352 24172 33392 24212
rect 33434 24172 33474 24212
rect 33516 24172 33556 24212
rect 33598 24172 33638 24212
rect 33680 24172 33720 24212
rect 48472 24172 48512 24212
rect 48554 24172 48594 24212
rect 48636 24172 48676 24212
rect 48718 24172 48758 24212
rect 48800 24172 48840 24212
rect 63592 24172 63632 24212
rect 63674 24172 63714 24212
rect 63756 24172 63796 24212
rect 63838 24172 63878 24212
rect 63920 24172 63960 24212
rect 78712 24172 78752 24212
rect 78794 24172 78834 24212
rect 78876 24172 78916 24212
rect 78958 24172 78998 24212
rect 79040 24172 79080 24212
rect 93832 24172 93872 24212
rect 93914 24172 93954 24212
rect 93996 24172 94036 24212
rect 94078 24172 94118 24212
rect 94160 24172 94200 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 19472 23416 19512 23456
rect 19554 23416 19594 23456
rect 19636 23416 19676 23456
rect 19718 23416 19758 23456
rect 19800 23416 19840 23456
rect 34592 23416 34632 23456
rect 34674 23416 34714 23456
rect 34756 23416 34796 23456
rect 34838 23416 34878 23456
rect 34920 23416 34960 23456
rect 49712 23416 49752 23456
rect 49794 23416 49834 23456
rect 49876 23416 49916 23456
rect 49958 23416 49998 23456
rect 50040 23416 50080 23456
rect 64832 23416 64872 23456
rect 64914 23416 64954 23456
rect 64996 23416 65036 23456
rect 65078 23416 65118 23456
rect 65160 23416 65200 23456
rect 79952 23416 79992 23456
rect 80034 23416 80074 23456
rect 80116 23416 80156 23456
rect 80198 23416 80238 23456
rect 80280 23416 80320 23456
rect 95072 23416 95112 23456
rect 95154 23416 95194 23456
rect 95236 23416 95276 23456
rect 95318 23416 95358 23456
rect 95400 23416 95440 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 18232 22660 18272 22700
rect 18314 22660 18354 22700
rect 18396 22660 18436 22700
rect 18478 22660 18518 22700
rect 18560 22660 18600 22700
rect 33352 22660 33392 22700
rect 33434 22660 33474 22700
rect 33516 22660 33556 22700
rect 33598 22660 33638 22700
rect 33680 22660 33720 22700
rect 48472 22660 48512 22700
rect 48554 22660 48594 22700
rect 48636 22660 48676 22700
rect 48718 22660 48758 22700
rect 48800 22660 48840 22700
rect 63592 22660 63632 22700
rect 63674 22660 63714 22700
rect 63756 22660 63796 22700
rect 63838 22660 63878 22700
rect 63920 22660 63960 22700
rect 78712 22660 78752 22700
rect 78794 22660 78834 22700
rect 78876 22660 78916 22700
rect 78958 22660 78998 22700
rect 79040 22660 79080 22700
rect 93832 22660 93872 22700
rect 93914 22660 93954 22700
rect 93996 22660 94036 22700
rect 94078 22660 94118 22700
rect 94160 22660 94200 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 19472 21904 19512 21944
rect 19554 21904 19594 21944
rect 19636 21904 19676 21944
rect 19718 21904 19758 21944
rect 19800 21904 19840 21944
rect 34592 21904 34632 21944
rect 34674 21904 34714 21944
rect 34756 21904 34796 21944
rect 34838 21904 34878 21944
rect 34920 21904 34960 21944
rect 49712 21904 49752 21944
rect 49794 21904 49834 21944
rect 49876 21904 49916 21944
rect 49958 21904 49998 21944
rect 50040 21904 50080 21944
rect 64832 21904 64872 21944
rect 64914 21904 64954 21944
rect 64996 21904 65036 21944
rect 65078 21904 65118 21944
rect 65160 21904 65200 21944
rect 79952 21904 79992 21944
rect 80034 21904 80074 21944
rect 80116 21904 80156 21944
rect 80198 21904 80238 21944
rect 80280 21904 80320 21944
rect 95072 21904 95112 21944
rect 95154 21904 95194 21944
rect 95236 21904 95276 21944
rect 95318 21904 95358 21944
rect 95400 21904 95440 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 18232 21148 18272 21188
rect 18314 21148 18354 21188
rect 18396 21148 18436 21188
rect 18478 21148 18518 21188
rect 18560 21148 18600 21188
rect 33352 21148 33392 21188
rect 33434 21148 33474 21188
rect 33516 21148 33556 21188
rect 33598 21148 33638 21188
rect 33680 21148 33720 21188
rect 48472 21148 48512 21188
rect 48554 21148 48594 21188
rect 48636 21148 48676 21188
rect 48718 21148 48758 21188
rect 48800 21148 48840 21188
rect 63592 21148 63632 21188
rect 63674 21148 63714 21188
rect 63756 21148 63796 21188
rect 63838 21148 63878 21188
rect 63920 21148 63960 21188
rect 78712 21148 78752 21188
rect 78794 21148 78834 21188
rect 78876 21148 78916 21188
rect 78958 21148 78998 21188
rect 79040 21148 79080 21188
rect 93832 21148 93872 21188
rect 93914 21148 93954 21188
rect 93996 21148 94036 21188
rect 94078 21148 94118 21188
rect 94160 21148 94200 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 19472 20392 19512 20432
rect 19554 20392 19594 20432
rect 19636 20392 19676 20432
rect 19718 20392 19758 20432
rect 19800 20392 19840 20432
rect 34592 20392 34632 20432
rect 34674 20392 34714 20432
rect 34756 20392 34796 20432
rect 34838 20392 34878 20432
rect 34920 20392 34960 20432
rect 49712 20392 49752 20432
rect 49794 20392 49834 20432
rect 49876 20392 49916 20432
rect 49958 20392 49998 20432
rect 50040 20392 50080 20432
rect 64832 20392 64872 20432
rect 64914 20392 64954 20432
rect 64996 20392 65036 20432
rect 65078 20392 65118 20432
rect 65160 20392 65200 20432
rect 79952 20392 79992 20432
rect 80034 20392 80074 20432
rect 80116 20392 80156 20432
rect 80198 20392 80238 20432
rect 80280 20392 80320 20432
rect 95072 20392 95112 20432
rect 95154 20392 95194 20432
rect 95236 20392 95276 20432
rect 95318 20392 95358 20432
rect 95400 20392 95440 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 18232 19636 18272 19676
rect 18314 19636 18354 19676
rect 18396 19636 18436 19676
rect 18478 19636 18518 19676
rect 18560 19636 18600 19676
rect 33352 19636 33392 19676
rect 33434 19636 33474 19676
rect 33516 19636 33556 19676
rect 33598 19636 33638 19676
rect 33680 19636 33720 19676
rect 48472 19636 48512 19676
rect 48554 19636 48594 19676
rect 48636 19636 48676 19676
rect 48718 19636 48758 19676
rect 48800 19636 48840 19676
rect 63592 19636 63632 19676
rect 63674 19636 63714 19676
rect 63756 19636 63796 19676
rect 63838 19636 63878 19676
rect 63920 19636 63960 19676
rect 78712 19636 78752 19676
rect 78794 19636 78834 19676
rect 78876 19636 78916 19676
rect 78958 19636 78998 19676
rect 79040 19636 79080 19676
rect 93832 19636 93872 19676
rect 93914 19636 93954 19676
rect 93996 19636 94036 19676
rect 94078 19636 94118 19676
rect 94160 19636 94200 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 19472 18880 19512 18920
rect 19554 18880 19594 18920
rect 19636 18880 19676 18920
rect 19718 18880 19758 18920
rect 19800 18880 19840 18920
rect 34592 18880 34632 18920
rect 34674 18880 34714 18920
rect 34756 18880 34796 18920
rect 34838 18880 34878 18920
rect 34920 18880 34960 18920
rect 49712 18880 49752 18920
rect 49794 18880 49834 18920
rect 49876 18880 49916 18920
rect 49958 18880 49998 18920
rect 50040 18880 50080 18920
rect 64832 18880 64872 18920
rect 64914 18880 64954 18920
rect 64996 18880 65036 18920
rect 65078 18880 65118 18920
rect 65160 18880 65200 18920
rect 79952 18880 79992 18920
rect 80034 18880 80074 18920
rect 80116 18880 80156 18920
rect 80198 18880 80238 18920
rect 80280 18880 80320 18920
rect 95072 18880 95112 18920
rect 95154 18880 95194 18920
rect 95236 18880 95276 18920
rect 95318 18880 95358 18920
rect 95400 18880 95440 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 18232 18124 18272 18164
rect 18314 18124 18354 18164
rect 18396 18124 18436 18164
rect 18478 18124 18518 18164
rect 18560 18124 18600 18164
rect 33352 18124 33392 18164
rect 33434 18124 33474 18164
rect 33516 18124 33556 18164
rect 33598 18124 33638 18164
rect 33680 18124 33720 18164
rect 48472 18124 48512 18164
rect 48554 18124 48594 18164
rect 48636 18124 48676 18164
rect 48718 18124 48758 18164
rect 48800 18124 48840 18164
rect 63592 18124 63632 18164
rect 63674 18124 63714 18164
rect 63756 18124 63796 18164
rect 63838 18124 63878 18164
rect 63920 18124 63960 18164
rect 78712 18124 78752 18164
rect 78794 18124 78834 18164
rect 78876 18124 78916 18164
rect 78958 18124 78998 18164
rect 79040 18124 79080 18164
rect 93832 18124 93872 18164
rect 93914 18124 93954 18164
rect 93996 18124 94036 18164
rect 94078 18124 94118 18164
rect 94160 18124 94200 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 19472 17368 19512 17408
rect 19554 17368 19594 17408
rect 19636 17368 19676 17408
rect 19718 17368 19758 17408
rect 19800 17368 19840 17408
rect 34592 17368 34632 17408
rect 34674 17368 34714 17408
rect 34756 17368 34796 17408
rect 34838 17368 34878 17408
rect 34920 17368 34960 17408
rect 49712 17368 49752 17408
rect 49794 17368 49834 17408
rect 49876 17368 49916 17408
rect 49958 17368 49998 17408
rect 50040 17368 50080 17408
rect 64832 17368 64872 17408
rect 64914 17368 64954 17408
rect 64996 17368 65036 17408
rect 65078 17368 65118 17408
rect 65160 17368 65200 17408
rect 79952 17368 79992 17408
rect 80034 17368 80074 17408
rect 80116 17368 80156 17408
rect 80198 17368 80238 17408
rect 80280 17368 80320 17408
rect 95072 17368 95112 17408
rect 95154 17368 95194 17408
rect 95236 17368 95276 17408
rect 95318 17368 95358 17408
rect 95400 17368 95440 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 18232 16612 18272 16652
rect 18314 16612 18354 16652
rect 18396 16612 18436 16652
rect 18478 16612 18518 16652
rect 18560 16612 18600 16652
rect 33352 16612 33392 16652
rect 33434 16612 33474 16652
rect 33516 16612 33556 16652
rect 33598 16612 33638 16652
rect 33680 16612 33720 16652
rect 48472 16612 48512 16652
rect 48554 16612 48594 16652
rect 48636 16612 48676 16652
rect 48718 16612 48758 16652
rect 48800 16612 48840 16652
rect 63592 16612 63632 16652
rect 63674 16612 63714 16652
rect 63756 16612 63796 16652
rect 63838 16612 63878 16652
rect 63920 16612 63960 16652
rect 78712 16612 78752 16652
rect 78794 16612 78834 16652
rect 78876 16612 78916 16652
rect 78958 16612 78998 16652
rect 79040 16612 79080 16652
rect 93832 16612 93872 16652
rect 93914 16612 93954 16652
rect 93996 16612 94036 16652
rect 94078 16612 94118 16652
rect 94160 16612 94200 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 19472 15856 19512 15896
rect 19554 15856 19594 15896
rect 19636 15856 19676 15896
rect 19718 15856 19758 15896
rect 19800 15856 19840 15896
rect 34592 15856 34632 15896
rect 34674 15856 34714 15896
rect 34756 15856 34796 15896
rect 34838 15856 34878 15896
rect 34920 15856 34960 15896
rect 49712 15856 49752 15896
rect 49794 15856 49834 15896
rect 49876 15856 49916 15896
rect 49958 15856 49998 15896
rect 50040 15856 50080 15896
rect 64832 15856 64872 15896
rect 64914 15856 64954 15896
rect 64996 15856 65036 15896
rect 65078 15856 65118 15896
rect 65160 15856 65200 15896
rect 79952 15856 79992 15896
rect 80034 15856 80074 15896
rect 80116 15856 80156 15896
rect 80198 15856 80238 15896
rect 80280 15856 80320 15896
rect 95072 15856 95112 15896
rect 95154 15856 95194 15896
rect 95236 15856 95276 15896
rect 95318 15856 95358 15896
rect 95400 15856 95440 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 18232 15100 18272 15140
rect 18314 15100 18354 15140
rect 18396 15100 18436 15140
rect 18478 15100 18518 15140
rect 18560 15100 18600 15140
rect 33352 15100 33392 15140
rect 33434 15100 33474 15140
rect 33516 15100 33556 15140
rect 33598 15100 33638 15140
rect 33680 15100 33720 15140
rect 48472 15100 48512 15140
rect 48554 15100 48594 15140
rect 48636 15100 48676 15140
rect 48718 15100 48758 15140
rect 48800 15100 48840 15140
rect 63592 15100 63632 15140
rect 63674 15100 63714 15140
rect 63756 15100 63796 15140
rect 63838 15100 63878 15140
rect 63920 15100 63960 15140
rect 78712 15100 78752 15140
rect 78794 15100 78834 15140
rect 78876 15100 78916 15140
rect 78958 15100 78998 15140
rect 79040 15100 79080 15140
rect 93832 15100 93872 15140
rect 93914 15100 93954 15140
rect 93996 15100 94036 15140
rect 94078 15100 94118 15140
rect 94160 15100 94200 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 19472 14344 19512 14384
rect 19554 14344 19594 14384
rect 19636 14344 19676 14384
rect 19718 14344 19758 14384
rect 19800 14344 19840 14384
rect 34592 14344 34632 14384
rect 34674 14344 34714 14384
rect 34756 14344 34796 14384
rect 34838 14344 34878 14384
rect 34920 14344 34960 14384
rect 49712 14344 49752 14384
rect 49794 14344 49834 14384
rect 49876 14344 49916 14384
rect 49958 14344 49998 14384
rect 50040 14344 50080 14384
rect 64832 14344 64872 14384
rect 64914 14344 64954 14384
rect 64996 14344 65036 14384
rect 65078 14344 65118 14384
rect 65160 14344 65200 14384
rect 79952 14344 79992 14384
rect 80034 14344 80074 14384
rect 80116 14344 80156 14384
rect 80198 14344 80238 14384
rect 80280 14344 80320 14384
rect 95072 14344 95112 14384
rect 95154 14344 95194 14384
rect 95236 14344 95276 14384
rect 95318 14344 95358 14384
rect 95400 14344 95440 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 18232 13588 18272 13628
rect 18314 13588 18354 13628
rect 18396 13588 18436 13628
rect 18478 13588 18518 13628
rect 18560 13588 18600 13628
rect 33352 13588 33392 13628
rect 33434 13588 33474 13628
rect 33516 13588 33556 13628
rect 33598 13588 33638 13628
rect 33680 13588 33720 13628
rect 48472 13588 48512 13628
rect 48554 13588 48594 13628
rect 48636 13588 48676 13628
rect 48718 13588 48758 13628
rect 48800 13588 48840 13628
rect 63592 13588 63632 13628
rect 63674 13588 63714 13628
rect 63756 13588 63796 13628
rect 63838 13588 63878 13628
rect 63920 13588 63960 13628
rect 78712 13588 78752 13628
rect 78794 13588 78834 13628
rect 78876 13588 78916 13628
rect 78958 13588 78998 13628
rect 79040 13588 79080 13628
rect 93832 13588 93872 13628
rect 93914 13588 93954 13628
rect 93996 13588 94036 13628
rect 94078 13588 94118 13628
rect 94160 13588 94200 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 19472 12832 19512 12872
rect 19554 12832 19594 12872
rect 19636 12832 19676 12872
rect 19718 12832 19758 12872
rect 19800 12832 19840 12872
rect 34592 12832 34632 12872
rect 34674 12832 34714 12872
rect 34756 12832 34796 12872
rect 34838 12832 34878 12872
rect 34920 12832 34960 12872
rect 49712 12832 49752 12872
rect 49794 12832 49834 12872
rect 49876 12832 49916 12872
rect 49958 12832 49998 12872
rect 50040 12832 50080 12872
rect 64832 12832 64872 12872
rect 64914 12832 64954 12872
rect 64996 12832 65036 12872
rect 65078 12832 65118 12872
rect 65160 12832 65200 12872
rect 79952 12832 79992 12872
rect 80034 12832 80074 12872
rect 80116 12832 80156 12872
rect 80198 12832 80238 12872
rect 80280 12832 80320 12872
rect 95072 12832 95112 12872
rect 95154 12832 95194 12872
rect 95236 12832 95276 12872
rect 95318 12832 95358 12872
rect 95400 12832 95440 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 18232 12076 18272 12116
rect 18314 12076 18354 12116
rect 18396 12076 18436 12116
rect 18478 12076 18518 12116
rect 18560 12076 18600 12116
rect 33352 12076 33392 12116
rect 33434 12076 33474 12116
rect 33516 12076 33556 12116
rect 33598 12076 33638 12116
rect 33680 12076 33720 12116
rect 48472 12076 48512 12116
rect 48554 12076 48594 12116
rect 48636 12076 48676 12116
rect 48718 12076 48758 12116
rect 48800 12076 48840 12116
rect 63592 12076 63632 12116
rect 63674 12076 63714 12116
rect 63756 12076 63796 12116
rect 63838 12076 63878 12116
rect 63920 12076 63960 12116
rect 78712 12076 78752 12116
rect 78794 12076 78834 12116
rect 78876 12076 78916 12116
rect 78958 12076 78998 12116
rect 79040 12076 79080 12116
rect 93832 12076 93872 12116
rect 93914 12076 93954 12116
rect 93996 12076 94036 12116
rect 94078 12076 94118 12116
rect 94160 12076 94200 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 19472 11320 19512 11360
rect 19554 11320 19594 11360
rect 19636 11320 19676 11360
rect 19718 11320 19758 11360
rect 19800 11320 19840 11360
rect 34592 11320 34632 11360
rect 34674 11320 34714 11360
rect 34756 11320 34796 11360
rect 34838 11320 34878 11360
rect 34920 11320 34960 11360
rect 49712 11320 49752 11360
rect 49794 11320 49834 11360
rect 49876 11320 49916 11360
rect 49958 11320 49998 11360
rect 50040 11320 50080 11360
rect 64832 11320 64872 11360
rect 64914 11320 64954 11360
rect 64996 11320 65036 11360
rect 65078 11320 65118 11360
rect 65160 11320 65200 11360
rect 79952 11320 79992 11360
rect 80034 11320 80074 11360
rect 80116 11320 80156 11360
rect 80198 11320 80238 11360
rect 80280 11320 80320 11360
rect 95072 11320 95112 11360
rect 95154 11320 95194 11360
rect 95236 11320 95276 11360
rect 95318 11320 95358 11360
rect 95400 11320 95440 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 18232 10564 18272 10604
rect 18314 10564 18354 10604
rect 18396 10564 18436 10604
rect 18478 10564 18518 10604
rect 18560 10564 18600 10604
rect 33352 10564 33392 10604
rect 33434 10564 33474 10604
rect 33516 10564 33556 10604
rect 33598 10564 33638 10604
rect 33680 10564 33720 10604
rect 48472 10564 48512 10604
rect 48554 10564 48594 10604
rect 48636 10564 48676 10604
rect 48718 10564 48758 10604
rect 48800 10564 48840 10604
rect 63592 10564 63632 10604
rect 63674 10564 63714 10604
rect 63756 10564 63796 10604
rect 63838 10564 63878 10604
rect 63920 10564 63960 10604
rect 78712 10564 78752 10604
rect 78794 10564 78834 10604
rect 78876 10564 78916 10604
rect 78958 10564 78998 10604
rect 79040 10564 79080 10604
rect 93832 10564 93872 10604
rect 93914 10564 93954 10604
rect 93996 10564 94036 10604
rect 94078 10564 94118 10604
rect 94160 10564 94200 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 19472 9808 19512 9848
rect 19554 9808 19594 9848
rect 19636 9808 19676 9848
rect 19718 9808 19758 9848
rect 19800 9808 19840 9848
rect 34592 9808 34632 9848
rect 34674 9808 34714 9848
rect 34756 9808 34796 9848
rect 34838 9808 34878 9848
rect 34920 9808 34960 9848
rect 49712 9808 49752 9848
rect 49794 9808 49834 9848
rect 49876 9808 49916 9848
rect 49958 9808 49998 9848
rect 50040 9808 50080 9848
rect 64832 9808 64872 9848
rect 64914 9808 64954 9848
rect 64996 9808 65036 9848
rect 65078 9808 65118 9848
rect 65160 9808 65200 9848
rect 79952 9808 79992 9848
rect 80034 9808 80074 9848
rect 80116 9808 80156 9848
rect 80198 9808 80238 9848
rect 80280 9808 80320 9848
rect 95072 9808 95112 9848
rect 95154 9808 95194 9848
rect 95236 9808 95276 9848
rect 95318 9808 95358 9848
rect 95400 9808 95440 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 18232 9052 18272 9092
rect 18314 9052 18354 9092
rect 18396 9052 18436 9092
rect 18478 9052 18518 9092
rect 18560 9052 18600 9092
rect 33352 9052 33392 9092
rect 33434 9052 33474 9092
rect 33516 9052 33556 9092
rect 33598 9052 33638 9092
rect 33680 9052 33720 9092
rect 48472 9052 48512 9092
rect 48554 9052 48594 9092
rect 48636 9052 48676 9092
rect 48718 9052 48758 9092
rect 48800 9052 48840 9092
rect 63592 9052 63632 9092
rect 63674 9052 63714 9092
rect 63756 9052 63796 9092
rect 63838 9052 63878 9092
rect 63920 9052 63960 9092
rect 78712 9052 78752 9092
rect 78794 9052 78834 9092
rect 78876 9052 78916 9092
rect 78958 9052 78998 9092
rect 79040 9052 79080 9092
rect 93832 9052 93872 9092
rect 93914 9052 93954 9092
rect 93996 9052 94036 9092
rect 94078 9052 94118 9092
rect 94160 9052 94200 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 19472 8296 19512 8336
rect 19554 8296 19594 8336
rect 19636 8296 19676 8336
rect 19718 8296 19758 8336
rect 19800 8296 19840 8336
rect 34592 8296 34632 8336
rect 34674 8296 34714 8336
rect 34756 8296 34796 8336
rect 34838 8296 34878 8336
rect 34920 8296 34960 8336
rect 49712 8296 49752 8336
rect 49794 8296 49834 8336
rect 49876 8296 49916 8336
rect 49958 8296 49998 8336
rect 50040 8296 50080 8336
rect 64832 8296 64872 8336
rect 64914 8296 64954 8336
rect 64996 8296 65036 8336
rect 65078 8296 65118 8336
rect 65160 8296 65200 8336
rect 79952 8296 79992 8336
rect 80034 8296 80074 8336
rect 80116 8296 80156 8336
rect 80198 8296 80238 8336
rect 80280 8296 80320 8336
rect 95072 8296 95112 8336
rect 95154 8296 95194 8336
rect 95236 8296 95276 8336
rect 95318 8296 95358 8336
rect 95400 8296 95440 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 18232 7540 18272 7580
rect 18314 7540 18354 7580
rect 18396 7540 18436 7580
rect 18478 7540 18518 7580
rect 18560 7540 18600 7580
rect 33352 7540 33392 7580
rect 33434 7540 33474 7580
rect 33516 7540 33556 7580
rect 33598 7540 33638 7580
rect 33680 7540 33720 7580
rect 48472 7540 48512 7580
rect 48554 7540 48594 7580
rect 48636 7540 48676 7580
rect 48718 7540 48758 7580
rect 48800 7540 48840 7580
rect 63592 7540 63632 7580
rect 63674 7540 63714 7580
rect 63756 7540 63796 7580
rect 63838 7540 63878 7580
rect 63920 7540 63960 7580
rect 78712 7540 78752 7580
rect 78794 7540 78834 7580
rect 78876 7540 78916 7580
rect 78958 7540 78998 7580
rect 79040 7540 79080 7580
rect 93832 7540 93872 7580
rect 93914 7540 93954 7580
rect 93996 7540 94036 7580
rect 94078 7540 94118 7580
rect 94160 7540 94200 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 19472 6784 19512 6824
rect 19554 6784 19594 6824
rect 19636 6784 19676 6824
rect 19718 6784 19758 6824
rect 19800 6784 19840 6824
rect 34592 6784 34632 6824
rect 34674 6784 34714 6824
rect 34756 6784 34796 6824
rect 34838 6784 34878 6824
rect 34920 6784 34960 6824
rect 49712 6784 49752 6824
rect 49794 6784 49834 6824
rect 49876 6784 49916 6824
rect 49958 6784 49998 6824
rect 50040 6784 50080 6824
rect 64832 6784 64872 6824
rect 64914 6784 64954 6824
rect 64996 6784 65036 6824
rect 65078 6784 65118 6824
rect 65160 6784 65200 6824
rect 79952 6784 79992 6824
rect 80034 6784 80074 6824
rect 80116 6784 80156 6824
rect 80198 6784 80238 6824
rect 80280 6784 80320 6824
rect 95072 6784 95112 6824
rect 95154 6784 95194 6824
rect 95236 6784 95276 6824
rect 95318 6784 95358 6824
rect 95400 6784 95440 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 18232 6028 18272 6068
rect 18314 6028 18354 6068
rect 18396 6028 18436 6068
rect 18478 6028 18518 6068
rect 18560 6028 18600 6068
rect 33352 6028 33392 6068
rect 33434 6028 33474 6068
rect 33516 6028 33556 6068
rect 33598 6028 33638 6068
rect 33680 6028 33720 6068
rect 48472 6028 48512 6068
rect 48554 6028 48594 6068
rect 48636 6028 48676 6068
rect 48718 6028 48758 6068
rect 48800 6028 48840 6068
rect 63592 6028 63632 6068
rect 63674 6028 63714 6068
rect 63756 6028 63796 6068
rect 63838 6028 63878 6068
rect 63920 6028 63960 6068
rect 78712 6028 78752 6068
rect 78794 6028 78834 6068
rect 78876 6028 78916 6068
rect 78958 6028 78998 6068
rect 79040 6028 79080 6068
rect 93832 6028 93872 6068
rect 93914 6028 93954 6068
rect 93996 6028 94036 6068
rect 94078 6028 94118 6068
rect 94160 6028 94200 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 19472 5272 19512 5312
rect 19554 5272 19594 5312
rect 19636 5272 19676 5312
rect 19718 5272 19758 5312
rect 19800 5272 19840 5312
rect 34592 5272 34632 5312
rect 34674 5272 34714 5312
rect 34756 5272 34796 5312
rect 34838 5272 34878 5312
rect 34920 5272 34960 5312
rect 49712 5272 49752 5312
rect 49794 5272 49834 5312
rect 49876 5272 49916 5312
rect 49958 5272 49998 5312
rect 50040 5272 50080 5312
rect 64832 5272 64872 5312
rect 64914 5272 64954 5312
rect 64996 5272 65036 5312
rect 65078 5272 65118 5312
rect 65160 5272 65200 5312
rect 79952 5272 79992 5312
rect 80034 5272 80074 5312
rect 80116 5272 80156 5312
rect 80198 5272 80238 5312
rect 80280 5272 80320 5312
rect 95072 5272 95112 5312
rect 95154 5272 95194 5312
rect 95236 5272 95276 5312
rect 95318 5272 95358 5312
rect 95400 5272 95440 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 18232 4516 18272 4556
rect 18314 4516 18354 4556
rect 18396 4516 18436 4556
rect 18478 4516 18518 4556
rect 18560 4516 18600 4556
rect 33352 4516 33392 4556
rect 33434 4516 33474 4556
rect 33516 4516 33556 4556
rect 33598 4516 33638 4556
rect 33680 4516 33720 4556
rect 48472 4516 48512 4556
rect 48554 4516 48594 4556
rect 48636 4516 48676 4556
rect 48718 4516 48758 4556
rect 48800 4516 48840 4556
rect 63592 4516 63632 4556
rect 63674 4516 63714 4556
rect 63756 4516 63796 4556
rect 63838 4516 63878 4556
rect 63920 4516 63960 4556
rect 78712 4516 78752 4556
rect 78794 4516 78834 4556
rect 78876 4516 78916 4556
rect 78958 4516 78998 4556
rect 79040 4516 79080 4556
rect 93832 4516 93872 4556
rect 93914 4516 93954 4556
rect 93996 4516 94036 4556
rect 94078 4516 94118 4556
rect 94160 4516 94200 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 19472 3760 19512 3800
rect 19554 3760 19594 3800
rect 19636 3760 19676 3800
rect 19718 3760 19758 3800
rect 19800 3760 19840 3800
rect 34592 3760 34632 3800
rect 34674 3760 34714 3800
rect 34756 3760 34796 3800
rect 34838 3760 34878 3800
rect 34920 3760 34960 3800
rect 49712 3760 49752 3800
rect 49794 3760 49834 3800
rect 49876 3760 49916 3800
rect 49958 3760 49998 3800
rect 50040 3760 50080 3800
rect 64832 3760 64872 3800
rect 64914 3760 64954 3800
rect 64996 3760 65036 3800
rect 65078 3760 65118 3800
rect 65160 3760 65200 3800
rect 79952 3760 79992 3800
rect 80034 3760 80074 3800
rect 80116 3760 80156 3800
rect 80198 3760 80238 3800
rect 80280 3760 80320 3800
rect 95072 3760 95112 3800
rect 95154 3760 95194 3800
rect 95236 3760 95276 3800
rect 95318 3760 95358 3800
rect 95400 3760 95440 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 18232 3004 18272 3044
rect 18314 3004 18354 3044
rect 18396 3004 18436 3044
rect 18478 3004 18518 3044
rect 18560 3004 18600 3044
rect 33352 3004 33392 3044
rect 33434 3004 33474 3044
rect 33516 3004 33556 3044
rect 33598 3004 33638 3044
rect 33680 3004 33720 3044
rect 48472 3004 48512 3044
rect 48554 3004 48594 3044
rect 48636 3004 48676 3044
rect 48718 3004 48758 3044
rect 48800 3004 48840 3044
rect 63592 3004 63632 3044
rect 63674 3004 63714 3044
rect 63756 3004 63796 3044
rect 63838 3004 63878 3044
rect 63920 3004 63960 3044
rect 78712 3004 78752 3044
rect 78794 3004 78834 3044
rect 78876 3004 78916 3044
rect 78958 3004 78998 3044
rect 79040 3004 79080 3044
rect 93832 3004 93872 3044
rect 93914 3004 93954 3044
rect 93996 3004 94036 3044
rect 94078 3004 94118 3044
rect 94160 3004 94200 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 19472 2248 19512 2288
rect 19554 2248 19594 2288
rect 19636 2248 19676 2288
rect 19718 2248 19758 2288
rect 19800 2248 19840 2288
rect 34592 2248 34632 2288
rect 34674 2248 34714 2288
rect 34756 2248 34796 2288
rect 34838 2248 34878 2288
rect 34920 2248 34960 2288
rect 49712 2248 49752 2288
rect 49794 2248 49834 2288
rect 49876 2248 49916 2288
rect 49958 2248 49998 2288
rect 50040 2248 50080 2288
rect 64832 2248 64872 2288
rect 64914 2248 64954 2288
rect 64996 2248 65036 2288
rect 65078 2248 65118 2288
rect 65160 2248 65200 2288
rect 79952 2248 79992 2288
rect 80034 2248 80074 2288
rect 80116 2248 80156 2288
rect 80198 2248 80238 2288
rect 80280 2248 80320 2288
rect 95072 2248 95112 2288
rect 95154 2248 95194 2288
rect 95236 2248 95276 2288
rect 95318 2248 95358 2288
rect 95400 2248 95440 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 18232 1492 18272 1532
rect 18314 1492 18354 1532
rect 18396 1492 18436 1532
rect 18478 1492 18518 1532
rect 18560 1492 18600 1532
rect 33352 1492 33392 1532
rect 33434 1492 33474 1532
rect 33516 1492 33556 1532
rect 33598 1492 33638 1532
rect 33680 1492 33720 1532
rect 48472 1492 48512 1532
rect 48554 1492 48594 1532
rect 48636 1492 48676 1532
rect 48718 1492 48758 1532
rect 48800 1492 48840 1532
rect 63592 1492 63632 1532
rect 63674 1492 63714 1532
rect 63756 1492 63796 1532
rect 63838 1492 63878 1532
rect 63920 1492 63960 1532
rect 78712 1492 78752 1532
rect 78794 1492 78834 1532
rect 78876 1492 78916 1532
rect 78958 1492 78998 1532
rect 79040 1492 79080 1532
rect 93832 1492 93872 1532
rect 93914 1492 93954 1532
rect 93996 1492 94036 1532
rect 94078 1492 94118 1532
rect 94160 1492 94200 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 19472 736 19512 776
rect 19554 736 19594 776
rect 19636 736 19676 776
rect 19718 736 19758 776
rect 19800 736 19840 776
rect 34592 736 34632 776
rect 34674 736 34714 776
rect 34756 736 34796 776
rect 34838 736 34878 776
rect 34920 736 34960 776
rect 49712 736 49752 776
rect 49794 736 49834 776
rect 49876 736 49916 776
rect 49958 736 49998 776
rect 50040 736 50080 776
rect 64832 736 64872 776
rect 64914 736 64954 776
rect 64996 736 65036 776
rect 65078 736 65118 776
rect 65160 736 65200 776
rect 79952 736 79992 776
rect 80034 736 80074 776
rect 80116 736 80156 776
rect 80198 736 80238 776
rect 80280 736 80320 776
rect 95072 736 95112 776
rect 95154 736 95194 776
rect 95236 736 95276 776
rect 95318 736 95358 776
rect 95400 736 95440 776
<< metal5 >>
rect 4343 38599 4729 38618
rect 4343 38576 4409 38599
rect 4495 38576 4577 38599
rect 4663 38576 4729 38599
rect 4343 38536 4352 38576
rect 4392 38536 4409 38576
rect 4495 38536 4516 38576
rect 4556 38536 4577 38576
rect 4663 38536 4680 38576
rect 4720 38536 4729 38576
rect 4343 38513 4409 38536
rect 4495 38513 4577 38536
rect 4663 38513 4729 38536
rect 4343 38494 4729 38513
rect 19463 38599 19849 38618
rect 19463 38576 19529 38599
rect 19615 38576 19697 38599
rect 19783 38576 19849 38599
rect 19463 38536 19472 38576
rect 19512 38536 19529 38576
rect 19615 38536 19636 38576
rect 19676 38536 19697 38576
rect 19783 38536 19800 38576
rect 19840 38536 19849 38576
rect 19463 38513 19529 38536
rect 19615 38513 19697 38536
rect 19783 38513 19849 38536
rect 19463 38494 19849 38513
rect 34583 38599 34969 38618
rect 34583 38576 34649 38599
rect 34735 38576 34817 38599
rect 34903 38576 34969 38599
rect 34583 38536 34592 38576
rect 34632 38536 34649 38576
rect 34735 38536 34756 38576
rect 34796 38536 34817 38576
rect 34903 38536 34920 38576
rect 34960 38536 34969 38576
rect 34583 38513 34649 38536
rect 34735 38513 34817 38536
rect 34903 38513 34969 38536
rect 34583 38494 34969 38513
rect 49703 38599 50089 38618
rect 49703 38576 49769 38599
rect 49855 38576 49937 38599
rect 50023 38576 50089 38599
rect 49703 38536 49712 38576
rect 49752 38536 49769 38576
rect 49855 38536 49876 38576
rect 49916 38536 49937 38576
rect 50023 38536 50040 38576
rect 50080 38536 50089 38576
rect 49703 38513 49769 38536
rect 49855 38513 49937 38536
rect 50023 38513 50089 38536
rect 49703 38494 50089 38513
rect 64823 38599 65209 38618
rect 64823 38576 64889 38599
rect 64975 38576 65057 38599
rect 65143 38576 65209 38599
rect 64823 38536 64832 38576
rect 64872 38536 64889 38576
rect 64975 38536 64996 38576
rect 65036 38536 65057 38576
rect 65143 38536 65160 38576
rect 65200 38536 65209 38576
rect 64823 38513 64889 38536
rect 64975 38513 65057 38536
rect 65143 38513 65209 38536
rect 64823 38494 65209 38513
rect 79943 38599 80329 38618
rect 79943 38576 80009 38599
rect 80095 38576 80177 38599
rect 80263 38576 80329 38599
rect 79943 38536 79952 38576
rect 79992 38536 80009 38576
rect 80095 38536 80116 38576
rect 80156 38536 80177 38576
rect 80263 38536 80280 38576
rect 80320 38536 80329 38576
rect 79943 38513 80009 38536
rect 80095 38513 80177 38536
rect 80263 38513 80329 38536
rect 79943 38494 80329 38513
rect 95063 38599 95449 38618
rect 95063 38576 95129 38599
rect 95215 38576 95297 38599
rect 95383 38576 95449 38599
rect 95063 38536 95072 38576
rect 95112 38536 95129 38576
rect 95215 38536 95236 38576
rect 95276 38536 95297 38576
rect 95383 38536 95400 38576
rect 95440 38536 95449 38576
rect 95063 38513 95129 38536
rect 95215 38513 95297 38536
rect 95383 38513 95449 38536
rect 95063 38494 95449 38513
rect 3103 37843 3489 37862
rect 3103 37820 3169 37843
rect 3255 37820 3337 37843
rect 3423 37820 3489 37843
rect 3103 37780 3112 37820
rect 3152 37780 3169 37820
rect 3255 37780 3276 37820
rect 3316 37780 3337 37820
rect 3423 37780 3440 37820
rect 3480 37780 3489 37820
rect 3103 37757 3169 37780
rect 3255 37757 3337 37780
rect 3423 37757 3489 37780
rect 3103 37738 3489 37757
rect 18223 37843 18609 37862
rect 18223 37820 18289 37843
rect 18375 37820 18457 37843
rect 18543 37820 18609 37843
rect 18223 37780 18232 37820
rect 18272 37780 18289 37820
rect 18375 37780 18396 37820
rect 18436 37780 18457 37820
rect 18543 37780 18560 37820
rect 18600 37780 18609 37820
rect 18223 37757 18289 37780
rect 18375 37757 18457 37780
rect 18543 37757 18609 37780
rect 18223 37738 18609 37757
rect 33343 37843 33729 37862
rect 33343 37820 33409 37843
rect 33495 37820 33577 37843
rect 33663 37820 33729 37843
rect 33343 37780 33352 37820
rect 33392 37780 33409 37820
rect 33495 37780 33516 37820
rect 33556 37780 33577 37820
rect 33663 37780 33680 37820
rect 33720 37780 33729 37820
rect 33343 37757 33409 37780
rect 33495 37757 33577 37780
rect 33663 37757 33729 37780
rect 33343 37738 33729 37757
rect 48463 37843 48849 37862
rect 48463 37820 48529 37843
rect 48615 37820 48697 37843
rect 48783 37820 48849 37843
rect 48463 37780 48472 37820
rect 48512 37780 48529 37820
rect 48615 37780 48636 37820
rect 48676 37780 48697 37820
rect 48783 37780 48800 37820
rect 48840 37780 48849 37820
rect 48463 37757 48529 37780
rect 48615 37757 48697 37780
rect 48783 37757 48849 37780
rect 48463 37738 48849 37757
rect 63583 37843 63969 37862
rect 63583 37820 63649 37843
rect 63735 37820 63817 37843
rect 63903 37820 63969 37843
rect 63583 37780 63592 37820
rect 63632 37780 63649 37820
rect 63735 37780 63756 37820
rect 63796 37780 63817 37820
rect 63903 37780 63920 37820
rect 63960 37780 63969 37820
rect 63583 37757 63649 37780
rect 63735 37757 63817 37780
rect 63903 37757 63969 37780
rect 63583 37738 63969 37757
rect 78703 37843 79089 37862
rect 78703 37820 78769 37843
rect 78855 37820 78937 37843
rect 79023 37820 79089 37843
rect 78703 37780 78712 37820
rect 78752 37780 78769 37820
rect 78855 37780 78876 37820
rect 78916 37780 78937 37820
rect 79023 37780 79040 37820
rect 79080 37780 79089 37820
rect 78703 37757 78769 37780
rect 78855 37757 78937 37780
rect 79023 37757 79089 37780
rect 78703 37738 79089 37757
rect 93823 37843 94209 37862
rect 93823 37820 93889 37843
rect 93975 37820 94057 37843
rect 94143 37820 94209 37843
rect 93823 37780 93832 37820
rect 93872 37780 93889 37820
rect 93975 37780 93996 37820
rect 94036 37780 94057 37820
rect 94143 37780 94160 37820
rect 94200 37780 94209 37820
rect 93823 37757 93889 37780
rect 93975 37757 94057 37780
rect 94143 37757 94209 37780
rect 93823 37738 94209 37757
rect 4343 37087 4729 37106
rect 4343 37064 4409 37087
rect 4495 37064 4577 37087
rect 4663 37064 4729 37087
rect 4343 37024 4352 37064
rect 4392 37024 4409 37064
rect 4495 37024 4516 37064
rect 4556 37024 4577 37064
rect 4663 37024 4680 37064
rect 4720 37024 4729 37064
rect 4343 37001 4409 37024
rect 4495 37001 4577 37024
rect 4663 37001 4729 37024
rect 4343 36982 4729 37001
rect 19463 37087 19849 37106
rect 19463 37064 19529 37087
rect 19615 37064 19697 37087
rect 19783 37064 19849 37087
rect 19463 37024 19472 37064
rect 19512 37024 19529 37064
rect 19615 37024 19636 37064
rect 19676 37024 19697 37064
rect 19783 37024 19800 37064
rect 19840 37024 19849 37064
rect 19463 37001 19529 37024
rect 19615 37001 19697 37024
rect 19783 37001 19849 37024
rect 19463 36982 19849 37001
rect 34583 37087 34969 37106
rect 34583 37064 34649 37087
rect 34735 37064 34817 37087
rect 34903 37064 34969 37087
rect 34583 37024 34592 37064
rect 34632 37024 34649 37064
rect 34735 37024 34756 37064
rect 34796 37024 34817 37064
rect 34903 37024 34920 37064
rect 34960 37024 34969 37064
rect 34583 37001 34649 37024
rect 34735 37001 34817 37024
rect 34903 37001 34969 37024
rect 34583 36982 34969 37001
rect 49703 37087 50089 37106
rect 49703 37064 49769 37087
rect 49855 37064 49937 37087
rect 50023 37064 50089 37087
rect 49703 37024 49712 37064
rect 49752 37024 49769 37064
rect 49855 37024 49876 37064
rect 49916 37024 49937 37064
rect 50023 37024 50040 37064
rect 50080 37024 50089 37064
rect 49703 37001 49769 37024
rect 49855 37001 49937 37024
rect 50023 37001 50089 37024
rect 49703 36982 50089 37001
rect 64823 37087 65209 37106
rect 64823 37064 64889 37087
rect 64975 37064 65057 37087
rect 65143 37064 65209 37087
rect 64823 37024 64832 37064
rect 64872 37024 64889 37064
rect 64975 37024 64996 37064
rect 65036 37024 65057 37064
rect 65143 37024 65160 37064
rect 65200 37024 65209 37064
rect 64823 37001 64889 37024
rect 64975 37001 65057 37024
rect 65143 37001 65209 37024
rect 64823 36982 65209 37001
rect 79943 37087 80329 37106
rect 79943 37064 80009 37087
rect 80095 37064 80177 37087
rect 80263 37064 80329 37087
rect 79943 37024 79952 37064
rect 79992 37024 80009 37064
rect 80095 37024 80116 37064
rect 80156 37024 80177 37064
rect 80263 37024 80280 37064
rect 80320 37024 80329 37064
rect 79943 37001 80009 37024
rect 80095 37001 80177 37024
rect 80263 37001 80329 37024
rect 79943 36982 80329 37001
rect 95063 37087 95449 37106
rect 95063 37064 95129 37087
rect 95215 37064 95297 37087
rect 95383 37064 95449 37087
rect 95063 37024 95072 37064
rect 95112 37024 95129 37064
rect 95215 37024 95236 37064
rect 95276 37024 95297 37064
rect 95383 37024 95400 37064
rect 95440 37024 95449 37064
rect 95063 37001 95129 37024
rect 95215 37001 95297 37024
rect 95383 37001 95449 37024
rect 95063 36982 95449 37001
rect 3103 36331 3489 36350
rect 3103 36308 3169 36331
rect 3255 36308 3337 36331
rect 3423 36308 3489 36331
rect 3103 36268 3112 36308
rect 3152 36268 3169 36308
rect 3255 36268 3276 36308
rect 3316 36268 3337 36308
rect 3423 36268 3440 36308
rect 3480 36268 3489 36308
rect 3103 36245 3169 36268
rect 3255 36245 3337 36268
rect 3423 36245 3489 36268
rect 3103 36226 3489 36245
rect 18223 36331 18609 36350
rect 18223 36308 18289 36331
rect 18375 36308 18457 36331
rect 18543 36308 18609 36331
rect 18223 36268 18232 36308
rect 18272 36268 18289 36308
rect 18375 36268 18396 36308
rect 18436 36268 18457 36308
rect 18543 36268 18560 36308
rect 18600 36268 18609 36308
rect 18223 36245 18289 36268
rect 18375 36245 18457 36268
rect 18543 36245 18609 36268
rect 18223 36226 18609 36245
rect 33343 36331 33729 36350
rect 33343 36308 33409 36331
rect 33495 36308 33577 36331
rect 33663 36308 33729 36331
rect 33343 36268 33352 36308
rect 33392 36268 33409 36308
rect 33495 36268 33516 36308
rect 33556 36268 33577 36308
rect 33663 36268 33680 36308
rect 33720 36268 33729 36308
rect 33343 36245 33409 36268
rect 33495 36245 33577 36268
rect 33663 36245 33729 36268
rect 33343 36226 33729 36245
rect 48463 36331 48849 36350
rect 48463 36308 48529 36331
rect 48615 36308 48697 36331
rect 48783 36308 48849 36331
rect 48463 36268 48472 36308
rect 48512 36268 48529 36308
rect 48615 36268 48636 36308
rect 48676 36268 48697 36308
rect 48783 36268 48800 36308
rect 48840 36268 48849 36308
rect 48463 36245 48529 36268
rect 48615 36245 48697 36268
rect 48783 36245 48849 36268
rect 48463 36226 48849 36245
rect 63583 36331 63969 36350
rect 63583 36308 63649 36331
rect 63735 36308 63817 36331
rect 63903 36308 63969 36331
rect 63583 36268 63592 36308
rect 63632 36268 63649 36308
rect 63735 36268 63756 36308
rect 63796 36268 63817 36308
rect 63903 36268 63920 36308
rect 63960 36268 63969 36308
rect 63583 36245 63649 36268
rect 63735 36245 63817 36268
rect 63903 36245 63969 36268
rect 63583 36226 63969 36245
rect 78703 36331 79089 36350
rect 78703 36308 78769 36331
rect 78855 36308 78937 36331
rect 79023 36308 79089 36331
rect 78703 36268 78712 36308
rect 78752 36268 78769 36308
rect 78855 36268 78876 36308
rect 78916 36268 78937 36308
rect 79023 36268 79040 36308
rect 79080 36268 79089 36308
rect 78703 36245 78769 36268
rect 78855 36245 78937 36268
rect 79023 36245 79089 36268
rect 78703 36226 79089 36245
rect 93823 36331 94209 36350
rect 93823 36308 93889 36331
rect 93975 36308 94057 36331
rect 94143 36308 94209 36331
rect 93823 36268 93832 36308
rect 93872 36268 93889 36308
rect 93975 36268 93996 36308
rect 94036 36268 94057 36308
rect 94143 36268 94160 36308
rect 94200 36268 94209 36308
rect 93823 36245 93889 36268
rect 93975 36245 94057 36268
rect 94143 36245 94209 36268
rect 93823 36226 94209 36245
rect 4343 35575 4729 35594
rect 4343 35552 4409 35575
rect 4495 35552 4577 35575
rect 4663 35552 4729 35575
rect 4343 35512 4352 35552
rect 4392 35512 4409 35552
rect 4495 35512 4516 35552
rect 4556 35512 4577 35552
rect 4663 35512 4680 35552
rect 4720 35512 4729 35552
rect 4343 35489 4409 35512
rect 4495 35489 4577 35512
rect 4663 35489 4729 35512
rect 4343 35470 4729 35489
rect 19463 35575 19849 35594
rect 19463 35552 19529 35575
rect 19615 35552 19697 35575
rect 19783 35552 19849 35575
rect 19463 35512 19472 35552
rect 19512 35512 19529 35552
rect 19615 35512 19636 35552
rect 19676 35512 19697 35552
rect 19783 35512 19800 35552
rect 19840 35512 19849 35552
rect 19463 35489 19529 35512
rect 19615 35489 19697 35512
rect 19783 35489 19849 35512
rect 19463 35470 19849 35489
rect 34583 35575 34969 35594
rect 34583 35552 34649 35575
rect 34735 35552 34817 35575
rect 34903 35552 34969 35575
rect 34583 35512 34592 35552
rect 34632 35512 34649 35552
rect 34735 35512 34756 35552
rect 34796 35512 34817 35552
rect 34903 35512 34920 35552
rect 34960 35512 34969 35552
rect 34583 35489 34649 35512
rect 34735 35489 34817 35512
rect 34903 35489 34969 35512
rect 34583 35470 34969 35489
rect 49703 35575 50089 35594
rect 49703 35552 49769 35575
rect 49855 35552 49937 35575
rect 50023 35552 50089 35575
rect 49703 35512 49712 35552
rect 49752 35512 49769 35552
rect 49855 35512 49876 35552
rect 49916 35512 49937 35552
rect 50023 35512 50040 35552
rect 50080 35512 50089 35552
rect 49703 35489 49769 35512
rect 49855 35489 49937 35512
rect 50023 35489 50089 35512
rect 49703 35470 50089 35489
rect 64823 35575 65209 35594
rect 64823 35552 64889 35575
rect 64975 35552 65057 35575
rect 65143 35552 65209 35575
rect 64823 35512 64832 35552
rect 64872 35512 64889 35552
rect 64975 35512 64996 35552
rect 65036 35512 65057 35552
rect 65143 35512 65160 35552
rect 65200 35512 65209 35552
rect 64823 35489 64889 35512
rect 64975 35489 65057 35512
rect 65143 35489 65209 35512
rect 64823 35470 65209 35489
rect 79943 35575 80329 35594
rect 79943 35552 80009 35575
rect 80095 35552 80177 35575
rect 80263 35552 80329 35575
rect 79943 35512 79952 35552
rect 79992 35512 80009 35552
rect 80095 35512 80116 35552
rect 80156 35512 80177 35552
rect 80263 35512 80280 35552
rect 80320 35512 80329 35552
rect 79943 35489 80009 35512
rect 80095 35489 80177 35512
rect 80263 35489 80329 35512
rect 79943 35470 80329 35489
rect 95063 35575 95449 35594
rect 95063 35552 95129 35575
rect 95215 35552 95297 35575
rect 95383 35552 95449 35575
rect 95063 35512 95072 35552
rect 95112 35512 95129 35552
rect 95215 35512 95236 35552
rect 95276 35512 95297 35552
rect 95383 35512 95400 35552
rect 95440 35512 95449 35552
rect 95063 35489 95129 35512
rect 95215 35489 95297 35512
rect 95383 35489 95449 35512
rect 95063 35470 95449 35489
rect 3103 34819 3489 34838
rect 3103 34796 3169 34819
rect 3255 34796 3337 34819
rect 3423 34796 3489 34819
rect 3103 34756 3112 34796
rect 3152 34756 3169 34796
rect 3255 34756 3276 34796
rect 3316 34756 3337 34796
rect 3423 34756 3440 34796
rect 3480 34756 3489 34796
rect 3103 34733 3169 34756
rect 3255 34733 3337 34756
rect 3423 34733 3489 34756
rect 3103 34714 3489 34733
rect 18223 34819 18609 34838
rect 18223 34796 18289 34819
rect 18375 34796 18457 34819
rect 18543 34796 18609 34819
rect 18223 34756 18232 34796
rect 18272 34756 18289 34796
rect 18375 34756 18396 34796
rect 18436 34756 18457 34796
rect 18543 34756 18560 34796
rect 18600 34756 18609 34796
rect 18223 34733 18289 34756
rect 18375 34733 18457 34756
rect 18543 34733 18609 34756
rect 18223 34714 18609 34733
rect 33343 34819 33729 34838
rect 33343 34796 33409 34819
rect 33495 34796 33577 34819
rect 33663 34796 33729 34819
rect 33343 34756 33352 34796
rect 33392 34756 33409 34796
rect 33495 34756 33516 34796
rect 33556 34756 33577 34796
rect 33663 34756 33680 34796
rect 33720 34756 33729 34796
rect 33343 34733 33409 34756
rect 33495 34733 33577 34756
rect 33663 34733 33729 34756
rect 33343 34714 33729 34733
rect 48463 34819 48849 34838
rect 48463 34796 48529 34819
rect 48615 34796 48697 34819
rect 48783 34796 48849 34819
rect 48463 34756 48472 34796
rect 48512 34756 48529 34796
rect 48615 34756 48636 34796
rect 48676 34756 48697 34796
rect 48783 34756 48800 34796
rect 48840 34756 48849 34796
rect 48463 34733 48529 34756
rect 48615 34733 48697 34756
rect 48783 34733 48849 34756
rect 48463 34714 48849 34733
rect 63583 34819 63969 34838
rect 63583 34796 63649 34819
rect 63735 34796 63817 34819
rect 63903 34796 63969 34819
rect 63583 34756 63592 34796
rect 63632 34756 63649 34796
rect 63735 34756 63756 34796
rect 63796 34756 63817 34796
rect 63903 34756 63920 34796
rect 63960 34756 63969 34796
rect 63583 34733 63649 34756
rect 63735 34733 63817 34756
rect 63903 34733 63969 34756
rect 63583 34714 63969 34733
rect 78703 34819 79089 34838
rect 78703 34796 78769 34819
rect 78855 34796 78937 34819
rect 79023 34796 79089 34819
rect 78703 34756 78712 34796
rect 78752 34756 78769 34796
rect 78855 34756 78876 34796
rect 78916 34756 78937 34796
rect 79023 34756 79040 34796
rect 79080 34756 79089 34796
rect 78703 34733 78769 34756
rect 78855 34733 78937 34756
rect 79023 34733 79089 34756
rect 78703 34714 79089 34733
rect 93823 34819 94209 34838
rect 93823 34796 93889 34819
rect 93975 34796 94057 34819
rect 94143 34796 94209 34819
rect 93823 34756 93832 34796
rect 93872 34756 93889 34796
rect 93975 34756 93996 34796
rect 94036 34756 94057 34796
rect 94143 34756 94160 34796
rect 94200 34756 94209 34796
rect 93823 34733 93889 34756
rect 93975 34733 94057 34756
rect 94143 34733 94209 34756
rect 93823 34714 94209 34733
rect 4343 34063 4729 34082
rect 4343 34040 4409 34063
rect 4495 34040 4577 34063
rect 4663 34040 4729 34063
rect 4343 34000 4352 34040
rect 4392 34000 4409 34040
rect 4495 34000 4516 34040
rect 4556 34000 4577 34040
rect 4663 34000 4680 34040
rect 4720 34000 4729 34040
rect 4343 33977 4409 34000
rect 4495 33977 4577 34000
rect 4663 33977 4729 34000
rect 4343 33958 4729 33977
rect 19463 34063 19849 34082
rect 19463 34040 19529 34063
rect 19615 34040 19697 34063
rect 19783 34040 19849 34063
rect 19463 34000 19472 34040
rect 19512 34000 19529 34040
rect 19615 34000 19636 34040
rect 19676 34000 19697 34040
rect 19783 34000 19800 34040
rect 19840 34000 19849 34040
rect 19463 33977 19529 34000
rect 19615 33977 19697 34000
rect 19783 33977 19849 34000
rect 19463 33958 19849 33977
rect 34583 34063 34969 34082
rect 34583 34040 34649 34063
rect 34735 34040 34817 34063
rect 34903 34040 34969 34063
rect 34583 34000 34592 34040
rect 34632 34000 34649 34040
rect 34735 34000 34756 34040
rect 34796 34000 34817 34040
rect 34903 34000 34920 34040
rect 34960 34000 34969 34040
rect 34583 33977 34649 34000
rect 34735 33977 34817 34000
rect 34903 33977 34969 34000
rect 34583 33958 34969 33977
rect 49703 34063 50089 34082
rect 49703 34040 49769 34063
rect 49855 34040 49937 34063
rect 50023 34040 50089 34063
rect 49703 34000 49712 34040
rect 49752 34000 49769 34040
rect 49855 34000 49876 34040
rect 49916 34000 49937 34040
rect 50023 34000 50040 34040
rect 50080 34000 50089 34040
rect 49703 33977 49769 34000
rect 49855 33977 49937 34000
rect 50023 33977 50089 34000
rect 49703 33958 50089 33977
rect 64823 34063 65209 34082
rect 64823 34040 64889 34063
rect 64975 34040 65057 34063
rect 65143 34040 65209 34063
rect 64823 34000 64832 34040
rect 64872 34000 64889 34040
rect 64975 34000 64996 34040
rect 65036 34000 65057 34040
rect 65143 34000 65160 34040
rect 65200 34000 65209 34040
rect 64823 33977 64889 34000
rect 64975 33977 65057 34000
rect 65143 33977 65209 34000
rect 64823 33958 65209 33977
rect 79943 34063 80329 34082
rect 79943 34040 80009 34063
rect 80095 34040 80177 34063
rect 80263 34040 80329 34063
rect 79943 34000 79952 34040
rect 79992 34000 80009 34040
rect 80095 34000 80116 34040
rect 80156 34000 80177 34040
rect 80263 34000 80280 34040
rect 80320 34000 80329 34040
rect 79943 33977 80009 34000
rect 80095 33977 80177 34000
rect 80263 33977 80329 34000
rect 79943 33958 80329 33977
rect 95063 34063 95449 34082
rect 95063 34040 95129 34063
rect 95215 34040 95297 34063
rect 95383 34040 95449 34063
rect 95063 34000 95072 34040
rect 95112 34000 95129 34040
rect 95215 34000 95236 34040
rect 95276 34000 95297 34040
rect 95383 34000 95400 34040
rect 95440 34000 95449 34040
rect 95063 33977 95129 34000
rect 95215 33977 95297 34000
rect 95383 33977 95449 34000
rect 95063 33958 95449 33977
rect 3103 33307 3489 33326
rect 3103 33284 3169 33307
rect 3255 33284 3337 33307
rect 3423 33284 3489 33307
rect 3103 33244 3112 33284
rect 3152 33244 3169 33284
rect 3255 33244 3276 33284
rect 3316 33244 3337 33284
rect 3423 33244 3440 33284
rect 3480 33244 3489 33284
rect 3103 33221 3169 33244
rect 3255 33221 3337 33244
rect 3423 33221 3489 33244
rect 3103 33202 3489 33221
rect 18223 33307 18609 33326
rect 18223 33284 18289 33307
rect 18375 33284 18457 33307
rect 18543 33284 18609 33307
rect 18223 33244 18232 33284
rect 18272 33244 18289 33284
rect 18375 33244 18396 33284
rect 18436 33244 18457 33284
rect 18543 33244 18560 33284
rect 18600 33244 18609 33284
rect 18223 33221 18289 33244
rect 18375 33221 18457 33244
rect 18543 33221 18609 33244
rect 18223 33202 18609 33221
rect 33343 33307 33729 33326
rect 33343 33284 33409 33307
rect 33495 33284 33577 33307
rect 33663 33284 33729 33307
rect 33343 33244 33352 33284
rect 33392 33244 33409 33284
rect 33495 33244 33516 33284
rect 33556 33244 33577 33284
rect 33663 33244 33680 33284
rect 33720 33244 33729 33284
rect 33343 33221 33409 33244
rect 33495 33221 33577 33244
rect 33663 33221 33729 33244
rect 33343 33202 33729 33221
rect 48463 33307 48849 33326
rect 48463 33284 48529 33307
rect 48615 33284 48697 33307
rect 48783 33284 48849 33307
rect 48463 33244 48472 33284
rect 48512 33244 48529 33284
rect 48615 33244 48636 33284
rect 48676 33244 48697 33284
rect 48783 33244 48800 33284
rect 48840 33244 48849 33284
rect 48463 33221 48529 33244
rect 48615 33221 48697 33244
rect 48783 33221 48849 33244
rect 48463 33202 48849 33221
rect 63583 33307 63969 33326
rect 63583 33284 63649 33307
rect 63735 33284 63817 33307
rect 63903 33284 63969 33307
rect 63583 33244 63592 33284
rect 63632 33244 63649 33284
rect 63735 33244 63756 33284
rect 63796 33244 63817 33284
rect 63903 33244 63920 33284
rect 63960 33244 63969 33284
rect 63583 33221 63649 33244
rect 63735 33221 63817 33244
rect 63903 33221 63969 33244
rect 63583 33202 63969 33221
rect 78703 33307 79089 33326
rect 78703 33284 78769 33307
rect 78855 33284 78937 33307
rect 79023 33284 79089 33307
rect 78703 33244 78712 33284
rect 78752 33244 78769 33284
rect 78855 33244 78876 33284
rect 78916 33244 78937 33284
rect 79023 33244 79040 33284
rect 79080 33244 79089 33284
rect 78703 33221 78769 33244
rect 78855 33221 78937 33244
rect 79023 33221 79089 33244
rect 78703 33202 79089 33221
rect 93823 33307 94209 33326
rect 93823 33284 93889 33307
rect 93975 33284 94057 33307
rect 94143 33284 94209 33307
rect 93823 33244 93832 33284
rect 93872 33244 93889 33284
rect 93975 33244 93996 33284
rect 94036 33244 94057 33284
rect 94143 33244 94160 33284
rect 94200 33244 94209 33284
rect 93823 33221 93889 33244
rect 93975 33221 94057 33244
rect 94143 33221 94209 33244
rect 93823 33202 94209 33221
rect 4343 32551 4729 32570
rect 4343 32528 4409 32551
rect 4495 32528 4577 32551
rect 4663 32528 4729 32551
rect 4343 32488 4352 32528
rect 4392 32488 4409 32528
rect 4495 32488 4516 32528
rect 4556 32488 4577 32528
rect 4663 32488 4680 32528
rect 4720 32488 4729 32528
rect 4343 32465 4409 32488
rect 4495 32465 4577 32488
rect 4663 32465 4729 32488
rect 4343 32446 4729 32465
rect 19463 32551 19849 32570
rect 19463 32528 19529 32551
rect 19615 32528 19697 32551
rect 19783 32528 19849 32551
rect 19463 32488 19472 32528
rect 19512 32488 19529 32528
rect 19615 32488 19636 32528
rect 19676 32488 19697 32528
rect 19783 32488 19800 32528
rect 19840 32488 19849 32528
rect 19463 32465 19529 32488
rect 19615 32465 19697 32488
rect 19783 32465 19849 32488
rect 19463 32446 19849 32465
rect 34583 32551 34969 32570
rect 34583 32528 34649 32551
rect 34735 32528 34817 32551
rect 34903 32528 34969 32551
rect 34583 32488 34592 32528
rect 34632 32488 34649 32528
rect 34735 32488 34756 32528
rect 34796 32488 34817 32528
rect 34903 32488 34920 32528
rect 34960 32488 34969 32528
rect 34583 32465 34649 32488
rect 34735 32465 34817 32488
rect 34903 32465 34969 32488
rect 34583 32446 34969 32465
rect 49703 32551 50089 32570
rect 49703 32528 49769 32551
rect 49855 32528 49937 32551
rect 50023 32528 50089 32551
rect 49703 32488 49712 32528
rect 49752 32488 49769 32528
rect 49855 32488 49876 32528
rect 49916 32488 49937 32528
rect 50023 32488 50040 32528
rect 50080 32488 50089 32528
rect 49703 32465 49769 32488
rect 49855 32465 49937 32488
rect 50023 32465 50089 32488
rect 49703 32446 50089 32465
rect 64823 32551 65209 32570
rect 64823 32528 64889 32551
rect 64975 32528 65057 32551
rect 65143 32528 65209 32551
rect 64823 32488 64832 32528
rect 64872 32488 64889 32528
rect 64975 32488 64996 32528
rect 65036 32488 65057 32528
rect 65143 32488 65160 32528
rect 65200 32488 65209 32528
rect 64823 32465 64889 32488
rect 64975 32465 65057 32488
rect 65143 32465 65209 32488
rect 64823 32446 65209 32465
rect 79943 32551 80329 32570
rect 79943 32528 80009 32551
rect 80095 32528 80177 32551
rect 80263 32528 80329 32551
rect 79943 32488 79952 32528
rect 79992 32488 80009 32528
rect 80095 32488 80116 32528
rect 80156 32488 80177 32528
rect 80263 32488 80280 32528
rect 80320 32488 80329 32528
rect 79943 32465 80009 32488
rect 80095 32465 80177 32488
rect 80263 32465 80329 32488
rect 79943 32446 80329 32465
rect 95063 32551 95449 32570
rect 95063 32528 95129 32551
rect 95215 32528 95297 32551
rect 95383 32528 95449 32551
rect 95063 32488 95072 32528
rect 95112 32488 95129 32528
rect 95215 32488 95236 32528
rect 95276 32488 95297 32528
rect 95383 32488 95400 32528
rect 95440 32488 95449 32528
rect 95063 32465 95129 32488
rect 95215 32465 95297 32488
rect 95383 32465 95449 32488
rect 95063 32446 95449 32465
rect 3103 31795 3489 31814
rect 3103 31772 3169 31795
rect 3255 31772 3337 31795
rect 3423 31772 3489 31795
rect 3103 31732 3112 31772
rect 3152 31732 3169 31772
rect 3255 31732 3276 31772
rect 3316 31732 3337 31772
rect 3423 31732 3440 31772
rect 3480 31732 3489 31772
rect 3103 31709 3169 31732
rect 3255 31709 3337 31732
rect 3423 31709 3489 31732
rect 3103 31690 3489 31709
rect 18223 31795 18609 31814
rect 18223 31772 18289 31795
rect 18375 31772 18457 31795
rect 18543 31772 18609 31795
rect 18223 31732 18232 31772
rect 18272 31732 18289 31772
rect 18375 31732 18396 31772
rect 18436 31732 18457 31772
rect 18543 31732 18560 31772
rect 18600 31732 18609 31772
rect 18223 31709 18289 31732
rect 18375 31709 18457 31732
rect 18543 31709 18609 31732
rect 18223 31690 18609 31709
rect 33343 31795 33729 31814
rect 33343 31772 33409 31795
rect 33495 31772 33577 31795
rect 33663 31772 33729 31795
rect 33343 31732 33352 31772
rect 33392 31732 33409 31772
rect 33495 31732 33516 31772
rect 33556 31732 33577 31772
rect 33663 31732 33680 31772
rect 33720 31732 33729 31772
rect 33343 31709 33409 31732
rect 33495 31709 33577 31732
rect 33663 31709 33729 31732
rect 33343 31690 33729 31709
rect 48463 31795 48849 31814
rect 48463 31772 48529 31795
rect 48615 31772 48697 31795
rect 48783 31772 48849 31795
rect 48463 31732 48472 31772
rect 48512 31732 48529 31772
rect 48615 31732 48636 31772
rect 48676 31732 48697 31772
rect 48783 31732 48800 31772
rect 48840 31732 48849 31772
rect 48463 31709 48529 31732
rect 48615 31709 48697 31732
rect 48783 31709 48849 31732
rect 48463 31690 48849 31709
rect 63583 31795 63969 31814
rect 63583 31772 63649 31795
rect 63735 31772 63817 31795
rect 63903 31772 63969 31795
rect 63583 31732 63592 31772
rect 63632 31732 63649 31772
rect 63735 31732 63756 31772
rect 63796 31732 63817 31772
rect 63903 31732 63920 31772
rect 63960 31732 63969 31772
rect 63583 31709 63649 31732
rect 63735 31709 63817 31732
rect 63903 31709 63969 31732
rect 63583 31690 63969 31709
rect 78703 31795 79089 31814
rect 78703 31772 78769 31795
rect 78855 31772 78937 31795
rect 79023 31772 79089 31795
rect 78703 31732 78712 31772
rect 78752 31732 78769 31772
rect 78855 31732 78876 31772
rect 78916 31732 78937 31772
rect 79023 31732 79040 31772
rect 79080 31732 79089 31772
rect 78703 31709 78769 31732
rect 78855 31709 78937 31732
rect 79023 31709 79089 31732
rect 78703 31690 79089 31709
rect 93823 31795 94209 31814
rect 93823 31772 93889 31795
rect 93975 31772 94057 31795
rect 94143 31772 94209 31795
rect 93823 31732 93832 31772
rect 93872 31732 93889 31772
rect 93975 31732 93996 31772
rect 94036 31732 94057 31772
rect 94143 31732 94160 31772
rect 94200 31732 94209 31772
rect 93823 31709 93889 31732
rect 93975 31709 94057 31732
rect 94143 31709 94209 31732
rect 93823 31690 94209 31709
rect 4343 31039 4729 31058
rect 4343 31016 4409 31039
rect 4495 31016 4577 31039
rect 4663 31016 4729 31039
rect 4343 30976 4352 31016
rect 4392 30976 4409 31016
rect 4495 30976 4516 31016
rect 4556 30976 4577 31016
rect 4663 30976 4680 31016
rect 4720 30976 4729 31016
rect 4343 30953 4409 30976
rect 4495 30953 4577 30976
rect 4663 30953 4729 30976
rect 4343 30934 4729 30953
rect 19463 31039 19849 31058
rect 19463 31016 19529 31039
rect 19615 31016 19697 31039
rect 19783 31016 19849 31039
rect 19463 30976 19472 31016
rect 19512 30976 19529 31016
rect 19615 30976 19636 31016
rect 19676 30976 19697 31016
rect 19783 30976 19800 31016
rect 19840 30976 19849 31016
rect 19463 30953 19529 30976
rect 19615 30953 19697 30976
rect 19783 30953 19849 30976
rect 19463 30934 19849 30953
rect 34583 31039 34969 31058
rect 34583 31016 34649 31039
rect 34735 31016 34817 31039
rect 34903 31016 34969 31039
rect 34583 30976 34592 31016
rect 34632 30976 34649 31016
rect 34735 30976 34756 31016
rect 34796 30976 34817 31016
rect 34903 30976 34920 31016
rect 34960 30976 34969 31016
rect 34583 30953 34649 30976
rect 34735 30953 34817 30976
rect 34903 30953 34969 30976
rect 34583 30934 34969 30953
rect 49703 31039 50089 31058
rect 49703 31016 49769 31039
rect 49855 31016 49937 31039
rect 50023 31016 50089 31039
rect 49703 30976 49712 31016
rect 49752 30976 49769 31016
rect 49855 30976 49876 31016
rect 49916 30976 49937 31016
rect 50023 30976 50040 31016
rect 50080 30976 50089 31016
rect 49703 30953 49769 30976
rect 49855 30953 49937 30976
rect 50023 30953 50089 30976
rect 49703 30934 50089 30953
rect 64823 31039 65209 31058
rect 64823 31016 64889 31039
rect 64975 31016 65057 31039
rect 65143 31016 65209 31039
rect 64823 30976 64832 31016
rect 64872 30976 64889 31016
rect 64975 30976 64996 31016
rect 65036 30976 65057 31016
rect 65143 30976 65160 31016
rect 65200 30976 65209 31016
rect 64823 30953 64889 30976
rect 64975 30953 65057 30976
rect 65143 30953 65209 30976
rect 64823 30934 65209 30953
rect 79943 31039 80329 31058
rect 79943 31016 80009 31039
rect 80095 31016 80177 31039
rect 80263 31016 80329 31039
rect 79943 30976 79952 31016
rect 79992 30976 80009 31016
rect 80095 30976 80116 31016
rect 80156 30976 80177 31016
rect 80263 30976 80280 31016
rect 80320 30976 80329 31016
rect 79943 30953 80009 30976
rect 80095 30953 80177 30976
rect 80263 30953 80329 30976
rect 79943 30934 80329 30953
rect 95063 31039 95449 31058
rect 95063 31016 95129 31039
rect 95215 31016 95297 31039
rect 95383 31016 95449 31039
rect 95063 30976 95072 31016
rect 95112 30976 95129 31016
rect 95215 30976 95236 31016
rect 95276 30976 95297 31016
rect 95383 30976 95400 31016
rect 95440 30976 95449 31016
rect 95063 30953 95129 30976
rect 95215 30953 95297 30976
rect 95383 30953 95449 30976
rect 95063 30934 95449 30953
rect 3103 30283 3489 30302
rect 3103 30260 3169 30283
rect 3255 30260 3337 30283
rect 3423 30260 3489 30283
rect 3103 30220 3112 30260
rect 3152 30220 3169 30260
rect 3255 30220 3276 30260
rect 3316 30220 3337 30260
rect 3423 30220 3440 30260
rect 3480 30220 3489 30260
rect 3103 30197 3169 30220
rect 3255 30197 3337 30220
rect 3423 30197 3489 30220
rect 3103 30178 3489 30197
rect 18223 30283 18609 30302
rect 18223 30260 18289 30283
rect 18375 30260 18457 30283
rect 18543 30260 18609 30283
rect 18223 30220 18232 30260
rect 18272 30220 18289 30260
rect 18375 30220 18396 30260
rect 18436 30220 18457 30260
rect 18543 30220 18560 30260
rect 18600 30220 18609 30260
rect 18223 30197 18289 30220
rect 18375 30197 18457 30220
rect 18543 30197 18609 30220
rect 18223 30178 18609 30197
rect 33343 30283 33729 30302
rect 33343 30260 33409 30283
rect 33495 30260 33577 30283
rect 33663 30260 33729 30283
rect 33343 30220 33352 30260
rect 33392 30220 33409 30260
rect 33495 30220 33516 30260
rect 33556 30220 33577 30260
rect 33663 30220 33680 30260
rect 33720 30220 33729 30260
rect 33343 30197 33409 30220
rect 33495 30197 33577 30220
rect 33663 30197 33729 30220
rect 33343 30178 33729 30197
rect 48463 30283 48849 30302
rect 48463 30260 48529 30283
rect 48615 30260 48697 30283
rect 48783 30260 48849 30283
rect 48463 30220 48472 30260
rect 48512 30220 48529 30260
rect 48615 30220 48636 30260
rect 48676 30220 48697 30260
rect 48783 30220 48800 30260
rect 48840 30220 48849 30260
rect 48463 30197 48529 30220
rect 48615 30197 48697 30220
rect 48783 30197 48849 30220
rect 48463 30178 48849 30197
rect 63583 30283 63969 30302
rect 63583 30260 63649 30283
rect 63735 30260 63817 30283
rect 63903 30260 63969 30283
rect 63583 30220 63592 30260
rect 63632 30220 63649 30260
rect 63735 30220 63756 30260
rect 63796 30220 63817 30260
rect 63903 30220 63920 30260
rect 63960 30220 63969 30260
rect 63583 30197 63649 30220
rect 63735 30197 63817 30220
rect 63903 30197 63969 30220
rect 63583 30178 63969 30197
rect 78703 30283 79089 30302
rect 78703 30260 78769 30283
rect 78855 30260 78937 30283
rect 79023 30260 79089 30283
rect 78703 30220 78712 30260
rect 78752 30220 78769 30260
rect 78855 30220 78876 30260
rect 78916 30220 78937 30260
rect 79023 30220 79040 30260
rect 79080 30220 79089 30260
rect 78703 30197 78769 30220
rect 78855 30197 78937 30220
rect 79023 30197 79089 30220
rect 78703 30178 79089 30197
rect 93823 30283 94209 30302
rect 93823 30260 93889 30283
rect 93975 30260 94057 30283
rect 94143 30260 94209 30283
rect 93823 30220 93832 30260
rect 93872 30220 93889 30260
rect 93975 30220 93996 30260
rect 94036 30220 94057 30260
rect 94143 30220 94160 30260
rect 94200 30220 94209 30260
rect 93823 30197 93889 30220
rect 93975 30197 94057 30220
rect 94143 30197 94209 30220
rect 93823 30178 94209 30197
rect 4343 29527 4729 29546
rect 4343 29504 4409 29527
rect 4495 29504 4577 29527
rect 4663 29504 4729 29527
rect 4343 29464 4352 29504
rect 4392 29464 4409 29504
rect 4495 29464 4516 29504
rect 4556 29464 4577 29504
rect 4663 29464 4680 29504
rect 4720 29464 4729 29504
rect 4343 29441 4409 29464
rect 4495 29441 4577 29464
rect 4663 29441 4729 29464
rect 4343 29422 4729 29441
rect 19463 29527 19849 29546
rect 19463 29504 19529 29527
rect 19615 29504 19697 29527
rect 19783 29504 19849 29527
rect 19463 29464 19472 29504
rect 19512 29464 19529 29504
rect 19615 29464 19636 29504
rect 19676 29464 19697 29504
rect 19783 29464 19800 29504
rect 19840 29464 19849 29504
rect 19463 29441 19529 29464
rect 19615 29441 19697 29464
rect 19783 29441 19849 29464
rect 19463 29422 19849 29441
rect 34583 29527 34969 29546
rect 34583 29504 34649 29527
rect 34735 29504 34817 29527
rect 34903 29504 34969 29527
rect 34583 29464 34592 29504
rect 34632 29464 34649 29504
rect 34735 29464 34756 29504
rect 34796 29464 34817 29504
rect 34903 29464 34920 29504
rect 34960 29464 34969 29504
rect 34583 29441 34649 29464
rect 34735 29441 34817 29464
rect 34903 29441 34969 29464
rect 34583 29422 34969 29441
rect 49703 29527 50089 29546
rect 49703 29504 49769 29527
rect 49855 29504 49937 29527
rect 50023 29504 50089 29527
rect 49703 29464 49712 29504
rect 49752 29464 49769 29504
rect 49855 29464 49876 29504
rect 49916 29464 49937 29504
rect 50023 29464 50040 29504
rect 50080 29464 50089 29504
rect 49703 29441 49769 29464
rect 49855 29441 49937 29464
rect 50023 29441 50089 29464
rect 49703 29422 50089 29441
rect 64823 29527 65209 29546
rect 64823 29504 64889 29527
rect 64975 29504 65057 29527
rect 65143 29504 65209 29527
rect 64823 29464 64832 29504
rect 64872 29464 64889 29504
rect 64975 29464 64996 29504
rect 65036 29464 65057 29504
rect 65143 29464 65160 29504
rect 65200 29464 65209 29504
rect 64823 29441 64889 29464
rect 64975 29441 65057 29464
rect 65143 29441 65209 29464
rect 64823 29422 65209 29441
rect 79943 29527 80329 29546
rect 79943 29504 80009 29527
rect 80095 29504 80177 29527
rect 80263 29504 80329 29527
rect 79943 29464 79952 29504
rect 79992 29464 80009 29504
rect 80095 29464 80116 29504
rect 80156 29464 80177 29504
rect 80263 29464 80280 29504
rect 80320 29464 80329 29504
rect 79943 29441 80009 29464
rect 80095 29441 80177 29464
rect 80263 29441 80329 29464
rect 79943 29422 80329 29441
rect 95063 29527 95449 29546
rect 95063 29504 95129 29527
rect 95215 29504 95297 29527
rect 95383 29504 95449 29527
rect 95063 29464 95072 29504
rect 95112 29464 95129 29504
rect 95215 29464 95236 29504
rect 95276 29464 95297 29504
rect 95383 29464 95400 29504
rect 95440 29464 95449 29504
rect 95063 29441 95129 29464
rect 95215 29441 95297 29464
rect 95383 29441 95449 29464
rect 95063 29422 95449 29441
rect 3103 28771 3489 28790
rect 3103 28748 3169 28771
rect 3255 28748 3337 28771
rect 3423 28748 3489 28771
rect 3103 28708 3112 28748
rect 3152 28708 3169 28748
rect 3255 28708 3276 28748
rect 3316 28708 3337 28748
rect 3423 28708 3440 28748
rect 3480 28708 3489 28748
rect 3103 28685 3169 28708
rect 3255 28685 3337 28708
rect 3423 28685 3489 28708
rect 3103 28666 3489 28685
rect 18223 28771 18609 28790
rect 18223 28748 18289 28771
rect 18375 28748 18457 28771
rect 18543 28748 18609 28771
rect 18223 28708 18232 28748
rect 18272 28708 18289 28748
rect 18375 28708 18396 28748
rect 18436 28708 18457 28748
rect 18543 28708 18560 28748
rect 18600 28708 18609 28748
rect 18223 28685 18289 28708
rect 18375 28685 18457 28708
rect 18543 28685 18609 28708
rect 18223 28666 18609 28685
rect 33343 28771 33729 28790
rect 33343 28748 33409 28771
rect 33495 28748 33577 28771
rect 33663 28748 33729 28771
rect 33343 28708 33352 28748
rect 33392 28708 33409 28748
rect 33495 28708 33516 28748
rect 33556 28708 33577 28748
rect 33663 28708 33680 28748
rect 33720 28708 33729 28748
rect 33343 28685 33409 28708
rect 33495 28685 33577 28708
rect 33663 28685 33729 28708
rect 33343 28666 33729 28685
rect 48463 28771 48849 28790
rect 48463 28748 48529 28771
rect 48615 28748 48697 28771
rect 48783 28748 48849 28771
rect 48463 28708 48472 28748
rect 48512 28708 48529 28748
rect 48615 28708 48636 28748
rect 48676 28708 48697 28748
rect 48783 28708 48800 28748
rect 48840 28708 48849 28748
rect 48463 28685 48529 28708
rect 48615 28685 48697 28708
rect 48783 28685 48849 28708
rect 48463 28666 48849 28685
rect 63583 28771 63969 28790
rect 63583 28748 63649 28771
rect 63735 28748 63817 28771
rect 63903 28748 63969 28771
rect 63583 28708 63592 28748
rect 63632 28708 63649 28748
rect 63735 28708 63756 28748
rect 63796 28708 63817 28748
rect 63903 28708 63920 28748
rect 63960 28708 63969 28748
rect 63583 28685 63649 28708
rect 63735 28685 63817 28708
rect 63903 28685 63969 28708
rect 63583 28666 63969 28685
rect 78703 28771 79089 28790
rect 78703 28748 78769 28771
rect 78855 28748 78937 28771
rect 79023 28748 79089 28771
rect 78703 28708 78712 28748
rect 78752 28708 78769 28748
rect 78855 28708 78876 28748
rect 78916 28708 78937 28748
rect 79023 28708 79040 28748
rect 79080 28708 79089 28748
rect 78703 28685 78769 28708
rect 78855 28685 78937 28708
rect 79023 28685 79089 28708
rect 78703 28666 79089 28685
rect 93823 28771 94209 28790
rect 93823 28748 93889 28771
rect 93975 28748 94057 28771
rect 94143 28748 94209 28771
rect 93823 28708 93832 28748
rect 93872 28708 93889 28748
rect 93975 28708 93996 28748
rect 94036 28708 94057 28748
rect 94143 28708 94160 28748
rect 94200 28708 94209 28748
rect 93823 28685 93889 28708
rect 93975 28685 94057 28708
rect 94143 28685 94209 28708
rect 93823 28666 94209 28685
rect 4343 28015 4729 28034
rect 4343 27992 4409 28015
rect 4495 27992 4577 28015
rect 4663 27992 4729 28015
rect 4343 27952 4352 27992
rect 4392 27952 4409 27992
rect 4495 27952 4516 27992
rect 4556 27952 4577 27992
rect 4663 27952 4680 27992
rect 4720 27952 4729 27992
rect 4343 27929 4409 27952
rect 4495 27929 4577 27952
rect 4663 27929 4729 27952
rect 4343 27910 4729 27929
rect 19463 28015 19849 28034
rect 19463 27992 19529 28015
rect 19615 27992 19697 28015
rect 19783 27992 19849 28015
rect 19463 27952 19472 27992
rect 19512 27952 19529 27992
rect 19615 27952 19636 27992
rect 19676 27952 19697 27992
rect 19783 27952 19800 27992
rect 19840 27952 19849 27992
rect 19463 27929 19529 27952
rect 19615 27929 19697 27952
rect 19783 27929 19849 27952
rect 19463 27910 19849 27929
rect 34583 28015 34969 28034
rect 34583 27992 34649 28015
rect 34735 27992 34817 28015
rect 34903 27992 34969 28015
rect 34583 27952 34592 27992
rect 34632 27952 34649 27992
rect 34735 27952 34756 27992
rect 34796 27952 34817 27992
rect 34903 27952 34920 27992
rect 34960 27952 34969 27992
rect 34583 27929 34649 27952
rect 34735 27929 34817 27952
rect 34903 27929 34969 27952
rect 34583 27910 34969 27929
rect 49703 28015 50089 28034
rect 49703 27992 49769 28015
rect 49855 27992 49937 28015
rect 50023 27992 50089 28015
rect 49703 27952 49712 27992
rect 49752 27952 49769 27992
rect 49855 27952 49876 27992
rect 49916 27952 49937 27992
rect 50023 27952 50040 27992
rect 50080 27952 50089 27992
rect 49703 27929 49769 27952
rect 49855 27929 49937 27952
rect 50023 27929 50089 27952
rect 49703 27910 50089 27929
rect 64823 28015 65209 28034
rect 64823 27992 64889 28015
rect 64975 27992 65057 28015
rect 65143 27992 65209 28015
rect 64823 27952 64832 27992
rect 64872 27952 64889 27992
rect 64975 27952 64996 27992
rect 65036 27952 65057 27992
rect 65143 27952 65160 27992
rect 65200 27952 65209 27992
rect 64823 27929 64889 27952
rect 64975 27929 65057 27952
rect 65143 27929 65209 27952
rect 64823 27910 65209 27929
rect 79943 28015 80329 28034
rect 79943 27992 80009 28015
rect 80095 27992 80177 28015
rect 80263 27992 80329 28015
rect 79943 27952 79952 27992
rect 79992 27952 80009 27992
rect 80095 27952 80116 27992
rect 80156 27952 80177 27992
rect 80263 27952 80280 27992
rect 80320 27952 80329 27992
rect 79943 27929 80009 27952
rect 80095 27929 80177 27952
rect 80263 27929 80329 27952
rect 79943 27910 80329 27929
rect 95063 28015 95449 28034
rect 95063 27992 95129 28015
rect 95215 27992 95297 28015
rect 95383 27992 95449 28015
rect 95063 27952 95072 27992
rect 95112 27952 95129 27992
rect 95215 27952 95236 27992
rect 95276 27952 95297 27992
rect 95383 27952 95400 27992
rect 95440 27952 95449 27992
rect 95063 27929 95129 27952
rect 95215 27929 95297 27952
rect 95383 27929 95449 27952
rect 95063 27910 95449 27929
rect 3103 27259 3489 27278
rect 3103 27236 3169 27259
rect 3255 27236 3337 27259
rect 3423 27236 3489 27259
rect 3103 27196 3112 27236
rect 3152 27196 3169 27236
rect 3255 27196 3276 27236
rect 3316 27196 3337 27236
rect 3423 27196 3440 27236
rect 3480 27196 3489 27236
rect 3103 27173 3169 27196
rect 3255 27173 3337 27196
rect 3423 27173 3489 27196
rect 3103 27154 3489 27173
rect 18223 27259 18609 27278
rect 18223 27236 18289 27259
rect 18375 27236 18457 27259
rect 18543 27236 18609 27259
rect 18223 27196 18232 27236
rect 18272 27196 18289 27236
rect 18375 27196 18396 27236
rect 18436 27196 18457 27236
rect 18543 27196 18560 27236
rect 18600 27196 18609 27236
rect 18223 27173 18289 27196
rect 18375 27173 18457 27196
rect 18543 27173 18609 27196
rect 18223 27154 18609 27173
rect 33343 27259 33729 27278
rect 33343 27236 33409 27259
rect 33495 27236 33577 27259
rect 33663 27236 33729 27259
rect 33343 27196 33352 27236
rect 33392 27196 33409 27236
rect 33495 27196 33516 27236
rect 33556 27196 33577 27236
rect 33663 27196 33680 27236
rect 33720 27196 33729 27236
rect 33343 27173 33409 27196
rect 33495 27173 33577 27196
rect 33663 27173 33729 27196
rect 33343 27154 33729 27173
rect 48463 27259 48849 27278
rect 48463 27236 48529 27259
rect 48615 27236 48697 27259
rect 48783 27236 48849 27259
rect 48463 27196 48472 27236
rect 48512 27196 48529 27236
rect 48615 27196 48636 27236
rect 48676 27196 48697 27236
rect 48783 27196 48800 27236
rect 48840 27196 48849 27236
rect 48463 27173 48529 27196
rect 48615 27173 48697 27196
rect 48783 27173 48849 27196
rect 48463 27154 48849 27173
rect 63583 27259 63969 27278
rect 63583 27236 63649 27259
rect 63735 27236 63817 27259
rect 63903 27236 63969 27259
rect 63583 27196 63592 27236
rect 63632 27196 63649 27236
rect 63735 27196 63756 27236
rect 63796 27196 63817 27236
rect 63903 27196 63920 27236
rect 63960 27196 63969 27236
rect 63583 27173 63649 27196
rect 63735 27173 63817 27196
rect 63903 27173 63969 27196
rect 63583 27154 63969 27173
rect 78703 27259 79089 27278
rect 78703 27236 78769 27259
rect 78855 27236 78937 27259
rect 79023 27236 79089 27259
rect 78703 27196 78712 27236
rect 78752 27196 78769 27236
rect 78855 27196 78876 27236
rect 78916 27196 78937 27236
rect 79023 27196 79040 27236
rect 79080 27196 79089 27236
rect 78703 27173 78769 27196
rect 78855 27173 78937 27196
rect 79023 27173 79089 27196
rect 78703 27154 79089 27173
rect 93823 27259 94209 27278
rect 93823 27236 93889 27259
rect 93975 27236 94057 27259
rect 94143 27236 94209 27259
rect 93823 27196 93832 27236
rect 93872 27196 93889 27236
rect 93975 27196 93996 27236
rect 94036 27196 94057 27236
rect 94143 27196 94160 27236
rect 94200 27196 94209 27236
rect 93823 27173 93889 27196
rect 93975 27173 94057 27196
rect 94143 27173 94209 27196
rect 93823 27154 94209 27173
rect 4343 26503 4729 26522
rect 4343 26480 4409 26503
rect 4495 26480 4577 26503
rect 4663 26480 4729 26503
rect 4343 26440 4352 26480
rect 4392 26440 4409 26480
rect 4495 26440 4516 26480
rect 4556 26440 4577 26480
rect 4663 26440 4680 26480
rect 4720 26440 4729 26480
rect 4343 26417 4409 26440
rect 4495 26417 4577 26440
rect 4663 26417 4729 26440
rect 4343 26398 4729 26417
rect 19463 26503 19849 26522
rect 19463 26480 19529 26503
rect 19615 26480 19697 26503
rect 19783 26480 19849 26503
rect 19463 26440 19472 26480
rect 19512 26440 19529 26480
rect 19615 26440 19636 26480
rect 19676 26440 19697 26480
rect 19783 26440 19800 26480
rect 19840 26440 19849 26480
rect 19463 26417 19529 26440
rect 19615 26417 19697 26440
rect 19783 26417 19849 26440
rect 19463 26398 19849 26417
rect 34583 26503 34969 26522
rect 34583 26480 34649 26503
rect 34735 26480 34817 26503
rect 34903 26480 34969 26503
rect 34583 26440 34592 26480
rect 34632 26440 34649 26480
rect 34735 26440 34756 26480
rect 34796 26440 34817 26480
rect 34903 26440 34920 26480
rect 34960 26440 34969 26480
rect 34583 26417 34649 26440
rect 34735 26417 34817 26440
rect 34903 26417 34969 26440
rect 34583 26398 34969 26417
rect 49703 26503 50089 26522
rect 49703 26480 49769 26503
rect 49855 26480 49937 26503
rect 50023 26480 50089 26503
rect 49703 26440 49712 26480
rect 49752 26440 49769 26480
rect 49855 26440 49876 26480
rect 49916 26440 49937 26480
rect 50023 26440 50040 26480
rect 50080 26440 50089 26480
rect 49703 26417 49769 26440
rect 49855 26417 49937 26440
rect 50023 26417 50089 26440
rect 49703 26398 50089 26417
rect 64823 26503 65209 26522
rect 64823 26480 64889 26503
rect 64975 26480 65057 26503
rect 65143 26480 65209 26503
rect 64823 26440 64832 26480
rect 64872 26440 64889 26480
rect 64975 26440 64996 26480
rect 65036 26440 65057 26480
rect 65143 26440 65160 26480
rect 65200 26440 65209 26480
rect 64823 26417 64889 26440
rect 64975 26417 65057 26440
rect 65143 26417 65209 26440
rect 64823 26398 65209 26417
rect 79943 26503 80329 26522
rect 79943 26480 80009 26503
rect 80095 26480 80177 26503
rect 80263 26480 80329 26503
rect 79943 26440 79952 26480
rect 79992 26440 80009 26480
rect 80095 26440 80116 26480
rect 80156 26440 80177 26480
rect 80263 26440 80280 26480
rect 80320 26440 80329 26480
rect 79943 26417 80009 26440
rect 80095 26417 80177 26440
rect 80263 26417 80329 26440
rect 79943 26398 80329 26417
rect 95063 26503 95449 26522
rect 95063 26480 95129 26503
rect 95215 26480 95297 26503
rect 95383 26480 95449 26503
rect 95063 26440 95072 26480
rect 95112 26440 95129 26480
rect 95215 26440 95236 26480
rect 95276 26440 95297 26480
rect 95383 26440 95400 26480
rect 95440 26440 95449 26480
rect 95063 26417 95129 26440
rect 95215 26417 95297 26440
rect 95383 26417 95449 26440
rect 95063 26398 95449 26417
rect 3103 25747 3489 25766
rect 3103 25724 3169 25747
rect 3255 25724 3337 25747
rect 3423 25724 3489 25747
rect 3103 25684 3112 25724
rect 3152 25684 3169 25724
rect 3255 25684 3276 25724
rect 3316 25684 3337 25724
rect 3423 25684 3440 25724
rect 3480 25684 3489 25724
rect 3103 25661 3169 25684
rect 3255 25661 3337 25684
rect 3423 25661 3489 25684
rect 3103 25642 3489 25661
rect 18223 25747 18609 25766
rect 18223 25724 18289 25747
rect 18375 25724 18457 25747
rect 18543 25724 18609 25747
rect 18223 25684 18232 25724
rect 18272 25684 18289 25724
rect 18375 25684 18396 25724
rect 18436 25684 18457 25724
rect 18543 25684 18560 25724
rect 18600 25684 18609 25724
rect 18223 25661 18289 25684
rect 18375 25661 18457 25684
rect 18543 25661 18609 25684
rect 18223 25642 18609 25661
rect 33343 25747 33729 25766
rect 33343 25724 33409 25747
rect 33495 25724 33577 25747
rect 33663 25724 33729 25747
rect 33343 25684 33352 25724
rect 33392 25684 33409 25724
rect 33495 25684 33516 25724
rect 33556 25684 33577 25724
rect 33663 25684 33680 25724
rect 33720 25684 33729 25724
rect 33343 25661 33409 25684
rect 33495 25661 33577 25684
rect 33663 25661 33729 25684
rect 33343 25642 33729 25661
rect 48463 25747 48849 25766
rect 48463 25724 48529 25747
rect 48615 25724 48697 25747
rect 48783 25724 48849 25747
rect 48463 25684 48472 25724
rect 48512 25684 48529 25724
rect 48615 25684 48636 25724
rect 48676 25684 48697 25724
rect 48783 25684 48800 25724
rect 48840 25684 48849 25724
rect 48463 25661 48529 25684
rect 48615 25661 48697 25684
rect 48783 25661 48849 25684
rect 48463 25642 48849 25661
rect 63583 25747 63969 25766
rect 63583 25724 63649 25747
rect 63735 25724 63817 25747
rect 63903 25724 63969 25747
rect 63583 25684 63592 25724
rect 63632 25684 63649 25724
rect 63735 25684 63756 25724
rect 63796 25684 63817 25724
rect 63903 25684 63920 25724
rect 63960 25684 63969 25724
rect 63583 25661 63649 25684
rect 63735 25661 63817 25684
rect 63903 25661 63969 25684
rect 63583 25642 63969 25661
rect 78703 25747 79089 25766
rect 78703 25724 78769 25747
rect 78855 25724 78937 25747
rect 79023 25724 79089 25747
rect 78703 25684 78712 25724
rect 78752 25684 78769 25724
rect 78855 25684 78876 25724
rect 78916 25684 78937 25724
rect 79023 25684 79040 25724
rect 79080 25684 79089 25724
rect 78703 25661 78769 25684
rect 78855 25661 78937 25684
rect 79023 25661 79089 25684
rect 78703 25642 79089 25661
rect 93823 25747 94209 25766
rect 93823 25724 93889 25747
rect 93975 25724 94057 25747
rect 94143 25724 94209 25747
rect 93823 25684 93832 25724
rect 93872 25684 93889 25724
rect 93975 25684 93996 25724
rect 94036 25684 94057 25724
rect 94143 25684 94160 25724
rect 94200 25684 94209 25724
rect 93823 25661 93889 25684
rect 93975 25661 94057 25684
rect 94143 25661 94209 25684
rect 93823 25642 94209 25661
rect 4343 24991 4729 25010
rect 4343 24968 4409 24991
rect 4495 24968 4577 24991
rect 4663 24968 4729 24991
rect 4343 24928 4352 24968
rect 4392 24928 4409 24968
rect 4495 24928 4516 24968
rect 4556 24928 4577 24968
rect 4663 24928 4680 24968
rect 4720 24928 4729 24968
rect 4343 24905 4409 24928
rect 4495 24905 4577 24928
rect 4663 24905 4729 24928
rect 4343 24886 4729 24905
rect 19463 24991 19849 25010
rect 19463 24968 19529 24991
rect 19615 24968 19697 24991
rect 19783 24968 19849 24991
rect 19463 24928 19472 24968
rect 19512 24928 19529 24968
rect 19615 24928 19636 24968
rect 19676 24928 19697 24968
rect 19783 24928 19800 24968
rect 19840 24928 19849 24968
rect 19463 24905 19529 24928
rect 19615 24905 19697 24928
rect 19783 24905 19849 24928
rect 19463 24886 19849 24905
rect 34583 24991 34969 25010
rect 34583 24968 34649 24991
rect 34735 24968 34817 24991
rect 34903 24968 34969 24991
rect 34583 24928 34592 24968
rect 34632 24928 34649 24968
rect 34735 24928 34756 24968
rect 34796 24928 34817 24968
rect 34903 24928 34920 24968
rect 34960 24928 34969 24968
rect 34583 24905 34649 24928
rect 34735 24905 34817 24928
rect 34903 24905 34969 24928
rect 34583 24886 34969 24905
rect 49703 24991 50089 25010
rect 49703 24968 49769 24991
rect 49855 24968 49937 24991
rect 50023 24968 50089 24991
rect 49703 24928 49712 24968
rect 49752 24928 49769 24968
rect 49855 24928 49876 24968
rect 49916 24928 49937 24968
rect 50023 24928 50040 24968
rect 50080 24928 50089 24968
rect 49703 24905 49769 24928
rect 49855 24905 49937 24928
rect 50023 24905 50089 24928
rect 49703 24886 50089 24905
rect 64823 24991 65209 25010
rect 64823 24968 64889 24991
rect 64975 24968 65057 24991
rect 65143 24968 65209 24991
rect 64823 24928 64832 24968
rect 64872 24928 64889 24968
rect 64975 24928 64996 24968
rect 65036 24928 65057 24968
rect 65143 24928 65160 24968
rect 65200 24928 65209 24968
rect 64823 24905 64889 24928
rect 64975 24905 65057 24928
rect 65143 24905 65209 24928
rect 64823 24886 65209 24905
rect 79943 24991 80329 25010
rect 79943 24968 80009 24991
rect 80095 24968 80177 24991
rect 80263 24968 80329 24991
rect 79943 24928 79952 24968
rect 79992 24928 80009 24968
rect 80095 24928 80116 24968
rect 80156 24928 80177 24968
rect 80263 24928 80280 24968
rect 80320 24928 80329 24968
rect 79943 24905 80009 24928
rect 80095 24905 80177 24928
rect 80263 24905 80329 24928
rect 79943 24886 80329 24905
rect 95063 24991 95449 25010
rect 95063 24968 95129 24991
rect 95215 24968 95297 24991
rect 95383 24968 95449 24991
rect 95063 24928 95072 24968
rect 95112 24928 95129 24968
rect 95215 24928 95236 24968
rect 95276 24928 95297 24968
rect 95383 24928 95400 24968
rect 95440 24928 95449 24968
rect 95063 24905 95129 24928
rect 95215 24905 95297 24928
rect 95383 24905 95449 24928
rect 95063 24886 95449 24905
rect 3103 24235 3489 24254
rect 3103 24212 3169 24235
rect 3255 24212 3337 24235
rect 3423 24212 3489 24235
rect 3103 24172 3112 24212
rect 3152 24172 3169 24212
rect 3255 24172 3276 24212
rect 3316 24172 3337 24212
rect 3423 24172 3440 24212
rect 3480 24172 3489 24212
rect 3103 24149 3169 24172
rect 3255 24149 3337 24172
rect 3423 24149 3489 24172
rect 3103 24130 3489 24149
rect 18223 24235 18609 24254
rect 18223 24212 18289 24235
rect 18375 24212 18457 24235
rect 18543 24212 18609 24235
rect 18223 24172 18232 24212
rect 18272 24172 18289 24212
rect 18375 24172 18396 24212
rect 18436 24172 18457 24212
rect 18543 24172 18560 24212
rect 18600 24172 18609 24212
rect 18223 24149 18289 24172
rect 18375 24149 18457 24172
rect 18543 24149 18609 24172
rect 18223 24130 18609 24149
rect 33343 24235 33729 24254
rect 33343 24212 33409 24235
rect 33495 24212 33577 24235
rect 33663 24212 33729 24235
rect 33343 24172 33352 24212
rect 33392 24172 33409 24212
rect 33495 24172 33516 24212
rect 33556 24172 33577 24212
rect 33663 24172 33680 24212
rect 33720 24172 33729 24212
rect 33343 24149 33409 24172
rect 33495 24149 33577 24172
rect 33663 24149 33729 24172
rect 33343 24130 33729 24149
rect 48463 24235 48849 24254
rect 48463 24212 48529 24235
rect 48615 24212 48697 24235
rect 48783 24212 48849 24235
rect 48463 24172 48472 24212
rect 48512 24172 48529 24212
rect 48615 24172 48636 24212
rect 48676 24172 48697 24212
rect 48783 24172 48800 24212
rect 48840 24172 48849 24212
rect 48463 24149 48529 24172
rect 48615 24149 48697 24172
rect 48783 24149 48849 24172
rect 48463 24130 48849 24149
rect 63583 24235 63969 24254
rect 63583 24212 63649 24235
rect 63735 24212 63817 24235
rect 63903 24212 63969 24235
rect 63583 24172 63592 24212
rect 63632 24172 63649 24212
rect 63735 24172 63756 24212
rect 63796 24172 63817 24212
rect 63903 24172 63920 24212
rect 63960 24172 63969 24212
rect 63583 24149 63649 24172
rect 63735 24149 63817 24172
rect 63903 24149 63969 24172
rect 63583 24130 63969 24149
rect 78703 24235 79089 24254
rect 78703 24212 78769 24235
rect 78855 24212 78937 24235
rect 79023 24212 79089 24235
rect 78703 24172 78712 24212
rect 78752 24172 78769 24212
rect 78855 24172 78876 24212
rect 78916 24172 78937 24212
rect 79023 24172 79040 24212
rect 79080 24172 79089 24212
rect 78703 24149 78769 24172
rect 78855 24149 78937 24172
rect 79023 24149 79089 24172
rect 78703 24130 79089 24149
rect 93823 24235 94209 24254
rect 93823 24212 93889 24235
rect 93975 24212 94057 24235
rect 94143 24212 94209 24235
rect 93823 24172 93832 24212
rect 93872 24172 93889 24212
rect 93975 24172 93996 24212
rect 94036 24172 94057 24212
rect 94143 24172 94160 24212
rect 94200 24172 94209 24212
rect 93823 24149 93889 24172
rect 93975 24149 94057 24172
rect 94143 24149 94209 24172
rect 93823 24130 94209 24149
rect 4343 23479 4729 23498
rect 4343 23456 4409 23479
rect 4495 23456 4577 23479
rect 4663 23456 4729 23479
rect 4343 23416 4352 23456
rect 4392 23416 4409 23456
rect 4495 23416 4516 23456
rect 4556 23416 4577 23456
rect 4663 23416 4680 23456
rect 4720 23416 4729 23456
rect 4343 23393 4409 23416
rect 4495 23393 4577 23416
rect 4663 23393 4729 23416
rect 4343 23374 4729 23393
rect 19463 23479 19849 23498
rect 19463 23456 19529 23479
rect 19615 23456 19697 23479
rect 19783 23456 19849 23479
rect 19463 23416 19472 23456
rect 19512 23416 19529 23456
rect 19615 23416 19636 23456
rect 19676 23416 19697 23456
rect 19783 23416 19800 23456
rect 19840 23416 19849 23456
rect 19463 23393 19529 23416
rect 19615 23393 19697 23416
rect 19783 23393 19849 23416
rect 19463 23374 19849 23393
rect 34583 23479 34969 23498
rect 34583 23456 34649 23479
rect 34735 23456 34817 23479
rect 34903 23456 34969 23479
rect 34583 23416 34592 23456
rect 34632 23416 34649 23456
rect 34735 23416 34756 23456
rect 34796 23416 34817 23456
rect 34903 23416 34920 23456
rect 34960 23416 34969 23456
rect 34583 23393 34649 23416
rect 34735 23393 34817 23416
rect 34903 23393 34969 23416
rect 34583 23374 34969 23393
rect 49703 23479 50089 23498
rect 49703 23456 49769 23479
rect 49855 23456 49937 23479
rect 50023 23456 50089 23479
rect 49703 23416 49712 23456
rect 49752 23416 49769 23456
rect 49855 23416 49876 23456
rect 49916 23416 49937 23456
rect 50023 23416 50040 23456
rect 50080 23416 50089 23456
rect 49703 23393 49769 23416
rect 49855 23393 49937 23416
rect 50023 23393 50089 23416
rect 49703 23374 50089 23393
rect 64823 23479 65209 23498
rect 64823 23456 64889 23479
rect 64975 23456 65057 23479
rect 65143 23456 65209 23479
rect 64823 23416 64832 23456
rect 64872 23416 64889 23456
rect 64975 23416 64996 23456
rect 65036 23416 65057 23456
rect 65143 23416 65160 23456
rect 65200 23416 65209 23456
rect 64823 23393 64889 23416
rect 64975 23393 65057 23416
rect 65143 23393 65209 23416
rect 64823 23374 65209 23393
rect 79943 23479 80329 23498
rect 79943 23456 80009 23479
rect 80095 23456 80177 23479
rect 80263 23456 80329 23479
rect 79943 23416 79952 23456
rect 79992 23416 80009 23456
rect 80095 23416 80116 23456
rect 80156 23416 80177 23456
rect 80263 23416 80280 23456
rect 80320 23416 80329 23456
rect 79943 23393 80009 23416
rect 80095 23393 80177 23416
rect 80263 23393 80329 23416
rect 79943 23374 80329 23393
rect 95063 23479 95449 23498
rect 95063 23456 95129 23479
rect 95215 23456 95297 23479
rect 95383 23456 95449 23479
rect 95063 23416 95072 23456
rect 95112 23416 95129 23456
rect 95215 23416 95236 23456
rect 95276 23416 95297 23456
rect 95383 23416 95400 23456
rect 95440 23416 95449 23456
rect 95063 23393 95129 23416
rect 95215 23393 95297 23416
rect 95383 23393 95449 23416
rect 95063 23374 95449 23393
rect 3103 22723 3489 22742
rect 3103 22700 3169 22723
rect 3255 22700 3337 22723
rect 3423 22700 3489 22723
rect 3103 22660 3112 22700
rect 3152 22660 3169 22700
rect 3255 22660 3276 22700
rect 3316 22660 3337 22700
rect 3423 22660 3440 22700
rect 3480 22660 3489 22700
rect 3103 22637 3169 22660
rect 3255 22637 3337 22660
rect 3423 22637 3489 22660
rect 3103 22618 3489 22637
rect 18223 22723 18609 22742
rect 18223 22700 18289 22723
rect 18375 22700 18457 22723
rect 18543 22700 18609 22723
rect 18223 22660 18232 22700
rect 18272 22660 18289 22700
rect 18375 22660 18396 22700
rect 18436 22660 18457 22700
rect 18543 22660 18560 22700
rect 18600 22660 18609 22700
rect 18223 22637 18289 22660
rect 18375 22637 18457 22660
rect 18543 22637 18609 22660
rect 18223 22618 18609 22637
rect 33343 22723 33729 22742
rect 33343 22700 33409 22723
rect 33495 22700 33577 22723
rect 33663 22700 33729 22723
rect 33343 22660 33352 22700
rect 33392 22660 33409 22700
rect 33495 22660 33516 22700
rect 33556 22660 33577 22700
rect 33663 22660 33680 22700
rect 33720 22660 33729 22700
rect 33343 22637 33409 22660
rect 33495 22637 33577 22660
rect 33663 22637 33729 22660
rect 33343 22618 33729 22637
rect 48463 22723 48849 22742
rect 48463 22700 48529 22723
rect 48615 22700 48697 22723
rect 48783 22700 48849 22723
rect 48463 22660 48472 22700
rect 48512 22660 48529 22700
rect 48615 22660 48636 22700
rect 48676 22660 48697 22700
rect 48783 22660 48800 22700
rect 48840 22660 48849 22700
rect 48463 22637 48529 22660
rect 48615 22637 48697 22660
rect 48783 22637 48849 22660
rect 48463 22618 48849 22637
rect 63583 22723 63969 22742
rect 63583 22700 63649 22723
rect 63735 22700 63817 22723
rect 63903 22700 63969 22723
rect 63583 22660 63592 22700
rect 63632 22660 63649 22700
rect 63735 22660 63756 22700
rect 63796 22660 63817 22700
rect 63903 22660 63920 22700
rect 63960 22660 63969 22700
rect 63583 22637 63649 22660
rect 63735 22637 63817 22660
rect 63903 22637 63969 22660
rect 63583 22618 63969 22637
rect 78703 22723 79089 22742
rect 78703 22700 78769 22723
rect 78855 22700 78937 22723
rect 79023 22700 79089 22723
rect 78703 22660 78712 22700
rect 78752 22660 78769 22700
rect 78855 22660 78876 22700
rect 78916 22660 78937 22700
rect 79023 22660 79040 22700
rect 79080 22660 79089 22700
rect 78703 22637 78769 22660
rect 78855 22637 78937 22660
rect 79023 22637 79089 22660
rect 78703 22618 79089 22637
rect 93823 22723 94209 22742
rect 93823 22700 93889 22723
rect 93975 22700 94057 22723
rect 94143 22700 94209 22723
rect 93823 22660 93832 22700
rect 93872 22660 93889 22700
rect 93975 22660 93996 22700
rect 94036 22660 94057 22700
rect 94143 22660 94160 22700
rect 94200 22660 94209 22700
rect 93823 22637 93889 22660
rect 93975 22637 94057 22660
rect 94143 22637 94209 22660
rect 93823 22618 94209 22637
rect 4343 21967 4729 21986
rect 4343 21944 4409 21967
rect 4495 21944 4577 21967
rect 4663 21944 4729 21967
rect 4343 21904 4352 21944
rect 4392 21904 4409 21944
rect 4495 21904 4516 21944
rect 4556 21904 4577 21944
rect 4663 21904 4680 21944
rect 4720 21904 4729 21944
rect 4343 21881 4409 21904
rect 4495 21881 4577 21904
rect 4663 21881 4729 21904
rect 4343 21862 4729 21881
rect 19463 21967 19849 21986
rect 19463 21944 19529 21967
rect 19615 21944 19697 21967
rect 19783 21944 19849 21967
rect 19463 21904 19472 21944
rect 19512 21904 19529 21944
rect 19615 21904 19636 21944
rect 19676 21904 19697 21944
rect 19783 21904 19800 21944
rect 19840 21904 19849 21944
rect 19463 21881 19529 21904
rect 19615 21881 19697 21904
rect 19783 21881 19849 21904
rect 19463 21862 19849 21881
rect 34583 21967 34969 21986
rect 34583 21944 34649 21967
rect 34735 21944 34817 21967
rect 34903 21944 34969 21967
rect 34583 21904 34592 21944
rect 34632 21904 34649 21944
rect 34735 21904 34756 21944
rect 34796 21904 34817 21944
rect 34903 21904 34920 21944
rect 34960 21904 34969 21944
rect 34583 21881 34649 21904
rect 34735 21881 34817 21904
rect 34903 21881 34969 21904
rect 34583 21862 34969 21881
rect 49703 21967 50089 21986
rect 49703 21944 49769 21967
rect 49855 21944 49937 21967
rect 50023 21944 50089 21967
rect 49703 21904 49712 21944
rect 49752 21904 49769 21944
rect 49855 21904 49876 21944
rect 49916 21904 49937 21944
rect 50023 21904 50040 21944
rect 50080 21904 50089 21944
rect 49703 21881 49769 21904
rect 49855 21881 49937 21904
rect 50023 21881 50089 21904
rect 49703 21862 50089 21881
rect 64823 21967 65209 21986
rect 64823 21944 64889 21967
rect 64975 21944 65057 21967
rect 65143 21944 65209 21967
rect 64823 21904 64832 21944
rect 64872 21904 64889 21944
rect 64975 21904 64996 21944
rect 65036 21904 65057 21944
rect 65143 21904 65160 21944
rect 65200 21904 65209 21944
rect 64823 21881 64889 21904
rect 64975 21881 65057 21904
rect 65143 21881 65209 21904
rect 64823 21862 65209 21881
rect 79943 21967 80329 21986
rect 79943 21944 80009 21967
rect 80095 21944 80177 21967
rect 80263 21944 80329 21967
rect 79943 21904 79952 21944
rect 79992 21904 80009 21944
rect 80095 21904 80116 21944
rect 80156 21904 80177 21944
rect 80263 21904 80280 21944
rect 80320 21904 80329 21944
rect 79943 21881 80009 21904
rect 80095 21881 80177 21904
rect 80263 21881 80329 21904
rect 79943 21862 80329 21881
rect 95063 21967 95449 21986
rect 95063 21944 95129 21967
rect 95215 21944 95297 21967
rect 95383 21944 95449 21967
rect 95063 21904 95072 21944
rect 95112 21904 95129 21944
rect 95215 21904 95236 21944
rect 95276 21904 95297 21944
rect 95383 21904 95400 21944
rect 95440 21904 95449 21944
rect 95063 21881 95129 21904
rect 95215 21881 95297 21904
rect 95383 21881 95449 21904
rect 95063 21862 95449 21881
rect 3103 21211 3489 21230
rect 3103 21188 3169 21211
rect 3255 21188 3337 21211
rect 3423 21188 3489 21211
rect 3103 21148 3112 21188
rect 3152 21148 3169 21188
rect 3255 21148 3276 21188
rect 3316 21148 3337 21188
rect 3423 21148 3440 21188
rect 3480 21148 3489 21188
rect 3103 21125 3169 21148
rect 3255 21125 3337 21148
rect 3423 21125 3489 21148
rect 3103 21106 3489 21125
rect 18223 21211 18609 21230
rect 18223 21188 18289 21211
rect 18375 21188 18457 21211
rect 18543 21188 18609 21211
rect 18223 21148 18232 21188
rect 18272 21148 18289 21188
rect 18375 21148 18396 21188
rect 18436 21148 18457 21188
rect 18543 21148 18560 21188
rect 18600 21148 18609 21188
rect 18223 21125 18289 21148
rect 18375 21125 18457 21148
rect 18543 21125 18609 21148
rect 18223 21106 18609 21125
rect 33343 21211 33729 21230
rect 33343 21188 33409 21211
rect 33495 21188 33577 21211
rect 33663 21188 33729 21211
rect 33343 21148 33352 21188
rect 33392 21148 33409 21188
rect 33495 21148 33516 21188
rect 33556 21148 33577 21188
rect 33663 21148 33680 21188
rect 33720 21148 33729 21188
rect 33343 21125 33409 21148
rect 33495 21125 33577 21148
rect 33663 21125 33729 21148
rect 33343 21106 33729 21125
rect 48463 21211 48849 21230
rect 48463 21188 48529 21211
rect 48615 21188 48697 21211
rect 48783 21188 48849 21211
rect 48463 21148 48472 21188
rect 48512 21148 48529 21188
rect 48615 21148 48636 21188
rect 48676 21148 48697 21188
rect 48783 21148 48800 21188
rect 48840 21148 48849 21188
rect 48463 21125 48529 21148
rect 48615 21125 48697 21148
rect 48783 21125 48849 21148
rect 48463 21106 48849 21125
rect 63583 21211 63969 21230
rect 63583 21188 63649 21211
rect 63735 21188 63817 21211
rect 63903 21188 63969 21211
rect 63583 21148 63592 21188
rect 63632 21148 63649 21188
rect 63735 21148 63756 21188
rect 63796 21148 63817 21188
rect 63903 21148 63920 21188
rect 63960 21148 63969 21188
rect 63583 21125 63649 21148
rect 63735 21125 63817 21148
rect 63903 21125 63969 21148
rect 63583 21106 63969 21125
rect 78703 21211 79089 21230
rect 78703 21188 78769 21211
rect 78855 21188 78937 21211
rect 79023 21188 79089 21211
rect 78703 21148 78712 21188
rect 78752 21148 78769 21188
rect 78855 21148 78876 21188
rect 78916 21148 78937 21188
rect 79023 21148 79040 21188
rect 79080 21148 79089 21188
rect 78703 21125 78769 21148
rect 78855 21125 78937 21148
rect 79023 21125 79089 21148
rect 78703 21106 79089 21125
rect 93823 21211 94209 21230
rect 93823 21188 93889 21211
rect 93975 21188 94057 21211
rect 94143 21188 94209 21211
rect 93823 21148 93832 21188
rect 93872 21148 93889 21188
rect 93975 21148 93996 21188
rect 94036 21148 94057 21188
rect 94143 21148 94160 21188
rect 94200 21148 94209 21188
rect 93823 21125 93889 21148
rect 93975 21125 94057 21148
rect 94143 21125 94209 21148
rect 93823 21106 94209 21125
rect 4343 20455 4729 20474
rect 4343 20432 4409 20455
rect 4495 20432 4577 20455
rect 4663 20432 4729 20455
rect 4343 20392 4352 20432
rect 4392 20392 4409 20432
rect 4495 20392 4516 20432
rect 4556 20392 4577 20432
rect 4663 20392 4680 20432
rect 4720 20392 4729 20432
rect 4343 20369 4409 20392
rect 4495 20369 4577 20392
rect 4663 20369 4729 20392
rect 4343 20350 4729 20369
rect 19463 20455 19849 20474
rect 19463 20432 19529 20455
rect 19615 20432 19697 20455
rect 19783 20432 19849 20455
rect 19463 20392 19472 20432
rect 19512 20392 19529 20432
rect 19615 20392 19636 20432
rect 19676 20392 19697 20432
rect 19783 20392 19800 20432
rect 19840 20392 19849 20432
rect 19463 20369 19529 20392
rect 19615 20369 19697 20392
rect 19783 20369 19849 20392
rect 19463 20350 19849 20369
rect 34583 20455 34969 20474
rect 34583 20432 34649 20455
rect 34735 20432 34817 20455
rect 34903 20432 34969 20455
rect 34583 20392 34592 20432
rect 34632 20392 34649 20432
rect 34735 20392 34756 20432
rect 34796 20392 34817 20432
rect 34903 20392 34920 20432
rect 34960 20392 34969 20432
rect 34583 20369 34649 20392
rect 34735 20369 34817 20392
rect 34903 20369 34969 20392
rect 34583 20350 34969 20369
rect 49703 20455 50089 20474
rect 49703 20432 49769 20455
rect 49855 20432 49937 20455
rect 50023 20432 50089 20455
rect 49703 20392 49712 20432
rect 49752 20392 49769 20432
rect 49855 20392 49876 20432
rect 49916 20392 49937 20432
rect 50023 20392 50040 20432
rect 50080 20392 50089 20432
rect 49703 20369 49769 20392
rect 49855 20369 49937 20392
rect 50023 20369 50089 20392
rect 49703 20350 50089 20369
rect 64823 20455 65209 20474
rect 64823 20432 64889 20455
rect 64975 20432 65057 20455
rect 65143 20432 65209 20455
rect 64823 20392 64832 20432
rect 64872 20392 64889 20432
rect 64975 20392 64996 20432
rect 65036 20392 65057 20432
rect 65143 20392 65160 20432
rect 65200 20392 65209 20432
rect 64823 20369 64889 20392
rect 64975 20369 65057 20392
rect 65143 20369 65209 20392
rect 64823 20350 65209 20369
rect 79943 20455 80329 20474
rect 79943 20432 80009 20455
rect 80095 20432 80177 20455
rect 80263 20432 80329 20455
rect 79943 20392 79952 20432
rect 79992 20392 80009 20432
rect 80095 20392 80116 20432
rect 80156 20392 80177 20432
rect 80263 20392 80280 20432
rect 80320 20392 80329 20432
rect 79943 20369 80009 20392
rect 80095 20369 80177 20392
rect 80263 20369 80329 20392
rect 79943 20350 80329 20369
rect 95063 20455 95449 20474
rect 95063 20432 95129 20455
rect 95215 20432 95297 20455
rect 95383 20432 95449 20455
rect 95063 20392 95072 20432
rect 95112 20392 95129 20432
rect 95215 20392 95236 20432
rect 95276 20392 95297 20432
rect 95383 20392 95400 20432
rect 95440 20392 95449 20432
rect 95063 20369 95129 20392
rect 95215 20369 95297 20392
rect 95383 20369 95449 20392
rect 95063 20350 95449 20369
rect 3103 19699 3489 19718
rect 3103 19676 3169 19699
rect 3255 19676 3337 19699
rect 3423 19676 3489 19699
rect 3103 19636 3112 19676
rect 3152 19636 3169 19676
rect 3255 19636 3276 19676
rect 3316 19636 3337 19676
rect 3423 19636 3440 19676
rect 3480 19636 3489 19676
rect 3103 19613 3169 19636
rect 3255 19613 3337 19636
rect 3423 19613 3489 19636
rect 3103 19594 3489 19613
rect 18223 19699 18609 19718
rect 18223 19676 18289 19699
rect 18375 19676 18457 19699
rect 18543 19676 18609 19699
rect 18223 19636 18232 19676
rect 18272 19636 18289 19676
rect 18375 19636 18396 19676
rect 18436 19636 18457 19676
rect 18543 19636 18560 19676
rect 18600 19636 18609 19676
rect 18223 19613 18289 19636
rect 18375 19613 18457 19636
rect 18543 19613 18609 19636
rect 18223 19594 18609 19613
rect 33343 19699 33729 19718
rect 33343 19676 33409 19699
rect 33495 19676 33577 19699
rect 33663 19676 33729 19699
rect 33343 19636 33352 19676
rect 33392 19636 33409 19676
rect 33495 19636 33516 19676
rect 33556 19636 33577 19676
rect 33663 19636 33680 19676
rect 33720 19636 33729 19676
rect 33343 19613 33409 19636
rect 33495 19613 33577 19636
rect 33663 19613 33729 19636
rect 33343 19594 33729 19613
rect 48463 19699 48849 19718
rect 48463 19676 48529 19699
rect 48615 19676 48697 19699
rect 48783 19676 48849 19699
rect 48463 19636 48472 19676
rect 48512 19636 48529 19676
rect 48615 19636 48636 19676
rect 48676 19636 48697 19676
rect 48783 19636 48800 19676
rect 48840 19636 48849 19676
rect 48463 19613 48529 19636
rect 48615 19613 48697 19636
rect 48783 19613 48849 19636
rect 48463 19594 48849 19613
rect 63583 19699 63969 19718
rect 63583 19676 63649 19699
rect 63735 19676 63817 19699
rect 63903 19676 63969 19699
rect 63583 19636 63592 19676
rect 63632 19636 63649 19676
rect 63735 19636 63756 19676
rect 63796 19636 63817 19676
rect 63903 19636 63920 19676
rect 63960 19636 63969 19676
rect 63583 19613 63649 19636
rect 63735 19613 63817 19636
rect 63903 19613 63969 19636
rect 63583 19594 63969 19613
rect 78703 19699 79089 19718
rect 78703 19676 78769 19699
rect 78855 19676 78937 19699
rect 79023 19676 79089 19699
rect 78703 19636 78712 19676
rect 78752 19636 78769 19676
rect 78855 19636 78876 19676
rect 78916 19636 78937 19676
rect 79023 19636 79040 19676
rect 79080 19636 79089 19676
rect 78703 19613 78769 19636
rect 78855 19613 78937 19636
rect 79023 19613 79089 19636
rect 78703 19594 79089 19613
rect 93823 19699 94209 19718
rect 93823 19676 93889 19699
rect 93975 19676 94057 19699
rect 94143 19676 94209 19699
rect 93823 19636 93832 19676
rect 93872 19636 93889 19676
rect 93975 19636 93996 19676
rect 94036 19636 94057 19676
rect 94143 19636 94160 19676
rect 94200 19636 94209 19676
rect 93823 19613 93889 19636
rect 93975 19613 94057 19636
rect 94143 19613 94209 19636
rect 93823 19594 94209 19613
rect 4343 18943 4729 18962
rect 4343 18920 4409 18943
rect 4495 18920 4577 18943
rect 4663 18920 4729 18943
rect 4343 18880 4352 18920
rect 4392 18880 4409 18920
rect 4495 18880 4516 18920
rect 4556 18880 4577 18920
rect 4663 18880 4680 18920
rect 4720 18880 4729 18920
rect 4343 18857 4409 18880
rect 4495 18857 4577 18880
rect 4663 18857 4729 18880
rect 4343 18838 4729 18857
rect 19463 18943 19849 18962
rect 19463 18920 19529 18943
rect 19615 18920 19697 18943
rect 19783 18920 19849 18943
rect 19463 18880 19472 18920
rect 19512 18880 19529 18920
rect 19615 18880 19636 18920
rect 19676 18880 19697 18920
rect 19783 18880 19800 18920
rect 19840 18880 19849 18920
rect 19463 18857 19529 18880
rect 19615 18857 19697 18880
rect 19783 18857 19849 18880
rect 19463 18838 19849 18857
rect 34583 18943 34969 18962
rect 34583 18920 34649 18943
rect 34735 18920 34817 18943
rect 34903 18920 34969 18943
rect 34583 18880 34592 18920
rect 34632 18880 34649 18920
rect 34735 18880 34756 18920
rect 34796 18880 34817 18920
rect 34903 18880 34920 18920
rect 34960 18880 34969 18920
rect 34583 18857 34649 18880
rect 34735 18857 34817 18880
rect 34903 18857 34969 18880
rect 34583 18838 34969 18857
rect 49703 18943 50089 18962
rect 49703 18920 49769 18943
rect 49855 18920 49937 18943
rect 50023 18920 50089 18943
rect 49703 18880 49712 18920
rect 49752 18880 49769 18920
rect 49855 18880 49876 18920
rect 49916 18880 49937 18920
rect 50023 18880 50040 18920
rect 50080 18880 50089 18920
rect 49703 18857 49769 18880
rect 49855 18857 49937 18880
rect 50023 18857 50089 18880
rect 49703 18838 50089 18857
rect 64823 18943 65209 18962
rect 64823 18920 64889 18943
rect 64975 18920 65057 18943
rect 65143 18920 65209 18943
rect 64823 18880 64832 18920
rect 64872 18880 64889 18920
rect 64975 18880 64996 18920
rect 65036 18880 65057 18920
rect 65143 18880 65160 18920
rect 65200 18880 65209 18920
rect 64823 18857 64889 18880
rect 64975 18857 65057 18880
rect 65143 18857 65209 18880
rect 64823 18838 65209 18857
rect 79943 18943 80329 18962
rect 79943 18920 80009 18943
rect 80095 18920 80177 18943
rect 80263 18920 80329 18943
rect 79943 18880 79952 18920
rect 79992 18880 80009 18920
rect 80095 18880 80116 18920
rect 80156 18880 80177 18920
rect 80263 18880 80280 18920
rect 80320 18880 80329 18920
rect 79943 18857 80009 18880
rect 80095 18857 80177 18880
rect 80263 18857 80329 18880
rect 79943 18838 80329 18857
rect 95063 18943 95449 18962
rect 95063 18920 95129 18943
rect 95215 18920 95297 18943
rect 95383 18920 95449 18943
rect 95063 18880 95072 18920
rect 95112 18880 95129 18920
rect 95215 18880 95236 18920
rect 95276 18880 95297 18920
rect 95383 18880 95400 18920
rect 95440 18880 95449 18920
rect 95063 18857 95129 18880
rect 95215 18857 95297 18880
rect 95383 18857 95449 18880
rect 95063 18838 95449 18857
rect 3103 18187 3489 18206
rect 3103 18164 3169 18187
rect 3255 18164 3337 18187
rect 3423 18164 3489 18187
rect 3103 18124 3112 18164
rect 3152 18124 3169 18164
rect 3255 18124 3276 18164
rect 3316 18124 3337 18164
rect 3423 18124 3440 18164
rect 3480 18124 3489 18164
rect 3103 18101 3169 18124
rect 3255 18101 3337 18124
rect 3423 18101 3489 18124
rect 3103 18082 3489 18101
rect 18223 18187 18609 18206
rect 18223 18164 18289 18187
rect 18375 18164 18457 18187
rect 18543 18164 18609 18187
rect 18223 18124 18232 18164
rect 18272 18124 18289 18164
rect 18375 18124 18396 18164
rect 18436 18124 18457 18164
rect 18543 18124 18560 18164
rect 18600 18124 18609 18164
rect 18223 18101 18289 18124
rect 18375 18101 18457 18124
rect 18543 18101 18609 18124
rect 18223 18082 18609 18101
rect 33343 18187 33729 18206
rect 33343 18164 33409 18187
rect 33495 18164 33577 18187
rect 33663 18164 33729 18187
rect 33343 18124 33352 18164
rect 33392 18124 33409 18164
rect 33495 18124 33516 18164
rect 33556 18124 33577 18164
rect 33663 18124 33680 18164
rect 33720 18124 33729 18164
rect 33343 18101 33409 18124
rect 33495 18101 33577 18124
rect 33663 18101 33729 18124
rect 33343 18082 33729 18101
rect 48463 18187 48849 18206
rect 48463 18164 48529 18187
rect 48615 18164 48697 18187
rect 48783 18164 48849 18187
rect 48463 18124 48472 18164
rect 48512 18124 48529 18164
rect 48615 18124 48636 18164
rect 48676 18124 48697 18164
rect 48783 18124 48800 18164
rect 48840 18124 48849 18164
rect 48463 18101 48529 18124
rect 48615 18101 48697 18124
rect 48783 18101 48849 18124
rect 48463 18082 48849 18101
rect 63583 18187 63969 18206
rect 63583 18164 63649 18187
rect 63735 18164 63817 18187
rect 63903 18164 63969 18187
rect 63583 18124 63592 18164
rect 63632 18124 63649 18164
rect 63735 18124 63756 18164
rect 63796 18124 63817 18164
rect 63903 18124 63920 18164
rect 63960 18124 63969 18164
rect 63583 18101 63649 18124
rect 63735 18101 63817 18124
rect 63903 18101 63969 18124
rect 63583 18082 63969 18101
rect 78703 18187 79089 18206
rect 78703 18164 78769 18187
rect 78855 18164 78937 18187
rect 79023 18164 79089 18187
rect 78703 18124 78712 18164
rect 78752 18124 78769 18164
rect 78855 18124 78876 18164
rect 78916 18124 78937 18164
rect 79023 18124 79040 18164
rect 79080 18124 79089 18164
rect 78703 18101 78769 18124
rect 78855 18101 78937 18124
rect 79023 18101 79089 18124
rect 78703 18082 79089 18101
rect 93823 18187 94209 18206
rect 93823 18164 93889 18187
rect 93975 18164 94057 18187
rect 94143 18164 94209 18187
rect 93823 18124 93832 18164
rect 93872 18124 93889 18164
rect 93975 18124 93996 18164
rect 94036 18124 94057 18164
rect 94143 18124 94160 18164
rect 94200 18124 94209 18164
rect 93823 18101 93889 18124
rect 93975 18101 94057 18124
rect 94143 18101 94209 18124
rect 93823 18082 94209 18101
rect 4343 17431 4729 17450
rect 4343 17408 4409 17431
rect 4495 17408 4577 17431
rect 4663 17408 4729 17431
rect 4343 17368 4352 17408
rect 4392 17368 4409 17408
rect 4495 17368 4516 17408
rect 4556 17368 4577 17408
rect 4663 17368 4680 17408
rect 4720 17368 4729 17408
rect 4343 17345 4409 17368
rect 4495 17345 4577 17368
rect 4663 17345 4729 17368
rect 4343 17326 4729 17345
rect 19463 17431 19849 17450
rect 19463 17408 19529 17431
rect 19615 17408 19697 17431
rect 19783 17408 19849 17431
rect 19463 17368 19472 17408
rect 19512 17368 19529 17408
rect 19615 17368 19636 17408
rect 19676 17368 19697 17408
rect 19783 17368 19800 17408
rect 19840 17368 19849 17408
rect 19463 17345 19529 17368
rect 19615 17345 19697 17368
rect 19783 17345 19849 17368
rect 19463 17326 19849 17345
rect 34583 17431 34969 17450
rect 34583 17408 34649 17431
rect 34735 17408 34817 17431
rect 34903 17408 34969 17431
rect 34583 17368 34592 17408
rect 34632 17368 34649 17408
rect 34735 17368 34756 17408
rect 34796 17368 34817 17408
rect 34903 17368 34920 17408
rect 34960 17368 34969 17408
rect 34583 17345 34649 17368
rect 34735 17345 34817 17368
rect 34903 17345 34969 17368
rect 34583 17326 34969 17345
rect 49703 17431 50089 17450
rect 49703 17408 49769 17431
rect 49855 17408 49937 17431
rect 50023 17408 50089 17431
rect 49703 17368 49712 17408
rect 49752 17368 49769 17408
rect 49855 17368 49876 17408
rect 49916 17368 49937 17408
rect 50023 17368 50040 17408
rect 50080 17368 50089 17408
rect 49703 17345 49769 17368
rect 49855 17345 49937 17368
rect 50023 17345 50089 17368
rect 49703 17326 50089 17345
rect 64823 17431 65209 17450
rect 64823 17408 64889 17431
rect 64975 17408 65057 17431
rect 65143 17408 65209 17431
rect 64823 17368 64832 17408
rect 64872 17368 64889 17408
rect 64975 17368 64996 17408
rect 65036 17368 65057 17408
rect 65143 17368 65160 17408
rect 65200 17368 65209 17408
rect 64823 17345 64889 17368
rect 64975 17345 65057 17368
rect 65143 17345 65209 17368
rect 64823 17326 65209 17345
rect 79943 17431 80329 17450
rect 79943 17408 80009 17431
rect 80095 17408 80177 17431
rect 80263 17408 80329 17431
rect 79943 17368 79952 17408
rect 79992 17368 80009 17408
rect 80095 17368 80116 17408
rect 80156 17368 80177 17408
rect 80263 17368 80280 17408
rect 80320 17368 80329 17408
rect 79943 17345 80009 17368
rect 80095 17345 80177 17368
rect 80263 17345 80329 17368
rect 79943 17326 80329 17345
rect 95063 17431 95449 17450
rect 95063 17408 95129 17431
rect 95215 17408 95297 17431
rect 95383 17408 95449 17431
rect 95063 17368 95072 17408
rect 95112 17368 95129 17408
rect 95215 17368 95236 17408
rect 95276 17368 95297 17408
rect 95383 17368 95400 17408
rect 95440 17368 95449 17408
rect 95063 17345 95129 17368
rect 95215 17345 95297 17368
rect 95383 17345 95449 17368
rect 95063 17326 95449 17345
rect 3103 16675 3489 16694
rect 3103 16652 3169 16675
rect 3255 16652 3337 16675
rect 3423 16652 3489 16675
rect 3103 16612 3112 16652
rect 3152 16612 3169 16652
rect 3255 16612 3276 16652
rect 3316 16612 3337 16652
rect 3423 16612 3440 16652
rect 3480 16612 3489 16652
rect 3103 16589 3169 16612
rect 3255 16589 3337 16612
rect 3423 16589 3489 16612
rect 3103 16570 3489 16589
rect 18223 16675 18609 16694
rect 18223 16652 18289 16675
rect 18375 16652 18457 16675
rect 18543 16652 18609 16675
rect 18223 16612 18232 16652
rect 18272 16612 18289 16652
rect 18375 16612 18396 16652
rect 18436 16612 18457 16652
rect 18543 16612 18560 16652
rect 18600 16612 18609 16652
rect 18223 16589 18289 16612
rect 18375 16589 18457 16612
rect 18543 16589 18609 16612
rect 18223 16570 18609 16589
rect 33343 16675 33729 16694
rect 33343 16652 33409 16675
rect 33495 16652 33577 16675
rect 33663 16652 33729 16675
rect 33343 16612 33352 16652
rect 33392 16612 33409 16652
rect 33495 16612 33516 16652
rect 33556 16612 33577 16652
rect 33663 16612 33680 16652
rect 33720 16612 33729 16652
rect 33343 16589 33409 16612
rect 33495 16589 33577 16612
rect 33663 16589 33729 16612
rect 33343 16570 33729 16589
rect 48463 16675 48849 16694
rect 48463 16652 48529 16675
rect 48615 16652 48697 16675
rect 48783 16652 48849 16675
rect 48463 16612 48472 16652
rect 48512 16612 48529 16652
rect 48615 16612 48636 16652
rect 48676 16612 48697 16652
rect 48783 16612 48800 16652
rect 48840 16612 48849 16652
rect 48463 16589 48529 16612
rect 48615 16589 48697 16612
rect 48783 16589 48849 16612
rect 48463 16570 48849 16589
rect 63583 16675 63969 16694
rect 63583 16652 63649 16675
rect 63735 16652 63817 16675
rect 63903 16652 63969 16675
rect 63583 16612 63592 16652
rect 63632 16612 63649 16652
rect 63735 16612 63756 16652
rect 63796 16612 63817 16652
rect 63903 16612 63920 16652
rect 63960 16612 63969 16652
rect 63583 16589 63649 16612
rect 63735 16589 63817 16612
rect 63903 16589 63969 16612
rect 63583 16570 63969 16589
rect 78703 16675 79089 16694
rect 78703 16652 78769 16675
rect 78855 16652 78937 16675
rect 79023 16652 79089 16675
rect 78703 16612 78712 16652
rect 78752 16612 78769 16652
rect 78855 16612 78876 16652
rect 78916 16612 78937 16652
rect 79023 16612 79040 16652
rect 79080 16612 79089 16652
rect 78703 16589 78769 16612
rect 78855 16589 78937 16612
rect 79023 16589 79089 16612
rect 78703 16570 79089 16589
rect 93823 16675 94209 16694
rect 93823 16652 93889 16675
rect 93975 16652 94057 16675
rect 94143 16652 94209 16675
rect 93823 16612 93832 16652
rect 93872 16612 93889 16652
rect 93975 16612 93996 16652
rect 94036 16612 94057 16652
rect 94143 16612 94160 16652
rect 94200 16612 94209 16652
rect 93823 16589 93889 16612
rect 93975 16589 94057 16612
rect 94143 16589 94209 16612
rect 93823 16570 94209 16589
rect 4343 15919 4729 15938
rect 4343 15896 4409 15919
rect 4495 15896 4577 15919
rect 4663 15896 4729 15919
rect 4343 15856 4352 15896
rect 4392 15856 4409 15896
rect 4495 15856 4516 15896
rect 4556 15856 4577 15896
rect 4663 15856 4680 15896
rect 4720 15856 4729 15896
rect 4343 15833 4409 15856
rect 4495 15833 4577 15856
rect 4663 15833 4729 15856
rect 4343 15814 4729 15833
rect 19463 15919 19849 15938
rect 19463 15896 19529 15919
rect 19615 15896 19697 15919
rect 19783 15896 19849 15919
rect 19463 15856 19472 15896
rect 19512 15856 19529 15896
rect 19615 15856 19636 15896
rect 19676 15856 19697 15896
rect 19783 15856 19800 15896
rect 19840 15856 19849 15896
rect 19463 15833 19529 15856
rect 19615 15833 19697 15856
rect 19783 15833 19849 15856
rect 19463 15814 19849 15833
rect 34583 15919 34969 15938
rect 34583 15896 34649 15919
rect 34735 15896 34817 15919
rect 34903 15896 34969 15919
rect 34583 15856 34592 15896
rect 34632 15856 34649 15896
rect 34735 15856 34756 15896
rect 34796 15856 34817 15896
rect 34903 15856 34920 15896
rect 34960 15856 34969 15896
rect 34583 15833 34649 15856
rect 34735 15833 34817 15856
rect 34903 15833 34969 15856
rect 34583 15814 34969 15833
rect 49703 15919 50089 15938
rect 49703 15896 49769 15919
rect 49855 15896 49937 15919
rect 50023 15896 50089 15919
rect 49703 15856 49712 15896
rect 49752 15856 49769 15896
rect 49855 15856 49876 15896
rect 49916 15856 49937 15896
rect 50023 15856 50040 15896
rect 50080 15856 50089 15896
rect 49703 15833 49769 15856
rect 49855 15833 49937 15856
rect 50023 15833 50089 15856
rect 49703 15814 50089 15833
rect 64823 15919 65209 15938
rect 64823 15896 64889 15919
rect 64975 15896 65057 15919
rect 65143 15896 65209 15919
rect 64823 15856 64832 15896
rect 64872 15856 64889 15896
rect 64975 15856 64996 15896
rect 65036 15856 65057 15896
rect 65143 15856 65160 15896
rect 65200 15856 65209 15896
rect 64823 15833 64889 15856
rect 64975 15833 65057 15856
rect 65143 15833 65209 15856
rect 64823 15814 65209 15833
rect 79943 15919 80329 15938
rect 79943 15896 80009 15919
rect 80095 15896 80177 15919
rect 80263 15896 80329 15919
rect 79943 15856 79952 15896
rect 79992 15856 80009 15896
rect 80095 15856 80116 15896
rect 80156 15856 80177 15896
rect 80263 15856 80280 15896
rect 80320 15856 80329 15896
rect 79943 15833 80009 15856
rect 80095 15833 80177 15856
rect 80263 15833 80329 15856
rect 79943 15814 80329 15833
rect 95063 15919 95449 15938
rect 95063 15896 95129 15919
rect 95215 15896 95297 15919
rect 95383 15896 95449 15919
rect 95063 15856 95072 15896
rect 95112 15856 95129 15896
rect 95215 15856 95236 15896
rect 95276 15856 95297 15896
rect 95383 15856 95400 15896
rect 95440 15856 95449 15896
rect 95063 15833 95129 15856
rect 95215 15833 95297 15856
rect 95383 15833 95449 15856
rect 95063 15814 95449 15833
rect 3103 15163 3489 15182
rect 3103 15140 3169 15163
rect 3255 15140 3337 15163
rect 3423 15140 3489 15163
rect 3103 15100 3112 15140
rect 3152 15100 3169 15140
rect 3255 15100 3276 15140
rect 3316 15100 3337 15140
rect 3423 15100 3440 15140
rect 3480 15100 3489 15140
rect 3103 15077 3169 15100
rect 3255 15077 3337 15100
rect 3423 15077 3489 15100
rect 3103 15058 3489 15077
rect 18223 15163 18609 15182
rect 18223 15140 18289 15163
rect 18375 15140 18457 15163
rect 18543 15140 18609 15163
rect 18223 15100 18232 15140
rect 18272 15100 18289 15140
rect 18375 15100 18396 15140
rect 18436 15100 18457 15140
rect 18543 15100 18560 15140
rect 18600 15100 18609 15140
rect 18223 15077 18289 15100
rect 18375 15077 18457 15100
rect 18543 15077 18609 15100
rect 18223 15058 18609 15077
rect 33343 15163 33729 15182
rect 33343 15140 33409 15163
rect 33495 15140 33577 15163
rect 33663 15140 33729 15163
rect 33343 15100 33352 15140
rect 33392 15100 33409 15140
rect 33495 15100 33516 15140
rect 33556 15100 33577 15140
rect 33663 15100 33680 15140
rect 33720 15100 33729 15140
rect 33343 15077 33409 15100
rect 33495 15077 33577 15100
rect 33663 15077 33729 15100
rect 33343 15058 33729 15077
rect 48463 15163 48849 15182
rect 48463 15140 48529 15163
rect 48615 15140 48697 15163
rect 48783 15140 48849 15163
rect 48463 15100 48472 15140
rect 48512 15100 48529 15140
rect 48615 15100 48636 15140
rect 48676 15100 48697 15140
rect 48783 15100 48800 15140
rect 48840 15100 48849 15140
rect 48463 15077 48529 15100
rect 48615 15077 48697 15100
rect 48783 15077 48849 15100
rect 48463 15058 48849 15077
rect 63583 15163 63969 15182
rect 63583 15140 63649 15163
rect 63735 15140 63817 15163
rect 63903 15140 63969 15163
rect 63583 15100 63592 15140
rect 63632 15100 63649 15140
rect 63735 15100 63756 15140
rect 63796 15100 63817 15140
rect 63903 15100 63920 15140
rect 63960 15100 63969 15140
rect 63583 15077 63649 15100
rect 63735 15077 63817 15100
rect 63903 15077 63969 15100
rect 63583 15058 63969 15077
rect 78703 15163 79089 15182
rect 78703 15140 78769 15163
rect 78855 15140 78937 15163
rect 79023 15140 79089 15163
rect 78703 15100 78712 15140
rect 78752 15100 78769 15140
rect 78855 15100 78876 15140
rect 78916 15100 78937 15140
rect 79023 15100 79040 15140
rect 79080 15100 79089 15140
rect 78703 15077 78769 15100
rect 78855 15077 78937 15100
rect 79023 15077 79089 15100
rect 78703 15058 79089 15077
rect 93823 15163 94209 15182
rect 93823 15140 93889 15163
rect 93975 15140 94057 15163
rect 94143 15140 94209 15163
rect 93823 15100 93832 15140
rect 93872 15100 93889 15140
rect 93975 15100 93996 15140
rect 94036 15100 94057 15140
rect 94143 15100 94160 15140
rect 94200 15100 94209 15140
rect 93823 15077 93889 15100
rect 93975 15077 94057 15100
rect 94143 15077 94209 15100
rect 93823 15058 94209 15077
rect 4343 14407 4729 14426
rect 4343 14384 4409 14407
rect 4495 14384 4577 14407
rect 4663 14384 4729 14407
rect 4343 14344 4352 14384
rect 4392 14344 4409 14384
rect 4495 14344 4516 14384
rect 4556 14344 4577 14384
rect 4663 14344 4680 14384
rect 4720 14344 4729 14384
rect 4343 14321 4409 14344
rect 4495 14321 4577 14344
rect 4663 14321 4729 14344
rect 4343 14302 4729 14321
rect 19463 14407 19849 14426
rect 19463 14384 19529 14407
rect 19615 14384 19697 14407
rect 19783 14384 19849 14407
rect 19463 14344 19472 14384
rect 19512 14344 19529 14384
rect 19615 14344 19636 14384
rect 19676 14344 19697 14384
rect 19783 14344 19800 14384
rect 19840 14344 19849 14384
rect 19463 14321 19529 14344
rect 19615 14321 19697 14344
rect 19783 14321 19849 14344
rect 19463 14302 19849 14321
rect 34583 14407 34969 14426
rect 34583 14384 34649 14407
rect 34735 14384 34817 14407
rect 34903 14384 34969 14407
rect 34583 14344 34592 14384
rect 34632 14344 34649 14384
rect 34735 14344 34756 14384
rect 34796 14344 34817 14384
rect 34903 14344 34920 14384
rect 34960 14344 34969 14384
rect 34583 14321 34649 14344
rect 34735 14321 34817 14344
rect 34903 14321 34969 14344
rect 34583 14302 34969 14321
rect 49703 14407 50089 14426
rect 49703 14384 49769 14407
rect 49855 14384 49937 14407
rect 50023 14384 50089 14407
rect 49703 14344 49712 14384
rect 49752 14344 49769 14384
rect 49855 14344 49876 14384
rect 49916 14344 49937 14384
rect 50023 14344 50040 14384
rect 50080 14344 50089 14384
rect 49703 14321 49769 14344
rect 49855 14321 49937 14344
rect 50023 14321 50089 14344
rect 49703 14302 50089 14321
rect 64823 14407 65209 14426
rect 64823 14384 64889 14407
rect 64975 14384 65057 14407
rect 65143 14384 65209 14407
rect 64823 14344 64832 14384
rect 64872 14344 64889 14384
rect 64975 14344 64996 14384
rect 65036 14344 65057 14384
rect 65143 14344 65160 14384
rect 65200 14344 65209 14384
rect 64823 14321 64889 14344
rect 64975 14321 65057 14344
rect 65143 14321 65209 14344
rect 64823 14302 65209 14321
rect 79943 14407 80329 14426
rect 79943 14384 80009 14407
rect 80095 14384 80177 14407
rect 80263 14384 80329 14407
rect 79943 14344 79952 14384
rect 79992 14344 80009 14384
rect 80095 14344 80116 14384
rect 80156 14344 80177 14384
rect 80263 14344 80280 14384
rect 80320 14344 80329 14384
rect 79943 14321 80009 14344
rect 80095 14321 80177 14344
rect 80263 14321 80329 14344
rect 79943 14302 80329 14321
rect 95063 14407 95449 14426
rect 95063 14384 95129 14407
rect 95215 14384 95297 14407
rect 95383 14384 95449 14407
rect 95063 14344 95072 14384
rect 95112 14344 95129 14384
rect 95215 14344 95236 14384
rect 95276 14344 95297 14384
rect 95383 14344 95400 14384
rect 95440 14344 95449 14384
rect 95063 14321 95129 14344
rect 95215 14321 95297 14344
rect 95383 14321 95449 14344
rect 95063 14302 95449 14321
rect 3103 13651 3489 13670
rect 3103 13628 3169 13651
rect 3255 13628 3337 13651
rect 3423 13628 3489 13651
rect 3103 13588 3112 13628
rect 3152 13588 3169 13628
rect 3255 13588 3276 13628
rect 3316 13588 3337 13628
rect 3423 13588 3440 13628
rect 3480 13588 3489 13628
rect 3103 13565 3169 13588
rect 3255 13565 3337 13588
rect 3423 13565 3489 13588
rect 3103 13546 3489 13565
rect 18223 13651 18609 13670
rect 18223 13628 18289 13651
rect 18375 13628 18457 13651
rect 18543 13628 18609 13651
rect 18223 13588 18232 13628
rect 18272 13588 18289 13628
rect 18375 13588 18396 13628
rect 18436 13588 18457 13628
rect 18543 13588 18560 13628
rect 18600 13588 18609 13628
rect 18223 13565 18289 13588
rect 18375 13565 18457 13588
rect 18543 13565 18609 13588
rect 18223 13546 18609 13565
rect 33343 13651 33729 13670
rect 33343 13628 33409 13651
rect 33495 13628 33577 13651
rect 33663 13628 33729 13651
rect 33343 13588 33352 13628
rect 33392 13588 33409 13628
rect 33495 13588 33516 13628
rect 33556 13588 33577 13628
rect 33663 13588 33680 13628
rect 33720 13588 33729 13628
rect 33343 13565 33409 13588
rect 33495 13565 33577 13588
rect 33663 13565 33729 13588
rect 33343 13546 33729 13565
rect 48463 13651 48849 13670
rect 48463 13628 48529 13651
rect 48615 13628 48697 13651
rect 48783 13628 48849 13651
rect 48463 13588 48472 13628
rect 48512 13588 48529 13628
rect 48615 13588 48636 13628
rect 48676 13588 48697 13628
rect 48783 13588 48800 13628
rect 48840 13588 48849 13628
rect 48463 13565 48529 13588
rect 48615 13565 48697 13588
rect 48783 13565 48849 13588
rect 48463 13546 48849 13565
rect 63583 13651 63969 13670
rect 63583 13628 63649 13651
rect 63735 13628 63817 13651
rect 63903 13628 63969 13651
rect 63583 13588 63592 13628
rect 63632 13588 63649 13628
rect 63735 13588 63756 13628
rect 63796 13588 63817 13628
rect 63903 13588 63920 13628
rect 63960 13588 63969 13628
rect 63583 13565 63649 13588
rect 63735 13565 63817 13588
rect 63903 13565 63969 13588
rect 63583 13546 63969 13565
rect 78703 13651 79089 13670
rect 78703 13628 78769 13651
rect 78855 13628 78937 13651
rect 79023 13628 79089 13651
rect 78703 13588 78712 13628
rect 78752 13588 78769 13628
rect 78855 13588 78876 13628
rect 78916 13588 78937 13628
rect 79023 13588 79040 13628
rect 79080 13588 79089 13628
rect 78703 13565 78769 13588
rect 78855 13565 78937 13588
rect 79023 13565 79089 13588
rect 78703 13546 79089 13565
rect 93823 13651 94209 13670
rect 93823 13628 93889 13651
rect 93975 13628 94057 13651
rect 94143 13628 94209 13651
rect 93823 13588 93832 13628
rect 93872 13588 93889 13628
rect 93975 13588 93996 13628
rect 94036 13588 94057 13628
rect 94143 13588 94160 13628
rect 94200 13588 94209 13628
rect 93823 13565 93889 13588
rect 93975 13565 94057 13588
rect 94143 13565 94209 13588
rect 93823 13546 94209 13565
rect 4343 12895 4729 12914
rect 4343 12872 4409 12895
rect 4495 12872 4577 12895
rect 4663 12872 4729 12895
rect 4343 12832 4352 12872
rect 4392 12832 4409 12872
rect 4495 12832 4516 12872
rect 4556 12832 4577 12872
rect 4663 12832 4680 12872
rect 4720 12832 4729 12872
rect 4343 12809 4409 12832
rect 4495 12809 4577 12832
rect 4663 12809 4729 12832
rect 4343 12790 4729 12809
rect 19463 12895 19849 12914
rect 19463 12872 19529 12895
rect 19615 12872 19697 12895
rect 19783 12872 19849 12895
rect 19463 12832 19472 12872
rect 19512 12832 19529 12872
rect 19615 12832 19636 12872
rect 19676 12832 19697 12872
rect 19783 12832 19800 12872
rect 19840 12832 19849 12872
rect 19463 12809 19529 12832
rect 19615 12809 19697 12832
rect 19783 12809 19849 12832
rect 19463 12790 19849 12809
rect 34583 12895 34969 12914
rect 34583 12872 34649 12895
rect 34735 12872 34817 12895
rect 34903 12872 34969 12895
rect 34583 12832 34592 12872
rect 34632 12832 34649 12872
rect 34735 12832 34756 12872
rect 34796 12832 34817 12872
rect 34903 12832 34920 12872
rect 34960 12832 34969 12872
rect 34583 12809 34649 12832
rect 34735 12809 34817 12832
rect 34903 12809 34969 12832
rect 34583 12790 34969 12809
rect 49703 12895 50089 12914
rect 49703 12872 49769 12895
rect 49855 12872 49937 12895
rect 50023 12872 50089 12895
rect 49703 12832 49712 12872
rect 49752 12832 49769 12872
rect 49855 12832 49876 12872
rect 49916 12832 49937 12872
rect 50023 12832 50040 12872
rect 50080 12832 50089 12872
rect 49703 12809 49769 12832
rect 49855 12809 49937 12832
rect 50023 12809 50089 12832
rect 49703 12790 50089 12809
rect 64823 12895 65209 12914
rect 64823 12872 64889 12895
rect 64975 12872 65057 12895
rect 65143 12872 65209 12895
rect 64823 12832 64832 12872
rect 64872 12832 64889 12872
rect 64975 12832 64996 12872
rect 65036 12832 65057 12872
rect 65143 12832 65160 12872
rect 65200 12832 65209 12872
rect 64823 12809 64889 12832
rect 64975 12809 65057 12832
rect 65143 12809 65209 12832
rect 64823 12790 65209 12809
rect 79943 12895 80329 12914
rect 79943 12872 80009 12895
rect 80095 12872 80177 12895
rect 80263 12872 80329 12895
rect 79943 12832 79952 12872
rect 79992 12832 80009 12872
rect 80095 12832 80116 12872
rect 80156 12832 80177 12872
rect 80263 12832 80280 12872
rect 80320 12832 80329 12872
rect 79943 12809 80009 12832
rect 80095 12809 80177 12832
rect 80263 12809 80329 12832
rect 79943 12790 80329 12809
rect 95063 12895 95449 12914
rect 95063 12872 95129 12895
rect 95215 12872 95297 12895
rect 95383 12872 95449 12895
rect 95063 12832 95072 12872
rect 95112 12832 95129 12872
rect 95215 12832 95236 12872
rect 95276 12832 95297 12872
rect 95383 12832 95400 12872
rect 95440 12832 95449 12872
rect 95063 12809 95129 12832
rect 95215 12809 95297 12832
rect 95383 12809 95449 12832
rect 95063 12790 95449 12809
rect 3103 12139 3489 12158
rect 3103 12116 3169 12139
rect 3255 12116 3337 12139
rect 3423 12116 3489 12139
rect 3103 12076 3112 12116
rect 3152 12076 3169 12116
rect 3255 12076 3276 12116
rect 3316 12076 3337 12116
rect 3423 12076 3440 12116
rect 3480 12076 3489 12116
rect 3103 12053 3169 12076
rect 3255 12053 3337 12076
rect 3423 12053 3489 12076
rect 3103 12034 3489 12053
rect 18223 12139 18609 12158
rect 18223 12116 18289 12139
rect 18375 12116 18457 12139
rect 18543 12116 18609 12139
rect 18223 12076 18232 12116
rect 18272 12076 18289 12116
rect 18375 12076 18396 12116
rect 18436 12076 18457 12116
rect 18543 12076 18560 12116
rect 18600 12076 18609 12116
rect 18223 12053 18289 12076
rect 18375 12053 18457 12076
rect 18543 12053 18609 12076
rect 18223 12034 18609 12053
rect 33343 12139 33729 12158
rect 33343 12116 33409 12139
rect 33495 12116 33577 12139
rect 33663 12116 33729 12139
rect 33343 12076 33352 12116
rect 33392 12076 33409 12116
rect 33495 12076 33516 12116
rect 33556 12076 33577 12116
rect 33663 12076 33680 12116
rect 33720 12076 33729 12116
rect 33343 12053 33409 12076
rect 33495 12053 33577 12076
rect 33663 12053 33729 12076
rect 33343 12034 33729 12053
rect 48463 12139 48849 12158
rect 48463 12116 48529 12139
rect 48615 12116 48697 12139
rect 48783 12116 48849 12139
rect 48463 12076 48472 12116
rect 48512 12076 48529 12116
rect 48615 12076 48636 12116
rect 48676 12076 48697 12116
rect 48783 12076 48800 12116
rect 48840 12076 48849 12116
rect 48463 12053 48529 12076
rect 48615 12053 48697 12076
rect 48783 12053 48849 12076
rect 48463 12034 48849 12053
rect 63583 12139 63969 12158
rect 63583 12116 63649 12139
rect 63735 12116 63817 12139
rect 63903 12116 63969 12139
rect 63583 12076 63592 12116
rect 63632 12076 63649 12116
rect 63735 12076 63756 12116
rect 63796 12076 63817 12116
rect 63903 12076 63920 12116
rect 63960 12076 63969 12116
rect 63583 12053 63649 12076
rect 63735 12053 63817 12076
rect 63903 12053 63969 12076
rect 63583 12034 63969 12053
rect 78703 12139 79089 12158
rect 78703 12116 78769 12139
rect 78855 12116 78937 12139
rect 79023 12116 79089 12139
rect 78703 12076 78712 12116
rect 78752 12076 78769 12116
rect 78855 12076 78876 12116
rect 78916 12076 78937 12116
rect 79023 12076 79040 12116
rect 79080 12076 79089 12116
rect 78703 12053 78769 12076
rect 78855 12053 78937 12076
rect 79023 12053 79089 12076
rect 78703 12034 79089 12053
rect 93823 12139 94209 12158
rect 93823 12116 93889 12139
rect 93975 12116 94057 12139
rect 94143 12116 94209 12139
rect 93823 12076 93832 12116
rect 93872 12076 93889 12116
rect 93975 12076 93996 12116
rect 94036 12076 94057 12116
rect 94143 12076 94160 12116
rect 94200 12076 94209 12116
rect 93823 12053 93889 12076
rect 93975 12053 94057 12076
rect 94143 12053 94209 12076
rect 93823 12034 94209 12053
rect 4343 11383 4729 11402
rect 4343 11360 4409 11383
rect 4495 11360 4577 11383
rect 4663 11360 4729 11383
rect 4343 11320 4352 11360
rect 4392 11320 4409 11360
rect 4495 11320 4516 11360
rect 4556 11320 4577 11360
rect 4663 11320 4680 11360
rect 4720 11320 4729 11360
rect 4343 11297 4409 11320
rect 4495 11297 4577 11320
rect 4663 11297 4729 11320
rect 4343 11278 4729 11297
rect 19463 11383 19849 11402
rect 19463 11360 19529 11383
rect 19615 11360 19697 11383
rect 19783 11360 19849 11383
rect 19463 11320 19472 11360
rect 19512 11320 19529 11360
rect 19615 11320 19636 11360
rect 19676 11320 19697 11360
rect 19783 11320 19800 11360
rect 19840 11320 19849 11360
rect 19463 11297 19529 11320
rect 19615 11297 19697 11320
rect 19783 11297 19849 11320
rect 19463 11278 19849 11297
rect 34583 11383 34969 11402
rect 34583 11360 34649 11383
rect 34735 11360 34817 11383
rect 34903 11360 34969 11383
rect 34583 11320 34592 11360
rect 34632 11320 34649 11360
rect 34735 11320 34756 11360
rect 34796 11320 34817 11360
rect 34903 11320 34920 11360
rect 34960 11320 34969 11360
rect 34583 11297 34649 11320
rect 34735 11297 34817 11320
rect 34903 11297 34969 11320
rect 34583 11278 34969 11297
rect 49703 11383 50089 11402
rect 49703 11360 49769 11383
rect 49855 11360 49937 11383
rect 50023 11360 50089 11383
rect 49703 11320 49712 11360
rect 49752 11320 49769 11360
rect 49855 11320 49876 11360
rect 49916 11320 49937 11360
rect 50023 11320 50040 11360
rect 50080 11320 50089 11360
rect 49703 11297 49769 11320
rect 49855 11297 49937 11320
rect 50023 11297 50089 11320
rect 49703 11278 50089 11297
rect 64823 11383 65209 11402
rect 64823 11360 64889 11383
rect 64975 11360 65057 11383
rect 65143 11360 65209 11383
rect 64823 11320 64832 11360
rect 64872 11320 64889 11360
rect 64975 11320 64996 11360
rect 65036 11320 65057 11360
rect 65143 11320 65160 11360
rect 65200 11320 65209 11360
rect 64823 11297 64889 11320
rect 64975 11297 65057 11320
rect 65143 11297 65209 11320
rect 64823 11278 65209 11297
rect 79943 11383 80329 11402
rect 79943 11360 80009 11383
rect 80095 11360 80177 11383
rect 80263 11360 80329 11383
rect 79943 11320 79952 11360
rect 79992 11320 80009 11360
rect 80095 11320 80116 11360
rect 80156 11320 80177 11360
rect 80263 11320 80280 11360
rect 80320 11320 80329 11360
rect 79943 11297 80009 11320
rect 80095 11297 80177 11320
rect 80263 11297 80329 11320
rect 79943 11278 80329 11297
rect 95063 11383 95449 11402
rect 95063 11360 95129 11383
rect 95215 11360 95297 11383
rect 95383 11360 95449 11383
rect 95063 11320 95072 11360
rect 95112 11320 95129 11360
rect 95215 11320 95236 11360
rect 95276 11320 95297 11360
rect 95383 11320 95400 11360
rect 95440 11320 95449 11360
rect 95063 11297 95129 11320
rect 95215 11297 95297 11320
rect 95383 11297 95449 11320
rect 95063 11278 95449 11297
rect 3103 10627 3489 10646
rect 3103 10604 3169 10627
rect 3255 10604 3337 10627
rect 3423 10604 3489 10627
rect 3103 10564 3112 10604
rect 3152 10564 3169 10604
rect 3255 10564 3276 10604
rect 3316 10564 3337 10604
rect 3423 10564 3440 10604
rect 3480 10564 3489 10604
rect 3103 10541 3169 10564
rect 3255 10541 3337 10564
rect 3423 10541 3489 10564
rect 3103 10522 3489 10541
rect 18223 10627 18609 10646
rect 18223 10604 18289 10627
rect 18375 10604 18457 10627
rect 18543 10604 18609 10627
rect 18223 10564 18232 10604
rect 18272 10564 18289 10604
rect 18375 10564 18396 10604
rect 18436 10564 18457 10604
rect 18543 10564 18560 10604
rect 18600 10564 18609 10604
rect 18223 10541 18289 10564
rect 18375 10541 18457 10564
rect 18543 10541 18609 10564
rect 18223 10522 18609 10541
rect 33343 10627 33729 10646
rect 33343 10604 33409 10627
rect 33495 10604 33577 10627
rect 33663 10604 33729 10627
rect 33343 10564 33352 10604
rect 33392 10564 33409 10604
rect 33495 10564 33516 10604
rect 33556 10564 33577 10604
rect 33663 10564 33680 10604
rect 33720 10564 33729 10604
rect 33343 10541 33409 10564
rect 33495 10541 33577 10564
rect 33663 10541 33729 10564
rect 33343 10522 33729 10541
rect 48463 10627 48849 10646
rect 48463 10604 48529 10627
rect 48615 10604 48697 10627
rect 48783 10604 48849 10627
rect 48463 10564 48472 10604
rect 48512 10564 48529 10604
rect 48615 10564 48636 10604
rect 48676 10564 48697 10604
rect 48783 10564 48800 10604
rect 48840 10564 48849 10604
rect 48463 10541 48529 10564
rect 48615 10541 48697 10564
rect 48783 10541 48849 10564
rect 48463 10522 48849 10541
rect 63583 10627 63969 10646
rect 63583 10604 63649 10627
rect 63735 10604 63817 10627
rect 63903 10604 63969 10627
rect 63583 10564 63592 10604
rect 63632 10564 63649 10604
rect 63735 10564 63756 10604
rect 63796 10564 63817 10604
rect 63903 10564 63920 10604
rect 63960 10564 63969 10604
rect 63583 10541 63649 10564
rect 63735 10541 63817 10564
rect 63903 10541 63969 10564
rect 63583 10522 63969 10541
rect 78703 10627 79089 10646
rect 78703 10604 78769 10627
rect 78855 10604 78937 10627
rect 79023 10604 79089 10627
rect 78703 10564 78712 10604
rect 78752 10564 78769 10604
rect 78855 10564 78876 10604
rect 78916 10564 78937 10604
rect 79023 10564 79040 10604
rect 79080 10564 79089 10604
rect 78703 10541 78769 10564
rect 78855 10541 78937 10564
rect 79023 10541 79089 10564
rect 78703 10522 79089 10541
rect 93823 10627 94209 10646
rect 93823 10604 93889 10627
rect 93975 10604 94057 10627
rect 94143 10604 94209 10627
rect 93823 10564 93832 10604
rect 93872 10564 93889 10604
rect 93975 10564 93996 10604
rect 94036 10564 94057 10604
rect 94143 10564 94160 10604
rect 94200 10564 94209 10604
rect 93823 10541 93889 10564
rect 93975 10541 94057 10564
rect 94143 10541 94209 10564
rect 93823 10522 94209 10541
rect 4343 9871 4729 9890
rect 4343 9848 4409 9871
rect 4495 9848 4577 9871
rect 4663 9848 4729 9871
rect 4343 9808 4352 9848
rect 4392 9808 4409 9848
rect 4495 9808 4516 9848
rect 4556 9808 4577 9848
rect 4663 9808 4680 9848
rect 4720 9808 4729 9848
rect 4343 9785 4409 9808
rect 4495 9785 4577 9808
rect 4663 9785 4729 9808
rect 4343 9766 4729 9785
rect 19463 9871 19849 9890
rect 19463 9848 19529 9871
rect 19615 9848 19697 9871
rect 19783 9848 19849 9871
rect 19463 9808 19472 9848
rect 19512 9808 19529 9848
rect 19615 9808 19636 9848
rect 19676 9808 19697 9848
rect 19783 9808 19800 9848
rect 19840 9808 19849 9848
rect 19463 9785 19529 9808
rect 19615 9785 19697 9808
rect 19783 9785 19849 9808
rect 19463 9766 19849 9785
rect 34583 9871 34969 9890
rect 34583 9848 34649 9871
rect 34735 9848 34817 9871
rect 34903 9848 34969 9871
rect 34583 9808 34592 9848
rect 34632 9808 34649 9848
rect 34735 9808 34756 9848
rect 34796 9808 34817 9848
rect 34903 9808 34920 9848
rect 34960 9808 34969 9848
rect 34583 9785 34649 9808
rect 34735 9785 34817 9808
rect 34903 9785 34969 9808
rect 34583 9766 34969 9785
rect 49703 9871 50089 9890
rect 49703 9848 49769 9871
rect 49855 9848 49937 9871
rect 50023 9848 50089 9871
rect 49703 9808 49712 9848
rect 49752 9808 49769 9848
rect 49855 9808 49876 9848
rect 49916 9808 49937 9848
rect 50023 9808 50040 9848
rect 50080 9808 50089 9848
rect 49703 9785 49769 9808
rect 49855 9785 49937 9808
rect 50023 9785 50089 9808
rect 49703 9766 50089 9785
rect 64823 9871 65209 9890
rect 64823 9848 64889 9871
rect 64975 9848 65057 9871
rect 65143 9848 65209 9871
rect 64823 9808 64832 9848
rect 64872 9808 64889 9848
rect 64975 9808 64996 9848
rect 65036 9808 65057 9848
rect 65143 9808 65160 9848
rect 65200 9808 65209 9848
rect 64823 9785 64889 9808
rect 64975 9785 65057 9808
rect 65143 9785 65209 9808
rect 64823 9766 65209 9785
rect 79943 9871 80329 9890
rect 79943 9848 80009 9871
rect 80095 9848 80177 9871
rect 80263 9848 80329 9871
rect 79943 9808 79952 9848
rect 79992 9808 80009 9848
rect 80095 9808 80116 9848
rect 80156 9808 80177 9848
rect 80263 9808 80280 9848
rect 80320 9808 80329 9848
rect 79943 9785 80009 9808
rect 80095 9785 80177 9808
rect 80263 9785 80329 9808
rect 79943 9766 80329 9785
rect 95063 9871 95449 9890
rect 95063 9848 95129 9871
rect 95215 9848 95297 9871
rect 95383 9848 95449 9871
rect 95063 9808 95072 9848
rect 95112 9808 95129 9848
rect 95215 9808 95236 9848
rect 95276 9808 95297 9848
rect 95383 9808 95400 9848
rect 95440 9808 95449 9848
rect 95063 9785 95129 9808
rect 95215 9785 95297 9808
rect 95383 9785 95449 9808
rect 95063 9766 95449 9785
rect 3103 9115 3489 9134
rect 3103 9092 3169 9115
rect 3255 9092 3337 9115
rect 3423 9092 3489 9115
rect 3103 9052 3112 9092
rect 3152 9052 3169 9092
rect 3255 9052 3276 9092
rect 3316 9052 3337 9092
rect 3423 9052 3440 9092
rect 3480 9052 3489 9092
rect 3103 9029 3169 9052
rect 3255 9029 3337 9052
rect 3423 9029 3489 9052
rect 3103 9010 3489 9029
rect 18223 9115 18609 9134
rect 18223 9092 18289 9115
rect 18375 9092 18457 9115
rect 18543 9092 18609 9115
rect 18223 9052 18232 9092
rect 18272 9052 18289 9092
rect 18375 9052 18396 9092
rect 18436 9052 18457 9092
rect 18543 9052 18560 9092
rect 18600 9052 18609 9092
rect 18223 9029 18289 9052
rect 18375 9029 18457 9052
rect 18543 9029 18609 9052
rect 18223 9010 18609 9029
rect 33343 9115 33729 9134
rect 33343 9092 33409 9115
rect 33495 9092 33577 9115
rect 33663 9092 33729 9115
rect 33343 9052 33352 9092
rect 33392 9052 33409 9092
rect 33495 9052 33516 9092
rect 33556 9052 33577 9092
rect 33663 9052 33680 9092
rect 33720 9052 33729 9092
rect 33343 9029 33409 9052
rect 33495 9029 33577 9052
rect 33663 9029 33729 9052
rect 33343 9010 33729 9029
rect 48463 9115 48849 9134
rect 48463 9092 48529 9115
rect 48615 9092 48697 9115
rect 48783 9092 48849 9115
rect 48463 9052 48472 9092
rect 48512 9052 48529 9092
rect 48615 9052 48636 9092
rect 48676 9052 48697 9092
rect 48783 9052 48800 9092
rect 48840 9052 48849 9092
rect 48463 9029 48529 9052
rect 48615 9029 48697 9052
rect 48783 9029 48849 9052
rect 48463 9010 48849 9029
rect 63583 9115 63969 9134
rect 63583 9092 63649 9115
rect 63735 9092 63817 9115
rect 63903 9092 63969 9115
rect 63583 9052 63592 9092
rect 63632 9052 63649 9092
rect 63735 9052 63756 9092
rect 63796 9052 63817 9092
rect 63903 9052 63920 9092
rect 63960 9052 63969 9092
rect 63583 9029 63649 9052
rect 63735 9029 63817 9052
rect 63903 9029 63969 9052
rect 63583 9010 63969 9029
rect 78703 9115 79089 9134
rect 78703 9092 78769 9115
rect 78855 9092 78937 9115
rect 79023 9092 79089 9115
rect 78703 9052 78712 9092
rect 78752 9052 78769 9092
rect 78855 9052 78876 9092
rect 78916 9052 78937 9092
rect 79023 9052 79040 9092
rect 79080 9052 79089 9092
rect 78703 9029 78769 9052
rect 78855 9029 78937 9052
rect 79023 9029 79089 9052
rect 78703 9010 79089 9029
rect 93823 9115 94209 9134
rect 93823 9092 93889 9115
rect 93975 9092 94057 9115
rect 94143 9092 94209 9115
rect 93823 9052 93832 9092
rect 93872 9052 93889 9092
rect 93975 9052 93996 9092
rect 94036 9052 94057 9092
rect 94143 9052 94160 9092
rect 94200 9052 94209 9092
rect 93823 9029 93889 9052
rect 93975 9029 94057 9052
rect 94143 9029 94209 9052
rect 93823 9010 94209 9029
rect 4343 8359 4729 8378
rect 4343 8336 4409 8359
rect 4495 8336 4577 8359
rect 4663 8336 4729 8359
rect 4343 8296 4352 8336
rect 4392 8296 4409 8336
rect 4495 8296 4516 8336
rect 4556 8296 4577 8336
rect 4663 8296 4680 8336
rect 4720 8296 4729 8336
rect 4343 8273 4409 8296
rect 4495 8273 4577 8296
rect 4663 8273 4729 8296
rect 4343 8254 4729 8273
rect 19463 8359 19849 8378
rect 19463 8336 19529 8359
rect 19615 8336 19697 8359
rect 19783 8336 19849 8359
rect 19463 8296 19472 8336
rect 19512 8296 19529 8336
rect 19615 8296 19636 8336
rect 19676 8296 19697 8336
rect 19783 8296 19800 8336
rect 19840 8296 19849 8336
rect 19463 8273 19529 8296
rect 19615 8273 19697 8296
rect 19783 8273 19849 8296
rect 19463 8254 19849 8273
rect 34583 8359 34969 8378
rect 34583 8336 34649 8359
rect 34735 8336 34817 8359
rect 34903 8336 34969 8359
rect 34583 8296 34592 8336
rect 34632 8296 34649 8336
rect 34735 8296 34756 8336
rect 34796 8296 34817 8336
rect 34903 8296 34920 8336
rect 34960 8296 34969 8336
rect 34583 8273 34649 8296
rect 34735 8273 34817 8296
rect 34903 8273 34969 8296
rect 34583 8254 34969 8273
rect 49703 8359 50089 8378
rect 49703 8336 49769 8359
rect 49855 8336 49937 8359
rect 50023 8336 50089 8359
rect 49703 8296 49712 8336
rect 49752 8296 49769 8336
rect 49855 8296 49876 8336
rect 49916 8296 49937 8336
rect 50023 8296 50040 8336
rect 50080 8296 50089 8336
rect 49703 8273 49769 8296
rect 49855 8273 49937 8296
rect 50023 8273 50089 8296
rect 49703 8254 50089 8273
rect 64823 8359 65209 8378
rect 64823 8336 64889 8359
rect 64975 8336 65057 8359
rect 65143 8336 65209 8359
rect 64823 8296 64832 8336
rect 64872 8296 64889 8336
rect 64975 8296 64996 8336
rect 65036 8296 65057 8336
rect 65143 8296 65160 8336
rect 65200 8296 65209 8336
rect 64823 8273 64889 8296
rect 64975 8273 65057 8296
rect 65143 8273 65209 8296
rect 64823 8254 65209 8273
rect 79943 8359 80329 8378
rect 79943 8336 80009 8359
rect 80095 8336 80177 8359
rect 80263 8336 80329 8359
rect 79943 8296 79952 8336
rect 79992 8296 80009 8336
rect 80095 8296 80116 8336
rect 80156 8296 80177 8336
rect 80263 8296 80280 8336
rect 80320 8296 80329 8336
rect 79943 8273 80009 8296
rect 80095 8273 80177 8296
rect 80263 8273 80329 8296
rect 79943 8254 80329 8273
rect 95063 8359 95449 8378
rect 95063 8336 95129 8359
rect 95215 8336 95297 8359
rect 95383 8336 95449 8359
rect 95063 8296 95072 8336
rect 95112 8296 95129 8336
rect 95215 8296 95236 8336
rect 95276 8296 95297 8336
rect 95383 8296 95400 8336
rect 95440 8296 95449 8336
rect 95063 8273 95129 8296
rect 95215 8273 95297 8296
rect 95383 8273 95449 8296
rect 95063 8254 95449 8273
rect 3103 7603 3489 7622
rect 3103 7580 3169 7603
rect 3255 7580 3337 7603
rect 3423 7580 3489 7603
rect 3103 7540 3112 7580
rect 3152 7540 3169 7580
rect 3255 7540 3276 7580
rect 3316 7540 3337 7580
rect 3423 7540 3440 7580
rect 3480 7540 3489 7580
rect 3103 7517 3169 7540
rect 3255 7517 3337 7540
rect 3423 7517 3489 7540
rect 3103 7498 3489 7517
rect 18223 7603 18609 7622
rect 18223 7580 18289 7603
rect 18375 7580 18457 7603
rect 18543 7580 18609 7603
rect 18223 7540 18232 7580
rect 18272 7540 18289 7580
rect 18375 7540 18396 7580
rect 18436 7540 18457 7580
rect 18543 7540 18560 7580
rect 18600 7540 18609 7580
rect 18223 7517 18289 7540
rect 18375 7517 18457 7540
rect 18543 7517 18609 7540
rect 18223 7498 18609 7517
rect 33343 7603 33729 7622
rect 33343 7580 33409 7603
rect 33495 7580 33577 7603
rect 33663 7580 33729 7603
rect 33343 7540 33352 7580
rect 33392 7540 33409 7580
rect 33495 7540 33516 7580
rect 33556 7540 33577 7580
rect 33663 7540 33680 7580
rect 33720 7540 33729 7580
rect 33343 7517 33409 7540
rect 33495 7517 33577 7540
rect 33663 7517 33729 7540
rect 33343 7498 33729 7517
rect 48463 7603 48849 7622
rect 48463 7580 48529 7603
rect 48615 7580 48697 7603
rect 48783 7580 48849 7603
rect 48463 7540 48472 7580
rect 48512 7540 48529 7580
rect 48615 7540 48636 7580
rect 48676 7540 48697 7580
rect 48783 7540 48800 7580
rect 48840 7540 48849 7580
rect 48463 7517 48529 7540
rect 48615 7517 48697 7540
rect 48783 7517 48849 7540
rect 48463 7498 48849 7517
rect 63583 7603 63969 7622
rect 63583 7580 63649 7603
rect 63735 7580 63817 7603
rect 63903 7580 63969 7603
rect 63583 7540 63592 7580
rect 63632 7540 63649 7580
rect 63735 7540 63756 7580
rect 63796 7540 63817 7580
rect 63903 7540 63920 7580
rect 63960 7540 63969 7580
rect 63583 7517 63649 7540
rect 63735 7517 63817 7540
rect 63903 7517 63969 7540
rect 63583 7498 63969 7517
rect 78703 7603 79089 7622
rect 78703 7580 78769 7603
rect 78855 7580 78937 7603
rect 79023 7580 79089 7603
rect 78703 7540 78712 7580
rect 78752 7540 78769 7580
rect 78855 7540 78876 7580
rect 78916 7540 78937 7580
rect 79023 7540 79040 7580
rect 79080 7540 79089 7580
rect 78703 7517 78769 7540
rect 78855 7517 78937 7540
rect 79023 7517 79089 7540
rect 78703 7498 79089 7517
rect 93823 7603 94209 7622
rect 93823 7580 93889 7603
rect 93975 7580 94057 7603
rect 94143 7580 94209 7603
rect 93823 7540 93832 7580
rect 93872 7540 93889 7580
rect 93975 7540 93996 7580
rect 94036 7540 94057 7580
rect 94143 7540 94160 7580
rect 94200 7540 94209 7580
rect 93823 7517 93889 7540
rect 93975 7517 94057 7540
rect 94143 7517 94209 7540
rect 93823 7498 94209 7517
rect 4343 6847 4729 6866
rect 4343 6824 4409 6847
rect 4495 6824 4577 6847
rect 4663 6824 4729 6847
rect 4343 6784 4352 6824
rect 4392 6784 4409 6824
rect 4495 6784 4516 6824
rect 4556 6784 4577 6824
rect 4663 6784 4680 6824
rect 4720 6784 4729 6824
rect 4343 6761 4409 6784
rect 4495 6761 4577 6784
rect 4663 6761 4729 6784
rect 4343 6742 4729 6761
rect 19463 6847 19849 6866
rect 19463 6824 19529 6847
rect 19615 6824 19697 6847
rect 19783 6824 19849 6847
rect 19463 6784 19472 6824
rect 19512 6784 19529 6824
rect 19615 6784 19636 6824
rect 19676 6784 19697 6824
rect 19783 6784 19800 6824
rect 19840 6784 19849 6824
rect 19463 6761 19529 6784
rect 19615 6761 19697 6784
rect 19783 6761 19849 6784
rect 19463 6742 19849 6761
rect 34583 6847 34969 6866
rect 34583 6824 34649 6847
rect 34735 6824 34817 6847
rect 34903 6824 34969 6847
rect 34583 6784 34592 6824
rect 34632 6784 34649 6824
rect 34735 6784 34756 6824
rect 34796 6784 34817 6824
rect 34903 6784 34920 6824
rect 34960 6784 34969 6824
rect 34583 6761 34649 6784
rect 34735 6761 34817 6784
rect 34903 6761 34969 6784
rect 34583 6742 34969 6761
rect 49703 6847 50089 6866
rect 49703 6824 49769 6847
rect 49855 6824 49937 6847
rect 50023 6824 50089 6847
rect 49703 6784 49712 6824
rect 49752 6784 49769 6824
rect 49855 6784 49876 6824
rect 49916 6784 49937 6824
rect 50023 6784 50040 6824
rect 50080 6784 50089 6824
rect 49703 6761 49769 6784
rect 49855 6761 49937 6784
rect 50023 6761 50089 6784
rect 49703 6742 50089 6761
rect 64823 6847 65209 6866
rect 64823 6824 64889 6847
rect 64975 6824 65057 6847
rect 65143 6824 65209 6847
rect 64823 6784 64832 6824
rect 64872 6784 64889 6824
rect 64975 6784 64996 6824
rect 65036 6784 65057 6824
rect 65143 6784 65160 6824
rect 65200 6784 65209 6824
rect 64823 6761 64889 6784
rect 64975 6761 65057 6784
rect 65143 6761 65209 6784
rect 64823 6742 65209 6761
rect 79943 6847 80329 6866
rect 79943 6824 80009 6847
rect 80095 6824 80177 6847
rect 80263 6824 80329 6847
rect 79943 6784 79952 6824
rect 79992 6784 80009 6824
rect 80095 6784 80116 6824
rect 80156 6784 80177 6824
rect 80263 6784 80280 6824
rect 80320 6784 80329 6824
rect 79943 6761 80009 6784
rect 80095 6761 80177 6784
rect 80263 6761 80329 6784
rect 79943 6742 80329 6761
rect 95063 6847 95449 6866
rect 95063 6824 95129 6847
rect 95215 6824 95297 6847
rect 95383 6824 95449 6847
rect 95063 6784 95072 6824
rect 95112 6784 95129 6824
rect 95215 6784 95236 6824
rect 95276 6784 95297 6824
rect 95383 6784 95400 6824
rect 95440 6784 95449 6824
rect 95063 6761 95129 6784
rect 95215 6761 95297 6784
rect 95383 6761 95449 6784
rect 95063 6742 95449 6761
rect 3103 6091 3489 6110
rect 3103 6068 3169 6091
rect 3255 6068 3337 6091
rect 3423 6068 3489 6091
rect 3103 6028 3112 6068
rect 3152 6028 3169 6068
rect 3255 6028 3276 6068
rect 3316 6028 3337 6068
rect 3423 6028 3440 6068
rect 3480 6028 3489 6068
rect 3103 6005 3169 6028
rect 3255 6005 3337 6028
rect 3423 6005 3489 6028
rect 3103 5986 3489 6005
rect 18223 6091 18609 6110
rect 18223 6068 18289 6091
rect 18375 6068 18457 6091
rect 18543 6068 18609 6091
rect 18223 6028 18232 6068
rect 18272 6028 18289 6068
rect 18375 6028 18396 6068
rect 18436 6028 18457 6068
rect 18543 6028 18560 6068
rect 18600 6028 18609 6068
rect 18223 6005 18289 6028
rect 18375 6005 18457 6028
rect 18543 6005 18609 6028
rect 18223 5986 18609 6005
rect 33343 6091 33729 6110
rect 33343 6068 33409 6091
rect 33495 6068 33577 6091
rect 33663 6068 33729 6091
rect 33343 6028 33352 6068
rect 33392 6028 33409 6068
rect 33495 6028 33516 6068
rect 33556 6028 33577 6068
rect 33663 6028 33680 6068
rect 33720 6028 33729 6068
rect 33343 6005 33409 6028
rect 33495 6005 33577 6028
rect 33663 6005 33729 6028
rect 33343 5986 33729 6005
rect 48463 6091 48849 6110
rect 48463 6068 48529 6091
rect 48615 6068 48697 6091
rect 48783 6068 48849 6091
rect 48463 6028 48472 6068
rect 48512 6028 48529 6068
rect 48615 6028 48636 6068
rect 48676 6028 48697 6068
rect 48783 6028 48800 6068
rect 48840 6028 48849 6068
rect 48463 6005 48529 6028
rect 48615 6005 48697 6028
rect 48783 6005 48849 6028
rect 48463 5986 48849 6005
rect 63583 6091 63969 6110
rect 63583 6068 63649 6091
rect 63735 6068 63817 6091
rect 63903 6068 63969 6091
rect 63583 6028 63592 6068
rect 63632 6028 63649 6068
rect 63735 6028 63756 6068
rect 63796 6028 63817 6068
rect 63903 6028 63920 6068
rect 63960 6028 63969 6068
rect 63583 6005 63649 6028
rect 63735 6005 63817 6028
rect 63903 6005 63969 6028
rect 63583 5986 63969 6005
rect 78703 6091 79089 6110
rect 78703 6068 78769 6091
rect 78855 6068 78937 6091
rect 79023 6068 79089 6091
rect 78703 6028 78712 6068
rect 78752 6028 78769 6068
rect 78855 6028 78876 6068
rect 78916 6028 78937 6068
rect 79023 6028 79040 6068
rect 79080 6028 79089 6068
rect 78703 6005 78769 6028
rect 78855 6005 78937 6028
rect 79023 6005 79089 6028
rect 78703 5986 79089 6005
rect 93823 6091 94209 6110
rect 93823 6068 93889 6091
rect 93975 6068 94057 6091
rect 94143 6068 94209 6091
rect 93823 6028 93832 6068
rect 93872 6028 93889 6068
rect 93975 6028 93996 6068
rect 94036 6028 94057 6068
rect 94143 6028 94160 6068
rect 94200 6028 94209 6068
rect 93823 6005 93889 6028
rect 93975 6005 94057 6028
rect 94143 6005 94209 6028
rect 93823 5986 94209 6005
rect 4343 5335 4729 5354
rect 4343 5312 4409 5335
rect 4495 5312 4577 5335
rect 4663 5312 4729 5335
rect 4343 5272 4352 5312
rect 4392 5272 4409 5312
rect 4495 5272 4516 5312
rect 4556 5272 4577 5312
rect 4663 5272 4680 5312
rect 4720 5272 4729 5312
rect 4343 5249 4409 5272
rect 4495 5249 4577 5272
rect 4663 5249 4729 5272
rect 4343 5230 4729 5249
rect 19463 5335 19849 5354
rect 19463 5312 19529 5335
rect 19615 5312 19697 5335
rect 19783 5312 19849 5335
rect 19463 5272 19472 5312
rect 19512 5272 19529 5312
rect 19615 5272 19636 5312
rect 19676 5272 19697 5312
rect 19783 5272 19800 5312
rect 19840 5272 19849 5312
rect 19463 5249 19529 5272
rect 19615 5249 19697 5272
rect 19783 5249 19849 5272
rect 19463 5230 19849 5249
rect 34583 5335 34969 5354
rect 34583 5312 34649 5335
rect 34735 5312 34817 5335
rect 34903 5312 34969 5335
rect 34583 5272 34592 5312
rect 34632 5272 34649 5312
rect 34735 5272 34756 5312
rect 34796 5272 34817 5312
rect 34903 5272 34920 5312
rect 34960 5272 34969 5312
rect 34583 5249 34649 5272
rect 34735 5249 34817 5272
rect 34903 5249 34969 5272
rect 34583 5230 34969 5249
rect 49703 5335 50089 5354
rect 49703 5312 49769 5335
rect 49855 5312 49937 5335
rect 50023 5312 50089 5335
rect 49703 5272 49712 5312
rect 49752 5272 49769 5312
rect 49855 5272 49876 5312
rect 49916 5272 49937 5312
rect 50023 5272 50040 5312
rect 50080 5272 50089 5312
rect 49703 5249 49769 5272
rect 49855 5249 49937 5272
rect 50023 5249 50089 5272
rect 49703 5230 50089 5249
rect 64823 5335 65209 5354
rect 64823 5312 64889 5335
rect 64975 5312 65057 5335
rect 65143 5312 65209 5335
rect 64823 5272 64832 5312
rect 64872 5272 64889 5312
rect 64975 5272 64996 5312
rect 65036 5272 65057 5312
rect 65143 5272 65160 5312
rect 65200 5272 65209 5312
rect 64823 5249 64889 5272
rect 64975 5249 65057 5272
rect 65143 5249 65209 5272
rect 64823 5230 65209 5249
rect 79943 5335 80329 5354
rect 79943 5312 80009 5335
rect 80095 5312 80177 5335
rect 80263 5312 80329 5335
rect 79943 5272 79952 5312
rect 79992 5272 80009 5312
rect 80095 5272 80116 5312
rect 80156 5272 80177 5312
rect 80263 5272 80280 5312
rect 80320 5272 80329 5312
rect 79943 5249 80009 5272
rect 80095 5249 80177 5272
rect 80263 5249 80329 5272
rect 79943 5230 80329 5249
rect 95063 5335 95449 5354
rect 95063 5312 95129 5335
rect 95215 5312 95297 5335
rect 95383 5312 95449 5335
rect 95063 5272 95072 5312
rect 95112 5272 95129 5312
rect 95215 5272 95236 5312
rect 95276 5272 95297 5312
rect 95383 5272 95400 5312
rect 95440 5272 95449 5312
rect 95063 5249 95129 5272
rect 95215 5249 95297 5272
rect 95383 5249 95449 5272
rect 95063 5230 95449 5249
rect 3103 4579 3489 4598
rect 3103 4556 3169 4579
rect 3255 4556 3337 4579
rect 3423 4556 3489 4579
rect 3103 4516 3112 4556
rect 3152 4516 3169 4556
rect 3255 4516 3276 4556
rect 3316 4516 3337 4556
rect 3423 4516 3440 4556
rect 3480 4516 3489 4556
rect 3103 4493 3169 4516
rect 3255 4493 3337 4516
rect 3423 4493 3489 4516
rect 3103 4474 3489 4493
rect 18223 4579 18609 4598
rect 18223 4556 18289 4579
rect 18375 4556 18457 4579
rect 18543 4556 18609 4579
rect 18223 4516 18232 4556
rect 18272 4516 18289 4556
rect 18375 4516 18396 4556
rect 18436 4516 18457 4556
rect 18543 4516 18560 4556
rect 18600 4516 18609 4556
rect 18223 4493 18289 4516
rect 18375 4493 18457 4516
rect 18543 4493 18609 4516
rect 18223 4474 18609 4493
rect 33343 4579 33729 4598
rect 33343 4556 33409 4579
rect 33495 4556 33577 4579
rect 33663 4556 33729 4579
rect 33343 4516 33352 4556
rect 33392 4516 33409 4556
rect 33495 4516 33516 4556
rect 33556 4516 33577 4556
rect 33663 4516 33680 4556
rect 33720 4516 33729 4556
rect 33343 4493 33409 4516
rect 33495 4493 33577 4516
rect 33663 4493 33729 4516
rect 33343 4474 33729 4493
rect 48463 4579 48849 4598
rect 48463 4556 48529 4579
rect 48615 4556 48697 4579
rect 48783 4556 48849 4579
rect 48463 4516 48472 4556
rect 48512 4516 48529 4556
rect 48615 4516 48636 4556
rect 48676 4516 48697 4556
rect 48783 4516 48800 4556
rect 48840 4516 48849 4556
rect 48463 4493 48529 4516
rect 48615 4493 48697 4516
rect 48783 4493 48849 4516
rect 48463 4474 48849 4493
rect 63583 4579 63969 4598
rect 63583 4556 63649 4579
rect 63735 4556 63817 4579
rect 63903 4556 63969 4579
rect 63583 4516 63592 4556
rect 63632 4516 63649 4556
rect 63735 4516 63756 4556
rect 63796 4516 63817 4556
rect 63903 4516 63920 4556
rect 63960 4516 63969 4556
rect 63583 4493 63649 4516
rect 63735 4493 63817 4516
rect 63903 4493 63969 4516
rect 63583 4474 63969 4493
rect 78703 4579 79089 4598
rect 78703 4556 78769 4579
rect 78855 4556 78937 4579
rect 79023 4556 79089 4579
rect 78703 4516 78712 4556
rect 78752 4516 78769 4556
rect 78855 4516 78876 4556
rect 78916 4516 78937 4556
rect 79023 4516 79040 4556
rect 79080 4516 79089 4556
rect 78703 4493 78769 4516
rect 78855 4493 78937 4516
rect 79023 4493 79089 4516
rect 78703 4474 79089 4493
rect 93823 4579 94209 4598
rect 93823 4556 93889 4579
rect 93975 4556 94057 4579
rect 94143 4556 94209 4579
rect 93823 4516 93832 4556
rect 93872 4516 93889 4556
rect 93975 4516 93996 4556
rect 94036 4516 94057 4556
rect 94143 4516 94160 4556
rect 94200 4516 94209 4556
rect 93823 4493 93889 4516
rect 93975 4493 94057 4516
rect 94143 4493 94209 4516
rect 93823 4474 94209 4493
rect 4343 3823 4729 3842
rect 4343 3800 4409 3823
rect 4495 3800 4577 3823
rect 4663 3800 4729 3823
rect 4343 3760 4352 3800
rect 4392 3760 4409 3800
rect 4495 3760 4516 3800
rect 4556 3760 4577 3800
rect 4663 3760 4680 3800
rect 4720 3760 4729 3800
rect 4343 3737 4409 3760
rect 4495 3737 4577 3760
rect 4663 3737 4729 3760
rect 4343 3718 4729 3737
rect 19463 3823 19849 3842
rect 19463 3800 19529 3823
rect 19615 3800 19697 3823
rect 19783 3800 19849 3823
rect 19463 3760 19472 3800
rect 19512 3760 19529 3800
rect 19615 3760 19636 3800
rect 19676 3760 19697 3800
rect 19783 3760 19800 3800
rect 19840 3760 19849 3800
rect 19463 3737 19529 3760
rect 19615 3737 19697 3760
rect 19783 3737 19849 3760
rect 19463 3718 19849 3737
rect 34583 3823 34969 3842
rect 34583 3800 34649 3823
rect 34735 3800 34817 3823
rect 34903 3800 34969 3823
rect 34583 3760 34592 3800
rect 34632 3760 34649 3800
rect 34735 3760 34756 3800
rect 34796 3760 34817 3800
rect 34903 3760 34920 3800
rect 34960 3760 34969 3800
rect 34583 3737 34649 3760
rect 34735 3737 34817 3760
rect 34903 3737 34969 3760
rect 34583 3718 34969 3737
rect 49703 3823 50089 3842
rect 49703 3800 49769 3823
rect 49855 3800 49937 3823
rect 50023 3800 50089 3823
rect 49703 3760 49712 3800
rect 49752 3760 49769 3800
rect 49855 3760 49876 3800
rect 49916 3760 49937 3800
rect 50023 3760 50040 3800
rect 50080 3760 50089 3800
rect 49703 3737 49769 3760
rect 49855 3737 49937 3760
rect 50023 3737 50089 3760
rect 49703 3718 50089 3737
rect 64823 3823 65209 3842
rect 64823 3800 64889 3823
rect 64975 3800 65057 3823
rect 65143 3800 65209 3823
rect 64823 3760 64832 3800
rect 64872 3760 64889 3800
rect 64975 3760 64996 3800
rect 65036 3760 65057 3800
rect 65143 3760 65160 3800
rect 65200 3760 65209 3800
rect 64823 3737 64889 3760
rect 64975 3737 65057 3760
rect 65143 3737 65209 3760
rect 64823 3718 65209 3737
rect 79943 3823 80329 3842
rect 79943 3800 80009 3823
rect 80095 3800 80177 3823
rect 80263 3800 80329 3823
rect 79943 3760 79952 3800
rect 79992 3760 80009 3800
rect 80095 3760 80116 3800
rect 80156 3760 80177 3800
rect 80263 3760 80280 3800
rect 80320 3760 80329 3800
rect 79943 3737 80009 3760
rect 80095 3737 80177 3760
rect 80263 3737 80329 3760
rect 79943 3718 80329 3737
rect 95063 3823 95449 3842
rect 95063 3800 95129 3823
rect 95215 3800 95297 3823
rect 95383 3800 95449 3823
rect 95063 3760 95072 3800
rect 95112 3760 95129 3800
rect 95215 3760 95236 3800
rect 95276 3760 95297 3800
rect 95383 3760 95400 3800
rect 95440 3760 95449 3800
rect 95063 3737 95129 3760
rect 95215 3737 95297 3760
rect 95383 3737 95449 3760
rect 95063 3718 95449 3737
rect 3103 3067 3489 3086
rect 3103 3044 3169 3067
rect 3255 3044 3337 3067
rect 3423 3044 3489 3067
rect 3103 3004 3112 3044
rect 3152 3004 3169 3044
rect 3255 3004 3276 3044
rect 3316 3004 3337 3044
rect 3423 3004 3440 3044
rect 3480 3004 3489 3044
rect 3103 2981 3169 3004
rect 3255 2981 3337 3004
rect 3423 2981 3489 3004
rect 3103 2962 3489 2981
rect 18223 3067 18609 3086
rect 18223 3044 18289 3067
rect 18375 3044 18457 3067
rect 18543 3044 18609 3067
rect 18223 3004 18232 3044
rect 18272 3004 18289 3044
rect 18375 3004 18396 3044
rect 18436 3004 18457 3044
rect 18543 3004 18560 3044
rect 18600 3004 18609 3044
rect 18223 2981 18289 3004
rect 18375 2981 18457 3004
rect 18543 2981 18609 3004
rect 18223 2962 18609 2981
rect 33343 3067 33729 3086
rect 33343 3044 33409 3067
rect 33495 3044 33577 3067
rect 33663 3044 33729 3067
rect 33343 3004 33352 3044
rect 33392 3004 33409 3044
rect 33495 3004 33516 3044
rect 33556 3004 33577 3044
rect 33663 3004 33680 3044
rect 33720 3004 33729 3044
rect 33343 2981 33409 3004
rect 33495 2981 33577 3004
rect 33663 2981 33729 3004
rect 33343 2962 33729 2981
rect 48463 3067 48849 3086
rect 48463 3044 48529 3067
rect 48615 3044 48697 3067
rect 48783 3044 48849 3067
rect 48463 3004 48472 3044
rect 48512 3004 48529 3044
rect 48615 3004 48636 3044
rect 48676 3004 48697 3044
rect 48783 3004 48800 3044
rect 48840 3004 48849 3044
rect 48463 2981 48529 3004
rect 48615 2981 48697 3004
rect 48783 2981 48849 3004
rect 48463 2962 48849 2981
rect 63583 3067 63969 3086
rect 63583 3044 63649 3067
rect 63735 3044 63817 3067
rect 63903 3044 63969 3067
rect 63583 3004 63592 3044
rect 63632 3004 63649 3044
rect 63735 3004 63756 3044
rect 63796 3004 63817 3044
rect 63903 3004 63920 3044
rect 63960 3004 63969 3044
rect 63583 2981 63649 3004
rect 63735 2981 63817 3004
rect 63903 2981 63969 3004
rect 63583 2962 63969 2981
rect 78703 3067 79089 3086
rect 78703 3044 78769 3067
rect 78855 3044 78937 3067
rect 79023 3044 79089 3067
rect 78703 3004 78712 3044
rect 78752 3004 78769 3044
rect 78855 3004 78876 3044
rect 78916 3004 78937 3044
rect 79023 3004 79040 3044
rect 79080 3004 79089 3044
rect 78703 2981 78769 3004
rect 78855 2981 78937 3004
rect 79023 2981 79089 3004
rect 78703 2962 79089 2981
rect 93823 3067 94209 3086
rect 93823 3044 93889 3067
rect 93975 3044 94057 3067
rect 94143 3044 94209 3067
rect 93823 3004 93832 3044
rect 93872 3004 93889 3044
rect 93975 3004 93996 3044
rect 94036 3004 94057 3044
rect 94143 3004 94160 3044
rect 94200 3004 94209 3044
rect 93823 2981 93889 3004
rect 93975 2981 94057 3004
rect 94143 2981 94209 3004
rect 93823 2962 94209 2981
rect 4343 2311 4729 2330
rect 4343 2288 4409 2311
rect 4495 2288 4577 2311
rect 4663 2288 4729 2311
rect 4343 2248 4352 2288
rect 4392 2248 4409 2288
rect 4495 2248 4516 2288
rect 4556 2248 4577 2288
rect 4663 2248 4680 2288
rect 4720 2248 4729 2288
rect 4343 2225 4409 2248
rect 4495 2225 4577 2248
rect 4663 2225 4729 2248
rect 4343 2206 4729 2225
rect 19463 2311 19849 2330
rect 19463 2288 19529 2311
rect 19615 2288 19697 2311
rect 19783 2288 19849 2311
rect 19463 2248 19472 2288
rect 19512 2248 19529 2288
rect 19615 2248 19636 2288
rect 19676 2248 19697 2288
rect 19783 2248 19800 2288
rect 19840 2248 19849 2288
rect 19463 2225 19529 2248
rect 19615 2225 19697 2248
rect 19783 2225 19849 2248
rect 19463 2206 19849 2225
rect 34583 2311 34969 2330
rect 34583 2288 34649 2311
rect 34735 2288 34817 2311
rect 34903 2288 34969 2311
rect 34583 2248 34592 2288
rect 34632 2248 34649 2288
rect 34735 2248 34756 2288
rect 34796 2248 34817 2288
rect 34903 2248 34920 2288
rect 34960 2248 34969 2288
rect 34583 2225 34649 2248
rect 34735 2225 34817 2248
rect 34903 2225 34969 2248
rect 34583 2206 34969 2225
rect 49703 2311 50089 2330
rect 49703 2288 49769 2311
rect 49855 2288 49937 2311
rect 50023 2288 50089 2311
rect 49703 2248 49712 2288
rect 49752 2248 49769 2288
rect 49855 2248 49876 2288
rect 49916 2248 49937 2288
rect 50023 2248 50040 2288
rect 50080 2248 50089 2288
rect 49703 2225 49769 2248
rect 49855 2225 49937 2248
rect 50023 2225 50089 2248
rect 49703 2206 50089 2225
rect 64823 2311 65209 2330
rect 64823 2288 64889 2311
rect 64975 2288 65057 2311
rect 65143 2288 65209 2311
rect 64823 2248 64832 2288
rect 64872 2248 64889 2288
rect 64975 2248 64996 2288
rect 65036 2248 65057 2288
rect 65143 2248 65160 2288
rect 65200 2248 65209 2288
rect 64823 2225 64889 2248
rect 64975 2225 65057 2248
rect 65143 2225 65209 2248
rect 64823 2206 65209 2225
rect 79943 2311 80329 2330
rect 79943 2288 80009 2311
rect 80095 2288 80177 2311
rect 80263 2288 80329 2311
rect 79943 2248 79952 2288
rect 79992 2248 80009 2288
rect 80095 2248 80116 2288
rect 80156 2248 80177 2288
rect 80263 2248 80280 2288
rect 80320 2248 80329 2288
rect 79943 2225 80009 2248
rect 80095 2225 80177 2248
rect 80263 2225 80329 2248
rect 79943 2206 80329 2225
rect 95063 2311 95449 2330
rect 95063 2288 95129 2311
rect 95215 2288 95297 2311
rect 95383 2288 95449 2311
rect 95063 2248 95072 2288
rect 95112 2248 95129 2288
rect 95215 2248 95236 2288
rect 95276 2248 95297 2288
rect 95383 2248 95400 2288
rect 95440 2248 95449 2288
rect 95063 2225 95129 2248
rect 95215 2225 95297 2248
rect 95383 2225 95449 2248
rect 95063 2206 95449 2225
rect 3103 1555 3489 1574
rect 3103 1532 3169 1555
rect 3255 1532 3337 1555
rect 3423 1532 3489 1555
rect 3103 1492 3112 1532
rect 3152 1492 3169 1532
rect 3255 1492 3276 1532
rect 3316 1492 3337 1532
rect 3423 1492 3440 1532
rect 3480 1492 3489 1532
rect 3103 1469 3169 1492
rect 3255 1469 3337 1492
rect 3423 1469 3489 1492
rect 3103 1450 3489 1469
rect 18223 1555 18609 1574
rect 18223 1532 18289 1555
rect 18375 1532 18457 1555
rect 18543 1532 18609 1555
rect 18223 1492 18232 1532
rect 18272 1492 18289 1532
rect 18375 1492 18396 1532
rect 18436 1492 18457 1532
rect 18543 1492 18560 1532
rect 18600 1492 18609 1532
rect 18223 1469 18289 1492
rect 18375 1469 18457 1492
rect 18543 1469 18609 1492
rect 18223 1450 18609 1469
rect 33343 1555 33729 1574
rect 33343 1532 33409 1555
rect 33495 1532 33577 1555
rect 33663 1532 33729 1555
rect 33343 1492 33352 1532
rect 33392 1492 33409 1532
rect 33495 1492 33516 1532
rect 33556 1492 33577 1532
rect 33663 1492 33680 1532
rect 33720 1492 33729 1532
rect 33343 1469 33409 1492
rect 33495 1469 33577 1492
rect 33663 1469 33729 1492
rect 33343 1450 33729 1469
rect 48463 1555 48849 1574
rect 48463 1532 48529 1555
rect 48615 1532 48697 1555
rect 48783 1532 48849 1555
rect 48463 1492 48472 1532
rect 48512 1492 48529 1532
rect 48615 1492 48636 1532
rect 48676 1492 48697 1532
rect 48783 1492 48800 1532
rect 48840 1492 48849 1532
rect 48463 1469 48529 1492
rect 48615 1469 48697 1492
rect 48783 1469 48849 1492
rect 48463 1450 48849 1469
rect 63583 1555 63969 1574
rect 63583 1532 63649 1555
rect 63735 1532 63817 1555
rect 63903 1532 63969 1555
rect 63583 1492 63592 1532
rect 63632 1492 63649 1532
rect 63735 1492 63756 1532
rect 63796 1492 63817 1532
rect 63903 1492 63920 1532
rect 63960 1492 63969 1532
rect 63583 1469 63649 1492
rect 63735 1469 63817 1492
rect 63903 1469 63969 1492
rect 63583 1450 63969 1469
rect 78703 1555 79089 1574
rect 78703 1532 78769 1555
rect 78855 1532 78937 1555
rect 79023 1532 79089 1555
rect 78703 1492 78712 1532
rect 78752 1492 78769 1532
rect 78855 1492 78876 1532
rect 78916 1492 78937 1532
rect 79023 1492 79040 1532
rect 79080 1492 79089 1532
rect 78703 1469 78769 1492
rect 78855 1469 78937 1492
rect 79023 1469 79089 1492
rect 78703 1450 79089 1469
rect 93823 1555 94209 1574
rect 93823 1532 93889 1555
rect 93975 1532 94057 1555
rect 94143 1532 94209 1555
rect 93823 1492 93832 1532
rect 93872 1492 93889 1532
rect 93975 1492 93996 1532
rect 94036 1492 94057 1532
rect 94143 1492 94160 1532
rect 94200 1492 94209 1532
rect 93823 1469 93889 1492
rect 93975 1469 94057 1492
rect 94143 1469 94209 1492
rect 93823 1450 94209 1469
rect 4343 799 4729 818
rect 4343 776 4409 799
rect 4495 776 4577 799
rect 4663 776 4729 799
rect 4343 736 4352 776
rect 4392 736 4409 776
rect 4495 736 4516 776
rect 4556 736 4577 776
rect 4663 736 4680 776
rect 4720 736 4729 776
rect 4343 713 4409 736
rect 4495 713 4577 736
rect 4663 713 4729 736
rect 4343 694 4729 713
rect 19463 799 19849 818
rect 19463 776 19529 799
rect 19615 776 19697 799
rect 19783 776 19849 799
rect 19463 736 19472 776
rect 19512 736 19529 776
rect 19615 736 19636 776
rect 19676 736 19697 776
rect 19783 736 19800 776
rect 19840 736 19849 776
rect 19463 713 19529 736
rect 19615 713 19697 736
rect 19783 713 19849 736
rect 19463 694 19849 713
rect 34583 799 34969 818
rect 34583 776 34649 799
rect 34735 776 34817 799
rect 34903 776 34969 799
rect 34583 736 34592 776
rect 34632 736 34649 776
rect 34735 736 34756 776
rect 34796 736 34817 776
rect 34903 736 34920 776
rect 34960 736 34969 776
rect 34583 713 34649 736
rect 34735 713 34817 736
rect 34903 713 34969 736
rect 34583 694 34969 713
rect 49703 799 50089 818
rect 49703 776 49769 799
rect 49855 776 49937 799
rect 50023 776 50089 799
rect 49703 736 49712 776
rect 49752 736 49769 776
rect 49855 736 49876 776
rect 49916 736 49937 776
rect 50023 736 50040 776
rect 50080 736 50089 776
rect 49703 713 49769 736
rect 49855 713 49937 736
rect 50023 713 50089 736
rect 49703 694 50089 713
rect 64823 799 65209 818
rect 64823 776 64889 799
rect 64975 776 65057 799
rect 65143 776 65209 799
rect 64823 736 64832 776
rect 64872 736 64889 776
rect 64975 736 64996 776
rect 65036 736 65057 776
rect 65143 736 65160 776
rect 65200 736 65209 776
rect 64823 713 64889 736
rect 64975 713 65057 736
rect 65143 713 65209 736
rect 64823 694 65209 713
rect 79943 799 80329 818
rect 79943 776 80009 799
rect 80095 776 80177 799
rect 80263 776 80329 799
rect 79943 736 79952 776
rect 79992 736 80009 776
rect 80095 736 80116 776
rect 80156 736 80177 776
rect 80263 736 80280 776
rect 80320 736 80329 776
rect 79943 713 80009 736
rect 80095 713 80177 736
rect 80263 713 80329 736
rect 79943 694 80329 713
rect 95063 799 95449 818
rect 95063 776 95129 799
rect 95215 776 95297 799
rect 95383 776 95449 799
rect 95063 736 95072 776
rect 95112 736 95129 776
rect 95215 736 95236 776
rect 95276 736 95297 776
rect 95383 736 95400 776
rect 95440 736 95449 776
rect 95063 713 95129 736
rect 95215 713 95297 736
rect 95383 713 95449 736
rect 95063 694 95449 713
<< via5 >>
rect 4409 38576 4495 38599
rect 4577 38576 4663 38599
rect 4409 38536 4434 38576
rect 4434 38536 4474 38576
rect 4474 38536 4495 38576
rect 4577 38536 4598 38576
rect 4598 38536 4638 38576
rect 4638 38536 4663 38576
rect 4409 38513 4495 38536
rect 4577 38513 4663 38536
rect 19529 38576 19615 38599
rect 19697 38576 19783 38599
rect 19529 38536 19554 38576
rect 19554 38536 19594 38576
rect 19594 38536 19615 38576
rect 19697 38536 19718 38576
rect 19718 38536 19758 38576
rect 19758 38536 19783 38576
rect 19529 38513 19615 38536
rect 19697 38513 19783 38536
rect 34649 38576 34735 38599
rect 34817 38576 34903 38599
rect 34649 38536 34674 38576
rect 34674 38536 34714 38576
rect 34714 38536 34735 38576
rect 34817 38536 34838 38576
rect 34838 38536 34878 38576
rect 34878 38536 34903 38576
rect 34649 38513 34735 38536
rect 34817 38513 34903 38536
rect 49769 38576 49855 38599
rect 49937 38576 50023 38599
rect 49769 38536 49794 38576
rect 49794 38536 49834 38576
rect 49834 38536 49855 38576
rect 49937 38536 49958 38576
rect 49958 38536 49998 38576
rect 49998 38536 50023 38576
rect 49769 38513 49855 38536
rect 49937 38513 50023 38536
rect 64889 38576 64975 38599
rect 65057 38576 65143 38599
rect 64889 38536 64914 38576
rect 64914 38536 64954 38576
rect 64954 38536 64975 38576
rect 65057 38536 65078 38576
rect 65078 38536 65118 38576
rect 65118 38536 65143 38576
rect 64889 38513 64975 38536
rect 65057 38513 65143 38536
rect 80009 38576 80095 38599
rect 80177 38576 80263 38599
rect 80009 38536 80034 38576
rect 80034 38536 80074 38576
rect 80074 38536 80095 38576
rect 80177 38536 80198 38576
rect 80198 38536 80238 38576
rect 80238 38536 80263 38576
rect 80009 38513 80095 38536
rect 80177 38513 80263 38536
rect 95129 38576 95215 38599
rect 95297 38576 95383 38599
rect 95129 38536 95154 38576
rect 95154 38536 95194 38576
rect 95194 38536 95215 38576
rect 95297 38536 95318 38576
rect 95318 38536 95358 38576
rect 95358 38536 95383 38576
rect 95129 38513 95215 38536
rect 95297 38513 95383 38536
rect 3169 37820 3255 37843
rect 3337 37820 3423 37843
rect 3169 37780 3194 37820
rect 3194 37780 3234 37820
rect 3234 37780 3255 37820
rect 3337 37780 3358 37820
rect 3358 37780 3398 37820
rect 3398 37780 3423 37820
rect 3169 37757 3255 37780
rect 3337 37757 3423 37780
rect 18289 37820 18375 37843
rect 18457 37820 18543 37843
rect 18289 37780 18314 37820
rect 18314 37780 18354 37820
rect 18354 37780 18375 37820
rect 18457 37780 18478 37820
rect 18478 37780 18518 37820
rect 18518 37780 18543 37820
rect 18289 37757 18375 37780
rect 18457 37757 18543 37780
rect 33409 37820 33495 37843
rect 33577 37820 33663 37843
rect 33409 37780 33434 37820
rect 33434 37780 33474 37820
rect 33474 37780 33495 37820
rect 33577 37780 33598 37820
rect 33598 37780 33638 37820
rect 33638 37780 33663 37820
rect 33409 37757 33495 37780
rect 33577 37757 33663 37780
rect 48529 37820 48615 37843
rect 48697 37820 48783 37843
rect 48529 37780 48554 37820
rect 48554 37780 48594 37820
rect 48594 37780 48615 37820
rect 48697 37780 48718 37820
rect 48718 37780 48758 37820
rect 48758 37780 48783 37820
rect 48529 37757 48615 37780
rect 48697 37757 48783 37780
rect 63649 37820 63735 37843
rect 63817 37820 63903 37843
rect 63649 37780 63674 37820
rect 63674 37780 63714 37820
rect 63714 37780 63735 37820
rect 63817 37780 63838 37820
rect 63838 37780 63878 37820
rect 63878 37780 63903 37820
rect 63649 37757 63735 37780
rect 63817 37757 63903 37780
rect 78769 37820 78855 37843
rect 78937 37820 79023 37843
rect 78769 37780 78794 37820
rect 78794 37780 78834 37820
rect 78834 37780 78855 37820
rect 78937 37780 78958 37820
rect 78958 37780 78998 37820
rect 78998 37780 79023 37820
rect 78769 37757 78855 37780
rect 78937 37757 79023 37780
rect 93889 37820 93975 37843
rect 94057 37820 94143 37843
rect 93889 37780 93914 37820
rect 93914 37780 93954 37820
rect 93954 37780 93975 37820
rect 94057 37780 94078 37820
rect 94078 37780 94118 37820
rect 94118 37780 94143 37820
rect 93889 37757 93975 37780
rect 94057 37757 94143 37780
rect 4409 37064 4495 37087
rect 4577 37064 4663 37087
rect 4409 37024 4434 37064
rect 4434 37024 4474 37064
rect 4474 37024 4495 37064
rect 4577 37024 4598 37064
rect 4598 37024 4638 37064
rect 4638 37024 4663 37064
rect 4409 37001 4495 37024
rect 4577 37001 4663 37024
rect 19529 37064 19615 37087
rect 19697 37064 19783 37087
rect 19529 37024 19554 37064
rect 19554 37024 19594 37064
rect 19594 37024 19615 37064
rect 19697 37024 19718 37064
rect 19718 37024 19758 37064
rect 19758 37024 19783 37064
rect 19529 37001 19615 37024
rect 19697 37001 19783 37024
rect 34649 37064 34735 37087
rect 34817 37064 34903 37087
rect 34649 37024 34674 37064
rect 34674 37024 34714 37064
rect 34714 37024 34735 37064
rect 34817 37024 34838 37064
rect 34838 37024 34878 37064
rect 34878 37024 34903 37064
rect 34649 37001 34735 37024
rect 34817 37001 34903 37024
rect 49769 37064 49855 37087
rect 49937 37064 50023 37087
rect 49769 37024 49794 37064
rect 49794 37024 49834 37064
rect 49834 37024 49855 37064
rect 49937 37024 49958 37064
rect 49958 37024 49998 37064
rect 49998 37024 50023 37064
rect 49769 37001 49855 37024
rect 49937 37001 50023 37024
rect 64889 37064 64975 37087
rect 65057 37064 65143 37087
rect 64889 37024 64914 37064
rect 64914 37024 64954 37064
rect 64954 37024 64975 37064
rect 65057 37024 65078 37064
rect 65078 37024 65118 37064
rect 65118 37024 65143 37064
rect 64889 37001 64975 37024
rect 65057 37001 65143 37024
rect 80009 37064 80095 37087
rect 80177 37064 80263 37087
rect 80009 37024 80034 37064
rect 80034 37024 80074 37064
rect 80074 37024 80095 37064
rect 80177 37024 80198 37064
rect 80198 37024 80238 37064
rect 80238 37024 80263 37064
rect 80009 37001 80095 37024
rect 80177 37001 80263 37024
rect 95129 37064 95215 37087
rect 95297 37064 95383 37087
rect 95129 37024 95154 37064
rect 95154 37024 95194 37064
rect 95194 37024 95215 37064
rect 95297 37024 95318 37064
rect 95318 37024 95358 37064
rect 95358 37024 95383 37064
rect 95129 37001 95215 37024
rect 95297 37001 95383 37024
rect 3169 36308 3255 36331
rect 3337 36308 3423 36331
rect 3169 36268 3194 36308
rect 3194 36268 3234 36308
rect 3234 36268 3255 36308
rect 3337 36268 3358 36308
rect 3358 36268 3398 36308
rect 3398 36268 3423 36308
rect 3169 36245 3255 36268
rect 3337 36245 3423 36268
rect 18289 36308 18375 36331
rect 18457 36308 18543 36331
rect 18289 36268 18314 36308
rect 18314 36268 18354 36308
rect 18354 36268 18375 36308
rect 18457 36268 18478 36308
rect 18478 36268 18518 36308
rect 18518 36268 18543 36308
rect 18289 36245 18375 36268
rect 18457 36245 18543 36268
rect 33409 36308 33495 36331
rect 33577 36308 33663 36331
rect 33409 36268 33434 36308
rect 33434 36268 33474 36308
rect 33474 36268 33495 36308
rect 33577 36268 33598 36308
rect 33598 36268 33638 36308
rect 33638 36268 33663 36308
rect 33409 36245 33495 36268
rect 33577 36245 33663 36268
rect 48529 36308 48615 36331
rect 48697 36308 48783 36331
rect 48529 36268 48554 36308
rect 48554 36268 48594 36308
rect 48594 36268 48615 36308
rect 48697 36268 48718 36308
rect 48718 36268 48758 36308
rect 48758 36268 48783 36308
rect 48529 36245 48615 36268
rect 48697 36245 48783 36268
rect 63649 36308 63735 36331
rect 63817 36308 63903 36331
rect 63649 36268 63674 36308
rect 63674 36268 63714 36308
rect 63714 36268 63735 36308
rect 63817 36268 63838 36308
rect 63838 36268 63878 36308
rect 63878 36268 63903 36308
rect 63649 36245 63735 36268
rect 63817 36245 63903 36268
rect 78769 36308 78855 36331
rect 78937 36308 79023 36331
rect 78769 36268 78794 36308
rect 78794 36268 78834 36308
rect 78834 36268 78855 36308
rect 78937 36268 78958 36308
rect 78958 36268 78998 36308
rect 78998 36268 79023 36308
rect 78769 36245 78855 36268
rect 78937 36245 79023 36268
rect 93889 36308 93975 36331
rect 94057 36308 94143 36331
rect 93889 36268 93914 36308
rect 93914 36268 93954 36308
rect 93954 36268 93975 36308
rect 94057 36268 94078 36308
rect 94078 36268 94118 36308
rect 94118 36268 94143 36308
rect 93889 36245 93975 36268
rect 94057 36245 94143 36268
rect 4409 35552 4495 35575
rect 4577 35552 4663 35575
rect 4409 35512 4434 35552
rect 4434 35512 4474 35552
rect 4474 35512 4495 35552
rect 4577 35512 4598 35552
rect 4598 35512 4638 35552
rect 4638 35512 4663 35552
rect 4409 35489 4495 35512
rect 4577 35489 4663 35512
rect 19529 35552 19615 35575
rect 19697 35552 19783 35575
rect 19529 35512 19554 35552
rect 19554 35512 19594 35552
rect 19594 35512 19615 35552
rect 19697 35512 19718 35552
rect 19718 35512 19758 35552
rect 19758 35512 19783 35552
rect 19529 35489 19615 35512
rect 19697 35489 19783 35512
rect 34649 35552 34735 35575
rect 34817 35552 34903 35575
rect 34649 35512 34674 35552
rect 34674 35512 34714 35552
rect 34714 35512 34735 35552
rect 34817 35512 34838 35552
rect 34838 35512 34878 35552
rect 34878 35512 34903 35552
rect 34649 35489 34735 35512
rect 34817 35489 34903 35512
rect 49769 35552 49855 35575
rect 49937 35552 50023 35575
rect 49769 35512 49794 35552
rect 49794 35512 49834 35552
rect 49834 35512 49855 35552
rect 49937 35512 49958 35552
rect 49958 35512 49998 35552
rect 49998 35512 50023 35552
rect 49769 35489 49855 35512
rect 49937 35489 50023 35512
rect 64889 35552 64975 35575
rect 65057 35552 65143 35575
rect 64889 35512 64914 35552
rect 64914 35512 64954 35552
rect 64954 35512 64975 35552
rect 65057 35512 65078 35552
rect 65078 35512 65118 35552
rect 65118 35512 65143 35552
rect 64889 35489 64975 35512
rect 65057 35489 65143 35512
rect 80009 35552 80095 35575
rect 80177 35552 80263 35575
rect 80009 35512 80034 35552
rect 80034 35512 80074 35552
rect 80074 35512 80095 35552
rect 80177 35512 80198 35552
rect 80198 35512 80238 35552
rect 80238 35512 80263 35552
rect 80009 35489 80095 35512
rect 80177 35489 80263 35512
rect 95129 35552 95215 35575
rect 95297 35552 95383 35575
rect 95129 35512 95154 35552
rect 95154 35512 95194 35552
rect 95194 35512 95215 35552
rect 95297 35512 95318 35552
rect 95318 35512 95358 35552
rect 95358 35512 95383 35552
rect 95129 35489 95215 35512
rect 95297 35489 95383 35512
rect 3169 34796 3255 34819
rect 3337 34796 3423 34819
rect 3169 34756 3194 34796
rect 3194 34756 3234 34796
rect 3234 34756 3255 34796
rect 3337 34756 3358 34796
rect 3358 34756 3398 34796
rect 3398 34756 3423 34796
rect 3169 34733 3255 34756
rect 3337 34733 3423 34756
rect 18289 34796 18375 34819
rect 18457 34796 18543 34819
rect 18289 34756 18314 34796
rect 18314 34756 18354 34796
rect 18354 34756 18375 34796
rect 18457 34756 18478 34796
rect 18478 34756 18518 34796
rect 18518 34756 18543 34796
rect 18289 34733 18375 34756
rect 18457 34733 18543 34756
rect 33409 34796 33495 34819
rect 33577 34796 33663 34819
rect 33409 34756 33434 34796
rect 33434 34756 33474 34796
rect 33474 34756 33495 34796
rect 33577 34756 33598 34796
rect 33598 34756 33638 34796
rect 33638 34756 33663 34796
rect 33409 34733 33495 34756
rect 33577 34733 33663 34756
rect 48529 34796 48615 34819
rect 48697 34796 48783 34819
rect 48529 34756 48554 34796
rect 48554 34756 48594 34796
rect 48594 34756 48615 34796
rect 48697 34756 48718 34796
rect 48718 34756 48758 34796
rect 48758 34756 48783 34796
rect 48529 34733 48615 34756
rect 48697 34733 48783 34756
rect 63649 34796 63735 34819
rect 63817 34796 63903 34819
rect 63649 34756 63674 34796
rect 63674 34756 63714 34796
rect 63714 34756 63735 34796
rect 63817 34756 63838 34796
rect 63838 34756 63878 34796
rect 63878 34756 63903 34796
rect 63649 34733 63735 34756
rect 63817 34733 63903 34756
rect 78769 34796 78855 34819
rect 78937 34796 79023 34819
rect 78769 34756 78794 34796
rect 78794 34756 78834 34796
rect 78834 34756 78855 34796
rect 78937 34756 78958 34796
rect 78958 34756 78998 34796
rect 78998 34756 79023 34796
rect 78769 34733 78855 34756
rect 78937 34733 79023 34756
rect 93889 34796 93975 34819
rect 94057 34796 94143 34819
rect 93889 34756 93914 34796
rect 93914 34756 93954 34796
rect 93954 34756 93975 34796
rect 94057 34756 94078 34796
rect 94078 34756 94118 34796
rect 94118 34756 94143 34796
rect 93889 34733 93975 34756
rect 94057 34733 94143 34756
rect 4409 34040 4495 34063
rect 4577 34040 4663 34063
rect 4409 34000 4434 34040
rect 4434 34000 4474 34040
rect 4474 34000 4495 34040
rect 4577 34000 4598 34040
rect 4598 34000 4638 34040
rect 4638 34000 4663 34040
rect 4409 33977 4495 34000
rect 4577 33977 4663 34000
rect 19529 34040 19615 34063
rect 19697 34040 19783 34063
rect 19529 34000 19554 34040
rect 19554 34000 19594 34040
rect 19594 34000 19615 34040
rect 19697 34000 19718 34040
rect 19718 34000 19758 34040
rect 19758 34000 19783 34040
rect 19529 33977 19615 34000
rect 19697 33977 19783 34000
rect 34649 34040 34735 34063
rect 34817 34040 34903 34063
rect 34649 34000 34674 34040
rect 34674 34000 34714 34040
rect 34714 34000 34735 34040
rect 34817 34000 34838 34040
rect 34838 34000 34878 34040
rect 34878 34000 34903 34040
rect 34649 33977 34735 34000
rect 34817 33977 34903 34000
rect 49769 34040 49855 34063
rect 49937 34040 50023 34063
rect 49769 34000 49794 34040
rect 49794 34000 49834 34040
rect 49834 34000 49855 34040
rect 49937 34000 49958 34040
rect 49958 34000 49998 34040
rect 49998 34000 50023 34040
rect 49769 33977 49855 34000
rect 49937 33977 50023 34000
rect 64889 34040 64975 34063
rect 65057 34040 65143 34063
rect 64889 34000 64914 34040
rect 64914 34000 64954 34040
rect 64954 34000 64975 34040
rect 65057 34000 65078 34040
rect 65078 34000 65118 34040
rect 65118 34000 65143 34040
rect 64889 33977 64975 34000
rect 65057 33977 65143 34000
rect 80009 34040 80095 34063
rect 80177 34040 80263 34063
rect 80009 34000 80034 34040
rect 80034 34000 80074 34040
rect 80074 34000 80095 34040
rect 80177 34000 80198 34040
rect 80198 34000 80238 34040
rect 80238 34000 80263 34040
rect 80009 33977 80095 34000
rect 80177 33977 80263 34000
rect 95129 34040 95215 34063
rect 95297 34040 95383 34063
rect 95129 34000 95154 34040
rect 95154 34000 95194 34040
rect 95194 34000 95215 34040
rect 95297 34000 95318 34040
rect 95318 34000 95358 34040
rect 95358 34000 95383 34040
rect 95129 33977 95215 34000
rect 95297 33977 95383 34000
rect 3169 33284 3255 33307
rect 3337 33284 3423 33307
rect 3169 33244 3194 33284
rect 3194 33244 3234 33284
rect 3234 33244 3255 33284
rect 3337 33244 3358 33284
rect 3358 33244 3398 33284
rect 3398 33244 3423 33284
rect 3169 33221 3255 33244
rect 3337 33221 3423 33244
rect 18289 33284 18375 33307
rect 18457 33284 18543 33307
rect 18289 33244 18314 33284
rect 18314 33244 18354 33284
rect 18354 33244 18375 33284
rect 18457 33244 18478 33284
rect 18478 33244 18518 33284
rect 18518 33244 18543 33284
rect 18289 33221 18375 33244
rect 18457 33221 18543 33244
rect 33409 33284 33495 33307
rect 33577 33284 33663 33307
rect 33409 33244 33434 33284
rect 33434 33244 33474 33284
rect 33474 33244 33495 33284
rect 33577 33244 33598 33284
rect 33598 33244 33638 33284
rect 33638 33244 33663 33284
rect 33409 33221 33495 33244
rect 33577 33221 33663 33244
rect 48529 33284 48615 33307
rect 48697 33284 48783 33307
rect 48529 33244 48554 33284
rect 48554 33244 48594 33284
rect 48594 33244 48615 33284
rect 48697 33244 48718 33284
rect 48718 33244 48758 33284
rect 48758 33244 48783 33284
rect 48529 33221 48615 33244
rect 48697 33221 48783 33244
rect 63649 33284 63735 33307
rect 63817 33284 63903 33307
rect 63649 33244 63674 33284
rect 63674 33244 63714 33284
rect 63714 33244 63735 33284
rect 63817 33244 63838 33284
rect 63838 33244 63878 33284
rect 63878 33244 63903 33284
rect 63649 33221 63735 33244
rect 63817 33221 63903 33244
rect 78769 33284 78855 33307
rect 78937 33284 79023 33307
rect 78769 33244 78794 33284
rect 78794 33244 78834 33284
rect 78834 33244 78855 33284
rect 78937 33244 78958 33284
rect 78958 33244 78998 33284
rect 78998 33244 79023 33284
rect 78769 33221 78855 33244
rect 78937 33221 79023 33244
rect 93889 33284 93975 33307
rect 94057 33284 94143 33307
rect 93889 33244 93914 33284
rect 93914 33244 93954 33284
rect 93954 33244 93975 33284
rect 94057 33244 94078 33284
rect 94078 33244 94118 33284
rect 94118 33244 94143 33284
rect 93889 33221 93975 33244
rect 94057 33221 94143 33244
rect 4409 32528 4495 32551
rect 4577 32528 4663 32551
rect 4409 32488 4434 32528
rect 4434 32488 4474 32528
rect 4474 32488 4495 32528
rect 4577 32488 4598 32528
rect 4598 32488 4638 32528
rect 4638 32488 4663 32528
rect 4409 32465 4495 32488
rect 4577 32465 4663 32488
rect 19529 32528 19615 32551
rect 19697 32528 19783 32551
rect 19529 32488 19554 32528
rect 19554 32488 19594 32528
rect 19594 32488 19615 32528
rect 19697 32488 19718 32528
rect 19718 32488 19758 32528
rect 19758 32488 19783 32528
rect 19529 32465 19615 32488
rect 19697 32465 19783 32488
rect 34649 32528 34735 32551
rect 34817 32528 34903 32551
rect 34649 32488 34674 32528
rect 34674 32488 34714 32528
rect 34714 32488 34735 32528
rect 34817 32488 34838 32528
rect 34838 32488 34878 32528
rect 34878 32488 34903 32528
rect 34649 32465 34735 32488
rect 34817 32465 34903 32488
rect 49769 32528 49855 32551
rect 49937 32528 50023 32551
rect 49769 32488 49794 32528
rect 49794 32488 49834 32528
rect 49834 32488 49855 32528
rect 49937 32488 49958 32528
rect 49958 32488 49998 32528
rect 49998 32488 50023 32528
rect 49769 32465 49855 32488
rect 49937 32465 50023 32488
rect 64889 32528 64975 32551
rect 65057 32528 65143 32551
rect 64889 32488 64914 32528
rect 64914 32488 64954 32528
rect 64954 32488 64975 32528
rect 65057 32488 65078 32528
rect 65078 32488 65118 32528
rect 65118 32488 65143 32528
rect 64889 32465 64975 32488
rect 65057 32465 65143 32488
rect 80009 32528 80095 32551
rect 80177 32528 80263 32551
rect 80009 32488 80034 32528
rect 80034 32488 80074 32528
rect 80074 32488 80095 32528
rect 80177 32488 80198 32528
rect 80198 32488 80238 32528
rect 80238 32488 80263 32528
rect 80009 32465 80095 32488
rect 80177 32465 80263 32488
rect 95129 32528 95215 32551
rect 95297 32528 95383 32551
rect 95129 32488 95154 32528
rect 95154 32488 95194 32528
rect 95194 32488 95215 32528
rect 95297 32488 95318 32528
rect 95318 32488 95358 32528
rect 95358 32488 95383 32528
rect 95129 32465 95215 32488
rect 95297 32465 95383 32488
rect 3169 31772 3255 31795
rect 3337 31772 3423 31795
rect 3169 31732 3194 31772
rect 3194 31732 3234 31772
rect 3234 31732 3255 31772
rect 3337 31732 3358 31772
rect 3358 31732 3398 31772
rect 3398 31732 3423 31772
rect 3169 31709 3255 31732
rect 3337 31709 3423 31732
rect 18289 31772 18375 31795
rect 18457 31772 18543 31795
rect 18289 31732 18314 31772
rect 18314 31732 18354 31772
rect 18354 31732 18375 31772
rect 18457 31732 18478 31772
rect 18478 31732 18518 31772
rect 18518 31732 18543 31772
rect 18289 31709 18375 31732
rect 18457 31709 18543 31732
rect 33409 31772 33495 31795
rect 33577 31772 33663 31795
rect 33409 31732 33434 31772
rect 33434 31732 33474 31772
rect 33474 31732 33495 31772
rect 33577 31732 33598 31772
rect 33598 31732 33638 31772
rect 33638 31732 33663 31772
rect 33409 31709 33495 31732
rect 33577 31709 33663 31732
rect 48529 31772 48615 31795
rect 48697 31772 48783 31795
rect 48529 31732 48554 31772
rect 48554 31732 48594 31772
rect 48594 31732 48615 31772
rect 48697 31732 48718 31772
rect 48718 31732 48758 31772
rect 48758 31732 48783 31772
rect 48529 31709 48615 31732
rect 48697 31709 48783 31732
rect 63649 31772 63735 31795
rect 63817 31772 63903 31795
rect 63649 31732 63674 31772
rect 63674 31732 63714 31772
rect 63714 31732 63735 31772
rect 63817 31732 63838 31772
rect 63838 31732 63878 31772
rect 63878 31732 63903 31772
rect 63649 31709 63735 31732
rect 63817 31709 63903 31732
rect 78769 31772 78855 31795
rect 78937 31772 79023 31795
rect 78769 31732 78794 31772
rect 78794 31732 78834 31772
rect 78834 31732 78855 31772
rect 78937 31732 78958 31772
rect 78958 31732 78998 31772
rect 78998 31732 79023 31772
rect 78769 31709 78855 31732
rect 78937 31709 79023 31732
rect 93889 31772 93975 31795
rect 94057 31772 94143 31795
rect 93889 31732 93914 31772
rect 93914 31732 93954 31772
rect 93954 31732 93975 31772
rect 94057 31732 94078 31772
rect 94078 31732 94118 31772
rect 94118 31732 94143 31772
rect 93889 31709 93975 31732
rect 94057 31709 94143 31732
rect 4409 31016 4495 31039
rect 4577 31016 4663 31039
rect 4409 30976 4434 31016
rect 4434 30976 4474 31016
rect 4474 30976 4495 31016
rect 4577 30976 4598 31016
rect 4598 30976 4638 31016
rect 4638 30976 4663 31016
rect 4409 30953 4495 30976
rect 4577 30953 4663 30976
rect 19529 31016 19615 31039
rect 19697 31016 19783 31039
rect 19529 30976 19554 31016
rect 19554 30976 19594 31016
rect 19594 30976 19615 31016
rect 19697 30976 19718 31016
rect 19718 30976 19758 31016
rect 19758 30976 19783 31016
rect 19529 30953 19615 30976
rect 19697 30953 19783 30976
rect 34649 31016 34735 31039
rect 34817 31016 34903 31039
rect 34649 30976 34674 31016
rect 34674 30976 34714 31016
rect 34714 30976 34735 31016
rect 34817 30976 34838 31016
rect 34838 30976 34878 31016
rect 34878 30976 34903 31016
rect 34649 30953 34735 30976
rect 34817 30953 34903 30976
rect 49769 31016 49855 31039
rect 49937 31016 50023 31039
rect 49769 30976 49794 31016
rect 49794 30976 49834 31016
rect 49834 30976 49855 31016
rect 49937 30976 49958 31016
rect 49958 30976 49998 31016
rect 49998 30976 50023 31016
rect 49769 30953 49855 30976
rect 49937 30953 50023 30976
rect 64889 31016 64975 31039
rect 65057 31016 65143 31039
rect 64889 30976 64914 31016
rect 64914 30976 64954 31016
rect 64954 30976 64975 31016
rect 65057 30976 65078 31016
rect 65078 30976 65118 31016
rect 65118 30976 65143 31016
rect 64889 30953 64975 30976
rect 65057 30953 65143 30976
rect 80009 31016 80095 31039
rect 80177 31016 80263 31039
rect 80009 30976 80034 31016
rect 80034 30976 80074 31016
rect 80074 30976 80095 31016
rect 80177 30976 80198 31016
rect 80198 30976 80238 31016
rect 80238 30976 80263 31016
rect 80009 30953 80095 30976
rect 80177 30953 80263 30976
rect 95129 31016 95215 31039
rect 95297 31016 95383 31039
rect 95129 30976 95154 31016
rect 95154 30976 95194 31016
rect 95194 30976 95215 31016
rect 95297 30976 95318 31016
rect 95318 30976 95358 31016
rect 95358 30976 95383 31016
rect 95129 30953 95215 30976
rect 95297 30953 95383 30976
rect 3169 30260 3255 30283
rect 3337 30260 3423 30283
rect 3169 30220 3194 30260
rect 3194 30220 3234 30260
rect 3234 30220 3255 30260
rect 3337 30220 3358 30260
rect 3358 30220 3398 30260
rect 3398 30220 3423 30260
rect 3169 30197 3255 30220
rect 3337 30197 3423 30220
rect 18289 30260 18375 30283
rect 18457 30260 18543 30283
rect 18289 30220 18314 30260
rect 18314 30220 18354 30260
rect 18354 30220 18375 30260
rect 18457 30220 18478 30260
rect 18478 30220 18518 30260
rect 18518 30220 18543 30260
rect 18289 30197 18375 30220
rect 18457 30197 18543 30220
rect 33409 30260 33495 30283
rect 33577 30260 33663 30283
rect 33409 30220 33434 30260
rect 33434 30220 33474 30260
rect 33474 30220 33495 30260
rect 33577 30220 33598 30260
rect 33598 30220 33638 30260
rect 33638 30220 33663 30260
rect 33409 30197 33495 30220
rect 33577 30197 33663 30220
rect 48529 30260 48615 30283
rect 48697 30260 48783 30283
rect 48529 30220 48554 30260
rect 48554 30220 48594 30260
rect 48594 30220 48615 30260
rect 48697 30220 48718 30260
rect 48718 30220 48758 30260
rect 48758 30220 48783 30260
rect 48529 30197 48615 30220
rect 48697 30197 48783 30220
rect 63649 30260 63735 30283
rect 63817 30260 63903 30283
rect 63649 30220 63674 30260
rect 63674 30220 63714 30260
rect 63714 30220 63735 30260
rect 63817 30220 63838 30260
rect 63838 30220 63878 30260
rect 63878 30220 63903 30260
rect 63649 30197 63735 30220
rect 63817 30197 63903 30220
rect 78769 30260 78855 30283
rect 78937 30260 79023 30283
rect 78769 30220 78794 30260
rect 78794 30220 78834 30260
rect 78834 30220 78855 30260
rect 78937 30220 78958 30260
rect 78958 30220 78998 30260
rect 78998 30220 79023 30260
rect 78769 30197 78855 30220
rect 78937 30197 79023 30220
rect 93889 30260 93975 30283
rect 94057 30260 94143 30283
rect 93889 30220 93914 30260
rect 93914 30220 93954 30260
rect 93954 30220 93975 30260
rect 94057 30220 94078 30260
rect 94078 30220 94118 30260
rect 94118 30220 94143 30260
rect 93889 30197 93975 30220
rect 94057 30197 94143 30220
rect 4409 29504 4495 29527
rect 4577 29504 4663 29527
rect 4409 29464 4434 29504
rect 4434 29464 4474 29504
rect 4474 29464 4495 29504
rect 4577 29464 4598 29504
rect 4598 29464 4638 29504
rect 4638 29464 4663 29504
rect 4409 29441 4495 29464
rect 4577 29441 4663 29464
rect 19529 29504 19615 29527
rect 19697 29504 19783 29527
rect 19529 29464 19554 29504
rect 19554 29464 19594 29504
rect 19594 29464 19615 29504
rect 19697 29464 19718 29504
rect 19718 29464 19758 29504
rect 19758 29464 19783 29504
rect 19529 29441 19615 29464
rect 19697 29441 19783 29464
rect 34649 29504 34735 29527
rect 34817 29504 34903 29527
rect 34649 29464 34674 29504
rect 34674 29464 34714 29504
rect 34714 29464 34735 29504
rect 34817 29464 34838 29504
rect 34838 29464 34878 29504
rect 34878 29464 34903 29504
rect 34649 29441 34735 29464
rect 34817 29441 34903 29464
rect 49769 29504 49855 29527
rect 49937 29504 50023 29527
rect 49769 29464 49794 29504
rect 49794 29464 49834 29504
rect 49834 29464 49855 29504
rect 49937 29464 49958 29504
rect 49958 29464 49998 29504
rect 49998 29464 50023 29504
rect 49769 29441 49855 29464
rect 49937 29441 50023 29464
rect 64889 29504 64975 29527
rect 65057 29504 65143 29527
rect 64889 29464 64914 29504
rect 64914 29464 64954 29504
rect 64954 29464 64975 29504
rect 65057 29464 65078 29504
rect 65078 29464 65118 29504
rect 65118 29464 65143 29504
rect 64889 29441 64975 29464
rect 65057 29441 65143 29464
rect 80009 29504 80095 29527
rect 80177 29504 80263 29527
rect 80009 29464 80034 29504
rect 80034 29464 80074 29504
rect 80074 29464 80095 29504
rect 80177 29464 80198 29504
rect 80198 29464 80238 29504
rect 80238 29464 80263 29504
rect 80009 29441 80095 29464
rect 80177 29441 80263 29464
rect 95129 29504 95215 29527
rect 95297 29504 95383 29527
rect 95129 29464 95154 29504
rect 95154 29464 95194 29504
rect 95194 29464 95215 29504
rect 95297 29464 95318 29504
rect 95318 29464 95358 29504
rect 95358 29464 95383 29504
rect 95129 29441 95215 29464
rect 95297 29441 95383 29464
rect 3169 28748 3255 28771
rect 3337 28748 3423 28771
rect 3169 28708 3194 28748
rect 3194 28708 3234 28748
rect 3234 28708 3255 28748
rect 3337 28708 3358 28748
rect 3358 28708 3398 28748
rect 3398 28708 3423 28748
rect 3169 28685 3255 28708
rect 3337 28685 3423 28708
rect 18289 28748 18375 28771
rect 18457 28748 18543 28771
rect 18289 28708 18314 28748
rect 18314 28708 18354 28748
rect 18354 28708 18375 28748
rect 18457 28708 18478 28748
rect 18478 28708 18518 28748
rect 18518 28708 18543 28748
rect 18289 28685 18375 28708
rect 18457 28685 18543 28708
rect 33409 28748 33495 28771
rect 33577 28748 33663 28771
rect 33409 28708 33434 28748
rect 33434 28708 33474 28748
rect 33474 28708 33495 28748
rect 33577 28708 33598 28748
rect 33598 28708 33638 28748
rect 33638 28708 33663 28748
rect 33409 28685 33495 28708
rect 33577 28685 33663 28708
rect 48529 28748 48615 28771
rect 48697 28748 48783 28771
rect 48529 28708 48554 28748
rect 48554 28708 48594 28748
rect 48594 28708 48615 28748
rect 48697 28708 48718 28748
rect 48718 28708 48758 28748
rect 48758 28708 48783 28748
rect 48529 28685 48615 28708
rect 48697 28685 48783 28708
rect 63649 28748 63735 28771
rect 63817 28748 63903 28771
rect 63649 28708 63674 28748
rect 63674 28708 63714 28748
rect 63714 28708 63735 28748
rect 63817 28708 63838 28748
rect 63838 28708 63878 28748
rect 63878 28708 63903 28748
rect 63649 28685 63735 28708
rect 63817 28685 63903 28708
rect 78769 28748 78855 28771
rect 78937 28748 79023 28771
rect 78769 28708 78794 28748
rect 78794 28708 78834 28748
rect 78834 28708 78855 28748
rect 78937 28708 78958 28748
rect 78958 28708 78998 28748
rect 78998 28708 79023 28748
rect 78769 28685 78855 28708
rect 78937 28685 79023 28708
rect 93889 28748 93975 28771
rect 94057 28748 94143 28771
rect 93889 28708 93914 28748
rect 93914 28708 93954 28748
rect 93954 28708 93975 28748
rect 94057 28708 94078 28748
rect 94078 28708 94118 28748
rect 94118 28708 94143 28748
rect 93889 28685 93975 28708
rect 94057 28685 94143 28708
rect 4409 27992 4495 28015
rect 4577 27992 4663 28015
rect 4409 27952 4434 27992
rect 4434 27952 4474 27992
rect 4474 27952 4495 27992
rect 4577 27952 4598 27992
rect 4598 27952 4638 27992
rect 4638 27952 4663 27992
rect 4409 27929 4495 27952
rect 4577 27929 4663 27952
rect 19529 27992 19615 28015
rect 19697 27992 19783 28015
rect 19529 27952 19554 27992
rect 19554 27952 19594 27992
rect 19594 27952 19615 27992
rect 19697 27952 19718 27992
rect 19718 27952 19758 27992
rect 19758 27952 19783 27992
rect 19529 27929 19615 27952
rect 19697 27929 19783 27952
rect 34649 27992 34735 28015
rect 34817 27992 34903 28015
rect 34649 27952 34674 27992
rect 34674 27952 34714 27992
rect 34714 27952 34735 27992
rect 34817 27952 34838 27992
rect 34838 27952 34878 27992
rect 34878 27952 34903 27992
rect 34649 27929 34735 27952
rect 34817 27929 34903 27952
rect 49769 27992 49855 28015
rect 49937 27992 50023 28015
rect 49769 27952 49794 27992
rect 49794 27952 49834 27992
rect 49834 27952 49855 27992
rect 49937 27952 49958 27992
rect 49958 27952 49998 27992
rect 49998 27952 50023 27992
rect 49769 27929 49855 27952
rect 49937 27929 50023 27952
rect 64889 27992 64975 28015
rect 65057 27992 65143 28015
rect 64889 27952 64914 27992
rect 64914 27952 64954 27992
rect 64954 27952 64975 27992
rect 65057 27952 65078 27992
rect 65078 27952 65118 27992
rect 65118 27952 65143 27992
rect 64889 27929 64975 27952
rect 65057 27929 65143 27952
rect 80009 27992 80095 28015
rect 80177 27992 80263 28015
rect 80009 27952 80034 27992
rect 80034 27952 80074 27992
rect 80074 27952 80095 27992
rect 80177 27952 80198 27992
rect 80198 27952 80238 27992
rect 80238 27952 80263 27992
rect 80009 27929 80095 27952
rect 80177 27929 80263 27952
rect 95129 27992 95215 28015
rect 95297 27992 95383 28015
rect 95129 27952 95154 27992
rect 95154 27952 95194 27992
rect 95194 27952 95215 27992
rect 95297 27952 95318 27992
rect 95318 27952 95358 27992
rect 95358 27952 95383 27992
rect 95129 27929 95215 27952
rect 95297 27929 95383 27952
rect 3169 27236 3255 27259
rect 3337 27236 3423 27259
rect 3169 27196 3194 27236
rect 3194 27196 3234 27236
rect 3234 27196 3255 27236
rect 3337 27196 3358 27236
rect 3358 27196 3398 27236
rect 3398 27196 3423 27236
rect 3169 27173 3255 27196
rect 3337 27173 3423 27196
rect 18289 27236 18375 27259
rect 18457 27236 18543 27259
rect 18289 27196 18314 27236
rect 18314 27196 18354 27236
rect 18354 27196 18375 27236
rect 18457 27196 18478 27236
rect 18478 27196 18518 27236
rect 18518 27196 18543 27236
rect 18289 27173 18375 27196
rect 18457 27173 18543 27196
rect 33409 27236 33495 27259
rect 33577 27236 33663 27259
rect 33409 27196 33434 27236
rect 33434 27196 33474 27236
rect 33474 27196 33495 27236
rect 33577 27196 33598 27236
rect 33598 27196 33638 27236
rect 33638 27196 33663 27236
rect 33409 27173 33495 27196
rect 33577 27173 33663 27196
rect 48529 27236 48615 27259
rect 48697 27236 48783 27259
rect 48529 27196 48554 27236
rect 48554 27196 48594 27236
rect 48594 27196 48615 27236
rect 48697 27196 48718 27236
rect 48718 27196 48758 27236
rect 48758 27196 48783 27236
rect 48529 27173 48615 27196
rect 48697 27173 48783 27196
rect 63649 27236 63735 27259
rect 63817 27236 63903 27259
rect 63649 27196 63674 27236
rect 63674 27196 63714 27236
rect 63714 27196 63735 27236
rect 63817 27196 63838 27236
rect 63838 27196 63878 27236
rect 63878 27196 63903 27236
rect 63649 27173 63735 27196
rect 63817 27173 63903 27196
rect 78769 27236 78855 27259
rect 78937 27236 79023 27259
rect 78769 27196 78794 27236
rect 78794 27196 78834 27236
rect 78834 27196 78855 27236
rect 78937 27196 78958 27236
rect 78958 27196 78998 27236
rect 78998 27196 79023 27236
rect 78769 27173 78855 27196
rect 78937 27173 79023 27196
rect 93889 27236 93975 27259
rect 94057 27236 94143 27259
rect 93889 27196 93914 27236
rect 93914 27196 93954 27236
rect 93954 27196 93975 27236
rect 94057 27196 94078 27236
rect 94078 27196 94118 27236
rect 94118 27196 94143 27236
rect 93889 27173 93975 27196
rect 94057 27173 94143 27196
rect 4409 26480 4495 26503
rect 4577 26480 4663 26503
rect 4409 26440 4434 26480
rect 4434 26440 4474 26480
rect 4474 26440 4495 26480
rect 4577 26440 4598 26480
rect 4598 26440 4638 26480
rect 4638 26440 4663 26480
rect 4409 26417 4495 26440
rect 4577 26417 4663 26440
rect 19529 26480 19615 26503
rect 19697 26480 19783 26503
rect 19529 26440 19554 26480
rect 19554 26440 19594 26480
rect 19594 26440 19615 26480
rect 19697 26440 19718 26480
rect 19718 26440 19758 26480
rect 19758 26440 19783 26480
rect 19529 26417 19615 26440
rect 19697 26417 19783 26440
rect 34649 26480 34735 26503
rect 34817 26480 34903 26503
rect 34649 26440 34674 26480
rect 34674 26440 34714 26480
rect 34714 26440 34735 26480
rect 34817 26440 34838 26480
rect 34838 26440 34878 26480
rect 34878 26440 34903 26480
rect 34649 26417 34735 26440
rect 34817 26417 34903 26440
rect 49769 26480 49855 26503
rect 49937 26480 50023 26503
rect 49769 26440 49794 26480
rect 49794 26440 49834 26480
rect 49834 26440 49855 26480
rect 49937 26440 49958 26480
rect 49958 26440 49998 26480
rect 49998 26440 50023 26480
rect 49769 26417 49855 26440
rect 49937 26417 50023 26440
rect 64889 26480 64975 26503
rect 65057 26480 65143 26503
rect 64889 26440 64914 26480
rect 64914 26440 64954 26480
rect 64954 26440 64975 26480
rect 65057 26440 65078 26480
rect 65078 26440 65118 26480
rect 65118 26440 65143 26480
rect 64889 26417 64975 26440
rect 65057 26417 65143 26440
rect 80009 26480 80095 26503
rect 80177 26480 80263 26503
rect 80009 26440 80034 26480
rect 80034 26440 80074 26480
rect 80074 26440 80095 26480
rect 80177 26440 80198 26480
rect 80198 26440 80238 26480
rect 80238 26440 80263 26480
rect 80009 26417 80095 26440
rect 80177 26417 80263 26440
rect 95129 26480 95215 26503
rect 95297 26480 95383 26503
rect 95129 26440 95154 26480
rect 95154 26440 95194 26480
rect 95194 26440 95215 26480
rect 95297 26440 95318 26480
rect 95318 26440 95358 26480
rect 95358 26440 95383 26480
rect 95129 26417 95215 26440
rect 95297 26417 95383 26440
rect 3169 25724 3255 25747
rect 3337 25724 3423 25747
rect 3169 25684 3194 25724
rect 3194 25684 3234 25724
rect 3234 25684 3255 25724
rect 3337 25684 3358 25724
rect 3358 25684 3398 25724
rect 3398 25684 3423 25724
rect 3169 25661 3255 25684
rect 3337 25661 3423 25684
rect 18289 25724 18375 25747
rect 18457 25724 18543 25747
rect 18289 25684 18314 25724
rect 18314 25684 18354 25724
rect 18354 25684 18375 25724
rect 18457 25684 18478 25724
rect 18478 25684 18518 25724
rect 18518 25684 18543 25724
rect 18289 25661 18375 25684
rect 18457 25661 18543 25684
rect 33409 25724 33495 25747
rect 33577 25724 33663 25747
rect 33409 25684 33434 25724
rect 33434 25684 33474 25724
rect 33474 25684 33495 25724
rect 33577 25684 33598 25724
rect 33598 25684 33638 25724
rect 33638 25684 33663 25724
rect 33409 25661 33495 25684
rect 33577 25661 33663 25684
rect 48529 25724 48615 25747
rect 48697 25724 48783 25747
rect 48529 25684 48554 25724
rect 48554 25684 48594 25724
rect 48594 25684 48615 25724
rect 48697 25684 48718 25724
rect 48718 25684 48758 25724
rect 48758 25684 48783 25724
rect 48529 25661 48615 25684
rect 48697 25661 48783 25684
rect 63649 25724 63735 25747
rect 63817 25724 63903 25747
rect 63649 25684 63674 25724
rect 63674 25684 63714 25724
rect 63714 25684 63735 25724
rect 63817 25684 63838 25724
rect 63838 25684 63878 25724
rect 63878 25684 63903 25724
rect 63649 25661 63735 25684
rect 63817 25661 63903 25684
rect 78769 25724 78855 25747
rect 78937 25724 79023 25747
rect 78769 25684 78794 25724
rect 78794 25684 78834 25724
rect 78834 25684 78855 25724
rect 78937 25684 78958 25724
rect 78958 25684 78998 25724
rect 78998 25684 79023 25724
rect 78769 25661 78855 25684
rect 78937 25661 79023 25684
rect 93889 25724 93975 25747
rect 94057 25724 94143 25747
rect 93889 25684 93914 25724
rect 93914 25684 93954 25724
rect 93954 25684 93975 25724
rect 94057 25684 94078 25724
rect 94078 25684 94118 25724
rect 94118 25684 94143 25724
rect 93889 25661 93975 25684
rect 94057 25661 94143 25684
rect 4409 24968 4495 24991
rect 4577 24968 4663 24991
rect 4409 24928 4434 24968
rect 4434 24928 4474 24968
rect 4474 24928 4495 24968
rect 4577 24928 4598 24968
rect 4598 24928 4638 24968
rect 4638 24928 4663 24968
rect 4409 24905 4495 24928
rect 4577 24905 4663 24928
rect 19529 24968 19615 24991
rect 19697 24968 19783 24991
rect 19529 24928 19554 24968
rect 19554 24928 19594 24968
rect 19594 24928 19615 24968
rect 19697 24928 19718 24968
rect 19718 24928 19758 24968
rect 19758 24928 19783 24968
rect 19529 24905 19615 24928
rect 19697 24905 19783 24928
rect 34649 24968 34735 24991
rect 34817 24968 34903 24991
rect 34649 24928 34674 24968
rect 34674 24928 34714 24968
rect 34714 24928 34735 24968
rect 34817 24928 34838 24968
rect 34838 24928 34878 24968
rect 34878 24928 34903 24968
rect 34649 24905 34735 24928
rect 34817 24905 34903 24928
rect 49769 24968 49855 24991
rect 49937 24968 50023 24991
rect 49769 24928 49794 24968
rect 49794 24928 49834 24968
rect 49834 24928 49855 24968
rect 49937 24928 49958 24968
rect 49958 24928 49998 24968
rect 49998 24928 50023 24968
rect 49769 24905 49855 24928
rect 49937 24905 50023 24928
rect 64889 24968 64975 24991
rect 65057 24968 65143 24991
rect 64889 24928 64914 24968
rect 64914 24928 64954 24968
rect 64954 24928 64975 24968
rect 65057 24928 65078 24968
rect 65078 24928 65118 24968
rect 65118 24928 65143 24968
rect 64889 24905 64975 24928
rect 65057 24905 65143 24928
rect 80009 24968 80095 24991
rect 80177 24968 80263 24991
rect 80009 24928 80034 24968
rect 80034 24928 80074 24968
rect 80074 24928 80095 24968
rect 80177 24928 80198 24968
rect 80198 24928 80238 24968
rect 80238 24928 80263 24968
rect 80009 24905 80095 24928
rect 80177 24905 80263 24928
rect 95129 24968 95215 24991
rect 95297 24968 95383 24991
rect 95129 24928 95154 24968
rect 95154 24928 95194 24968
rect 95194 24928 95215 24968
rect 95297 24928 95318 24968
rect 95318 24928 95358 24968
rect 95358 24928 95383 24968
rect 95129 24905 95215 24928
rect 95297 24905 95383 24928
rect 3169 24212 3255 24235
rect 3337 24212 3423 24235
rect 3169 24172 3194 24212
rect 3194 24172 3234 24212
rect 3234 24172 3255 24212
rect 3337 24172 3358 24212
rect 3358 24172 3398 24212
rect 3398 24172 3423 24212
rect 3169 24149 3255 24172
rect 3337 24149 3423 24172
rect 18289 24212 18375 24235
rect 18457 24212 18543 24235
rect 18289 24172 18314 24212
rect 18314 24172 18354 24212
rect 18354 24172 18375 24212
rect 18457 24172 18478 24212
rect 18478 24172 18518 24212
rect 18518 24172 18543 24212
rect 18289 24149 18375 24172
rect 18457 24149 18543 24172
rect 33409 24212 33495 24235
rect 33577 24212 33663 24235
rect 33409 24172 33434 24212
rect 33434 24172 33474 24212
rect 33474 24172 33495 24212
rect 33577 24172 33598 24212
rect 33598 24172 33638 24212
rect 33638 24172 33663 24212
rect 33409 24149 33495 24172
rect 33577 24149 33663 24172
rect 48529 24212 48615 24235
rect 48697 24212 48783 24235
rect 48529 24172 48554 24212
rect 48554 24172 48594 24212
rect 48594 24172 48615 24212
rect 48697 24172 48718 24212
rect 48718 24172 48758 24212
rect 48758 24172 48783 24212
rect 48529 24149 48615 24172
rect 48697 24149 48783 24172
rect 63649 24212 63735 24235
rect 63817 24212 63903 24235
rect 63649 24172 63674 24212
rect 63674 24172 63714 24212
rect 63714 24172 63735 24212
rect 63817 24172 63838 24212
rect 63838 24172 63878 24212
rect 63878 24172 63903 24212
rect 63649 24149 63735 24172
rect 63817 24149 63903 24172
rect 78769 24212 78855 24235
rect 78937 24212 79023 24235
rect 78769 24172 78794 24212
rect 78794 24172 78834 24212
rect 78834 24172 78855 24212
rect 78937 24172 78958 24212
rect 78958 24172 78998 24212
rect 78998 24172 79023 24212
rect 78769 24149 78855 24172
rect 78937 24149 79023 24172
rect 93889 24212 93975 24235
rect 94057 24212 94143 24235
rect 93889 24172 93914 24212
rect 93914 24172 93954 24212
rect 93954 24172 93975 24212
rect 94057 24172 94078 24212
rect 94078 24172 94118 24212
rect 94118 24172 94143 24212
rect 93889 24149 93975 24172
rect 94057 24149 94143 24172
rect 4409 23456 4495 23479
rect 4577 23456 4663 23479
rect 4409 23416 4434 23456
rect 4434 23416 4474 23456
rect 4474 23416 4495 23456
rect 4577 23416 4598 23456
rect 4598 23416 4638 23456
rect 4638 23416 4663 23456
rect 4409 23393 4495 23416
rect 4577 23393 4663 23416
rect 19529 23456 19615 23479
rect 19697 23456 19783 23479
rect 19529 23416 19554 23456
rect 19554 23416 19594 23456
rect 19594 23416 19615 23456
rect 19697 23416 19718 23456
rect 19718 23416 19758 23456
rect 19758 23416 19783 23456
rect 19529 23393 19615 23416
rect 19697 23393 19783 23416
rect 34649 23456 34735 23479
rect 34817 23456 34903 23479
rect 34649 23416 34674 23456
rect 34674 23416 34714 23456
rect 34714 23416 34735 23456
rect 34817 23416 34838 23456
rect 34838 23416 34878 23456
rect 34878 23416 34903 23456
rect 34649 23393 34735 23416
rect 34817 23393 34903 23416
rect 49769 23456 49855 23479
rect 49937 23456 50023 23479
rect 49769 23416 49794 23456
rect 49794 23416 49834 23456
rect 49834 23416 49855 23456
rect 49937 23416 49958 23456
rect 49958 23416 49998 23456
rect 49998 23416 50023 23456
rect 49769 23393 49855 23416
rect 49937 23393 50023 23416
rect 64889 23456 64975 23479
rect 65057 23456 65143 23479
rect 64889 23416 64914 23456
rect 64914 23416 64954 23456
rect 64954 23416 64975 23456
rect 65057 23416 65078 23456
rect 65078 23416 65118 23456
rect 65118 23416 65143 23456
rect 64889 23393 64975 23416
rect 65057 23393 65143 23416
rect 80009 23456 80095 23479
rect 80177 23456 80263 23479
rect 80009 23416 80034 23456
rect 80034 23416 80074 23456
rect 80074 23416 80095 23456
rect 80177 23416 80198 23456
rect 80198 23416 80238 23456
rect 80238 23416 80263 23456
rect 80009 23393 80095 23416
rect 80177 23393 80263 23416
rect 95129 23456 95215 23479
rect 95297 23456 95383 23479
rect 95129 23416 95154 23456
rect 95154 23416 95194 23456
rect 95194 23416 95215 23456
rect 95297 23416 95318 23456
rect 95318 23416 95358 23456
rect 95358 23416 95383 23456
rect 95129 23393 95215 23416
rect 95297 23393 95383 23416
rect 3169 22700 3255 22723
rect 3337 22700 3423 22723
rect 3169 22660 3194 22700
rect 3194 22660 3234 22700
rect 3234 22660 3255 22700
rect 3337 22660 3358 22700
rect 3358 22660 3398 22700
rect 3398 22660 3423 22700
rect 3169 22637 3255 22660
rect 3337 22637 3423 22660
rect 18289 22700 18375 22723
rect 18457 22700 18543 22723
rect 18289 22660 18314 22700
rect 18314 22660 18354 22700
rect 18354 22660 18375 22700
rect 18457 22660 18478 22700
rect 18478 22660 18518 22700
rect 18518 22660 18543 22700
rect 18289 22637 18375 22660
rect 18457 22637 18543 22660
rect 33409 22700 33495 22723
rect 33577 22700 33663 22723
rect 33409 22660 33434 22700
rect 33434 22660 33474 22700
rect 33474 22660 33495 22700
rect 33577 22660 33598 22700
rect 33598 22660 33638 22700
rect 33638 22660 33663 22700
rect 33409 22637 33495 22660
rect 33577 22637 33663 22660
rect 48529 22700 48615 22723
rect 48697 22700 48783 22723
rect 48529 22660 48554 22700
rect 48554 22660 48594 22700
rect 48594 22660 48615 22700
rect 48697 22660 48718 22700
rect 48718 22660 48758 22700
rect 48758 22660 48783 22700
rect 48529 22637 48615 22660
rect 48697 22637 48783 22660
rect 63649 22700 63735 22723
rect 63817 22700 63903 22723
rect 63649 22660 63674 22700
rect 63674 22660 63714 22700
rect 63714 22660 63735 22700
rect 63817 22660 63838 22700
rect 63838 22660 63878 22700
rect 63878 22660 63903 22700
rect 63649 22637 63735 22660
rect 63817 22637 63903 22660
rect 78769 22700 78855 22723
rect 78937 22700 79023 22723
rect 78769 22660 78794 22700
rect 78794 22660 78834 22700
rect 78834 22660 78855 22700
rect 78937 22660 78958 22700
rect 78958 22660 78998 22700
rect 78998 22660 79023 22700
rect 78769 22637 78855 22660
rect 78937 22637 79023 22660
rect 93889 22700 93975 22723
rect 94057 22700 94143 22723
rect 93889 22660 93914 22700
rect 93914 22660 93954 22700
rect 93954 22660 93975 22700
rect 94057 22660 94078 22700
rect 94078 22660 94118 22700
rect 94118 22660 94143 22700
rect 93889 22637 93975 22660
rect 94057 22637 94143 22660
rect 4409 21944 4495 21967
rect 4577 21944 4663 21967
rect 4409 21904 4434 21944
rect 4434 21904 4474 21944
rect 4474 21904 4495 21944
rect 4577 21904 4598 21944
rect 4598 21904 4638 21944
rect 4638 21904 4663 21944
rect 4409 21881 4495 21904
rect 4577 21881 4663 21904
rect 19529 21944 19615 21967
rect 19697 21944 19783 21967
rect 19529 21904 19554 21944
rect 19554 21904 19594 21944
rect 19594 21904 19615 21944
rect 19697 21904 19718 21944
rect 19718 21904 19758 21944
rect 19758 21904 19783 21944
rect 19529 21881 19615 21904
rect 19697 21881 19783 21904
rect 34649 21944 34735 21967
rect 34817 21944 34903 21967
rect 34649 21904 34674 21944
rect 34674 21904 34714 21944
rect 34714 21904 34735 21944
rect 34817 21904 34838 21944
rect 34838 21904 34878 21944
rect 34878 21904 34903 21944
rect 34649 21881 34735 21904
rect 34817 21881 34903 21904
rect 49769 21944 49855 21967
rect 49937 21944 50023 21967
rect 49769 21904 49794 21944
rect 49794 21904 49834 21944
rect 49834 21904 49855 21944
rect 49937 21904 49958 21944
rect 49958 21904 49998 21944
rect 49998 21904 50023 21944
rect 49769 21881 49855 21904
rect 49937 21881 50023 21904
rect 64889 21944 64975 21967
rect 65057 21944 65143 21967
rect 64889 21904 64914 21944
rect 64914 21904 64954 21944
rect 64954 21904 64975 21944
rect 65057 21904 65078 21944
rect 65078 21904 65118 21944
rect 65118 21904 65143 21944
rect 64889 21881 64975 21904
rect 65057 21881 65143 21904
rect 80009 21944 80095 21967
rect 80177 21944 80263 21967
rect 80009 21904 80034 21944
rect 80034 21904 80074 21944
rect 80074 21904 80095 21944
rect 80177 21904 80198 21944
rect 80198 21904 80238 21944
rect 80238 21904 80263 21944
rect 80009 21881 80095 21904
rect 80177 21881 80263 21904
rect 95129 21944 95215 21967
rect 95297 21944 95383 21967
rect 95129 21904 95154 21944
rect 95154 21904 95194 21944
rect 95194 21904 95215 21944
rect 95297 21904 95318 21944
rect 95318 21904 95358 21944
rect 95358 21904 95383 21944
rect 95129 21881 95215 21904
rect 95297 21881 95383 21904
rect 3169 21188 3255 21211
rect 3337 21188 3423 21211
rect 3169 21148 3194 21188
rect 3194 21148 3234 21188
rect 3234 21148 3255 21188
rect 3337 21148 3358 21188
rect 3358 21148 3398 21188
rect 3398 21148 3423 21188
rect 3169 21125 3255 21148
rect 3337 21125 3423 21148
rect 18289 21188 18375 21211
rect 18457 21188 18543 21211
rect 18289 21148 18314 21188
rect 18314 21148 18354 21188
rect 18354 21148 18375 21188
rect 18457 21148 18478 21188
rect 18478 21148 18518 21188
rect 18518 21148 18543 21188
rect 18289 21125 18375 21148
rect 18457 21125 18543 21148
rect 33409 21188 33495 21211
rect 33577 21188 33663 21211
rect 33409 21148 33434 21188
rect 33434 21148 33474 21188
rect 33474 21148 33495 21188
rect 33577 21148 33598 21188
rect 33598 21148 33638 21188
rect 33638 21148 33663 21188
rect 33409 21125 33495 21148
rect 33577 21125 33663 21148
rect 48529 21188 48615 21211
rect 48697 21188 48783 21211
rect 48529 21148 48554 21188
rect 48554 21148 48594 21188
rect 48594 21148 48615 21188
rect 48697 21148 48718 21188
rect 48718 21148 48758 21188
rect 48758 21148 48783 21188
rect 48529 21125 48615 21148
rect 48697 21125 48783 21148
rect 63649 21188 63735 21211
rect 63817 21188 63903 21211
rect 63649 21148 63674 21188
rect 63674 21148 63714 21188
rect 63714 21148 63735 21188
rect 63817 21148 63838 21188
rect 63838 21148 63878 21188
rect 63878 21148 63903 21188
rect 63649 21125 63735 21148
rect 63817 21125 63903 21148
rect 78769 21188 78855 21211
rect 78937 21188 79023 21211
rect 78769 21148 78794 21188
rect 78794 21148 78834 21188
rect 78834 21148 78855 21188
rect 78937 21148 78958 21188
rect 78958 21148 78998 21188
rect 78998 21148 79023 21188
rect 78769 21125 78855 21148
rect 78937 21125 79023 21148
rect 93889 21188 93975 21211
rect 94057 21188 94143 21211
rect 93889 21148 93914 21188
rect 93914 21148 93954 21188
rect 93954 21148 93975 21188
rect 94057 21148 94078 21188
rect 94078 21148 94118 21188
rect 94118 21148 94143 21188
rect 93889 21125 93975 21148
rect 94057 21125 94143 21148
rect 4409 20432 4495 20455
rect 4577 20432 4663 20455
rect 4409 20392 4434 20432
rect 4434 20392 4474 20432
rect 4474 20392 4495 20432
rect 4577 20392 4598 20432
rect 4598 20392 4638 20432
rect 4638 20392 4663 20432
rect 4409 20369 4495 20392
rect 4577 20369 4663 20392
rect 19529 20432 19615 20455
rect 19697 20432 19783 20455
rect 19529 20392 19554 20432
rect 19554 20392 19594 20432
rect 19594 20392 19615 20432
rect 19697 20392 19718 20432
rect 19718 20392 19758 20432
rect 19758 20392 19783 20432
rect 19529 20369 19615 20392
rect 19697 20369 19783 20392
rect 34649 20432 34735 20455
rect 34817 20432 34903 20455
rect 34649 20392 34674 20432
rect 34674 20392 34714 20432
rect 34714 20392 34735 20432
rect 34817 20392 34838 20432
rect 34838 20392 34878 20432
rect 34878 20392 34903 20432
rect 34649 20369 34735 20392
rect 34817 20369 34903 20392
rect 49769 20432 49855 20455
rect 49937 20432 50023 20455
rect 49769 20392 49794 20432
rect 49794 20392 49834 20432
rect 49834 20392 49855 20432
rect 49937 20392 49958 20432
rect 49958 20392 49998 20432
rect 49998 20392 50023 20432
rect 49769 20369 49855 20392
rect 49937 20369 50023 20392
rect 64889 20432 64975 20455
rect 65057 20432 65143 20455
rect 64889 20392 64914 20432
rect 64914 20392 64954 20432
rect 64954 20392 64975 20432
rect 65057 20392 65078 20432
rect 65078 20392 65118 20432
rect 65118 20392 65143 20432
rect 64889 20369 64975 20392
rect 65057 20369 65143 20392
rect 80009 20432 80095 20455
rect 80177 20432 80263 20455
rect 80009 20392 80034 20432
rect 80034 20392 80074 20432
rect 80074 20392 80095 20432
rect 80177 20392 80198 20432
rect 80198 20392 80238 20432
rect 80238 20392 80263 20432
rect 80009 20369 80095 20392
rect 80177 20369 80263 20392
rect 95129 20432 95215 20455
rect 95297 20432 95383 20455
rect 95129 20392 95154 20432
rect 95154 20392 95194 20432
rect 95194 20392 95215 20432
rect 95297 20392 95318 20432
rect 95318 20392 95358 20432
rect 95358 20392 95383 20432
rect 95129 20369 95215 20392
rect 95297 20369 95383 20392
rect 3169 19676 3255 19699
rect 3337 19676 3423 19699
rect 3169 19636 3194 19676
rect 3194 19636 3234 19676
rect 3234 19636 3255 19676
rect 3337 19636 3358 19676
rect 3358 19636 3398 19676
rect 3398 19636 3423 19676
rect 3169 19613 3255 19636
rect 3337 19613 3423 19636
rect 18289 19676 18375 19699
rect 18457 19676 18543 19699
rect 18289 19636 18314 19676
rect 18314 19636 18354 19676
rect 18354 19636 18375 19676
rect 18457 19636 18478 19676
rect 18478 19636 18518 19676
rect 18518 19636 18543 19676
rect 18289 19613 18375 19636
rect 18457 19613 18543 19636
rect 33409 19676 33495 19699
rect 33577 19676 33663 19699
rect 33409 19636 33434 19676
rect 33434 19636 33474 19676
rect 33474 19636 33495 19676
rect 33577 19636 33598 19676
rect 33598 19636 33638 19676
rect 33638 19636 33663 19676
rect 33409 19613 33495 19636
rect 33577 19613 33663 19636
rect 48529 19676 48615 19699
rect 48697 19676 48783 19699
rect 48529 19636 48554 19676
rect 48554 19636 48594 19676
rect 48594 19636 48615 19676
rect 48697 19636 48718 19676
rect 48718 19636 48758 19676
rect 48758 19636 48783 19676
rect 48529 19613 48615 19636
rect 48697 19613 48783 19636
rect 63649 19676 63735 19699
rect 63817 19676 63903 19699
rect 63649 19636 63674 19676
rect 63674 19636 63714 19676
rect 63714 19636 63735 19676
rect 63817 19636 63838 19676
rect 63838 19636 63878 19676
rect 63878 19636 63903 19676
rect 63649 19613 63735 19636
rect 63817 19613 63903 19636
rect 78769 19676 78855 19699
rect 78937 19676 79023 19699
rect 78769 19636 78794 19676
rect 78794 19636 78834 19676
rect 78834 19636 78855 19676
rect 78937 19636 78958 19676
rect 78958 19636 78998 19676
rect 78998 19636 79023 19676
rect 78769 19613 78855 19636
rect 78937 19613 79023 19636
rect 93889 19676 93975 19699
rect 94057 19676 94143 19699
rect 93889 19636 93914 19676
rect 93914 19636 93954 19676
rect 93954 19636 93975 19676
rect 94057 19636 94078 19676
rect 94078 19636 94118 19676
rect 94118 19636 94143 19676
rect 93889 19613 93975 19636
rect 94057 19613 94143 19636
rect 4409 18920 4495 18943
rect 4577 18920 4663 18943
rect 4409 18880 4434 18920
rect 4434 18880 4474 18920
rect 4474 18880 4495 18920
rect 4577 18880 4598 18920
rect 4598 18880 4638 18920
rect 4638 18880 4663 18920
rect 4409 18857 4495 18880
rect 4577 18857 4663 18880
rect 19529 18920 19615 18943
rect 19697 18920 19783 18943
rect 19529 18880 19554 18920
rect 19554 18880 19594 18920
rect 19594 18880 19615 18920
rect 19697 18880 19718 18920
rect 19718 18880 19758 18920
rect 19758 18880 19783 18920
rect 19529 18857 19615 18880
rect 19697 18857 19783 18880
rect 34649 18920 34735 18943
rect 34817 18920 34903 18943
rect 34649 18880 34674 18920
rect 34674 18880 34714 18920
rect 34714 18880 34735 18920
rect 34817 18880 34838 18920
rect 34838 18880 34878 18920
rect 34878 18880 34903 18920
rect 34649 18857 34735 18880
rect 34817 18857 34903 18880
rect 49769 18920 49855 18943
rect 49937 18920 50023 18943
rect 49769 18880 49794 18920
rect 49794 18880 49834 18920
rect 49834 18880 49855 18920
rect 49937 18880 49958 18920
rect 49958 18880 49998 18920
rect 49998 18880 50023 18920
rect 49769 18857 49855 18880
rect 49937 18857 50023 18880
rect 64889 18920 64975 18943
rect 65057 18920 65143 18943
rect 64889 18880 64914 18920
rect 64914 18880 64954 18920
rect 64954 18880 64975 18920
rect 65057 18880 65078 18920
rect 65078 18880 65118 18920
rect 65118 18880 65143 18920
rect 64889 18857 64975 18880
rect 65057 18857 65143 18880
rect 80009 18920 80095 18943
rect 80177 18920 80263 18943
rect 80009 18880 80034 18920
rect 80034 18880 80074 18920
rect 80074 18880 80095 18920
rect 80177 18880 80198 18920
rect 80198 18880 80238 18920
rect 80238 18880 80263 18920
rect 80009 18857 80095 18880
rect 80177 18857 80263 18880
rect 95129 18920 95215 18943
rect 95297 18920 95383 18943
rect 95129 18880 95154 18920
rect 95154 18880 95194 18920
rect 95194 18880 95215 18920
rect 95297 18880 95318 18920
rect 95318 18880 95358 18920
rect 95358 18880 95383 18920
rect 95129 18857 95215 18880
rect 95297 18857 95383 18880
rect 3169 18164 3255 18187
rect 3337 18164 3423 18187
rect 3169 18124 3194 18164
rect 3194 18124 3234 18164
rect 3234 18124 3255 18164
rect 3337 18124 3358 18164
rect 3358 18124 3398 18164
rect 3398 18124 3423 18164
rect 3169 18101 3255 18124
rect 3337 18101 3423 18124
rect 18289 18164 18375 18187
rect 18457 18164 18543 18187
rect 18289 18124 18314 18164
rect 18314 18124 18354 18164
rect 18354 18124 18375 18164
rect 18457 18124 18478 18164
rect 18478 18124 18518 18164
rect 18518 18124 18543 18164
rect 18289 18101 18375 18124
rect 18457 18101 18543 18124
rect 33409 18164 33495 18187
rect 33577 18164 33663 18187
rect 33409 18124 33434 18164
rect 33434 18124 33474 18164
rect 33474 18124 33495 18164
rect 33577 18124 33598 18164
rect 33598 18124 33638 18164
rect 33638 18124 33663 18164
rect 33409 18101 33495 18124
rect 33577 18101 33663 18124
rect 48529 18164 48615 18187
rect 48697 18164 48783 18187
rect 48529 18124 48554 18164
rect 48554 18124 48594 18164
rect 48594 18124 48615 18164
rect 48697 18124 48718 18164
rect 48718 18124 48758 18164
rect 48758 18124 48783 18164
rect 48529 18101 48615 18124
rect 48697 18101 48783 18124
rect 63649 18164 63735 18187
rect 63817 18164 63903 18187
rect 63649 18124 63674 18164
rect 63674 18124 63714 18164
rect 63714 18124 63735 18164
rect 63817 18124 63838 18164
rect 63838 18124 63878 18164
rect 63878 18124 63903 18164
rect 63649 18101 63735 18124
rect 63817 18101 63903 18124
rect 78769 18164 78855 18187
rect 78937 18164 79023 18187
rect 78769 18124 78794 18164
rect 78794 18124 78834 18164
rect 78834 18124 78855 18164
rect 78937 18124 78958 18164
rect 78958 18124 78998 18164
rect 78998 18124 79023 18164
rect 78769 18101 78855 18124
rect 78937 18101 79023 18124
rect 93889 18164 93975 18187
rect 94057 18164 94143 18187
rect 93889 18124 93914 18164
rect 93914 18124 93954 18164
rect 93954 18124 93975 18164
rect 94057 18124 94078 18164
rect 94078 18124 94118 18164
rect 94118 18124 94143 18164
rect 93889 18101 93975 18124
rect 94057 18101 94143 18124
rect 4409 17408 4495 17431
rect 4577 17408 4663 17431
rect 4409 17368 4434 17408
rect 4434 17368 4474 17408
rect 4474 17368 4495 17408
rect 4577 17368 4598 17408
rect 4598 17368 4638 17408
rect 4638 17368 4663 17408
rect 4409 17345 4495 17368
rect 4577 17345 4663 17368
rect 19529 17408 19615 17431
rect 19697 17408 19783 17431
rect 19529 17368 19554 17408
rect 19554 17368 19594 17408
rect 19594 17368 19615 17408
rect 19697 17368 19718 17408
rect 19718 17368 19758 17408
rect 19758 17368 19783 17408
rect 19529 17345 19615 17368
rect 19697 17345 19783 17368
rect 34649 17408 34735 17431
rect 34817 17408 34903 17431
rect 34649 17368 34674 17408
rect 34674 17368 34714 17408
rect 34714 17368 34735 17408
rect 34817 17368 34838 17408
rect 34838 17368 34878 17408
rect 34878 17368 34903 17408
rect 34649 17345 34735 17368
rect 34817 17345 34903 17368
rect 49769 17408 49855 17431
rect 49937 17408 50023 17431
rect 49769 17368 49794 17408
rect 49794 17368 49834 17408
rect 49834 17368 49855 17408
rect 49937 17368 49958 17408
rect 49958 17368 49998 17408
rect 49998 17368 50023 17408
rect 49769 17345 49855 17368
rect 49937 17345 50023 17368
rect 64889 17408 64975 17431
rect 65057 17408 65143 17431
rect 64889 17368 64914 17408
rect 64914 17368 64954 17408
rect 64954 17368 64975 17408
rect 65057 17368 65078 17408
rect 65078 17368 65118 17408
rect 65118 17368 65143 17408
rect 64889 17345 64975 17368
rect 65057 17345 65143 17368
rect 80009 17408 80095 17431
rect 80177 17408 80263 17431
rect 80009 17368 80034 17408
rect 80034 17368 80074 17408
rect 80074 17368 80095 17408
rect 80177 17368 80198 17408
rect 80198 17368 80238 17408
rect 80238 17368 80263 17408
rect 80009 17345 80095 17368
rect 80177 17345 80263 17368
rect 95129 17408 95215 17431
rect 95297 17408 95383 17431
rect 95129 17368 95154 17408
rect 95154 17368 95194 17408
rect 95194 17368 95215 17408
rect 95297 17368 95318 17408
rect 95318 17368 95358 17408
rect 95358 17368 95383 17408
rect 95129 17345 95215 17368
rect 95297 17345 95383 17368
rect 3169 16652 3255 16675
rect 3337 16652 3423 16675
rect 3169 16612 3194 16652
rect 3194 16612 3234 16652
rect 3234 16612 3255 16652
rect 3337 16612 3358 16652
rect 3358 16612 3398 16652
rect 3398 16612 3423 16652
rect 3169 16589 3255 16612
rect 3337 16589 3423 16612
rect 18289 16652 18375 16675
rect 18457 16652 18543 16675
rect 18289 16612 18314 16652
rect 18314 16612 18354 16652
rect 18354 16612 18375 16652
rect 18457 16612 18478 16652
rect 18478 16612 18518 16652
rect 18518 16612 18543 16652
rect 18289 16589 18375 16612
rect 18457 16589 18543 16612
rect 33409 16652 33495 16675
rect 33577 16652 33663 16675
rect 33409 16612 33434 16652
rect 33434 16612 33474 16652
rect 33474 16612 33495 16652
rect 33577 16612 33598 16652
rect 33598 16612 33638 16652
rect 33638 16612 33663 16652
rect 33409 16589 33495 16612
rect 33577 16589 33663 16612
rect 48529 16652 48615 16675
rect 48697 16652 48783 16675
rect 48529 16612 48554 16652
rect 48554 16612 48594 16652
rect 48594 16612 48615 16652
rect 48697 16612 48718 16652
rect 48718 16612 48758 16652
rect 48758 16612 48783 16652
rect 48529 16589 48615 16612
rect 48697 16589 48783 16612
rect 63649 16652 63735 16675
rect 63817 16652 63903 16675
rect 63649 16612 63674 16652
rect 63674 16612 63714 16652
rect 63714 16612 63735 16652
rect 63817 16612 63838 16652
rect 63838 16612 63878 16652
rect 63878 16612 63903 16652
rect 63649 16589 63735 16612
rect 63817 16589 63903 16612
rect 78769 16652 78855 16675
rect 78937 16652 79023 16675
rect 78769 16612 78794 16652
rect 78794 16612 78834 16652
rect 78834 16612 78855 16652
rect 78937 16612 78958 16652
rect 78958 16612 78998 16652
rect 78998 16612 79023 16652
rect 78769 16589 78855 16612
rect 78937 16589 79023 16612
rect 93889 16652 93975 16675
rect 94057 16652 94143 16675
rect 93889 16612 93914 16652
rect 93914 16612 93954 16652
rect 93954 16612 93975 16652
rect 94057 16612 94078 16652
rect 94078 16612 94118 16652
rect 94118 16612 94143 16652
rect 93889 16589 93975 16612
rect 94057 16589 94143 16612
rect 4409 15896 4495 15919
rect 4577 15896 4663 15919
rect 4409 15856 4434 15896
rect 4434 15856 4474 15896
rect 4474 15856 4495 15896
rect 4577 15856 4598 15896
rect 4598 15856 4638 15896
rect 4638 15856 4663 15896
rect 4409 15833 4495 15856
rect 4577 15833 4663 15856
rect 19529 15896 19615 15919
rect 19697 15896 19783 15919
rect 19529 15856 19554 15896
rect 19554 15856 19594 15896
rect 19594 15856 19615 15896
rect 19697 15856 19718 15896
rect 19718 15856 19758 15896
rect 19758 15856 19783 15896
rect 19529 15833 19615 15856
rect 19697 15833 19783 15856
rect 34649 15896 34735 15919
rect 34817 15896 34903 15919
rect 34649 15856 34674 15896
rect 34674 15856 34714 15896
rect 34714 15856 34735 15896
rect 34817 15856 34838 15896
rect 34838 15856 34878 15896
rect 34878 15856 34903 15896
rect 34649 15833 34735 15856
rect 34817 15833 34903 15856
rect 49769 15896 49855 15919
rect 49937 15896 50023 15919
rect 49769 15856 49794 15896
rect 49794 15856 49834 15896
rect 49834 15856 49855 15896
rect 49937 15856 49958 15896
rect 49958 15856 49998 15896
rect 49998 15856 50023 15896
rect 49769 15833 49855 15856
rect 49937 15833 50023 15856
rect 64889 15896 64975 15919
rect 65057 15896 65143 15919
rect 64889 15856 64914 15896
rect 64914 15856 64954 15896
rect 64954 15856 64975 15896
rect 65057 15856 65078 15896
rect 65078 15856 65118 15896
rect 65118 15856 65143 15896
rect 64889 15833 64975 15856
rect 65057 15833 65143 15856
rect 80009 15896 80095 15919
rect 80177 15896 80263 15919
rect 80009 15856 80034 15896
rect 80034 15856 80074 15896
rect 80074 15856 80095 15896
rect 80177 15856 80198 15896
rect 80198 15856 80238 15896
rect 80238 15856 80263 15896
rect 80009 15833 80095 15856
rect 80177 15833 80263 15856
rect 95129 15896 95215 15919
rect 95297 15896 95383 15919
rect 95129 15856 95154 15896
rect 95154 15856 95194 15896
rect 95194 15856 95215 15896
rect 95297 15856 95318 15896
rect 95318 15856 95358 15896
rect 95358 15856 95383 15896
rect 95129 15833 95215 15856
rect 95297 15833 95383 15856
rect 3169 15140 3255 15163
rect 3337 15140 3423 15163
rect 3169 15100 3194 15140
rect 3194 15100 3234 15140
rect 3234 15100 3255 15140
rect 3337 15100 3358 15140
rect 3358 15100 3398 15140
rect 3398 15100 3423 15140
rect 3169 15077 3255 15100
rect 3337 15077 3423 15100
rect 18289 15140 18375 15163
rect 18457 15140 18543 15163
rect 18289 15100 18314 15140
rect 18314 15100 18354 15140
rect 18354 15100 18375 15140
rect 18457 15100 18478 15140
rect 18478 15100 18518 15140
rect 18518 15100 18543 15140
rect 18289 15077 18375 15100
rect 18457 15077 18543 15100
rect 33409 15140 33495 15163
rect 33577 15140 33663 15163
rect 33409 15100 33434 15140
rect 33434 15100 33474 15140
rect 33474 15100 33495 15140
rect 33577 15100 33598 15140
rect 33598 15100 33638 15140
rect 33638 15100 33663 15140
rect 33409 15077 33495 15100
rect 33577 15077 33663 15100
rect 48529 15140 48615 15163
rect 48697 15140 48783 15163
rect 48529 15100 48554 15140
rect 48554 15100 48594 15140
rect 48594 15100 48615 15140
rect 48697 15100 48718 15140
rect 48718 15100 48758 15140
rect 48758 15100 48783 15140
rect 48529 15077 48615 15100
rect 48697 15077 48783 15100
rect 63649 15140 63735 15163
rect 63817 15140 63903 15163
rect 63649 15100 63674 15140
rect 63674 15100 63714 15140
rect 63714 15100 63735 15140
rect 63817 15100 63838 15140
rect 63838 15100 63878 15140
rect 63878 15100 63903 15140
rect 63649 15077 63735 15100
rect 63817 15077 63903 15100
rect 78769 15140 78855 15163
rect 78937 15140 79023 15163
rect 78769 15100 78794 15140
rect 78794 15100 78834 15140
rect 78834 15100 78855 15140
rect 78937 15100 78958 15140
rect 78958 15100 78998 15140
rect 78998 15100 79023 15140
rect 78769 15077 78855 15100
rect 78937 15077 79023 15100
rect 93889 15140 93975 15163
rect 94057 15140 94143 15163
rect 93889 15100 93914 15140
rect 93914 15100 93954 15140
rect 93954 15100 93975 15140
rect 94057 15100 94078 15140
rect 94078 15100 94118 15140
rect 94118 15100 94143 15140
rect 93889 15077 93975 15100
rect 94057 15077 94143 15100
rect 4409 14384 4495 14407
rect 4577 14384 4663 14407
rect 4409 14344 4434 14384
rect 4434 14344 4474 14384
rect 4474 14344 4495 14384
rect 4577 14344 4598 14384
rect 4598 14344 4638 14384
rect 4638 14344 4663 14384
rect 4409 14321 4495 14344
rect 4577 14321 4663 14344
rect 19529 14384 19615 14407
rect 19697 14384 19783 14407
rect 19529 14344 19554 14384
rect 19554 14344 19594 14384
rect 19594 14344 19615 14384
rect 19697 14344 19718 14384
rect 19718 14344 19758 14384
rect 19758 14344 19783 14384
rect 19529 14321 19615 14344
rect 19697 14321 19783 14344
rect 34649 14384 34735 14407
rect 34817 14384 34903 14407
rect 34649 14344 34674 14384
rect 34674 14344 34714 14384
rect 34714 14344 34735 14384
rect 34817 14344 34838 14384
rect 34838 14344 34878 14384
rect 34878 14344 34903 14384
rect 34649 14321 34735 14344
rect 34817 14321 34903 14344
rect 49769 14384 49855 14407
rect 49937 14384 50023 14407
rect 49769 14344 49794 14384
rect 49794 14344 49834 14384
rect 49834 14344 49855 14384
rect 49937 14344 49958 14384
rect 49958 14344 49998 14384
rect 49998 14344 50023 14384
rect 49769 14321 49855 14344
rect 49937 14321 50023 14344
rect 64889 14384 64975 14407
rect 65057 14384 65143 14407
rect 64889 14344 64914 14384
rect 64914 14344 64954 14384
rect 64954 14344 64975 14384
rect 65057 14344 65078 14384
rect 65078 14344 65118 14384
rect 65118 14344 65143 14384
rect 64889 14321 64975 14344
rect 65057 14321 65143 14344
rect 80009 14384 80095 14407
rect 80177 14384 80263 14407
rect 80009 14344 80034 14384
rect 80034 14344 80074 14384
rect 80074 14344 80095 14384
rect 80177 14344 80198 14384
rect 80198 14344 80238 14384
rect 80238 14344 80263 14384
rect 80009 14321 80095 14344
rect 80177 14321 80263 14344
rect 95129 14384 95215 14407
rect 95297 14384 95383 14407
rect 95129 14344 95154 14384
rect 95154 14344 95194 14384
rect 95194 14344 95215 14384
rect 95297 14344 95318 14384
rect 95318 14344 95358 14384
rect 95358 14344 95383 14384
rect 95129 14321 95215 14344
rect 95297 14321 95383 14344
rect 3169 13628 3255 13651
rect 3337 13628 3423 13651
rect 3169 13588 3194 13628
rect 3194 13588 3234 13628
rect 3234 13588 3255 13628
rect 3337 13588 3358 13628
rect 3358 13588 3398 13628
rect 3398 13588 3423 13628
rect 3169 13565 3255 13588
rect 3337 13565 3423 13588
rect 18289 13628 18375 13651
rect 18457 13628 18543 13651
rect 18289 13588 18314 13628
rect 18314 13588 18354 13628
rect 18354 13588 18375 13628
rect 18457 13588 18478 13628
rect 18478 13588 18518 13628
rect 18518 13588 18543 13628
rect 18289 13565 18375 13588
rect 18457 13565 18543 13588
rect 33409 13628 33495 13651
rect 33577 13628 33663 13651
rect 33409 13588 33434 13628
rect 33434 13588 33474 13628
rect 33474 13588 33495 13628
rect 33577 13588 33598 13628
rect 33598 13588 33638 13628
rect 33638 13588 33663 13628
rect 33409 13565 33495 13588
rect 33577 13565 33663 13588
rect 48529 13628 48615 13651
rect 48697 13628 48783 13651
rect 48529 13588 48554 13628
rect 48554 13588 48594 13628
rect 48594 13588 48615 13628
rect 48697 13588 48718 13628
rect 48718 13588 48758 13628
rect 48758 13588 48783 13628
rect 48529 13565 48615 13588
rect 48697 13565 48783 13588
rect 63649 13628 63735 13651
rect 63817 13628 63903 13651
rect 63649 13588 63674 13628
rect 63674 13588 63714 13628
rect 63714 13588 63735 13628
rect 63817 13588 63838 13628
rect 63838 13588 63878 13628
rect 63878 13588 63903 13628
rect 63649 13565 63735 13588
rect 63817 13565 63903 13588
rect 78769 13628 78855 13651
rect 78937 13628 79023 13651
rect 78769 13588 78794 13628
rect 78794 13588 78834 13628
rect 78834 13588 78855 13628
rect 78937 13588 78958 13628
rect 78958 13588 78998 13628
rect 78998 13588 79023 13628
rect 78769 13565 78855 13588
rect 78937 13565 79023 13588
rect 93889 13628 93975 13651
rect 94057 13628 94143 13651
rect 93889 13588 93914 13628
rect 93914 13588 93954 13628
rect 93954 13588 93975 13628
rect 94057 13588 94078 13628
rect 94078 13588 94118 13628
rect 94118 13588 94143 13628
rect 93889 13565 93975 13588
rect 94057 13565 94143 13588
rect 4409 12872 4495 12895
rect 4577 12872 4663 12895
rect 4409 12832 4434 12872
rect 4434 12832 4474 12872
rect 4474 12832 4495 12872
rect 4577 12832 4598 12872
rect 4598 12832 4638 12872
rect 4638 12832 4663 12872
rect 4409 12809 4495 12832
rect 4577 12809 4663 12832
rect 19529 12872 19615 12895
rect 19697 12872 19783 12895
rect 19529 12832 19554 12872
rect 19554 12832 19594 12872
rect 19594 12832 19615 12872
rect 19697 12832 19718 12872
rect 19718 12832 19758 12872
rect 19758 12832 19783 12872
rect 19529 12809 19615 12832
rect 19697 12809 19783 12832
rect 34649 12872 34735 12895
rect 34817 12872 34903 12895
rect 34649 12832 34674 12872
rect 34674 12832 34714 12872
rect 34714 12832 34735 12872
rect 34817 12832 34838 12872
rect 34838 12832 34878 12872
rect 34878 12832 34903 12872
rect 34649 12809 34735 12832
rect 34817 12809 34903 12832
rect 49769 12872 49855 12895
rect 49937 12872 50023 12895
rect 49769 12832 49794 12872
rect 49794 12832 49834 12872
rect 49834 12832 49855 12872
rect 49937 12832 49958 12872
rect 49958 12832 49998 12872
rect 49998 12832 50023 12872
rect 49769 12809 49855 12832
rect 49937 12809 50023 12832
rect 64889 12872 64975 12895
rect 65057 12872 65143 12895
rect 64889 12832 64914 12872
rect 64914 12832 64954 12872
rect 64954 12832 64975 12872
rect 65057 12832 65078 12872
rect 65078 12832 65118 12872
rect 65118 12832 65143 12872
rect 64889 12809 64975 12832
rect 65057 12809 65143 12832
rect 80009 12872 80095 12895
rect 80177 12872 80263 12895
rect 80009 12832 80034 12872
rect 80034 12832 80074 12872
rect 80074 12832 80095 12872
rect 80177 12832 80198 12872
rect 80198 12832 80238 12872
rect 80238 12832 80263 12872
rect 80009 12809 80095 12832
rect 80177 12809 80263 12832
rect 95129 12872 95215 12895
rect 95297 12872 95383 12895
rect 95129 12832 95154 12872
rect 95154 12832 95194 12872
rect 95194 12832 95215 12872
rect 95297 12832 95318 12872
rect 95318 12832 95358 12872
rect 95358 12832 95383 12872
rect 95129 12809 95215 12832
rect 95297 12809 95383 12832
rect 3169 12116 3255 12139
rect 3337 12116 3423 12139
rect 3169 12076 3194 12116
rect 3194 12076 3234 12116
rect 3234 12076 3255 12116
rect 3337 12076 3358 12116
rect 3358 12076 3398 12116
rect 3398 12076 3423 12116
rect 3169 12053 3255 12076
rect 3337 12053 3423 12076
rect 18289 12116 18375 12139
rect 18457 12116 18543 12139
rect 18289 12076 18314 12116
rect 18314 12076 18354 12116
rect 18354 12076 18375 12116
rect 18457 12076 18478 12116
rect 18478 12076 18518 12116
rect 18518 12076 18543 12116
rect 18289 12053 18375 12076
rect 18457 12053 18543 12076
rect 33409 12116 33495 12139
rect 33577 12116 33663 12139
rect 33409 12076 33434 12116
rect 33434 12076 33474 12116
rect 33474 12076 33495 12116
rect 33577 12076 33598 12116
rect 33598 12076 33638 12116
rect 33638 12076 33663 12116
rect 33409 12053 33495 12076
rect 33577 12053 33663 12076
rect 48529 12116 48615 12139
rect 48697 12116 48783 12139
rect 48529 12076 48554 12116
rect 48554 12076 48594 12116
rect 48594 12076 48615 12116
rect 48697 12076 48718 12116
rect 48718 12076 48758 12116
rect 48758 12076 48783 12116
rect 48529 12053 48615 12076
rect 48697 12053 48783 12076
rect 63649 12116 63735 12139
rect 63817 12116 63903 12139
rect 63649 12076 63674 12116
rect 63674 12076 63714 12116
rect 63714 12076 63735 12116
rect 63817 12076 63838 12116
rect 63838 12076 63878 12116
rect 63878 12076 63903 12116
rect 63649 12053 63735 12076
rect 63817 12053 63903 12076
rect 78769 12116 78855 12139
rect 78937 12116 79023 12139
rect 78769 12076 78794 12116
rect 78794 12076 78834 12116
rect 78834 12076 78855 12116
rect 78937 12076 78958 12116
rect 78958 12076 78998 12116
rect 78998 12076 79023 12116
rect 78769 12053 78855 12076
rect 78937 12053 79023 12076
rect 93889 12116 93975 12139
rect 94057 12116 94143 12139
rect 93889 12076 93914 12116
rect 93914 12076 93954 12116
rect 93954 12076 93975 12116
rect 94057 12076 94078 12116
rect 94078 12076 94118 12116
rect 94118 12076 94143 12116
rect 93889 12053 93975 12076
rect 94057 12053 94143 12076
rect 4409 11360 4495 11383
rect 4577 11360 4663 11383
rect 4409 11320 4434 11360
rect 4434 11320 4474 11360
rect 4474 11320 4495 11360
rect 4577 11320 4598 11360
rect 4598 11320 4638 11360
rect 4638 11320 4663 11360
rect 4409 11297 4495 11320
rect 4577 11297 4663 11320
rect 19529 11360 19615 11383
rect 19697 11360 19783 11383
rect 19529 11320 19554 11360
rect 19554 11320 19594 11360
rect 19594 11320 19615 11360
rect 19697 11320 19718 11360
rect 19718 11320 19758 11360
rect 19758 11320 19783 11360
rect 19529 11297 19615 11320
rect 19697 11297 19783 11320
rect 34649 11360 34735 11383
rect 34817 11360 34903 11383
rect 34649 11320 34674 11360
rect 34674 11320 34714 11360
rect 34714 11320 34735 11360
rect 34817 11320 34838 11360
rect 34838 11320 34878 11360
rect 34878 11320 34903 11360
rect 34649 11297 34735 11320
rect 34817 11297 34903 11320
rect 49769 11360 49855 11383
rect 49937 11360 50023 11383
rect 49769 11320 49794 11360
rect 49794 11320 49834 11360
rect 49834 11320 49855 11360
rect 49937 11320 49958 11360
rect 49958 11320 49998 11360
rect 49998 11320 50023 11360
rect 49769 11297 49855 11320
rect 49937 11297 50023 11320
rect 64889 11360 64975 11383
rect 65057 11360 65143 11383
rect 64889 11320 64914 11360
rect 64914 11320 64954 11360
rect 64954 11320 64975 11360
rect 65057 11320 65078 11360
rect 65078 11320 65118 11360
rect 65118 11320 65143 11360
rect 64889 11297 64975 11320
rect 65057 11297 65143 11320
rect 80009 11360 80095 11383
rect 80177 11360 80263 11383
rect 80009 11320 80034 11360
rect 80034 11320 80074 11360
rect 80074 11320 80095 11360
rect 80177 11320 80198 11360
rect 80198 11320 80238 11360
rect 80238 11320 80263 11360
rect 80009 11297 80095 11320
rect 80177 11297 80263 11320
rect 95129 11360 95215 11383
rect 95297 11360 95383 11383
rect 95129 11320 95154 11360
rect 95154 11320 95194 11360
rect 95194 11320 95215 11360
rect 95297 11320 95318 11360
rect 95318 11320 95358 11360
rect 95358 11320 95383 11360
rect 95129 11297 95215 11320
rect 95297 11297 95383 11320
rect 3169 10604 3255 10627
rect 3337 10604 3423 10627
rect 3169 10564 3194 10604
rect 3194 10564 3234 10604
rect 3234 10564 3255 10604
rect 3337 10564 3358 10604
rect 3358 10564 3398 10604
rect 3398 10564 3423 10604
rect 3169 10541 3255 10564
rect 3337 10541 3423 10564
rect 18289 10604 18375 10627
rect 18457 10604 18543 10627
rect 18289 10564 18314 10604
rect 18314 10564 18354 10604
rect 18354 10564 18375 10604
rect 18457 10564 18478 10604
rect 18478 10564 18518 10604
rect 18518 10564 18543 10604
rect 18289 10541 18375 10564
rect 18457 10541 18543 10564
rect 33409 10604 33495 10627
rect 33577 10604 33663 10627
rect 33409 10564 33434 10604
rect 33434 10564 33474 10604
rect 33474 10564 33495 10604
rect 33577 10564 33598 10604
rect 33598 10564 33638 10604
rect 33638 10564 33663 10604
rect 33409 10541 33495 10564
rect 33577 10541 33663 10564
rect 48529 10604 48615 10627
rect 48697 10604 48783 10627
rect 48529 10564 48554 10604
rect 48554 10564 48594 10604
rect 48594 10564 48615 10604
rect 48697 10564 48718 10604
rect 48718 10564 48758 10604
rect 48758 10564 48783 10604
rect 48529 10541 48615 10564
rect 48697 10541 48783 10564
rect 63649 10604 63735 10627
rect 63817 10604 63903 10627
rect 63649 10564 63674 10604
rect 63674 10564 63714 10604
rect 63714 10564 63735 10604
rect 63817 10564 63838 10604
rect 63838 10564 63878 10604
rect 63878 10564 63903 10604
rect 63649 10541 63735 10564
rect 63817 10541 63903 10564
rect 78769 10604 78855 10627
rect 78937 10604 79023 10627
rect 78769 10564 78794 10604
rect 78794 10564 78834 10604
rect 78834 10564 78855 10604
rect 78937 10564 78958 10604
rect 78958 10564 78998 10604
rect 78998 10564 79023 10604
rect 78769 10541 78855 10564
rect 78937 10541 79023 10564
rect 93889 10604 93975 10627
rect 94057 10604 94143 10627
rect 93889 10564 93914 10604
rect 93914 10564 93954 10604
rect 93954 10564 93975 10604
rect 94057 10564 94078 10604
rect 94078 10564 94118 10604
rect 94118 10564 94143 10604
rect 93889 10541 93975 10564
rect 94057 10541 94143 10564
rect 4409 9848 4495 9871
rect 4577 9848 4663 9871
rect 4409 9808 4434 9848
rect 4434 9808 4474 9848
rect 4474 9808 4495 9848
rect 4577 9808 4598 9848
rect 4598 9808 4638 9848
rect 4638 9808 4663 9848
rect 4409 9785 4495 9808
rect 4577 9785 4663 9808
rect 19529 9848 19615 9871
rect 19697 9848 19783 9871
rect 19529 9808 19554 9848
rect 19554 9808 19594 9848
rect 19594 9808 19615 9848
rect 19697 9808 19718 9848
rect 19718 9808 19758 9848
rect 19758 9808 19783 9848
rect 19529 9785 19615 9808
rect 19697 9785 19783 9808
rect 34649 9848 34735 9871
rect 34817 9848 34903 9871
rect 34649 9808 34674 9848
rect 34674 9808 34714 9848
rect 34714 9808 34735 9848
rect 34817 9808 34838 9848
rect 34838 9808 34878 9848
rect 34878 9808 34903 9848
rect 34649 9785 34735 9808
rect 34817 9785 34903 9808
rect 49769 9848 49855 9871
rect 49937 9848 50023 9871
rect 49769 9808 49794 9848
rect 49794 9808 49834 9848
rect 49834 9808 49855 9848
rect 49937 9808 49958 9848
rect 49958 9808 49998 9848
rect 49998 9808 50023 9848
rect 49769 9785 49855 9808
rect 49937 9785 50023 9808
rect 64889 9848 64975 9871
rect 65057 9848 65143 9871
rect 64889 9808 64914 9848
rect 64914 9808 64954 9848
rect 64954 9808 64975 9848
rect 65057 9808 65078 9848
rect 65078 9808 65118 9848
rect 65118 9808 65143 9848
rect 64889 9785 64975 9808
rect 65057 9785 65143 9808
rect 80009 9848 80095 9871
rect 80177 9848 80263 9871
rect 80009 9808 80034 9848
rect 80034 9808 80074 9848
rect 80074 9808 80095 9848
rect 80177 9808 80198 9848
rect 80198 9808 80238 9848
rect 80238 9808 80263 9848
rect 80009 9785 80095 9808
rect 80177 9785 80263 9808
rect 95129 9848 95215 9871
rect 95297 9848 95383 9871
rect 95129 9808 95154 9848
rect 95154 9808 95194 9848
rect 95194 9808 95215 9848
rect 95297 9808 95318 9848
rect 95318 9808 95358 9848
rect 95358 9808 95383 9848
rect 95129 9785 95215 9808
rect 95297 9785 95383 9808
rect 3169 9092 3255 9115
rect 3337 9092 3423 9115
rect 3169 9052 3194 9092
rect 3194 9052 3234 9092
rect 3234 9052 3255 9092
rect 3337 9052 3358 9092
rect 3358 9052 3398 9092
rect 3398 9052 3423 9092
rect 3169 9029 3255 9052
rect 3337 9029 3423 9052
rect 18289 9092 18375 9115
rect 18457 9092 18543 9115
rect 18289 9052 18314 9092
rect 18314 9052 18354 9092
rect 18354 9052 18375 9092
rect 18457 9052 18478 9092
rect 18478 9052 18518 9092
rect 18518 9052 18543 9092
rect 18289 9029 18375 9052
rect 18457 9029 18543 9052
rect 33409 9092 33495 9115
rect 33577 9092 33663 9115
rect 33409 9052 33434 9092
rect 33434 9052 33474 9092
rect 33474 9052 33495 9092
rect 33577 9052 33598 9092
rect 33598 9052 33638 9092
rect 33638 9052 33663 9092
rect 33409 9029 33495 9052
rect 33577 9029 33663 9052
rect 48529 9092 48615 9115
rect 48697 9092 48783 9115
rect 48529 9052 48554 9092
rect 48554 9052 48594 9092
rect 48594 9052 48615 9092
rect 48697 9052 48718 9092
rect 48718 9052 48758 9092
rect 48758 9052 48783 9092
rect 48529 9029 48615 9052
rect 48697 9029 48783 9052
rect 63649 9092 63735 9115
rect 63817 9092 63903 9115
rect 63649 9052 63674 9092
rect 63674 9052 63714 9092
rect 63714 9052 63735 9092
rect 63817 9052 63838 9092
rect 63838 9052 63878 9092
rect 63878 9052 63903 9092
rect 63649 9029 63735 9052
rect 63817 9029 63903 9052
rect 78769 9092 78855 9115
rect 78937 9092 79023 9115
rect 78769 9052 78794 9092
rect 78794 9052 78834 9092
rect 78834 9052 78855 9092
rect 78937 9052 78958 9092
rect 78958 9052 78998 9092
rect 78998 9052 79023 9092
rect 78769 9029 78855 9052
rect 78937 9029 79023 9052
rect 93889 9092 93975 9115
rect 94057 9092 94143 9115
rect 93889 9052 93914 9092
rect 93914 9052 93954 9092
rect 93954 9052 93975 9092
rect 94057 9052 94078 9092
rect 94078 9052 94118 9092
rect 94118 9052 94143 9092
rect 93889 9029 93975 9052
rect 94057 9029 94143 9052
rect 4409 8336 4495 8359
rect 4577 8336 4663 8359
rect 4409 8296 4434 8336
rect 4434 8296 4474 8336
rect 4474 8296 4495 8336
rect 4577 8296 4598 8336
rect 4598 8296 4638 8336
rect 4638 8296 4663 8336
rect 4409 8273 4495 8296
rect 4577 8273 4663 8296
rect 19529 8336 19615 8359
rect 19697 8336 19783 8359
rect 19529 8296 19554 8336
rect 19554 8296 19594 8336
rect 19594 8296 19615 8336
rect 19697 8296 19718 8336
rect 19718 8296 19758 8336
rect 19758 8296 19783 8336
rect 19529 8273 19615 8296
rect 19697 8273 19783 8296
rect 34649 8336 34735 8359
rect 34817 8336 34903 8359
rect 34649 8296 34674 8336
rect 34674 8296 34714 8336
rect 34714 8296 34735 8336
rect 34817 8296 34838 8336
rect 34838 8296 34878 8336
rect 34878 8296 34903 8336
rect 34649 8273 34735 8296
rect 34817 8273 34903 8296
rect 49769 8336 49855 8359
rect 49937 8336 50023 8359
rect 49769 8296 49794 8336
rect 49794 8296 49834 8336
rect 49834 8296 49855 8336
rect 49937 8296 49958 8336
rect 49958 8296 49998 8336
rect 49998 8296 50023 8336
rect 49769 8273 49855 8296
rect 49937 8273 50023 8296
rect 64889 8336 64975 8359
rect 65057 8336 65143 8359
rect 64889 8296 64914 8336
rect 64914 8296 64954 8336
rect 64954 8296 64975 8336
rect 65057 8296 65078 8336
rect 65078 8296 65118 8336
rect 65118 8296 65143 8336
rect 64889 8273 64975 8296
rect 65057 8273 65143 8296
rect 80009 8336 80095 8359
rect 80177 8336 80263 8359
rect 80009 8296 80034 8336
rect 80034 8296 80074 8336
rect 80074 8296 80095 8336
rect 80177 8296 80198 8336
rect 80198 8296 80238 8336
rect 80238 8296 80263 8336
rect 80009 8273 80095 8296
rect 80177 8273 80263 8296
rect 95129 8336 95215 8359
rect 95297 8336 95383 8359
rect 95129 8296 95154 8336
rect 95154 8296 95194 8336
rect 95194 8296 95215 8336
rect 95297 8296 95318 8336
rect 95318 8296 95358 8336
rect 95358 8296 95383 8336
rect 95129 8273 95215 8296
rect 95297 8273 95383 8296
rect 3169 7580 3255 7603
rect 3337 7580 3423 7603
rect 3169 7540 3194 7580
rect 3194 7540 3234 7580
rect 3234 7540 3255 7580
rect 3337 7540 3358 7580
rect 3358 7540 3398 7580
rect 3398 7540 3423 7580
rect 3169 7517 3255 7540
rect 3337 7517 3423 7540
rect 18289 7580 18375 7603
rect 18457 7580 18543 7603
rect 18289 7540 18314 7580
rect 18314 7540 18354 7580
rect 18354 7540 18375 7580
rect 18457 7540 18478 7580
rect 18478 7540 18518 7580
rect 18518 7540 18543 7580
rect 18289 7517 18375 7540
rect 18457 7517 18543 7540
rect 33409 7580 33495 7603
rect 33577 7580 33663 7603
rect 33409 7540 33434 7580
rect 33434 7540 33474 7580
rect 33474 7540 33495 7580
rect 33577 7540 33598 7580
rect 33598 7540 33638 7580
rect 33638 7540 33663 7580
rect 33409 7517 33495 7540
rect 33577 7517 33663 7540
rect 48529 7580 48615 7603
rect 48697 7580 48783 7603
rect 48529 7540 48554 7580
rect 48554 7540 48594 7580
rect 48594 7540 48615 7580
rect 48697 7540 48718 7580
rect 48718 7540 48758 7580
rect 48758 7540 48783 7580
rect 48529 7517 48615 7540
rect 48697 7517 48783 7540
rect 63649 7580 63735 7603
rect 63817 7580 63903 7603
rect 63649 7540 63674 7580
rect 63674 7540 63714 7580
rect 63714 7540 63735 7580
rect 63817 7540 63838 7580
rect 63838 7540 63878 7580
rect 63878 7540 63903 7580
rect 63649 7517 63735 7540
rect 63817 7517 63903 7540
rect 78769 7580 78855 7603
rect 78937 7580 79023 7603
rect 78769 7540 78794 7580
rect 78794 7540 78834 7580
rect 78834 7540 78855 7580
rect 78937 7540 78958 7580
rect 78958 7540 78998 7580
rect 78998 7540 79023 7580
rect 78769 7517 78855 7540
rect 78937 7517 79023 7540
rect 93889 7580 93975 7603
rect 94057 7580 94143 7603
rect 93889 7540 93914 7580
rect 93914 7540 93954 7580
rect 93954 7540 93975 7580
rect 94057 7540 94078 7580
rect 94078 7540 94118 7580
rect 94118 7540 94143 7580
rect 93889 7517 93975 7540
rect 94057 7517 94143 7540
rect 4409 6824 4495 6847
rect 4577 6824 4663 6847
rect 4409 6784 4434 6824
rect 4434 6784 4474 6824
rect 4474 6784 4495 6824
rect 4577 6784 4598 6824
rect 4598 6784 4638 6824
rect 4638 6784 4663 6824
rect 4409 6761 4495 6784
rect 4577 6761 4663 6784
rect 19529 6824 19615 6847
rect 19697 6824 19783 6847
rect 19529 6784 19554 6824
rect 19554 6784 19594 6824
rect 19594 6784 19615 6824
rect 19697 6784 19718 6824
rect 19718 6784 19758 6824
rect 19758 6784 19783 6824
rect 19529 6761 19615 6784
rect 19697 6761 19783 6784
rect 34649 6824 34735 6847
rect 34817 6824 34903 6847
rect 34649 6784 34674 6824
rect 34674 6784 34714 6824
rect 34714 6784 34735 6824
rect 34817 6784 34838 6824
rect 34838 6784 34878 6824
rect 34878 6784 34903 6824
rect 34649 6761 34735 6784
rect 34817 6761 34903 6784
rect 49769 6824 49855 6847
rect 49937 6824 50023 6847
rect 49769 6784 49794 6824
rect 49794 6784 49834 6824
rect 49834 6784 49855 6824
rect 49937 6784 49958 6824
rect 49958 6784 49998 6824
rect 49998 6784 50023 6824
rect 49769 6761 49855 6784
rect 49937 6761 50023 6784
rect 64889 6824 64975 6847
rect 65057 6824 65143 6847
rect 64889 6784 64914 6824
rect 64914 6784 64954 6824
rect 64954 6784 64975 6824
rect 65057 6784 65078 6824
rect 65078 6784 65118 6824
rect 65118 6784 65143 6824
rect 64889 6761 64975 6784
rect 65057 6761 65143 6784
rect 80009 6824 80095 6847
rect 80177 6824 80263 6847
rect 80009 6784 80034 6824
rect 80034 6784 80074 6824
rect 80074 6784 80095 6824
rect 80177 6784 80198 6824
rect 80198 6784 80238 6824
rect 80238 6784 80263 6824
rect 80009 6761 80095 6784
rect 80177 6761 80263 6784
rect 95129 6824 95215 6847
rect 95297 6824 95383 6847
rect 95129 6784 95154 6824
rect 95154 6784 95194 6824
rect 95194 6784 95215 6824
rect 95297 6784 95318 6824
rect 95318 6784 95358 6824
rect 95358 6784 95383 6824
rect 95129 6761 95215 6784
rect 95297 6761 95383 6784
rect 3169 6068 3255 6091
rect 3337 6068 3423 6091
rect 3169 6028 3194 6068
rect 3194 6028 3234 6068
rect 3234 6028 3255 6068
rect 3337 6028 3358 6068
rect 3358 6028 3398 6068
rect 3398 6028 3423 6068
rect 3169 6005 3255 6028
rect 3337 6005 3423 6028
rect 18289 6068 18375 6091
rect 18457 6068 18543 6091
rect 18289 6028 18314 6068
rect 18314 6028 18354 6068
rect 18354 6028 18375 6068
rect 18457 6028 18478 6068
rect 18478 6028 18518 6068
rect 18518 6028 18543 6068
rect 18289 6005 18375 6028
rect 18457 6005 18543 6028
rect 33409 6068 33495 6091
rect 33577 6068 33663 6091
rect 33409 6028 33434 6068
rect 33434 6028 33474 6068
rect 33474 6028 33495 6068
rect 33577 6028 33598 6068
rect 33598 6028 33638 6068
rect 33638 6028 33663 6068
rect 33409 6005 33495 6028
rect 33577 6005 33663 6028
rect 48529 6068 48615 6091
rect 48697 6068 48783 6091
rect 48529 6028 48554 6068
rect 48554 6028 48594 6068
rect 48594 6028 48615 6068
rect 48697 6028 48718 6068
rect 48718 6028 48758 6068
rect 48758 6028 48783 6068
rect 48529 6005 48615 6028
rect 48697 6005 48783 6028
rect 63649 6068 63735 6091
rect 63817 6068 63903 6091
rect 63649 6028 63674 6068
rect 63674 6028 63714 6068
rect 63714 6028 63735 6068
rect 63817 6028 63838 6068
rect 63838 6028 63878 6068
rect 63878 6028 63903 6068
rect 63649 6005 63735 6028
rect 63817 6005 63903 6028
rect 78769 6068 78855 6091
rect 78937 6068 79023 6091
rect 78769 6028 78794 6068
rect 78794 6028 78834 6068
rect 78834 6028 78855 6068
rect 78937 6028 78958 6068
rect 78958 6028 78998 6068
rect 78998 6028 79023 6068
rect 78769 6005 78855 6028
rect 78937 6005 79023 6028
rect 93889 6068 93975 6091
rect 94057 6068 94143 6091
rect 93889 6028 93914 6068
rect 93914 6028 93954 6068
rect 93954 6028 93975 6068
rect 94057 6028 94078 6068
rect 94078 6028 94118 6068
rect 94118 6028 94143 6068
rect 93889 6005 93975 6028
rect 94057 6005 94143 6028
rect 4409 5312 4495 5335
rect 4577 5312 4663 5335
rect 4409 5272 4434 5312
rect 4434 5272 4474 5312
rect 4474 5272 4495 5312
rect 4577 5272 4598 5312
rect 4598 5272 4638 5312
rect 4638 5272 4663 5312
rect 4409 5249 4495 5272
rect 4577 5249 4663 5272
rect 19529 5312 19615 5335
rect 19697 5312 19783 5335
rect 19529 5272 19554 5312
rect 19554 5272 19594 5312
rect 19594 5272 19615 5312
rect 19697 5272 19718 5312
rect 19718 5272 19758 5312
rect 19758 5272 19783 5312
rect 19529 5249 19615 5272
rect 19697 5249 19783 5272
rect 34649 5312 34735 5335
rect 34817 5312 34903 5335
rect 34649 5272 34674 5312
rect 34674 5272 34714 5312
rect 34714 5272 34735 5312
rect 34817 5272 34838 5312
rect 34838 5272 34878 5312
rect 34878 5272 34903 5312
rect 34649 5249 34735 5272
rect 34817 5249 34903 5272
rect 49769 5312 49855 5335
rect 49937 5312 50023 5335
rect 49769 5272 49794 5312
rect 49794 5272 49834 5312
rect 49834 5272 49855 5312
rect 49937 5272 49958 5312
rect 49958 5272 49998 5312
rect 49998 5272 50023 5312
rect 49769 5249 49855 5272
rect 49937 5249 50023 5272
rect 64889 5312 64975 5335
rect 65057 5312 65143 5335
rect 64889 5272 64914 5312
rect 64914 5272 64954 5312
rect 64954 5272 64975 5312
rect 65057 5272 65078 5312
rect 65078 5272 65118 5312
rect 65118 5272 65143 5312
rect 64889 5249 64975 5272
rect 65057 5249 65143 5272
rect 80009 5312 80095 5335
rect 80177 5312 80263 5335
rect 80009 5272 80034 5312
rect 80034 5272 80074 5312
rect 80074 5272 80095 5312
rect 80177 5272 80198 5312
rect 80198 5272 80238 5312
rect 80238 5272 80263 5312
rect 80009 5249 80095 5272
rect 80177 5249 80263 5272
rect 95129 5312 95215 5335
rect 95297 5312 95383 5335
rect 95129 5272 95154 5312
rect 95154 5272 95194 5312
rect 95194 5272 95215 5312
rect 95297 5272 95318 5312
rect 95318 5272 95358 5312
rect 95358 5272 95383 5312
rect 95129 5249 95215 5272
rect 95297 5249 95383 5272
rect 3169 4556 3255 4579
rect 3337 4556 3423 4579
rect 3169 4516 3194 4556
rect 3194 4516 3234 4556
rect 3234 4516 3255 4556
rect 3337 4516 3358 4556
rect 3358 4516 3398 4556
rect 3398 4516 3423 4556
rect 3169 4493 3255 4516
rect 3337 4493 3423 4516
rect 18289 4556 18375 4579
rect 18457 4556 18543 4579
rect 18289 4516 18314 4556
rect 18314 4516 18354 4556
rect 18354 4516 18375 4556
rect 18457 4516 18478 4556
rect 18478 4516 18518 4556
rect 18518 4516 18543 4556
rect 18289 4493 18375 4516
rect 18457 4493 18543 4516
rect 33409 4556 33495 4579
rect 33577 4556 33663 4579
rect 33409 4516 33434 4556
rect 33434 4516 33474 4556
rect 33474 4516 33495 4556
rect 33577 4516 33598 4556
rect 33598 4516 33638 4556
rect 33638 4516 33663 4556
rect 33409 4493 33495 4516
rect 33577 4493 33663 4516
rect 48529 4556 48615 4579
rect 48697 4556 48783 4579
rect 48529 4516 48554 4556
rect 48554 4516 48594 4556
rect 48594 4516 48615 4556
rect 48697 4516 48718 4556
rect 48718 4516 48758 4556
rect 48758 4516 48783 4556
rect 48529 4493 48615 4516
rect 48697 4493 48783 4516
rect 63649 4556 63735 4579
rect 63817 4556 63903 4579
rect 63649 4516 63674 4556
rect 63674 4516 63714 4556
rect 63714 4516 63735 4556
rect 63817 4516 63838 4556
rect 63838 4516 63878 4556
rect 63878 4516 63903 4556
rect 63649 4493 63735 4516
rect 63817 4493 63903 4516
rect 78769 4556 78855 4579
rect 78937 4556 79023 4579
rect 78769 4516 78794 4556
rect 78794 4516 78834 4556
rect 78834 4516 78855 4556
rect 78937 4516 78958 4556
rect 78958 4516 78998 4556
rect 78998 4516 79023 4556
rect 78769 4493 78855 4516
rect 78937 4493 79023 4516
rect 93889 4556 93975 4579
rect 94057 4556 94143 4579
rect 93889 4516 93914 4556
rect 93914 4516 93954 4556
rect 93954 4516 93975 4556
rect 94057 4516 94078 4556
rect 94078 4516 94118 4556
rect 94118 4516 94143 4556
rect 93889 4493 93975 4516
rect 94057 4493 94143 4516
rect 4409 3800 4495 3823
rect 4577 3800 4663 3823
rect 4409 3760 4434 3800
rect 4434 3760 4474 3800
rect 4474 3760 4495 3800
rect 4577 3760 4598 3800
rect 4598 3760 4638 3800
rect 4638 3760 4663 3800
rect 4409 3737 4495 3760
rect 4577 3737 4663 3760
rect 19529 3800 19615 3823
rect 19697 3800 19783 3823
rect 19529 3760 19554 3800
rect 19554 3760 19594 3800
rect 19594 3760 19615 3800
rect 19697 3760 19718 3800
rect 19718 3760 19758 3800
rect 19758 3760 19783 3800
rect 19529 3737 19615 3760
rect 19697 3737 19783 3760
rect 34649 3800 34735 3823
rect 34817 3800 34903 3823
rect 34649 3760 34674 3800
rect 34674 3760 34714 3800
rect 34714 3760 34735 3800
rect 34817 3760 34838 3800
rect 34838 3760 34878 3800
rect 34878 3760 34903 3800
rect 34649 3737 34735 3760
rect 34817 3737 34903 3760
rect 49769 3800 49855 3823
rect 49937 3800 50023 3823
rect 49769 3760 49794 3800
rect 49794 3760 49834 3800
rect 49834 3760 49855 3800
rect 49937 3760 49958 3800
rect 49958 3760 49998 3800
rect 49998 3760 50023 3800
rect 49769 3737 49855 3760
rect 49937 3737 50023 3760
rect 64889 3800 64975 3823
rect 65057 3800 65143 3823
rect 64889 3760 64914 3800
rect 64914 3760 64954 3800
rect 64954 3760 64975 3800
rect 65057 3760 65078 3800
rect 65078 3760 65118 3800
rect 65118 3760 65143 3800
rect 64889 3737 64975 3760
rect 65057 3737 65143 3760
rect 80009 3800 80095 3823
rect 80177 3800 80263 3823
rect 80009 3760 80034 3800
rect 80034 3760 80074 3800
rect 80074 3760 80095 3800
rect 80177 3760 80198 3800
rect 80198 3760 80238 3800
rect 80238 3760 80263 3800
rect 80009 3737 80095 3760
rect 80177 3737 80263 3760
rect 95129 3800 95215 3823
rect 95297 3800 95383 3823
rect 95129 3760 95154 3800
rect 95154 3760 95194 3800
rect 95194 3760 95215 3800
rect 95297 3760 95318 3800
rect 95318 3760 95358 3800
rect 95358 3760 95383 3800
rect 95129 3737 95215 3760
rect 95297 3737 95383 3760
rect 3169 3044 3255 3067
rect 3337 3044 3423 3067
rect 3169 3004 3194 3044
rect 3194 3004 3234 3044
rect 3234 3004 3255 3044
rect 3337 3004 3358 3044
rect 3358 3004 3398 3044
rect 3398 3004 3423 3044
rect 3169 2981 3255 3004
rect 3337 2981 3423 3004
rect 18289 3044 18375 3067
rect 18457 3044 18543 3067
rect 18289 3004 18314 3044
rect 18314 3004 18354 3044
rect 18354 3004 18375 3044
rect 18457 3004 18478 3044
rect 18478 3004 18518 3044
rect 18518 3004 18543 3044
rect 18289 2981 18375 3004
rect 18457 2981 18543 3004
rect 33409 3044 33495 3067
rect 33577 3044 33663 3067
rect 33409 3004 33434 3044
rect 33434 3004 33474 3044
rect 33474 3004 33495 3044
rect 33577 3004 33598 3044
rect 33598 3004 33638 3044
rect 33638 3004 33663 3044
rect 33409 2981 33495 3004
rect 33577 2981 33663 3004
rect 48529 3044 48615 3067
rect 48697 3044 48783 3067
rect 48529 3004 48554 3044
rect 48554 3004 48594 3044
rect 48594 3004 48615 3044
rect 48697 3004 48718 3044
rect 48718 3004 48758 3044
rect 48758 3004 48783 3044
rect 48529 2981 48615 3004
rect 48697 2981 48783 3004
rect 63649 3044 63735 3067
rect 63817 3044 63903 3067
rect 63649 3004 63674 3044
rect 63674 3004 63714 3044
rect 63714 3004 63735 3044
rect 63817 3004 63838 3044
rect 63838 3004 63878 3044
rect 63878 3004 63903 3044
rect 63649 2981 63735 3004
rect 63817 2981 63903 3004
rect 78769 3044 78855 3067
rect 78937 3044 79023 3067
rect 78769 3004 78794 3044
rect 78794 3004 78834 3044
rect 78834 3004 78855 3044
rect 78937 3004 78958 3044
rect 78958 3004 78998 3044
rect 78998 3004 79023 3044
rect 78769 2981 78855 3004
rect 78937 2981 79023 3004
rect 93889 3044 93975 3067
rect 94057 3044 94143 3067
rect 93889 3004 93914 3044
rect 93914 3004 93954 3044
rect 93954 3004 93975 3044
rect 94057 3004 94078 3044
rect 94078 3004 94118 3044
rect 94118 3004 94143 3044
rect 93889 2981 93975 3004
rect 94057 2981 94143 3004
rect 4409 2288 4495 2311
rect 4577 2288 4663 2311
rect 4409 2248 4434 2288
rect 4434 2248 4474 2288
rect 4474 2248 4495 2288
rect 4577 2248 4598 2288
rect 4598 2248 4638 2288
rect 4638 2248 4663 2288
rect 4409 2225 4495 2248
rect 4577 2225 4663 2248
rect 19529 2288 19615 2311
rect 19697 2288 19783 2311
rect 19529 2248 19554 2288
rect 19554 2248 19594 2288
rect 19594 2248 19615 2288
rect 19697 2248 19718 2288
rect 19718 2248 19758 2288
rect 19758 2248 19783 2288
rect 19529 2225 19615 2248
rect 19697 2225 19783 2248
rect 34649 2288 34735 2311
rect 34817 2288 34903 2311
rect 34649 2248 34674 2288
rect 34674 2248 34714 2288
rect 34714 2248 34735 2288
rect 34817 2248 34838 2288
rect 34838 2248 34878 2288
rect 34878 2248 34903 2288
rect 34649 2225 34735 2248
rect 34817 2225 34903 2248
rect 49769 2288 49855 2311
rect 49937 2288 50023 2311
rect 49769 2248 49794 2288
rect 49794 2248 49834 2288
rect 49834 2248 49855 2288
rect 49937 2248 49958 2288
rect 49958 2248 49998 2288
rect 49998 2248 50023 2288
rect 49769 2225 49855 2248
rect 49937 2225 50023 2248
rect 64889 2288 64975 2311
rect 65057 2288 65143 2311
rect 64889 2248 64914 2288
rect 64914 2248 64954 2288
rect 64954 2248 64975 2288
rect 65057 2248 65078 2288
rect 65078 2248 65118 2288
rect 65118 2248 65143 2288
rect 64889 2225 64975 2248
rect 65057 2225 65143 2248
rect 80009 2288 80095 2311
rect 80177 2288 80263 2311
rect 80009 2248 80034 2288
rect 80034 2248 80074 2288
rect 80074 2248 80095 2288
rect 80177 2248 80198 2288
rect 80198 2248 80238 2288
rect 80238 2248 80263 2288
rect 80009 2225 80095 2248
rect 80177 2225 80263 2248
rect 95129 2288 95215 2311
rect 95297 2288 95383 2311
rect 95129 2248 95154 2288
rect 95154 2248 95194 2288
rect 95194 2248 95215 2288
rect 95297 2248 95318 2288
rect 95318 2248 95358 2288
rect 95358 2248 95383 2288
rect 95129 2225 95215 2248
rect 95297 2225 95383 2248
rect 3169 1532 3255 1555
rect 3337 1532 3423 1555
rect 3169 1492 3194 1532
rect 3194 1492 3234 1532
rect 3234 1492 3255 1532
rect 3337 1492 3358 1532
rect 3358 1492 3398 1532
rect 3398 1492 3423 1532
rect 3169 1469 3255 1492
rect 3337 1469 3423 1492
rect 18289 1532 18375 1555
rect 18457 1532 18543 1555
rect 18289 1492 18314 1532
rect 18314 1492 18354 1532
rect 18354 1492 18375 1532
rect 18457 1492 18478 1532
rect 18478 1492 18518 1532
rect 18518 1492 18543 1532
rect 18289 1469 18375 1492
rect 18457 1469 18543 1492
rect 33409 1532 33495 1555
rect 33577 1532 33663 1555
rect 33409 1492 33434 1532
rect 33434 1492 33474 1532
rect 33474 1492 33495 1532
rect 33577 1492 33598 1532
rect 33598 1492 33638 1532
rect 33638 1492 33663 1532
rect 33409 1469 33495 1492
rect 33577 1469 33663 1492
rect 48529 1532 48615 1555
rect 48697 1532 48783 1555
rect 48529 1492 48554 1532
rect 48554 1492 48594 1532
rect 48594 1492 48615 1532
rect 48697 1492 48718 1532
rect 48718 1492 48758 1532
rect 48758 1492 48783 1532
rect 48529 1469 48615 1492
rect 48697 1469 48783 1492
rect 63649 1532 63735 1555
rect 63817 1532 63903 1555
rect 63649 1492 63674 1532
rect 63674 1492 63714 1532
rect 63714 1492 63735 1532
rect 63817 1492 63838 1532
rect 63838 1492 63878 1532
rect 63878 1492 63903 1532
rect 63649 1469 63735 1492
rect 63817 1469 63903 1492
rect 78769 1532 78855 1555
rect 78937 1532 79023 1555
rect 78769 1492 78794 1532
rect 78794 1492 78834 1532
rect 78834 1492 78855 1532
rect 78937 1492 78958 1532
rect 78958 1492 78998 1532
rect 78998 1492 79023 1532
rect 78769 1469 78855 1492
rect 78937 1469 79023 1492
rect 93889 1532 93975 1555
rect 94057 1532 94143 1555
rect 93889 1492 93914 1532
rect 93914 1492 93954 1532
rect 93954 1492 93975 1532
rect 94057 1492 94078 1532
rect 94078 1492 94118 1532
rect 94118 1492 94143 1532
rect 93889 1469 93975 1492
rect 94057 1469 94143 1492
rect 4409 776 4495 799
rect 4577 776 4663 799
rect 4409 736 4434 776
rect 4434 736 4474 776
rect 4474 736 4495 776
rect 4577 736 4598 776
rect 4598 736 4638 776
rect 4638 736 4663 776
rect 4409 713 4495 736
rect 4577 713 4663 736
rect 19529 776 19615 799
rect 19697 776 19783 799
rect 19529 736 19554 776
rect 19554 736 19594 776
rect 19594 736 19615 776
rect 19697 736 19718 776
rect 19718 736 19758 776
rect 19758 736 19783 776
rect 19529 713 19615 736
rect 19697 713 19783 736
rect 34649 776 34735 799
rect 34817 776 34903 799
rect 34649 736 34674 776
rect 34674 736 34714 776
rect 34714 736 34735 776
rect 34817 736 34838 776
rect 34838 736 34878 776
rect 34878 736 34903 776
rect 34649 713 34735 736
rect 34817 713 34903 736
rect 49769 776 49855 799
rect 49937 776 50023 799
rect 49769 736 49794 776
rect 49794 736 49834 776
rect 49834 736 49855 776
rect 49937 736 49958 776
rect 49958 736 49998 776
rect 49998 736 50023 776
rect 49769 713 49855 736
rect 49937 713 50023 736
rect 64889 776 64975 799
rect 65057 776 65143 799
rect 64889 736 64914 776
rect 64914 736 64954 776
rect 64954 736 64975 776
rect 65057 736 65078 776
rect 65078 736 65118 776
rect 65118 736 65143 776
rect 64889 713 64975 736
rect 65057 713 65143 736
rect 80009 776 80095 799
rect 80177 776 80263 799
rect 80009 736 80034 776
rect 80034 736 80074 776
rect 80074 736 80095 776
rect 80177 736 80198 776
rect 80198 736 80238 776
rect 80238 736 80263 776
rect 80009 713 80095 736
rect 80177 713 80263 736
rect 95129 776 95215 799
rect 95297 776 95383 799
rect 95129 736 95154 776
rect 95154 736 95194 776
rect 95194 736 95215 776
rect 95297 736 95318 776
rect 95318 736 95358 776
rect 95358 736 95383 776
rect 95129 713 95215 736
rect 95297 713 95383 736
<< metal6 >>
rect 3076 37843 3516 38600
rect 3076 37757 3169 37843
rect 3255 37757 3337 37843
rect 3423 37757 3516 37843
rect 3076 36331 3516 37757
rect 3076 36245 3169 36331
rect 3255 36245 3337 36331
rect 3423 36245 3516 36331
rect 3076 34819 3516 36245
rect 3076 34733 3169 34819
rect 3255 34733 3337 34819
rect 3423 34733 3516 34819
rect 3076 33307 3516 34733
rect 3076 33221 3169 33307
rect 3255 33221 3337 33307
rect 3423 33221 3516 33307
rect 3076 31795 3516 33221
rect 3076 31709 3169 31795
rect 3255 31709 3337 31795
rect 3423 31709 3516 31795
rect 3076 30283 3516 31709
rect 3076 30197 3169 30283
rect 3255 30197 3337 30283
rect 3423 30197 3516 30283
rect 3076 28771 3516 30197
rect 3076 28685 3169 28771
rect 3255 28685 3337 28771
rect 3423 28685 3516 28771
rect 3076 27259 3516 28685
rect 3076 27173 3169 27259
rect 3255 27173 3337 27259
rect 3423 27173 3516 27259
rect 3076 25747 3516 27173
rect 3076 25661 3169 25747
rect 3255 25661 3337 25747
rect 3423 25661 3516 25747
rect 3076 24235 3516 25661
rect 3076 24149 3169 24235
rect 3255 24149 3337 24235
rect 3423 24149 3516 24235
rect 3076 22723 3516 24149
rect 3076 22637 3169 22723
rect 3255 22637 3337 22723
rect 3423 22637 3516 22723
rect 3076 21211 3516 22637
rect 3076 21125 3169 21211
rect 3255 21125 3337 21211
rect 3423 21125 3516 21211
rect 3076 19699 3516 21125
rect 3076 19613 3169 19699
rect 3255 19613 3337 19699
rect 3423 19613 3516 19699
rect 3076 18187 3516 19613
rect 3076 18101 3169 18187
rect 3255 18101 3337 18187
rect 3423 18101 3516 18187
rect 3076 16675 3516 18101
rect 3076 16589 3169 16675
rect 3255 16589 3337 16675
rect 3423 16589 3516 16675
rect 3076 15163 3516 16589
rect 3076 15077 3169 15163
rect 3255 15077 3337 15163
rect 3423 15077 3516 15163
rect 3076 13651 3516 15077
rect 3076 13565 3169 13651
rect 3255 13565 3337 13651
rect 3423 13565 3516 13651
rect 3076 12139 3516 13565
rect 3076 12053 3169 12139
rect 3255 12053 3337 12139
rect 3423 12053 3516 12139
rect 3076 10627 3516 12053
rect 3076 10541 3169 10627
rect 3255 10541 3337 10627
rect 3423 10541 3516 10627
rect 3076 9115 3516 10541
rect 3076 9029 3169 9115
rect 3255 9029 3337 9115
rect 3423 9029 3516 9115
rect 3076 7603 3516 9029
rect 3076 7517 3169 7603
rect 3255 7517 3337 7603
rect 3423 7517 3516 7603
rect 3076 6091 3516 7517
rect 3076 6005 3169 6091
rect 3255 6005 3337 6091
rect 3423 6005 3516 6091
rect 3076 4579 3516 6005
rect 3076 4493 3169 4579
rect 3255 4493 3337 4579
rect 3423 4493 3516 4579
rect 3076 3067 3516 4493
rect 3076 2981 3169 3067
rect 3255 2981 3337 3067
rect 3423 2981 3516 3067
rect 3076 1555 3516 2981
rect 3076 1469 3169 1555
rect 3255 1469 3337 1555
rect 3423 1469 3516 1555
rect 3076 712 3516 1469
rect 4316 38599 4756 38682
rect 4316 38513 4409 38599
rect 4495 38513 4577 38599
rect 4663 38513 4756 38599
rect 4316 37087 4756 38513
rect 4316 37001 4409 37087
rect 4495 37001 4577 37087
rect 4663 37001 4756 37087
rect 4316 35575 4756 37001
rect 4316 35489 4409 35575
rect 4495 35489 4577 35575
rect 4663 35489 4756 35575
rect 4316 34063 4756 35489
rect 4316 33977 4409 34063
rect 4495 33977 4577 34063
rect 4663 33977 4756 34063
rect 4316 32551 4756 33977
rect 4316 32465 4409 32551
rect 4495 32465 4577 32551
rect 4663 32465 4756 32551
rect 4316 31039 4756 32465
rect 4316 30953 4409 31039
rect 4495 30953 4577 31039
rect 4663 30953 4756 31039
rect 4316 29527 4756 30953
rect 4316 29441 4409 29527
rect 4495 29441 4577 29527
rect 4663 29441 4756 29527
rect 4316 28015 4756 29441
rect 4316 27929 4409 28015
rect 4495 27929 4577 28015
rect 4663 27929 4756 28015
rect 4316 26503 4756 27929
rect 4316 26417 4409 26503
rect 4495 26417 4577 26503
rect 4663 26417 4756 26503
rect 4316 24991 4756 26417
rect 4316 24905 4409 24991
rect 4495 24905 4577 24991
rect 4663 24905 4756 24991
rect 4316 23479 4756 24905
rect 4316 23393 4409 23479
rect 4495 23393 4577 23479
rect 4663 23393 4756 23479
rect 4316 21967 4756 23393
rect 4316 21881 4409 21967
rect 4495 21881 4577 21967
rect 4663 21881 4756 21967
rect 4316 20455 4756 21881
rect 4316 20369 4409 20455
rect 4495 20369 4577 20455
rect 4663 20369 4756 20455
rect 4316 18943 4756 20369
rect 4316 18857 4409 18943
rect 4495 18857 4577 18943
rect 4663 18857 4756 18943
rect 4316 17431 4756 18857
rect 4316 17345 4409 17431
rect 4495 17345 4577 17431
rect 4663 17345 4756 17431
rect 4316 15919 4756 17345
rect 4316 15833 4409 15919
rect 4495 15833 4577 15919
rect 4663 15833 4756 15919
rect 4316 14407 4756 15833
rect 4316 14321 4409 14407
rect 4495 14321 4577 14407
rect 4663 14321 4756 14407
rect 4316 12895 4756 14321
rect 4316 12809 4409 12895
rect 4495 12809 4577 12895
rect 4663 12809 4756 12895
rect 4316 11383 4756 12809
rect 4316 11297 4409 11383
rect 4495 11297 4577 11383
rect 4663 11297 4756 11383
rect 4316 9871 4756 11297
rect 4316 9785 4409 9871
rect 4495 9785 4577 9871
rect 4663 9785 4756 9871
rect 4316 8359 4756 9785
rect 4316 8273 4409 8359
rect 4495 8273 4577 8359
rect 4663 8273 4756 8359
rect 4316 6847 4756 8273
rect 4316 6761 4409 6847
rect 4495 6761 4577 6847
rect 4663 6761 4756 6847
rect 4316 5335 4756 6761
rect 4316 5249 4409 5335
rect 4495 5249 4577 5335
rect 4663 5249 4756 5335
rect 4316 3823 4756 5249
rect 4316 3737 4409 3823
rect 4495 3737 4577 3823
rect 4663 3737 4756 3823
rect 4316 2311 4756 3737
rect 4316 2225 4409 2311
rect 4495 2225 4577 2311
rect 4663 2225 4756 2311
rect 4316 799 4756 2225
rect 4316 713 4409 799
rect 4495 713 4577 799
rect 4663 713 4756 799
rect 4316 630 4756 713
rect 18196 37843 18636 38600
rect 18196 37757 18289 37843
rect 18375 37757 18457 37843
rect 18543 37757 18636 37843
rect 18196 36331 18636 37757
rect 18196 36245 18289 36331
rect 18375 36245 18457 36331
rect 18543 36245 18636 36331
rect 18196 34819 18636 36245
rect 18196 34733 18289 34819
rect 18375 34733 18457 34819
rect 18543 34733 18636 34819
rect 18196 33307 18636 34733
rect 18196 33221 18289 33307
rect 18375 33221 18457 33307
rect 18543 33221 18636 33307
rect 18196 31795 18636 33221
rect 18196 31709 18289 31795
rect 18375 31709 18457 31795
rect 18543 31709 18636 31795
rect 18196 30283 18636 31709
rect 18196 30197 18289 30283
rect 18375 30197 18457 30283
rect 18543 30197 18636 30283
rect 18196 28771 18636 30197
rect 18196 28685 18289 28771
rect 18375 28685 18457 28771
rect 18543 28685 18636 28771
rect 18196 27259 18636 28685
rect 18196 27173 18289 27259
rect 18375 27173 18457 27259
rect 18543 27173 18636 27259
rect 18196 25747 18636 27173
rect 18196 25661 18289 25747
rect 18375 25661 18457 25747
rect 18543 25661 18636 25747
rect 18196 24235 18636 25661
rect 18196 24149 18289 24235
rect 18375 24149 18457 24235
rect 18543 24149 18636 24235
rect 18196 22723 18636 24149
rect 18196 22637 18289 22723
rect 18375 22637 18457 22723
rect 18543 22637 18636 22723
rect 18196 21211 18636 22637
rect 18196 21125 18289 21211
rect 18375 21125 18457 21211
rect 18543 21125 18636 21211
rect 18196 19699 18636 21125
rect 18196 19613 18289 19699
rect 18375 19613 18457 19699
rect 18543 19613 18636 19699
rect 18196 18187 18636 19613
rect 18196 18101 18289 18187
rect 18375 18101 18457 18187
rect 18543 18101 18636 18187
rect 18196 16675 18636 18101
rect 18196 16589 18289 16675
rect 18375 16589 18457 16675
rect 18543 16589 18636 16675
rect 18196 15163 18636 16589
rect 18196 15077 18289 15163
rect 18375 15077 18457 15163
rect 18543 15077 18636 15163
rect 18196 13651 18636 15077
rect 18196 13565 18289 13651
rect 18375 13565 18457 13651
rect 18543 13565 18636 13651
rect 18196 12139 18636 13565
rect 18196 12053 18289 12139
rect 18375 12053 18457 12139
rect 18543 12053 18636 12139
rect 18196 10627 18636 12053
rect 18196 10541 18289 10627
rect 18375 10541 18457 10627
rect 18543 10541 18636 10627
rect 18196 9115 18636 10541
rect 18196 9029 18289 9115
rect 18375 9029 18457 9115
rect 18543 9029 18636 9115
rect 18196 7603 18636 9029
rect 18196 7517 18289 7603
rect 18375 7517 18457 7603
rect 18543 7517 18636 7603
rect 18196 6091 18636 7517
rect 18196 6005 18289 6091
rect 18375 6005 18457 6091
rect 18543 6005 18636 6091
rect 18196 4579 18636 6005
rect 18196 4493 18289 4579
rect 18375 4493 18457 4579
rect 18543 4493 18636 4579
rect 18196 3067 18636 4493
rect 18196 2981 18289 3067
rect 18375 2981 18457 3067
rect 18543 2981 18636 3067
rect 18196 1555 18636 2981
rect 18196 1469 18289 1555
rect 18375 1469 18457 1555
rect 18543 1469 18636 1555
rect 18196 712 18636 1469
rect 19436 38599 19876 38682
rect 19436 38513 19529 38599
rect 19615 38513 19697 38599
rect 19783 38513 19876 38599
rect 19436 37087 19876 38513
rect 19436 37001 19529 37087
rect 19615 37001 19697 37087
rect 19783 37001 19876 37087
rect 19436 35575 19876 37001
rect 19436 35489 19529 35575
rect 19615 35489 19697 35575
rect 19783 35489 19876 35575
rect 19436 34063 19876 35489
rect 19436 33977 19529 34063
rect 19615 33977 19697 34063
rect 19783 33977 19876 34063
rect 19436 32551 19876 33977
rect 19436 32465 19529 32551
rect 19615 32465 19697 32551
rect 19783 32465 19876 32551
rect 19436 31039 19876 32465
rect 19436 30953 19529 31039
rect 19615 30953 19697 31039
rect 19783 30953 19876 31039
rect 19436 29527 19876 30953
rect 19436 29441 19529 29527
rect 19615 29441 19697 29527
rect 19783 29441 19876 29527
rect 19436 28015 19876 29441
rect 19436 27929 19529 28015
rect 19615 27929 19697 28015
rect 19783 27929 19876 28015
rect 19436 26503 19876 27929
rect 19436 26417 19529 26503
rect 19615 26417 19697 26503
rect 19783 26417 19876 26503
rect 19436 24991 19876 26417
rect 19436 24905 19529 24991
rect 19615 24905 19697 24991
rect 19783 24905 19876 24991
rect 19436 23479 19876 24905
rect 19436 23393 19529 23479
rect 19615 23393 19697 23479
rect 19783 23393 19876 23479
rect 19436 21967 19876 23393
rect 19436 21881 19529 21967
rect 19615 21881 19697 21967
rect 19783 21881 19876 21967
rect 19436 20455 19876 21881
rect 19436 20369 19529 20455
rect 19615 20369 19697 20455
rect 19783 20369 19876 20455
rect 19436 18943 19876 20369
rect 19436 18857 19529 18943
rect 19615 18857 19697 18943
rect 19783 18857 19876 18943
rect 19436 17431 19876 18857
rect 19436 17345 19529 17431
rect 19615 17345 19697 17431
rect 19783 17345 19876 17431
rect 19436 15919 19876 17345
rect 19436 15833 19529 15919
rect 19615 15833 19697 15919
rect 19783 15833 19876 15919
rect 19436 14407 19876 15833
rect 19436 14321 19529 14407
rect 19615 14321 19697 14407
rect 19783 14321 19876 14407
rect 19436 12895 19876 14321
rect 19436 12809 19529 12895
rect 19615 12809 19697 12895
rect 19783 12809 19876 12895
rect 19436 11383 19876 12809
rect 19436 11297 19529 11383
rect 19615 11297 19697 11383
rect 19783 11297 19876 11383
rect 19436 9871 19876 11297
rect 19436 9785 19529 9871
rect 19615 9785 19697 9871
rect 19783 9785 19876 9871
rect 19436 8359 19876 9785
rect 19436 8273 19529 8359
rect 19615 8273 19697 8359
rect 19783 8273 19876 8359
rect 19436 6847 19876 8273
rect 19436 6761 19529 6847
rect 19615 6761 19697 6847
rect 19783 6761 19876 6847
rect 19436 5335 19876 6761
rect 19436 5249 19529 5335
rect 19615 5249 19697 5335
rect 19783 5249 19876 5335
rect 19436 3823 19876 5249
rect 19436 3737 19529 3823
rect 19615 3737 19697 3823
rect 19783 3737 19876 3823
rect 19436 2311 19876 3737
rect 19436 2225 19529 2311
rect 19615 2225 19697 2311
rect 19783 2225 19876 2311
rect 19436 799 19876 2225
rect 19436 713 19529 799
rect 19615 713 19697 799
rect 19783 713 19876 799
rect 19436 630 19876 713
rect 33316 37843 33756 38600
rect 33316 37757 33409 37843
rect 33495 37757 33577 37843
rect 33663 37757 33756 37843
rect 33316 36331 33756 37757
rect 33316 36245 33409 36331
rect 33495 36245 33577 36331
rect 33663 36245 33756 36331
rect 33316 34819 33756 36245
rect 33316 34733 33409 34819
rect 33495 34733 33577 34819
rect 33663 34733 33756 34819
rect 33316 33307 33756 34733
rect 33316 33221 33409 33307
rect 33495 33221 33577 33307
rect 33663 33221 33756 33307
rect 33316 31795 33756 33221
rect 33316 31709 33409 31795
rect 33495 31709 33577 31795
rect 33663 31709 33756 31795
rect 33316 30283 33756 31709
rect 33316 30197 33409 30283
rect 33495 30197 33577 30283
rect 33663 30197 33756 30283
rect 33316 28771 33756 30197
rect 33316 28685 33409 28771
rect 33495 28685 33577 28771
rect 33663 28685 33756 28771
rect 33316 27259 33756 28685
rect 33316 27173 33409 27259
rect 33495 27173 33577 27259
rect 33663 27173 33756 27259
rect 33316 25747 33756 27173
rect 33316 25661 33409 25747
rect 33495 25661 33577 25747
rect 33663 25661 33756 25747
rect 33316 24235 33756 25661
rect 33316 24149 33409 24235
rect 33495 24149 33577 24235
rect 33663 24149 33756 24235
rect 33316 22723 33756 24149
rect 33316 22637 33409 22723
rect 33495 22637 33577 22723
rect 33663 22637 33756 22723
rect 33316 21211 33756 22637
rect 33316 21125 33409 21211
rect 33495 21125 33577 21211
rect 33663 21125 33756 21211
rect 33316 19699 33756 21125
rect 33316 19613 33409 19699
rect 33495 19613 33577 19699
rect 33663 19613 33756 19699
rect 33316 18187 33756 19613
rect 33316 18101 33409 18187
rect 33495 18101 33577 18187
rect 33663 18101 33756 18187
rect 33316 16675 33756 18101
rect 33316 16589 33409 16675
rect 33495 16589 33577 16675
rect 33663 16589 33756 16675
rect 33316 15163 33756 16589
rect 33316 15077 33409 15163
rect 33495 15077 33577 15163
rect 33663 15077 33756 15163
rect 33316 13651 33756 15077
rect 33316 13565 33409 13651
rect 33495 13565 33577 13651
rect 33663 13565 33756 13651
rect 33316 12139 33756 13565
rect 33316 12053 33409 12139
rect 33495 12053 33577 12139
rect 33663 12053 33756 12139
rect 33316 10627 33756 12053
rect 33316 10541 33409 10627
rect 33495 10541 33577 10627
rect 33663 10541 33756 10627
rect 33316 9115 33756 10541
rect 33316 9029 33409 9115
rect 33495 9029 33577 9115
rect 33663 9029 33756 9115
rect 33316 7603 33756 9029
rect 33316 7517 33409 7603
rect 33495 7517 33577 7603
rect 33663 7517 33756 7603
rect 33316 6091 33756 7517
rect 33316 6005 33409 6091
rect 33495 6005 33577 6091
rect 33663 6005 33756 6091
rect 33316 4579 33756 6005
rect 33316 4493 33409 4579
rect 33495 4493 33577 4579
rect 33663 4493 33756 4579
rect 33316 3067 33756 4493
rect 33316 2981 33409 3067
rect 33495 2981 33577 3067
rect 33663 2981 33756 3067
rect 33316 1555 33756 2981
rect 33316 1469 33409 1555
rect 33495 1469 33577 1555
rect 33663 1469 33756 1555
rect 33316 712 33756 1469
rect 34556 38599 34996 38682
rect 34556 38513 34649 38599
rect 34735 38513 34817 38599
rect 34903 38513 34996 38599
rect 34556 37087 34996 38513
rect 34556 37001 34649 37087
rect 34735 37001 34817 37087
rect 34903 37001 34996 37087
rect 34556 35575 34996 37001
rect 34556 35489 34649 35575
rect 34735 35489 34817 35575
rect 34903 35489 34996 35575
rect 34556 34063 34996 35489
rect 34556 33977 34649 34063
rect 34735 33977 34817 34063
rect 34903 33977 34996 34063
rect 34556 32551 34996 33977
rect 34556 32465 34649 32551
rect 34735 32465 34817 32551
rect 34903 32465 34996 32551
rect 34556 31039 34996 32465
rect 34556 30953 34649 31039
rect 34735 30953 34817 31039
rect 34903 30953 34996 31039
rect 34556 29527 34996 30953
rect 34556 29441 34649 29527
rect 34735 29441 34817 29527
rect 34903 29441 34996 29527
rect 34556 28015 34996 29441
rect 34556 27929 34649 28015
rect 34735 27929 34817 28015
rect 34903 27929 34996 28015
rect 34556 26503 34996 27929
rect 34556 26417 34649 26503
rect 34735 26417 34817 26503
rect 34903 26417 34996 26503
rect 34556 24991 34996 26417
rect 34556 24905 34649 24991
rect 34735 24905 34817 24991
rect 34903 24905 34996 24991
rect 34556 23479 34996 24905
rect 34556 23393 34649 23479
rect 34735 23393 34817 23479
rect 34903 23393 34996 23479
rect 34556 21967 34996 23393
rect 34556 21881 34649 21967
rect 34735 21881 34817 21967
rect 34903 21881 34996 21967
rect 34556 20455 34996 21881
rect 34556 20369 34649 20455
rect 34735 20369 34817 20455
rect 34903 20369 34996 20455
rect 34556 18943 34996 20369
rect 34556 18857 34649 18943
rect 34735 18857 34817 18943
rect 34903 18857 34996 18943
rect 34556 17431 34996 18857
rect 34556 17345 34649 17431
rect 34735 17345 34817 17431
rect 34903 17345 34996 17431
rect 34556 15919 34996 17345
rect 34556 15833 34649 15919
rect 34735 15833 34817 15919
rect 34903 15833 34996 15919
rect 34556 14407 34996 15833
rect 34556 14321 34649 14407
rect 34735 14321 34817 14407
rect 34903 14321 34996 14407
rect 34556 12895 34996 14321
rect 34556 12809 34649 12895
rect 34735 12809 34817 12895
rect 34903 12809 34996 12895
rect 34556 11383 34996 12809
rect 34556 11297 34649 11383
rect 34735 11297 34817 11383
rect 34903 11297 34996 11383
rect 34556 9871 34996 11297
rect 34556 9785 34649 9871
rect 34735 9785 34817 9871
rect 34903 9785 34996 9871
rect 34556 8359 34996 9785
rect 34556 8273 34649 8359
rect 34735 8273 34817 8359
rect 34903 8273 34996 8359
rect 34556 6847 34996 8273
rect 34556 6761 34649 6847
rect 34735 6761 34817 6847
rect 34903 6761 34996 6847
rect 34556 5335 34996 6761
rect 34556 5249 34649 5335
rect 34735 5249 34817 5335
rect 34903 5249 34996 5335
rect 34556 3823 34996 5249
rect 34556 3737 34649 3823
rect 34735 3737 34817 3823
rect 34903 3737 34996 3823
rect 34556 2311 34996 3737
rect 34556 2225 34649 2311
rect 34735 2225 34817 2311
rect 34903 2225 34996 2311
rect 34556 799 34996 2225
rect 34556 713 34649 799
rect 34735 713 34817 799
rect 34903 713 34996 799
rect 34556 630 34996 713
rect 48436 37843 48876 38600
rect 48436 37757 48529 37843
rect 48615 37757 48697 37843
rect 48783 37757 48876 37843
rect 48436 36331 48876 37757
rect 48436 36245 48529 36331
rect 48615 36245 48697 36331
rect 48783 36245 48876 36331
rect 48436 34819 48876 36245
rect 48436 34733 48529 34819
rect 48615 34733 48697 34819
rect 48783 34733 48876 34819
rect 48436 33307 48876 34733
rect 48436 33221 48529 33307
rect 48615 33221 48697 33307
rect 48783 33221 48876 33307
rect 48436 31795 48876 33221
rect 48436 31709 48529 31795
rect 48615 31709 48697 31795
rect 48783 31709 48876 31795
rect 48436 30283 48876 31709
rect 48436 30197 48529 30283
rect 48615 30197 48697 30283
rect 48783 30197 48876 30283
rect 48436 28771 48876 30197
rect 48436 28685 48529 28771
rect 48615 28685 48697 28771
rect 48783 28685 48876 28771
rect 48436 27259 48876 28685
rect 48436 27173 48529 27259
rect 48615 27173 48697 27259
rect 48783 27173 48876 27259
rect 48436 25747 48876 27173
rect 48436 25661 48529 25747
rect 48615 25661 48697 25747
rect 48783 25661 48876 25747
rect 48436 24235 48876 25661
rect 48436 24149 48529 24235
rect 48615 24149 48697 24235
rect 48783 24149 48876 24235
rect 48436 22723 48876 24149
rect 48436 22637 48529 22723
rect 48615 22637 48697 22723
rect 48783 22637 48876 22723
rect 48436 21211 48876 22637
rect 48436 21125 48529 21211
rect 48615 21125 48697 21211
rect 48783 21125 48876 21211
rect 48436 19699 48876 21125
rect 48436 19613 48529 19699
rect 48615 19613 48697 19699
rect 48783 19613 48876 19699
rect 48436 18187 48876 19613
rect 48436 18101 48529 18187
rect 48615 18101 48697 18187
rect 48783 18101 48876 18187
rect 48436 16675 48876 18101
rect 48436 16589 48529 16675
rect 48615 16589 48697 16675
rect 48783 16589 48876 16675
rect 48436 15163 48876 16589
rect 48436 15077 48529 15163
rect 48615 15077 48697 15163
rect 48783 15077 48876 15163
rect 48436 13651 48876 15077
rect 48436 13565 48529 13651
rect 48615 13565 48697 13651
rect 48783 13565 48876 13651
rect 48436 12139 48876 13565
rect 48436 12053 48529 12139
rect 48615 12053 48697 12139
rect 48783 12053 48876 12139
rect 48436 10627 48876 12053
rect 48436 10541 48529 10627
rect 48615 10541 48697 10627
rect 48783 10541 48876 10627
rect 48436 9115 48876 10541
rect 48436 9029 48529 9115
rect 48615 9029 48697 9115
rect 48783 9029 48876 9115
rect 48436 7603 48876 9029
rect 48436 7517 48529 7603
rect 48615 7517 48697 7603
rect 48783 7517 48876 7603
rect 48436 6091 48876 7517
rect 48436 6005 48529 6091
rect 48615 6005 48697 6091
rect 48783 6005 48876 6091
rect 48436 4579 48876 6005
rect 48436 4493 48529 4579
rect 48615 4493 48697 4579
rect 48783 4493 48876 4579
rect 48436 3067 48876 4493
rect 48436 2981 48529 3067
rect 48615 2981 48697 3067
rect 48783 2981 48876 3067
rect 48436 1555 48876 2981
rect 48436 1469 48529 1555
rect 48615 1469 48697 1555
rect 48783 1469 48876 1555
rect 48436 712 48876 1469
rect 49676 38599 50116 38682
rect 49676 38513 49769 38599
rect 49855 38513 49937 38599
rect 50023 38513 50116 38599
rect 49676 37087 50116 38513
rect 49676 37001 49769 37087
rect 49855 37001 49937 37087
rect 50023 37001 50116 37087
rect 49676 35575 50116 37001
rect 49676 35489 49769 35575
rect 49855 35489 49937 35575
rect 50023 35489 50116 35575
rect 49676 34063 50116 35489
rect 49676 33977 49769 34063
rect 49855 33977 49937 34063
rect 50023 33977 50116 34063
rect 49676 32551 50116 33977
rect 49676 32465 49769 32551
rect 49855 32465 49937 32551
rect 50023 32465 50116 32551
rect 49676 31039 50116 32465
rect 49676 30953 49769 31039
rect 49855 30953 49937 31039
rect 50023 30953 50116 31039
rect 49676 29527 50116 30953
rect 49676 29441 49769 29527
rect 49855 29441 49937 29527
rect 50023 29441 50116 29527
rect 49676 28015 50116 29441
rect 49676 27929 49769 28015
rect 49855 27929 49937 28015
rect 50023 27929 50116 28015
rect 49676 26503 50116 27929
rect 49676 26417 49769 26503
rect 49855 26417 49937 26503
rect 50023 26417 50116 26503
rect 49676 24991 50116 26417
rect 49676 24905 49769 24991
rect 49855 24905 49937 24991
rect 50023 24905 50116 24991
rect 49676 23479 50116 24905
rect 49676 23393 49769 23479
rect 49855 23393 49937 23479
rect 50023 23393 50116 23479
rect 49676 21967 50116 23393
rect 49676 21881 49769 21967
rect 49855 21881 49937 21967
rect 50023 21881 50116 21967
rect 49676 20455 50116 21881
rect 49676 20369 49769 20455
rect 49855 20369 49937 20455
rect 50023 20369 50116 20455
rect 49676 18943 50116 20369
rect 49676 18857 49769 18943
rect 49855 18857 49937 18943
rect 50023 18857 50116 18943
rect 49676 17431 50116 18857
rect 49676 17345 49769 17431
rect 49855 17345 49937 17431
rect 50023 17345 50116 17431
rect 49676 15919 50116 17345
rect 49676 15833 49769 15919
rect 49855 15833 49937 15919
rect 50023 15833 50116 15919
rect 49676 14407 50116 15833
rect 49676 14321 49769 14407
rect 49855 14321 49937 14407
rect 50023 14321 50116 14407
rect 49676 12895 50116 14321
rect 49676 12809 49769 12895
rect 49855 12809 49937 12895
rect 50023 12809 50116 12895
rect 49676 11383 50116 12809
rect 49676 11297 49769 11383
rect 49855 11297 49937 11383
rect 50023 11297 50116 11383
rect 49676 9871 50116 11297
rect 49676 9785 49769 9871
rect 49855 9785 49937 9871
rect 50023 9785 50116 9871
rect 49676 8359 50116 9785
rect 49676 8273 49769 8359
rect 49855 8273 49937 8359
rect 50023 8273 50116 8359
rect 49676 6847 50116 8273
rect 49676 6761 49769 6847
rect 49855 6761 49937 6847
rect 50023 6761 50116 6847
rect 49676 5335 50116 6761
rect 49676 5249 49769 5335
rect 49855 5249 49937 5335
rect 50023 5249 50116 5335
rect 49676 3823 50116 5249
rect 49676 3737 49769 3823
rect 49855 3737 49937 3823
rect 50023 3737 50116 3823
rect 49676 2311 50116 3737
rect 49676 2225 49769 2311
rect 49855 2225 49937 2311
rect 50023 2225 50116 2311
rect 49676 799 50116 2225
rect 49676 713 49769 799
rect 49855 713 49937 799
rect 50023 713 50116 799
rect 49676 630 50116 713
rect 63556 37843 63996 38600
rect 63556 37757 63649 37843
rect 63735 37757 63817 37843
rect 63903 37757 63996 37843
rect 63556 36331 63996 37757
rect 63556 36245 63649 36331
rect 63735 36245 63817 36331
rect 63903 36245 63996 36331
rect 63556 34819 63996 36245
rect 63556 34733 63649 34819
rect 63735 34733 63817 34819
rect 63903 34733 63996 34819
rect 63556 33307 63996 34733
rect 63556 33221 63649 33307
rect 63735 33221 63817 33307
rect 63903 33221 63996 33307
rect 63556 31795 63996 33221
rect 63556 31709 63649 31795
rect 63735 31709 63817 31795
rect 63903 31709 63996 31795
rect 63556 30283 63996 31709
rect 63556 30197 63649 30283
rect 63735 30197 63817 30283
rect 63903 30197 63996 30283
rect 63556 28771 63996 30197
rect 63556 28685 63649 28771
rect 63735 28685 63817 28771
rect 63903 28685 63996 28771
rect 63556 27259 63996 28685
rect 63556 27173 63649 27259
rect 63735 27173 63817 27259
rect 63903 27173 63996 27259
rect 63556 25747 63996 27173
rect 63556 25661 63649 25747
rect 63735 25661 63817 25747
rect 63903 25661 63996 25747
rect 63556 24235 63996 25661
rect 63556 24149 63649 24235
rect 63735 24149 63817 24235
rect 63903 24149 63996 24235
rect 63556 22723 63996 24149
rect 63556 22637 63649 22723
rect 63735 22637 63817 22723
rect 63903 22637 63996 22723
rect 63556 21211 63996 22637
rect 63556 21125 63649 21211
rect 63735 21125 63817 21211
rect 63903 21125 63996 21211
rect 63556 19699 63996 21125
rect 63556 19613 63649 19699
rect 63735 19613 63817 19699
rect 63903 19613 63996 19699
rect 63556 18187 63996 19613
rect 63556 18101 63649 18187
rect 63735 18101 63817 18187
rect 63903 18101 63996 18187
rect 63556 16675 63996 18101
rect 63556 16589 63649 16675
rect 63735 16589 63817 16675
rect 63903 16589 63996 16675
rect 63556 15163 63996 16589
rect 63556 15077 63649 15163
rect 63735 15077 63817 15163
rect 63903 15077 63996 15163
rect 63556 13651 63996 15077
rect 63556 13565 63649 13651
rect 63735 13565 63817 13651
rect 63903 13565 63996 13651
rect 63556 12139 63996 13565
rect 63556 12053 63649 12139
rect 63735 12053 63817 12139
rect 63903 12053 63996 12139
rect 63556 10627 63996 12053
rect 63556 10541 63649 10627
rect 63735 10541 63817 10627
rect 63903 10541 63996 10627
rect 63556 9115 63996 10541
rect 63556 9029 63649 9115
rect 63735 9029 63817 9115
rect 63903 9029 63996 9115
rect 63556 7603 63996 9029
rect 63556 7517 63649 7603
rect 63735 7517 63817 7603
rect 63903 7517 63996 7603
rect 63556 6091 63996 7517
rect 63556 6005 63649 6091
rect 63735 6005 63817 6091
rect 63903 6005 63996 6091
rect 63556 4579 63996 6005
rect 63556 4493 63649 4579
rect 63735 4493 63817 4579
rect 63903 4493 63996 4579
rect 63556 3067 63996 4493
rect 63556 2981 63649 3067
rect 63735 2981 63817 3067
rect 63903 2981 63996 3067
rect 63556 1555 63996 2981
rect 63556 1469 63649 1555
rect 63735 1469 63817 1555
rect 63903 1469 63996 1555
rect 63556 712 63996 1469
rect 64796 38599 65236 38682
rect 64796 38513 64889 38599
rect 64975 38513 65057 38599
rect 65143 38513 65236 38599
rect 64796 37087 65236 38513
rect 64796 37001 64889 37087
rect 64975 37001 65057 37087
rect 65143 37001 65236 37087
rect 64796 35575 65236 37001
rect 64796 35489 64889 35575
rect 64975 35489 65057 35575
rect 65143 35489 65236 35575
rect 64796 34063 65236 35489
rect 64796 33977 64889 34063
rect 64975 33977 65057 34063
rect 65143 33977 65236 34063
rect 64796 32551 65236 33977
rect 64796 32465 64889 32551
rect 64975 32465 65057 32551
rect 65143 32465 65236 32551
rect 64796 31039 65236 32465
rect 64796 30953 64889 31039
rect 64975 30953 65057 31039
rect 65143 30953 65236 31039
rect 64796 29527 65236 30953
rect 64796 29441 64889 29527
rect 64975 29441 65057 29527
rect 65143 29441 65236 29527
rect 64796 28015 65236 29441
rect 64796 27929 64889 28015
rect 64975 27929 65057 28015
rect 65143 27929 65236 28015
rect 64796 26503 65236 27929
rect 64796 26417 64889 26503
rect 64975 26417 65057 26503
rect 65143 26417 65236 26503
rect 64796 24991 65236 26417
rect 64796 24905 64889 24991
rect 64975 24905 65057 24991
rect 65143 24905 65236 24991
rect 64796 23479 65236 24905
rect 64796 23393 64889 23479
rect 64975 23393 65057 23479
rect 65143 23393 65236 23479
rect 64796 21967 65236 23393
rect 64796 21881 64889 21967
rect 64975 21881 65057 21967
rect 65143 21881 65236 21967
rect 64796 20455 65236 21881
rect 64796 20369 64889 20455
rect 64975 20369 65057 20455
rect 65143 20369 65236 20455
rect 64796 18943 65236 20369
rect 64796 18857 64889 18943
rect 64975 18857 65057 18943
rect 65143 18857 65236 18943
rect 64796 17431 65236 18857
rect 64796 17345 64889 17431
rect 64975 17345 65057 17431
rect 65143 17345 65236 17431
rect 64796 15919 65236 17345
rect 64796 15833 64889 15919
rect 64975 15833 65057 15919
rect 65143 15833 65236 15919
rect 64796 14407 65236 15833
rect 64796 14321 64889 14407
rect 64975 14321 65057 14407
rect 65143 14321 65236 14407
rect 64796 12895 65236 14321
rect 64796 12809 64889 12895
rect 64975 12809 65057 12895
rect 65143 12809 65236 12895
rect 64796 11383 65236 12809
rect 64796 11297 64889 11383
rect 64975 11297 65057 11383
rect 65143 11297 65236 11383
rect 64796 9871 65236 11297
rect 64796 9785 64889 9871
rect 64975 9785 65057 9871
rect 65143 9785 65236 9871
rect 64796 8359 65236 9785
rect 64796 8273 64889 8359
rect 64975 8273 65057 8359
rect 65143 8273 65236 8359
rect 64796 6847 65236 8273
rect 64796 6761 64889 6847
rect 64975 6761 65057 6847
rect 65143 6761 65236 6847
rect 64796 5335 65236 6761
rect 64796 5249 64889 5335
rect 64975 5249 65057 5335
rect 65143 5249 65236 5335
rect 64796 3823 65236 5249
rect 64796 3737 64889 3823
rect 64975 3737 65057 3823
rect 65143 3737 65236 3823
rect 64796 2311 65236 3737
rect 64796 2225 64889 2311
rect 64975 2225 65057 2311
rect 65143 2225 65236 2311
rect 64796 799 65236 2225
rect 64796 713 64889 799
rect 64975 713 65057 799
rect 65143 713 65236 799
rect 64796 630 65236 713
rect 78676 37843 79116 38600
rect 78676 37757 78769 37843
rect 78855 37757 78937 37843
rect 79023 37757 79116 37843
rect 78676 36331 79116 37757
rect 78676 36245 78769 36331
rect 78855 36245 78937 36331
rect 79023 36245 79116 36331
rect 78676 34819 79116 36245
rect 78676 34733 78769 34819
rect 78855 34733 78937 34819
rect 79023 34733 79116 34819
rect 78676 33307 79116 34733
rect 78676 33221 78769 33307
rect 78855 33221 78937 33307
rect 79023 33221 79116 33307
rect 78676 31795 79116 33221
rect 78676 31709 78769 31795
rect 78855 31709 78937 31795
rect 79023 31709 79116 31795
rect 78676 30283 79116 31709
rect 78676 30197 78769 30283
rect 78855 30197 78937 30283
rect 79023 30197 79116 30283
rect 78676 28771 79116 30197
rect 78676 28685 78769 28771
rect 78855 28685 78937 28771
rect 79023 28685 79116 28771
rect 78676 27259 79116 28685
rect 78676 27173 78769 27259
rect 78855 27173 78937 27259
rect 79023 27173 79116 27259
rect 78676 25747 79116 27173
rect 78676 25661 78769 25747
rect 78855 25661 78937 25747
rect 79023 25661 79116 25747
rect 78676 24235 79116 25661
rect 78676 24149 78769 24235
rect 78855 24149 78937 24235
rect 79023 24149 79116 24235
rect 78676 22723 79116 24149
rect 78676 22637 78769 22723
rect 78855 22637 78937 22723
rect 79023 22637 79116 22723
rect 78676 21211 79116 22637
rect 78676 21125 78769 21211
rect 78855 21125 78937 21211
rect 79023 21125 79116 21211
rect 78676 19699 79116 21125
rect 78676 19613 78769 19699
rect 78855 19613 78937 19699
rect 79023 19613 79116 19699
rect 78676 18187 79116 19613
rect 78676 18101 78769 18187
rect 78855 18101 78937 18187
rect 79023 18101 79116 18187
rect 78676 16675 79116 18101
rect 78676 16589 78769 16675
rect 78855 16589 78937 16675
rect 79023 16589 79116 16675
rect 78676 15163 79116 16589
rect 78676 15077 78769 15163
rect 78855 15077 78937 15163
rect 79023 15077 79116 15163
rect 78676 13651 79116 15077
rect 78676 13565 78769 13651
rect 78855 13565 78937 13651
rect 79023 13565 79116 13651
rect 78676 12139 79116 13565
rect 78676 12053 78769 12139
rect 78855 12053 78937 12139
rect 79023 12053 79116 12139
rect 78676 10627 79116 12053
rect 78676 10541 78769 10627
rect 78855 10541 78937 10627
rect 79023 10541 79116 10627
rect 78676 9115 79116 10541
rect 78676 9029 78769 9115
rect 78855 9029 78937 9115
rect 79023 9029 79116 9115
rect 78676 7603 79116 9029
rect 78676 7517 78769 7603
rect 78855 7517 78937 7603
rect 79023 7517 79116 7603
rect 78676 6091 79116 7517
rect 78676 6005 78769 6091
rect 78855 6005 78937 6091
rect 79023 6005 79116 6091
rect 78676 4579 79116 6005
rect 78676 4493 78769 4579
rect 78855 4493 78937 4579
rect 79023 4493 79116 4579
rect 78676 3067 79116 4493
rect 78676 2981 78769 3067
rect 78855 2981 78937 3067
rect 79023 2981 79116 3067
rect 78676 1555 79116 2981
rect 78676 1469 78769 1555
rect 78855 1469 78937 1555
rect 79023 1469 79116 1555
rect 78676 712 79116 1469
rect 79916 38599 80356 38682
rect 79916 38513 80009 38599
rect 80095 38513 80177 38599
rect 80263 38513 80356 38599
rect 79916 37087 80356 38513
rect 79916 37001 80009 37087
rect 80095 37001 80177 37087
rect 80263 37001 80356 37087
rect 79916 35575 80356 37001
rect 79916 35489 80009 35575
rect 80095 35489 80177 35575
rect 80263 35489 80356 35575
rect 79916 34063 80356 35489
rect 79916 33977 80009 34063
rect 80095 33977 80177 34063
rect 80263 33977 80356 34063
rect 79916 32551 80356 33977
rect 79916 32465 80009 32551
rect 80095 32465 80177 32551
rect 80263 32465 80356 32551
rect 79916 31039 80356 32465
rect 79916 30953 80009 31039
rect 80095 30953 80177 31039
rect 80263 30953 80356 31039
rect 79916 29527 80356 30953
rect 79916 29441 80009 29527
rect 80095 29441 80177 29527
rect 80263 29441 80356 29527
rect 79916 28015 80356 29441
rect 79916 27929 80009 28015
rect 80095 27929 80177 28015
rect 80263 27929 80356 28015
rect 79916 26503 80356 27929
rect 79916 26417 80009 26503
rect 80095 26417 80177 26503
rect 80263 26417 80356 26503
rect 79916 24991 80356 26417
rect 79916 24905 80009 24991
rect 80095 24905 80177 24991
rect 80263 24905 80356 24991
rect 79916 23479 80356 24905
rect 79916 23393 80009 23479
rect 80095 23393 80177 23479
rect 80263 23393 80356 23479
rect 79916 21967 80356 23393
rect 79916 21881 80009 21967
rect 80095 21881 80177 21967
rect 80263 21881 80356 21967
rect 79916 20455 80356 21881
rect 79916 20369 80009 20455
rect 80095 20369 80177 20455
rect 80263 20369 80356 20455
rect 79916 18943 80356 20369
rect 79916 18857 80009 18943
rect 80095 18857 80177 18943
rect 80263 18857 80356 18943
rect 79916 17431 80356 18857
rect 79916 17345 80009 17431
rect 80095 17345 80177 17431
rect 80263 17345 80356 17431
rect 79916 15919 80356 17345
rect 79916 15833 80009 15919
rect 80095 15833 80177 15919
rect 80263 15833 80356 15919
rect 79916 14407 80356 15833
rect 79916 14321 80009 14407
rect 80095 14321 80177 14407
rect 80263 14321 80356 14407
rect 79916 12895 80356 14321
rect 79916 12809 80009 12895
rect 80095 12809 80177 12895
rect 80263 12809 80356 12895
rect 79916 11383 80356 12809
rect 79916 11297 80009 11383
rect 80095 11297 80177 11383
rect 80263 11297 80356 11383
rect 79916 9871 80356 11297
rect 79916 9785 80009 9871
rect 80095 9785 80177 9871
rect 80263 9785 80356 9871
rect 79916 8359 80356 9785
rect 79916 8273 80009 8359
rect 80095 8273 80177 8359
rect 80263 8273 80356 8359
rect 79916 6847 80356 8273
rect 79916 6761 80009 6847
rect 80095 6761 80177 6847
rect 80263 6761 80356 6847
rect 79916 5335 80356 6761
rect 79916 5249 80009 5335
rect 80095 5249 80177 5335
rect 80263 5249 80356 5335
rect 79916 3823 80356 5249
rect 79916 3737 80009 3823
rect 80095 3737 80177 3823
rect 80263 3737 80356 3823
rect 79916 2311 80356 3737
rect 79916 2225 80009 2311
rect 80095 2225 80177 2311
rect 80263 2225 80356 2311
rect 79916 799 80356 2225
rect 79916 713 80009 799
rect 80095 713 80177 799
rect 80263 713 80356 799
rect 79916 630 80356 713
rect 93796 37843 94236 38600
rect 93796 37757 93889 37843
rect 93975 37757 94057 37843
rect 94143 37757 94236 37843
rect 93796 36331 94236 37757
rect 93796 36245 93889 36331
rect 93975 36245 94057 36331
rect 94143 36245 94236 36331
rect 93796 34819 94236 36245
rect 93796 34733 93889 34819
rect 93975 34733 94057 34819
rect 94143 34733 94236 34819
rect 93796 33307 94236 34733
rect 93796 33221 93889 33307
rect 93975 33221 94057 33307
rect 94143 33221 94236 33307
rect 93796 31795 94236 33221
rect 93796 31709 93889 31795
rect 93975 31709 94057 31795
rect 94143 31709 94236 31795
rect 93796 30283 94236 31709
rect 93796 30197 93889 30283
rect 93975 30197 94057 30283
rect 94143 30197 94236 30283
rect 93796 28771 94236 30197
rect 93796 28685 93889 28771
rect 93975 28685 94057 28771
rect 94143 28685 94236 28771
rect 93796 27259 94236 28685
rect 93796 27173 93889 27259
rect 93975 27173 94057 27259
rect 94143 27173 94236 27259
rect 93796 25747 94236 27173
rect 93796 25661 93889 25747
rect 93975 25661 94057 25747
rect 94143 25661 94236 25747
rect 93796 24235 94236 25661
rect 93796 24149 93889 24235
rect 93975 24149 94057 24235
rect 94143 24149 94236 24235
rect 93796 22723 94236 24149
rect 93796 22637 93889 22723
rect 93975 22637 94057 22723
rect 94143 22637 94236 22723
rect 93796 21211 94236 22637
rect 93796 21125 93889 21211
rect 93975 21125 94057 21211
rect 94143 21125 94236 21211
rect 93796 19699 94236 21125
rect 93796 19613 93889 19699
rect 93975 19613 94057 19699
rect 94143 19613 94236 19699
rect 93796 18187 94236 19613
rect 93796 18101 93889 18187
rect 93975 18101 94057 18187
rect 94143 18101 94236 18187
rect 93796 16675 94236 18101
rect 93796 16589 93889 16675
rect 93975 16589 94057 16675
rect 94143 16589 94236 16675
rect 93796 15163 94236 16589
rect 93796 15077 93889 15163
rect 93975 15077 94057 15163
rect 94143 15077 94236 15163
rect 93796 13651 94236 15077
rect 93796 13565 93889 13651
rect 93975 13565 94057 13651
rect 94143 13565 94236 13651
rect 93796 12139 94236 13565
rect 93796 12053 93889 12139
rect 93975 12053 94057 12139
rect 94143 12053 94236 12139
rect 93796 10627 94236 12053
rect 93796 10541 93889 10627
rect 93975 10541 94057 10627
rect 94143 10541 94236 10627
rect 93796 9115 94236 10541
rect 93796 9029 93889 9115
rect 93975 9029 94057 9115
rect 94143 9029 94236 9115
rect 93796 7603 94236 9029
rect 93796 7517 93889 7603
rect 93975 7517 94057 7603
rect 94143 7517 94236 7603
rect 93796 6091 94236 7517
rect 93796 6005 93889 6091
rect 93975 6005 94057 6091
rect 94143 6005 94236 6091
rect 93796 4579 94236 6005
rect 93796 4493 93889 4579
rect 93975 4493 94057 4579
rect 94143 4493 94236 4579
rect 93796 3067 94236 4493
rect 93796 2981 93889 3067
rect 93975 2981 94057 3067
rect 94143 2981 94236 3067
rect 93796 1555 94236 2981
rect 93796 1469 93889 1555
rect 93975 1469 94057 1555
rect 94143 1469 94236 1555
rect 93796 712 94236 1469
rect 95036 38599 95476 38682
rect 95036 38513 95129 38599
rect 95215 38513 95297 38599
rect 95383 38513 95476 38599
rect 95036 37087 95476 38513
rect 95036 37001 95129 37087
rect 95215 37001 95297 37087
rect 95383 37001 95476 37087
rect 95036 35575 95476 37001
rect 95036 35489 95129 35575
rect 95215 35489 95297 35575
rect 95383 35489 95476 35575
rect 95036 34063 95476 35489
rect 95036 33977 95129 34063
rect 95215 33977 95297 34063
rect 95383 33977 95476 34063
rect 95036 32551 95476 33977
rect 95036 32465 95129 32551
rect 95215 32465 95297 32551
rect 95383 32465 95476 32551
rect 95036 31039 95476 32465
rect 95036 30953 95129 31039
rect 95215 30953 95297 31039
rect 95383 30953 95476 31039
rect 95036 29527 95476 30953
rect 95036 29441 95129 29527
rect 95215 29441 95297 29527
rect 95383 29441 95476 29527
rect 95036 28015 95476 29441
rect 95036 27929 95129 28015
rect 95215 27929 95297 28015
rect 95383 27929 95476 28015
rect 95036 26503 95476 27929
rect 95036 26417 95129 26503
rect 95215 26417 95297 26503
rect 95383 26417 95476 26503
rect 95036 24991 95476 26417
rect 95036 24905 95129 24991
rect 95215 24905 95297 24991
rect 95383 24905 95476 24991
rect 95036 23479 95476 24905
rect 95036 23393 95129 23479
rect 95215 23393 95297 23479
rect 95383 23393 95476 23479
rect 95036 21967 95476 23393
rect 95036 21881 95129 21967
rect 95215 21881 95297 21967
rect 95383 21881 95476 21967
rect 95036 20455 95476 21881
rect 95036 20369 95129 20455
rect 95215 20369 95297 20455
rect 95383 20369 95476 20455
rect 95036 18943 95476 20369
rect 95036 18857 95129 18943
rect 95215 18857 95297 18943
rect 95383 18857 95476 18943
rect 95036 17431 95476 18857
rect 95036 17345 95129 17431
rect 95215 17345 95297 17431
rect 95383 17345 95476 17431
rect 95036 15919 95476 17345
rect 95036 15833 95129 15919
rect 95215 15833 95297 15919
rect 95383 15833 95476 15919
rect 95036 14407 95476 15833
rect 95036 14321 95129 14407
rect 95215 14321 95297 14407
rect 95383 14321 95476 14407
rect 95036 12895 95476 14321
rect 95036 12809 95129 12895
rect 95215 12809 95297 12895
rect 95383 12809 95476 12895
rect 95036 11383 95476 12809
rect 95036 11297 95129 11383
rect 95215 11297 95297 11383
rect 95383 11297 95476 11383
rect 95036 9871 95476 11297
rect 95036 9785 95129 9871
rect 95215 9785 95297 9871
rect 95383 9785 95476 9871
rect 95036 8359 95476 9785
rect 95036 8273 95129 8359
rect 95215 8273 95297 8359
rect 95383 8273 95476 8359
rect 95036 6847 95476 8273
rect 95036 6761 95129 6847
rect 95215 6761 95297 6847
rect 95383 6761 95476 6847
rect 95036 5335 95476 6761
rect 95036 5249 95129 5335
rect 95215 5249 95297 5335
rect 95383 5249 95476 5335
rect 95036 3823 95476 5249
rect 95036 3737 95129 3823
rect 95215 3737 95297 3823
rect 95383 3737 95476 3823
rect 95036 2311 95476 3737
rect 95036 2225 95129 2311
rect 95215 2225 95297 2311
rect 95383 2225 95476 2311
rect 95036 799 95476 2225
rect 95036 713 95129 799
rect 95215 713 95297 799
rect 95383 713 95476 799
rect 95036 630 95476 713
use sg13g2_and2_1  _222_
timestamp 1676905363
transform 1 0 8736 0 1 14364
box -48 -56 528 834
use sg13g2_and2_1  _223_
timestamp 1676905363
transform 1 0 4992 0 1 5292
box -48 -56 528 834
use sg13g2_and2_1  _224_
timestamp 1676905363
transform 1 0 7872 0 1 34020
box -48 -56 528 834
use sg13g2_and2_1  _225_
timestamp 1676905363
transform 1 0 5472 0 1 20412
box -48 -56 528 834
use sg13g2_and2_1  _226_
timestamp 1676905363
transform -1 0 55584 0 1 9828
box -48 -56 528 834
use sg13g2_and2_1  _227_
timestamp 1676905363
transform -1 0 44736 0 1 30996
box -48 -56 528 834
use sg13g2_and2_1  _228_
timestamp 1676905363
transform 1 0 29088 0 1 17388
box -48 -56 528 834
use sg13g2_and2_1  _229_
timestamp 1676905363
transform 1 0 44832 0 1 21924
box -48 -56 528 834
use sg13g2_and2_1  _230_
timestamp 1676905363
transform 1 0 35040 0 1 21924
box -48 -56 528 834
use sg13g2_and2_1  _231_
timestamp 1676905363
transform 1 0 50016 0 -1 5292
box -48 -56 528 834
use sg13g2_and2_1  _232_
timestamp 1676905363
transform 1 0 40608 0 -1 6804
box -48 -56 528 834
use sg13g2_and2_1  _233_
timestamp 1676905363
transform 1 0 52224 0 1 17388
box -48 -56 528 834
use sg13g2_and2_1  _234_
timestamp 1676905363
transform 1 0 17472 0 1 3780
box -48 -56 528 834
use sg13g2_and2_1  _235_
timestamp 1676905363
transform 1 0 4896 0 -1 27972
box -48 -56 528 834
use sg13g2_and2_1  _236_
timestamp 1676905363
transform 1 0 19872 0 -1 15876
box -48 -56 528 834
use sg13g2_and2_1  _237_
timestamp 1676905363
transform 1 0 18144 0 -1 30996
box -48 -56 528 834
use sg13g2_and2_1  _238_
timestamp 1676905363
transform 1 0 25152 0 -1 35532
box -48 -56 528 834
use sg13g2_and2_1  _239_
timestamp 1676905363
transform 1 0 33696 0 1 34020
box -48 -56 528 834
use sg13g2_nand2_1  _240_
timestamp 1676560849
transform 1 0 25824 0 1 8316
box -48 -56 432 834
use sg13g2_nand2_1  _241_
timestamp 1676560849
transform 1 0 28128 0 1 9828
box -48 -56 432 834
use sg13g2_nor2_1  _242_
timestamp 1676630787
transform 1 0 27744 0 1 9828
box -48 -56 432 834
use sg13g2_xor2_1  _243_
timestamp 1677581577
transform -1 0 28416 0 1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _244_
timestamp 1677520200
transform -1 0 27648 0 1 8316
box -48 -56 816 834
use sg13g2_o21ai_1  _245_
timestamp 1685179043
transform 1 0 29472 0 1 8316
box -48 -56 538 834
use sg13g2_and2_1  _246_
timestamp 1676905363
transform 1 0 31584 0 -1 12852
box -48 -56 528 834
use sg13g2_or2_1  _247_
timestamp 1684239771
transform 1 0 29760 0 1 11340
box -48 -56 528 834
use sg13g2_nand2b_1  _248_
timestamp 1676570795
transform 1 0 31872 0 -1 11340
box -48 -56 528 834
use sg13g2_xnor2_1  _249_
timestamp 1677520200
transform -1 0 31584 0 -1 12852
box -48 -56 816 834
use sg13g2_xor2_1  _250_
timestamp 1677581577
transform -1 0 25920 0 -1 8316
box -48 -56 816 834
use sg13g2_nand2_1  _251_
timestamp 1676560849
transform 1 0 55296 0 1 14364
box -48 -56 432 834
use sg13g2_xor2_1  _252_
timestamp 1677581577
transform -1 0 59904 0 1 14364
box -48 -56 816 834
use sg13g2_xnor2_1  _253_
timestamp 1677520200
transform 1 0 55680 0 1 14364
box -48 -56 816 834
use sg13g2_xor2_1  _254_
timestamp 1677581577
transform -1 0 55776 0 -1 14364
box -48 -56 816 834
use sg13g2_nand2_1  _255_
timestamp 1676560849
transform 1 0 42528 0 -1 12852
box -48 -56 432 834
use sg13g2_xor2_1  _256_
timestamp 1677581577
transform -1 0 44160 0 -1 14364
box -48 -56 816 834
use sg13g2_xnor2_1  _257_
timestamp 1677520200
transform -1 0 43488 0 1 11340
box -48 -56 816 834
use sg13g2_xor2_1  _258_
timestamp 1677581577
transform -1 0 41856 0 1 9828
box -48 -56 816 834
use sg13g2_nand2_1  _259_
timestamp 1676560849
transform 1 0 39456 0 -1 15876
box -48 -56 432 834
use sg13g2_xor2_1  _260_
timestamp 1677581577
transform 1 0 40320 0 -1 17388
box -48 -56 816 834
use sg13g2_xnor2_1  _261_
timestamp 1677520200
transform 1 0 40320 0 -1 15876
box -48 -56 816 834
use sg13g2_xor2_1  _262_
timestamp 1677581577
transform 1 0 38208 0 1 14364
box -48 -56 816 834
use sg13g2_nand2_1  _263_
timestamp 1676560849
transform 1 0 49248 0 -1 12852
box -48 -56 432 834
use sg13g2_xor2_1  _264_
timestamp 1677581577
transform -1 0 51072 0 -1 12852
box -48 -56 816 834
use sg13g2_xnor2_1  _265_
timestamp 1677520200
transform -1 0 50208 0 1 12852
box -48 -56 816 834
use sg13g2_xor2_1  _266_
timestamp 1677581577
transform -1 0 49440 0 1 11340
box -48 -56 816 834
use sg13g2_nand2_1  _267_
timestamp 1676560849
transform -1 0 33792 0 -1 15876
box -48 -56 432 834
use sg13g2_xor2_1  _268_
timestamp 1677581577
transform 1 0 32640 0 -1 17388
box -48 -56 816 834
use sg13g2_xnor2_1  _269_
timestamp 1677520200
transform 1 0 33696 0 1 15876
box -48 -56 816 834
use sg13g2_xor2_1  _270_
timestamp 1677581577
transform 1 0 33600 0 1 14364
box -48 -56 816 834
use sg13g2_nand2_1  _271_
timestamp 1676560849
transform 1 0 39648 0 1 20412
box -48 -56 432 834
use sg13g2_xor2_1  _272_
timestamp 1677581577
transform -1 0 40896 0 -1 23436
box -48 -56 816 834
use sg13g2_xnor2_1  _273_
timestamp 1677520200
transform 1 0 40032 0 1 20412
box -48 -56 816 834
use sg13g2_xor2_1  _274_
timestamp 1677581577
transform 1 0 38592 0 -1 20412
box -48 -56 816 834
use sg13g2_nand2_1  _275_
timestamp 1676560849
transform -1 0 46848 0 -1 8316
box -48 -56 432 834
use sg13g2_xor2_1  _276_
timestamp 1677581577
transform 1 0 46368 0 -1 6804
box -48 -56 816 834
use sg13g2_xnor2_1  _277_
timestamp 1677520200
transform 1 0 46848 0 -1 8316
box -48 -56 816 834
use sg13g2_xor2_1  _278_
timestamp 1677581577
transform -1 0 47232 0 1 8316
box -48 -56 816 834
use sg13g2_nand2_1  _279_
timestamp 1676560849
transform 1 0 37152 0 -1 32508
box -48 -56 432 834
use sg13g2_xor2_1  _280_
timestamp 1677581577
transform -1 0 40512 0 -1 32508
box -48 -56 816 834
use sg13g2_xnor2_1  _281_
timestamp 1677520200
transform -1 0 39168 0 1 30996
box -48 -56 816 834
use sg13g2_xor2_1  _282_
timestamp 1677581577
transform 1 0 37536 0 -1 32508
box -48 -56 816 834
use sg13g2_nand2_1  _283_
timestamp 1676560849
transform -1 0 33504 0 1 6804
box -48 -56 432 834
use sg13g2_nand2_1  _284_
timestamp 1676560849
transform 1 0 33120 0 1 8316
box -48 -56 432 834
use sg13g2_nor2_1  _285_
timestamp 1676630787
transform 1 0 34272 0 1 8316
box -48 -56 432 834
use sg13g2_xor2_1  _286_
timestamp 1677581577
transform -1 0 34272 0 1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _287_
timestamp 1677520200
transform -1 0 33792 0 -1 8316
box -48 -56 816 834
use sg13g2_xor2_1  _288_
timestamp 1677581577
transform -1 0 34560 0 -1 8316
box -48 -56 816 834
use sg13g2_nand2_1  _289_
timestamp 1676560849
transform 1 0 20832 0 -1 24948
box -48 -56 432 834
use sg13g2_xor2_1  _290_
timestamp 1677581577
transform 1 0 21696 0 1 24948
box -48 -56 816 834
use sg13g2_xnor2_1  _291_
timestamp 1677520200
transform -1 0 22368 0 1 23436
box -48 -56 816 834
use sg13g2_xor2_1  _292_
timestamp 1677581577
transform -1 0 21312 0 -1 23436
box -48 -56 816 834
use sg13g2_nand2_1  _293_
timestamp 1676560849
transform -1 0 17184 0 -1 24948
box -48 -56 432 834
use sg13g2_xor2_1  _294_
timestamp 1677581577
transform 1 0 16032 0 -1 24948
box -48 -56 816 834
use sg13g2_xnor2_1  _295_
timestamp 1677520200
transform 1 0 16320 0 1 24948
box -48 -56 816 834
use sg13g2_xor2_1  _296_
timestamp 1677581577
transform 1 0 15360 0 1 23436
box -48 -56 816 834
use sg13g2_nand2_1  _297_
timestamp 1676560849
transform 1 0 28608 0 1 26460
box -48 -56 432 834
use sg13g2_xor2_1  _298_
timestamp 1677581577
transform 1 0 29952 0 1 29484
box -48 -56 816 834
use sg13g2_xnor2_1  _299_
timestamp 1677520200
transform -1 0 29472 0 1 27972
box -48 -56 816 834
use sg13g2_xor2_1  _300_
timestamp 1677581577
transform -1 0 29280 0 -1 26460
box -48 -56 816 834
use sg13g2_nand2_1  _301_
timestamp 1676560849
transform 1 0 11328 0 1 20412
box -48 -56 432 834
use sg13g2_xor2_1  _302_
timestamp 1677581577
transform 1 0 10656 0 -1 18900
box -48 -56 816 834
use sg13g2_xnor2_1  _303_
timestamp 1677520200
transform 1 0 11808 0 -1 20412
box -48 -56 816 834
use sg13g2_xor2_1  _304_
timestamp 1677581577
transform 1 0 11712 0 1 20412
box -48 -56 816 834
use sg13g2_nand2_1  _305_
timestamp 1676560849
transform -1 0 11328 0 1 26460
box -48 -56 432 834
use sg13g2_xor2_1  _306_
timestamp 1677581577
transform 1 0 10464 0 1 29484
box -48 -56 816 834
use sg13g2_xnor2_1  _307_
timestamp 1677520200
transform 1 0 10752 0 -1 27972
box -48 -56 816 834
use sg13g2_xor2_1  _308_
timestamp 1677581577
transform 1 0 9984 0 -1 26460
box -48 -56 816 834
use sg13g2_nand2_1  _309_
timestamp 1676560849
transform -1 0 25440 0 -1 30996
box -48 -56 432 834
use sg13g2_xor2_1  _310_
timestamp 1677581577
transform 1 0 23808 0 1 30996
box -48 -56 816 834
use sg13g2_xnor2_1  _311_
timestamp 1677520200
transform 1 0 25440 0 -1 30996
box -48 -56 816 834
use sg13g2_xor2_1  _312_
timestamp 1677581577
transform 1 0 25248 0 1 29484
box -48 -56 816 834
use sg13g2_nand2_1  _313_
timestamp 1676560849
transform 1 0 21792 0 1 9828
box -48 -56 432 834
use sg13g2_nand2_1  _314_
timestamp 1676560849
transform 1 0 22944 0 1 12852
box -48 -56 432 834
use sg13g2_nor2_1  _315_
timestamp 1676630787
transform -1 0 24288 0 -1 12852
box -48 -56 432 834
use sg13g2_xor2_1  _316_
timestamp 1677581577
transform 1 0 22656 0 -1 12852
box -48 -56 816 834
use sg13g2_xnor2_1  _317_
timestamp 1677520200
transform 1 0 23040 0 1 11340
box -48 -56 816 834
use sg13g2_xor2_1  _318_
timestamp 1677581577
transform 1 0 21024 0 1 9828
box -48 -56 816 834
use sg13g2_nand2_1  _319_
timestamp 1676560849
transform 1 0 7008 0 -1 14364
box -48 -56 432 834
use sg13g2_nand2_1  _320_
timestamp 1676560849
transform -1 0 9408 0 -1 14364
box -48 -56 432 834
use sg13g2_xor2_1  _321_
timestamp 1677581577
transform 1 0 7968 0 1 14364
box -48 -56 816 834
use sg13g2_nand2_1  _322_
timestamp 1676560849
transform 1 0 4416 0 1 5292
box -48 -56 432 834
use sg13g2_nand2_1  _323_
timestamp 1676560849
transform 1 0 4320 0 -1 8316
box -48 -56 432 834
use sg13g2_xor2_1  _324_
timestamp 1677581577
transform 1 0 5568 0 -1 8316
box -48 -56 816 834
use sg13g2_a21o_2  _325_
timestamp 1683999997
transform 1 0 30720 0 -1 11340
box -48 -56 816 834
use sg13g2_nand2_1  _326_
timestamp 1676560849
transform 1 0 7200 0 -1 35532
box -48 -56 432 834
use sg13g2_nand2_1  _327_
timestamp 1676560849
transform -1 0 9504 0 1 35532
box -48 -56 432 834
use sg13g2_xor2_1  _328_
timestamp 1677581577
transform 1 0 8352 0 1 34020
box -48 -56 816 834
use sg13g2_nand2_1  _329_
timestamp 1676560849
transform 1 0 4416 0 -1 20412
box -48 -56 432 834
use sg13g2_nand2_1  _330_
timestamp 1676560849
transform 1 0 4416 0 -1 21924
box -48 -56 432 834
use sg13g2_xor2_1  _331_
timestamp 1677581577
transform 1 0 4800 0 -1 20412
box -48 -56 816 834
use sg13g2_nand2_1  _332_
timestamp 1676560849
transform 1 0 58368 0 1 9828
box -48 -56 432 834
use sg13g2_nand2_1  _333_
timestamp 1676560849
transform -1 0 59136 0 1 9828
box -48 -56 432 834
use sg13g2_xor2_1  _334_
timestamp 1677581577
transform 1 0 58656 0 -1 11340
box -48 -56 816 834
use sg13g2_nand2_1  _335_
timestamp 1676560849
transform 1 0 44736 0 1 29484
box -48 -56 432 834
use sg13g2_nand2_1  _336_
timestamp 1676560849
transform -1 0 46752 0 -1 30996
box -48 -56 432 834
use sg13g2_xor2_1  _337_
timestamp 1677581577
transform 1 0 44928 0 -1 30996
box -48 -56 816 834
use sg13g2_nand2_1  _338_
timestamp 1676560849
transform 1 0 27840 0 -1 20412
box -48 -56 432 834
use sg13g2_nand2_1  _339_
timestamp 1676560849
transform 1 0 28224 0 -1 20412
box -48 -56 432 834
use sg13g2_xor2_1  _340_
timestamp 1677581577
transform 1 0 28800 0 1 18900
box -48 -56 816 834
use sg13g2_nand2_1  _341_
timestamp 1676560849
transform -1 0 43680 0 -1 24948
box -48 -56 432 834
use sg13g2_nand2_1  _342_
timestamp 1676560849
transform -1 0 45792 0 1 23436
box -48 -56 432 834
use sg13g2_xor2_1  _343_
timestamp 1677581577
transform 1 0 43392 0 1 23436
box -48 -56 816 834
use sg13g2_nand2_1  _344_
timestamp 1676560849
transform -1 0 34176 0 -1 24948
box -48 -56 432 834
use sg13g2_nand2_1  _345_
timestamp 1676560849
transform 1 0 34752 0 1 23436
box -48 -56 432 834
use sg13g2_xor2_1  _346_
timestamp 1677581577
transform 1 0 35136 0 1 23436
box -48 -56 816 834
use sg13g2_nand2_1  _347_
timestamp 1676560849
transform 1 0 50304 0 -1 3780
box -48 -56 432 834
use sg13g2_nand2_1  _348_
timestamp 1676560849
transform 1 0 49056 0 -1 3780
box -48 -56 432 834
use sg13g2_xor2_1  _349_
timestamp 1677581577
transform -1 0 49728 0 1 3780
box -48 -56 816 834
use sg13g2_nand2_1  _350_
timestamp 1676560849
transform -1 0 39648 0 1 5292
box -48 -56 432 834
use sg13g2_nand2_1  _351_
timestamp 1676560849
transform -1 0 41376 0 1 3780
box -48 -56 432 834
use sg13g2_xor2_1  _352_
timestamp 1677581577
transform 1 0 40992 0 -1 5292
box -48 -56 816 834
use sg13g2_nand2_1  _353_
timestamp 1676560849
transform 1 0 55104 0 -1 18900
box -48 -56 432 834
use sg13g2_nand2_1  _354_
timestamp 1676560849
transform 1 0 51072 0 1 17388
box -48 -56 432 834
use sg13g2_xor2_1  _355_
timestamp 1677581577
transform 1 0 55104 0 1 17388
box -48 -56 816 834
use sg13g2_o21ai_1  _356_
timestamp 1685179043
transform -1 0 33408 0 -1 9828
box -48 -56 538 834
use sg13g2_nand2_1  _357_
timestamp 1676560849
transform 1 0 17952 0 1 2268
box -48 -56 432 834
use sg13g2_nand2_1  _358_
timestamp 1676560849
transform 1 0 17376 0 1 2268
box -48 -56 432 834
use sg13g2_xor2_1  _359_
timestamp 1677581577
transform 1 0 18624 0 1 2268
box -48 -56 816 834
use sg13g2_nand2_1  _360_
timestamp 1676560849
transform 1 0 4128 0 -1 27972
box -48 -56 432 834
use sg13g2_nand2_1  _361_
timestamp 1676560849
transform 1 0 4512 0 -1 27972
box -48 -56 432 834
use sg13g2_xor2_1  _362_
timestamp 1677581577
transform 1 0 5376 0 -1 27972
box -48 -56 816 834
use sg13g2_nand2_1  _363_
timestamp 1676560849
transform -1 0 18144 0 -1 15876
box -48 -56 432 834
use sg13g2_nand2_1  _364_
timestamp 1676560849
transform 1 0 17376 0 -1 15876
box -48 -56 432 834
use sg13g2_xor2_1  _365_
timestamp 1677581577
transform 1 0 18144 0 -1 15876
box -48 -56 816 834
use sg13g2_nand2_1  _366_
timestamp 1676560849
transform 1 0 16992 0 -1 30996
box -48 -56 432 834
use sg13g2_nand2_1  _367_
timestamp 1676560849
transform 1 0 16896 0 -1 32508
box -48 -56 432 834
use sg13g2_xor2_1  _368_
timestamp 1677581577
transform 1 0 17376 0 -1 30996
box -48 -56 816 834
use sg13g2_nand2_1  _369_
timestamp 1676560849
transform 1 0 21216 0 -1 35532
box -48 -56 432 834
use sg13g2_nand2_1  _370_
timestamp 1676560849
transform 1 0 22080 0 1 35532
box -48 -56 432 834
use sg13g2_xor2_1  _371_
timestamp 1677581577
transform 1 0 21600 0 -1 35532
box -48 -56 816 834
use sg13g2_nand2_1  _372_
timestamp 1676560849
transform 1 0 33024 0 -1 35532
box -48 -56 432 834
use sg13g2_nand2_1  _373_
timestamp 1676560849
transform -1 0 36384 0 1 35532
box -48 -56 432 834
use sg13g2_xor2_1  _374_
timestamp 1677581577
transform 1 0 35712 0 -1 35532
box -48 -56 816 834
use sg13g2_o21ai_1  _375_
timestamp 1685179043
transform 1 0 23424 0 -1 12852
box -48 -56 538 834
use sg13g2_buf_1  _376_
timestamp 1676385511
transform -1 0 55008 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _377_
timestamp 1676385511
transform 1 0 59136 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _378_
timestamp 1676385511
transform -1 0 49632 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  _379_
timestamp 1676385511
transform 1 0 55200 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  _380_
timestamp 1676385511
transform -1 0 39552 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _381_
timestamp 1676385511
transform 1 0 37344 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _382_
timestamp 1676385511
transform -1 0 52224 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _383_
timestamp 1676385511
transform 1 0 51744 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _384_
timestamp 1676385511
transform -1 0 33600 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  _385_
timestamp 1676385511
transform 1 0 33312 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  _386_
timestamp 1676385511
transform -1 0 45120 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  _387_
timestamp 1676385511
transform -1 0 41760 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  _388_
timestamp 1676385511
transform -1 0 27360 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  _389_
timestamp 1676385511
transform -1 0 27168 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  _390_
timestamp 1676385511
transform -1 0 17664 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  _391_
timestamp 1676385511
transform -1 0 15936 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  _392_
timestamp 1676385511
transform -1 0 17184 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _393_
timestamp 1676385511
transform -1 0 17760 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _394_
timestamp 1676385511
transform -1 0 55872 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _395_
timestamp 1676385511
transform -1 0 60096 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  _396_
timestamp 1676385511
transform -1 0 52800 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  _397_
timestamp 1676385511
transform -1 0 49152 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  _398_
timestamp 1676385511
transform -1 0 38976 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _399_
timestamp 1676385511
transform 1 0 41760 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _400_
timestamp 1676385511
transform -1 0 48864 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _401_
timestamp 1676385511
transform 1 0 46560 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _402_
timestamp 1676385511
transform -1 0 31584 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  _403_
timestamp 1676385511
transform -1 0 34368 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  _404_
timestamp 1676385511
transform 1 0 44832 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  _405_
timestamp 1676385511
transform 1 0 46080 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  _406_
timestamp 1676385511
transform -1 0 26976 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  _407_
timestamp 1676385511
transform -1 0 26784 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  _408_
timestamp 1676385511
transform 1 0 18432 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  _409_
timestamp 1676385511
transform -1 0 16128 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  _410_
timestamp 1676385511
transform -1 0 13056 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _411_
timestamp 1676385511
transform -1 0 13632 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _412_
timestamp 1676385511
transform -1 0 45792 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  _413_
timestamp 1676385511
transform -1 0 44736 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  _414_
timestamp 1676385511
transform -1 0 35520 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _415_
timestamp 1676385511
transform -1 0 31488 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _416_
timestamp 1676385511
transform -1 0 24960 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _417_
timestamp 1676385511
transform -1 0 19584 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _418_
timestamp 1676385511
transform -1 0 16224 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  _419_
timestamp 1676385511
transform -1 0 15552 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  _420_
timestamp 1676385511
transform -1 0 4224 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  _421_
timestamp 1676385511
transform -1 0 3552 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  _422_
timestamp 1676385511
transform 1 0 9216 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _423_
timestamp 1676385511
transform -1 0 5952 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _424_
timestamp 1676385511
transform -1 0 4608 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  _425_
timestamp 1676385511
transform -1 0 3360 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  _426_
timestamp 1676385511
transform 1 0 9024 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  _427_
timestamp 1676385511
transform -1 0 5856 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  _428_
timestamp 1676385511
transform -1 0 4032 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _429_
timestamp 1676385511
transform 1 0 2880 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _430_
timestamp 1676385511
transform -1 0 43680 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  _431_
timestamp 1676385511
transform -1 0 47616 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  _432_
timestamp 1676385511
transform -1 0 31584 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _433_
timestamp 1676385511
transform -1 0 36768 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _434_
timestamp 1676385511
transform 1 0 23136 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _435_
timestamp 1676385511
transform -1 0 20160 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _436_
timestamp 1676385511
transform -1 0 16512 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  _437_
timestamp 1676385511
transform -1 0 15744 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  _438_
timestamp 1676385511
transform -1 0 3840 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  _439_
timestamp 1676385511
transform -1 0 3936 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  _440_
timestamp 1676385511
transform -1 0 5184 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _441_
timestamp 1676385511
transform -1 0 9600 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _442_
timestamp 1676385511
transform -1 0 3264 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  _443_
timestamp 1676385511
transform 1 0 2880 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  _444_
timestamp 1676385511
transform -1 0 4128 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  _445_
timestamp 1676385511
transform 1 0 9408 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  _446_
timestamp 1676385511
transform -1 0 4704 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _447_
timestamp 1676385511
transform -1 0 3456 0 1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _448_
timestamp 1746538728
transform 1 0 54048 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _449_
timestamp 1746538728
transform 1 0 59520 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _450_
timestamp 1746538728
transform 1 0 48672 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _451_
timestamp 1746538728
transform 1 0 55584 0 1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _452_
timestamp 1746538728
transform 1 0 38016 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _453_
timestamp 1746538728
transform -1 0 38496 0 -1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _454_
timestamp 1746538728
transform 1 0 51840 0 -1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _455_
timestamp 1746538728
transform 1 0 52128 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _456_
timestamp 1746538728
transform 1 0 32352 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _457_
timestamp 1746538728
transform -1 0 35040 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _458_
timestamp 1746538728
transform 1 0 44352 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _459_
timestamp 1746538728
transform 1 0 40224 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _460_
timestamp 1746538728
transform 1 0 26112 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _461_
timestamp 1746538728
transform 1 0 25728 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _462_
timestamp 1746538728
transform 1 0 16800 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _463_
timestamp 1746538728
transform 1 0 14496 0 1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _464_
timestamp 1746538728
transform 1 0 16224 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _465_
timestamp 1746538728
transform 1 0 16608 0 1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _466_
timestamp 1746538728
transform 1 0 55200 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _467_
timestamp 1746538728
transform 1 0 59520 0 -1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _468_
timestamp 1746538728
transform 1 0 52032 0 -1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _469_
timestamp 1746538728
transform 1 0 47712 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _470_
timestamp 1746538728
transform 1 0 37824 0 -1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _471_
timestamp 1746538728
transform -1 0 43200 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _472_
timestamp 1746538728
transform 1 0 47520 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _473_
timestamp 1746538728
transform -1 0 47520 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _474_
timestamp 1746538728
transform 1 0 30144 0 1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _475_
timestamp 1746538728
transform 1 0 33984 0 1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _476_
timestamp 1746538728
transform 1 0 45120 0 1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _477_
timestamp 1746538728
transform 1 0 46464 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _478_
timestamp 1746538728
transform 1 0 25632 0 1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _479_
timestamp 1746538728
transform 1 0 25632 0 1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _480_
timestamp 1746538728
transform 1 0 18816 0 1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _481_
timestamp 1746538728
transform 1 0 14784 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _482_
timestamp 1746538728
transform 1 0 11712 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _483_
timestamp 1746538728
transform 1 0 12192 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _484_
timestamp 1746538728
transform 1 0 45312 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _485_
timestamp 1746538728
transform 1 0 44448 0 1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _486_
timestamp 1746538728
transform 1 0 35136 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _487_
timestamp 1746538728
transform 1 0 30144 0 1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _488_
timestamp 1746538728
transform 1 0 24480 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _489_
timestamp 1746538728
transform 1 0 18240 0 1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _490_
timestamp 1746538728
transform 1 0 14880 0 -1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _491_
timestamp 1746538728
transform 1 0 14304 0 1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _492_
timestamp 1746538728
transform 1 0 2784 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _493_
timestamp 1746538728
transform 1 0 2304 0 1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _494_
timestamp 1746538728
transform 1 0 9504 0 1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _495_
timestamp 1746538728
transform 1 0 4608 0 1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _496_
timestamp 1746538728
transform 1 0 3744 0 1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _497_
timestamp 1746538728
transform 1 0 2112 0 1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _498_
timestamp 1746538728
transform 1 0 9408 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _499_
timestamp 1746538728
transform 1 0 3936 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _500_
timestamp 1746538728
transform 1 0 2880 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _501_
timestamp 1746538728
transform -1 0 3840 0 -1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _502_
timestamp 1746538728
transform 1 0 42432 0 -1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _503_
timestamp 1746538728
transform 1 0 46848 0 1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _504_
timestamp 1746538728
transform 1 0 30240 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _505_
timestamp 1746538728
transform 1 0 36480 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _506_
timestamp 1746538728
transform 1 0 23520 0 1 35532
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _507_
timestamp 1746538728
transform 1 0 18720 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _508_
timestamp 1746538728
transform 1 0 15360 0 -1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _509_
timestamp 1746538728
transform 1 0 14400 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _510_
timestamp 1746538728
transform 1 0 2688 0 -1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _511_
timestamp 1746538728
transform 1 0 2400 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _512_
timestamp 1746538728
transform 1 0 3840 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _513_
timestamp 1746538728
transform 1 0 9312 0 -1 37044
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _514_
timestamp 1746538728
transform 1 0 2208 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _515_
timestamp 1746538728
transform -1 0 3744 0 1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _516_
timestamp 1746538728
transform 1 0 2880 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _517_
timestamp 1746538728
transform 1 0 9792 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _518_
timestamp 1746538728
transform 1 0 3840 0 -1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _519_
timestamp 1746538728
transform 1 0 2208 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _520_
timestamp 1746538728
transform -1 0 46944 0 1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _521_
timestamp 1746538728
transform -1 0 43392 0 1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _522_
timestamp 1746538728
transform 1 0 36192 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _523_
timestamp 1746538728
transform 1 0 36768 0 -1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _524_
timestamp 1746538728
transform -1 0 50688 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _525_
timestamp 1746538728
transform -1 0 56160 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _526_
timestamp 1746538728
transform 1 0 46752 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _527_
timestamp 1746538728
transform 1 0 48000 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _528_
timestamp 1746538728
transform 1 0 19296 0 -1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _529_
timestamp 1746538728
transform 1 0 20832 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _530_
timestamp 1746538728
transform -1 0 39552 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _531_
timestamp 1746538728
transform -1 0 43200 0 -1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _532_
timestamp 1746538728
transform -1 0 52896 0 1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _533_
timestamp 1746538728
transform -1 0 48864 0 1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _534_
timestamp 1746538728
transform 1 0 35328 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _535_
timestamp 1746538728
transform 1 0 36192 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _536_
timestamp 1746538728
transform 1 0 23712 0 1 3780
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _537_
timestamp 1746538728
transform 1 0 24576 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _538_
timestamp 1746538728
transform 1 0 21216 0 1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _539_
timestamp 1746538728
transform 1 0 25248 0 -1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _540_
timestamp 1746538728
transform 1 0 42048 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _541_
timestamp 1746538728
transform 1 0 42144 0 1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _542_
timestamp 1746538728
transform -1 0 44448 0 -1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _543_
timestamp 1746538728
transform -1 0 46752 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _544_
timestamp 1746538728
transform 1 0 52704 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _545_
timestamp 1746538728
transform 1 0 56544 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _546_
timestamp 1746538728
transform 1 0 38400 0 1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _547_
timestamp 1746538728
transform 1 0 41664 0 -1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _548_
timestamp 1746538728
transform 1 0 27648 0 -1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _549_
timestamp 1746538728
transform 1 0 28128 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _550_
timestamp 1746538728
transform 1 0 54336 0 -1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _551_
timestamp 1746538728
transform 1 0 58944 0 -1 14364
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _552_
timestamp 1746538728
transform 1 0 31008 0 1 15876
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _553_
timestamp 1746538728
transform 1 0 31008 0 1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _554_
timestamp 1746538728
transform 1 0 22944 0 1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _555_
timestamp 1746538728
transform -1 0 30144 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _556_
timestamp 1746538728
transform -1 0 32832 0 1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _557_
timestamp 1746538728
transform -1 0 39648 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_2  _558_
timestamp 1746538784
transform -1 0 38400 0 -1 11340
box -48 -56 2736 834
use sg13g2_dfrbpq_1  _559_
timestamp 1746538728
transform 1 0 31008 0 1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_2  _560_
timestamp 1746538784
transform 1 0 31008 0 -1 3780
box -48 -56 2736 834
use sg13g2_dfrbpq_1  _561_
timestamp 1746538728
transform 1 0 8736 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _562_
timestamp 1746538728
transform 1 0 8736 0 -1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _563_
timestamp 1746538728
transform 1 0 7008 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _564_
timestamp 1746538728
transform 1 0 7776 0 -1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_2  _565_
timestamp 1746538784
transform -1 0 40992 0 -1 27972
box -48 -56 2736 834
use sg13g2_dfrbpq_1  _566_
timestamp 1746538728
transform -1 0 32928 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _567_
timestamp 1746538728
transform 1 0 26112 0 -1 27972
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _568_
timestamp 1746538728
transform 1 0 27264 0 1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _569_
timestamp 1746538728
transform 1 0 6912 0 -1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _570_
timestamp 1746538728
transform 1 0 6720 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _571_
timestamp 1746538728
transform 1 0 11328 0 1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _572_
timestamp 1746538728
transform 1 0 11616 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _573_
timestamp 1746538728
transform 1 0 20736 0 1 29484
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _574_
timestamp 1746538728
transform 1 0 20064 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _575_
timestamp 1746538728
transform 1 0 13536 0 1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _576_
timestamp 1746538728
transform 1 0 13536 0 1 20412
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _577_
timestamp 1746538728
transform 1 0 9696 0 1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _578_
timestamp 1746538728
transform 1 0 10272 0 -1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _579_
timestamp 1746538728
transform 1 0 9504 0 -1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _580_
timestamp 1746538728
transform 1 0 8544 0 1 17388
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _581_
timestamp 1746538728
transform 1 0 25536 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _582_
timestamp 1746538728
transform 1 0 21696 0 1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _583_
timestamp 1746538728
transform -1 0 27264 0 -1 24948
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _584_
timestamp 1746538728
transform -1 0 24096 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _585_
timestamp 1746538728
transform 1 0 33792 0 -1 32508
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _586_
timestamp 1746538728
transform 1 0 37248 0 1 34020
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _587_
timestamp 1746538728
transform 1 0 17856 0 1 23436
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _588_
timestamp 1746538728
transform 1 0 18624 0 -1 26460
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _589_
timestamp 1746538728
transform 1 0 12288 0 1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _590_
timestamp 1746538728
transform 1 0 12864 0 1 9828
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _591_
timestamp 1746538728
transform -1 0 38496 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _592_
timestamp 1746538728
transform -1 0 41952 0 -1 30996
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _593_
timestamp 1746538728
transform 1 0 7968 0 -1 21924
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _594_
timestamp 1746538728
transform 1 0 7296 0 1 18900
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _595_
timestamp 1746538728
transform 1 0 21888 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _596_
timestamp 1746538728
transform 1 0 24384 0 -1 11340
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _597_
timestamp 1746538728
transform 1 0 28224 0 -1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_2  _598_
timestamp 1746538784
transform 1 0 19872 0 1 18900
box -48 -56 2736 834
use sg13g2_dfrbpq_2  _599_
timestamp 1746538784
transform 1 0 20928 0 -1 20412
box -48 -56 2736 834
use sg13g2_dfrbpq_1  _600_
timestamp 1746538728
transform 1 0 16608 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _601_
timestamp 1746538728
transform 1 0 16224 0 -1 11340
box -48 -56 2640 834
use sg13g2_buf_8  clkbuf_0_clk
timestamp 1676454965
transform 1 0 31008 0 -1 20412
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_0_0_clk
timestamp 1676454965
transform -1 0 10464 0 -1 11340
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_1_0_clk
timestamp 1676454965
transform -1 0 9696 0 -1 12852
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_2_0_clk
timestamp 1676454965
transform -1 0 21888 0 -1 11340
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_3_0_clk
timestamp 1676454965
transform -1 0 19680 0 -1 12852
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_4_0_clk
timestamp 1676454965
transform -1 0 9984 0 -1 27972
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_5_0_clk
timestamp 1676454965
transform -1 0 10368 0 1 29484
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_6_0_clk
timestamp 1676454965
transform -1 0 23328 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_7_0_clk
timestamp 1676454965
transform -1 0 22848 0 1 30996
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_8_0_clk
timestamp 1676454965
transform -1 0 38688 0 1 8316
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_9_0_clk
timestamp 1676454965
transform -1 0 39360 0 1 9828
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_10_0_clk
timestamp 1676454965
transform -1 0 53760 0 -1 9828
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_11_0_clk
timestamp 1676454965
transform 1 0 53376 0 1 11340
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_12_0_clk
timestamp 1676454965
transform -1 0 35424 0 -1 24948
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_13_0_clk
timestamp 1676454965
transform -1 0 36768 0 -1 26460
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_14_0_clk
timestamp 1676454965
transform -1 0 46464 0 -1 24948
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_4_15_0_clk
timestamp 1676454965
transform -1 0 44640 0 -1 26460
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_0__f_clk
timestamp 1676454965
transform -1 0 7776 0 -1 8316
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_1__f_clk
timestamp 1676454965
transform 1 0 11040 0 1 6804
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_2__f_clk
timestamp 1676454965
transform -1 0 6528 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_3__f_clk
timestamp 1676454965
transform 1 0 10080 0 1 15876
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_4__f_clk
timestamp 1676454965
transform -1 0 20832 0 1 5292
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_5__f_clk
timestamp 1676454965
transform 1 0 23328 0 1 8316
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_6__f_clk
timestamp 1676454965
transform -1 0 17184 0 -1 15876
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_7__f_clk
timestamp 1676454965
transform 1 0 20256 0 -1 17388
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_8__f_clk
timestamp 1676454965
transform -1 0 7008 0 1 24948
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_9__f_clk
timestamp 1676454965
transform 1 0 11712 0 -1 24948
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_10__f_clk
timestamp 1676454965
transform -1 0 7680 0 1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_11__f_clk
timestamp 1676454965
transform 1 0 10944 0 -1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_12__f_clk
timestamp 1676454965
transform -1 0 20832 0 1 27972
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_13__f_clk
timestamp 1676454965
transform 1 0 24096 0 1 24948
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_14__f_clk
timestamp 1676454965
transform -1 0 21024 0 1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_15__f_clk
timestamp 1676454965
transform 1 0 24384 0 -1 34020
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_16__f_clk
timestamp 1676454965
transform -1 0 35520 0 -1 6804
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_17__f_clk
timestamp 1676454965
transform 1 0 39744 0 -1 5292
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_18__f_clk
timestamp 1676454965
transform -1 0 36096 0 -1 12852
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_19__f_clk
timestamp 1676454965
transform 1 0 41472 0 1 11340
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_20__f_clk
timestamp 1676454965
transform -1 0 50016 0 1 6804
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_21__f_clk
timestamp 1676454965
transform 1 0 56256 0 1 6804
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_22__f_clk
timestamp 1676454965
transform -1 0 52416 0 1 14364
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_23__f_clk
timestamp 1676454965
transform 1 0 56832 0 -1 14364
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_24__f_clk
timestamp 1676454965
transform -1 0 32352 0 -1 21924
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_25__f_clk
timestamp 1676454965
transform 1 0 34752 0 1 18900
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_26__f_clk
timestamp 1676454965
transform -1 0 35328 0 -1 30996
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_27__f_clk
timestamp 1676454965
transform 1 0 36288 0 1 30996
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_28__f_clk
timestamp 1676454965
transform -1 0 44256 0 -1 21924
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_29__f_clk
timestamp 1676454965
transform 1 0 49152 0 1 21924
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_30__f_clk
timestamp 1676454965
transform -1 0 41184 0 1 27972
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_5_31__f_clk
timestamp 1676454965
transform 1 0 45120 0 1 29484
box -48 -56 1296 834
use sg13g2_inv_1  clkload0
timestamp 1676386529
transform 1 0 20352 0 -1 15876
box -48 -56 336 834
use sg13g2_inv_1  clkload1
timestamp 1676386529
transform 1 0 10656 0 -1 34020
box -48 -56 336 834
use sg13g2_buf_1  clkload2
timestamp 1676385511
transform 1 0 19200 0 1 27972
box -48 -56 432 834
use sg13g2_inv_1  clkload3
timestamp 1676386529
transform -1 0 24384 0 -1 34020
box -48 -56 336 834
use sg13g2_buf_1  clkload4
timestamp 1676385511
transform 1 0 39360 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  clkload5
timestamp 1676385511
transform 1 0 41088 0 -1 12852
box -48 -56 432 834
use sg13g2_inv_1  clkload6
timestamp 1676386529
transform 1 0 56544 0 1 12852
box -48 -56 336 834
use sg13g2_inv_1  clkload7
timestamp 1676386529
transform -1 0 35904 0 -1 30996
box -48 -56 336 834
use sg13g2_inv_1  clkload8
timestamp 1676386529
transform 1 0 44448 0 1 29484
box -48 -56 336 834
use sg13g2_buf_8  fanout56
timestamp 1676454965
transform 1 0 17856 0 -1 8316
box -48 -56 1296 834
use sg13g2_buf_8  fanout57
timestamp 1676454965
transform -1 0 13344 0 -1 6804
box -48 -56 1296 834
use sg13g2_buf_2  fanout58
timestamp 1676385467
transform 1 0 12384 0 1 9828
box -48 -56 528 834
use sg13g2_buf_8  fanout59
timestamp 1676454965
transform -1 0 19296 0 1 11340
box -48 -56 1296 834
use sg13g2_buf_8  fanout60
timestamp 1676454965
transform -1 0 28032 0 -1 14364
box -48 -56 1296 834
use sg13g2_buf_8  fanout61
timestamp 1676454965
transform 1 0 21120 0 -1 12852
box -48 -56 1296 834
use sg13g2_buf_8  fanout62
timestamp 1676454965
transform -1 0 20928 0 -1 20412
box -48 -56 1296 834
use sg13g2_buf_8  fanout63
timestamp 1676454965
transform 1 0 3264 0 1 18900
box -48 -56 1296 834
use sg13g2_buf_8  fanout64
timestamp 1676454965
transform -1 0 10176 0 1 21924
box -48 -56 1296 834
use sg13g2_buf_8  fanout65
timestamp 1676454965
transform 1 0 3744 0 1 30996
box -48 -56 1296 834
use sg13g2_buf_1  fanout66
timestamp 1676385511
transform -1 0 15360 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_8  fanout67
timestamp 1676454965
transform 1 0 14592 0 -1 21924
box -48 -56 1296 834
use sg13g2_buf_8  fanout68
timestamp 1676454965
transform -1 0 20736 0 1 20412
box -48 -56 1296 834
use sg13g2_buf_8  fanout69
timestamp 1676454965
transform 1 0 36864 0 1 9828
box -48 -56 1296 834
use sg13g2_buf_8  fanout70
timestamp 1676454965
transform -1 0 43872 0 1 17388
box -48 -56 1296 834
use sg13g2_buf_8  fanout71
timestamp 1676454965
transform -1 0 52800 0 -1 11340
box -48 -56 1296 834
use sg13g2_buf_8  fanout72
timestamp 1676454965
transform 1 0 52992 0 -1 12852
box -48 -56 1296 834
use sg13g2_buf_8  fanout73
timestamp 1676454965
transform 1 0 45696 0 1 15876
box -48 -56 1296 834
use sg13g2_buf_8  fanout74
timestamp 1676454965
transform 1 0 44928 0 -1 17388
box -48 -56 1296 834
use sg13g2_buf_8  fanout75
timestamp 1676454965
transform 1 0 32256 0 -1 20412
box -48 -56 1296 834
use sg13g2_buf_8  fanout76
timestamp 1676454965
transform -1 0 27264 0 1 29484
box -48 -56 1296 834
use sg13g2_buf_8  fanout77
timestamp 1676454965
transform 1 0 28512 0 1 24948
box -48 -56 1296 834
use sg13g2_buf_8  fanout78
timestamp 1676454965
transform 1 0 39744 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  fanout79
timestamp 1676454965
transform -1 0 34272 0 1 30996
box -48 -56 1296 834
use sg13g2_buf_8  fanout80
timestamp 1676454965
transform 1 0 32736 0 1 27972
box -48 -56 1296 834
use sg13g2_buf_8  fanout81
timestamp 1676454965
transform 1 0 20832 0 1 20412
box -48 -56 1296 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679585382
transform 1 0 576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679585382
transform 1 0 1248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679585382
transform 1 0 1920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679585382
transform 1 0 2592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679585382
transform 1 0 3264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679585382
transform 1 0 3936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679585382
transform 1 0 4608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679585382
transform 1 0 5280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679585382
transform 1 0 5952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679585382
transform 1 0 6624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679585382
transform 1 0 7296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679585382
transform 1 0 7968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679585382
transform 1 0 8640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679585382
transform 1 0 9312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679585382
transform 1 0 9984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679585382
transform 1 0 10656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679585382
transform 1 0 11328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679585382
transform 1 0 12000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679585382
transform 1 0 12672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679585382
transform 1 0 13344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679585382
transform 1 0 14016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679585382
transform 1 0 14688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679585382
transform 1 0 15360 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679585382
transform 1 0 16032 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679585382
transform 1 0 16704 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679585382
transform 1 0 17376 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679585382
transform 1 0 18048 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679585382
transform 1 0 18720 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1679585382
transform 1 0 19392 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1679585382
transform 1 0 20064 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1679585382
transform 1 0 20736 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1679585382
transform 1 0 21408 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_224
timestamp 1679585382
transform 1 0 22080 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_231
timestamp 1679585382
transform 1 0 22752 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_238
timestamp 1679585382
transform 1 0 23424 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_245
timestamp 1679585382
transform 1 0 24096 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_252
timestamp 1679585382
transform 1 0 24768 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_259
timestamp 1679585382
transform 1 0 25440 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_266
timestamp 1679585382
transform 1 0 26112 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_273
timestamp 1679585382
transform 1 0 26784 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_280
timestamp 1679585382
transform 1 0 27456 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_287
timestamp 1679585382
transform 1 0 28128 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_294
timestamp 1679585382
transform 1 0 28800 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_301
timestamp 1679585382
transform 1 0 29472 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_308
timestamp 1679585382
transform 1 0 30144 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_315
timestamp 1679585382
transform 1 0 30816 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_322
timestamp 1679585382
transform 1 0 31488 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_329
timestamp 1679585382
transform 1 0 32160 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_336
timestamp 1679585382
transform 1 0 32832 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_343
timestamp 1679585382
transform 1 0 33504 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_350
timestamp 1679585382
transform 1 0 34176 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_357
timestamp 1679585382
transform 1 0 34848 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_364
timestamp 1679585382
transform 1 0 35520 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_371
timestamp 1679585382
transform 1 0 36192 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_378
timestamp 1679585382
transform 1 0 36864 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_385
timestamp 1679585382
transform 1 0 37536 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_392
timestamp 1679585382
transform 1 0 38208 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_399
timestamp 1679585382
transform 1 0 38880 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_406
timestamp 1679585382
transform 1 0 39552 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_413
timestamp 1679585382
transform 1 0 40224 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_420
timestamp 1679585382
transform 1 0 40896 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_427
timestamp 1679585382
transform 1 0 41568 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_434
timestamp 1679585382
transform 1 0 42240 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_441
timestamp 1679585382
transform 1 0 42912 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_448
timestamp 1679585382
transform 1 0 43584 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_455
timestamp 1679585382
transform 1 0 44256 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_462
timestamp 1679585382
transform 1 0 44928 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_469
timestamp 1679585382
transform 1 0 45600 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_476
timestamp 1679585382
transform 1 0 46272 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_483
timestamp 1679585382
transform 1 0 46944 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_490
timestamp 1679585382
transform 1 0 47616 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_497
timestamp 1679585382
transform 1 0 48288 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_504
timestamp 1679585382
transform 1 0 48960 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_511
timestamp 1679585382
transform 1 0 49632 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_518
timestamp 1679585382
transform 1 0 50304 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_525
timestamp 1679585382
transform 1 0 50976 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_532
timestamp 1679585382
transform 1 0 51648 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_539
timestamp 1679585382
transform 1 0 52320 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_546
timestamp 1679585382
transform 1 0 52992 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_553
timestamp 1679585382
transform 1 0 53664 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_560
timestamp 1679585382
transform 1 0 54336 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_567
timestamp 1679585382
transform 1 0 55008 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_574
timestamp 1679585382
transform 1 0 55680 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_581
timestamp 1679585382
transform 1 0 56352 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_588
timestamp 1679585382
transform 1 0 57024 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_595
timestamp 1679585382
transform 1 0 57696 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_602
timestamp 1679585382
transform 1 0 58368 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_609
timestamp 1679585382
transform 1 0 59040 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_616
timestamp 1679585382
transform 1 0 59712 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_623
timestamp 1679585382
transform 1 0 60384 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_630
timestamp 1679585382
transform 1 0 61056 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_637
timestamp 1679585382
transform 1 0 61728 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_644
timestamp 1679585382
transform 1 0 62400 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_651
timestamp 1679585382
transform 1 0 63072 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_658
timestamp 1679585382
transform 1 0 63744 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_665
timestamp 1679585382
transform 1 0 64416 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_672
timestamp 1679585382
transform 1 0 65088 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_679
timestamp 1679585382
transform 1 0 65760 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_686
timestamp 1679585382
transform 1 0 66432 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_693
timestamp 1679585382
transform 1 0 67104 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_700
timestamp 1679585382
transform 1 0 67776 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_707
timestamp 1679585382
transform 1 0 68448 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_714
timestamp 1679585382
transform 1 0 69120 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_721
timestamp 1679585382
transform 1 0 69792 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_728
timestamp 1679585382
transform 1 0 70464 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_735
timestamp 1679585382
transform 1 0 71136 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_742
timestamp 1679585382
transform 1 0 71808 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_749
timestamp 1679585382
transform 1 0 72480 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_756
timestamp 1679585382
transform 1 0 73152 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_763
timestamp 1679585382
transform 1 0 73824 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_770
timestamp 1679585382
transform 1 0 74496 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_777
timestamp 1679585382
transform 1 0 75168 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_784
timestamp 1679585382
transform 1 0 75840 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_791
timestamp 1679585382
transform 1 0 76512 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_798
timestamp 1679585382
transform 1 0 77184 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_805
timestamp 1679585382
transform 1 0 77856 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_812
timestamp 1679585382
transform 1 0 78528 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_819
timestamp 1679585382
transform 1 0 79200 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_826
timestamp 1679585382
transform 1 0 79872 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_833
timestamp 1679585382
transform 1 0 80544 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_840
timestamp 1679585382
transform 1 0 81216 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_847
timestamp 1679585382
transform 1 0 81888 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_854
timestamp 1679585382
transform 1 0 82560 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_861
timestamp 1679585382
transform 1 0 83232 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_868
timestamp 1679585382
transform 1 0 83904 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_875
timestamp 1679585382
transform 1 0 84576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_882
timestamp 1679585382
transform 1 0 85248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_889
timestamp 1679585382
transform 1 0 85920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_896
timestamp 1679585382
transform 1 0 86592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_903
timestamp 1679585382
transform 1 0 87264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_910
timestamp 1679585382
transform 1 0 87936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_917
timestamp 1679585382
transform 1 0 88608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_924
timestamp 1679585382
transform 1 0 89280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_931
timestamp 1679585382
transform 1 0 89952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_938
timestamp 1679585382
transform 1 0 90624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_945
timestamp 1679585382
transform 1 0 91296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_952
timestamp 1679585382
transform 1 0 91968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_959
timestamp 1679585382
transform 1 0 92640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_966
timestamp 1679585382
transform 1 0 93312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_973
timestamp 1679585382
transform 1 0 93984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_980
timestamp 1679585382
transform 1 0 94656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_987
timestamp 1679585382
transform 1 0 95328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_994
timestamp 1679585382
transform 1 0 96000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1001
timestamp 1679585382
transform 1 0 96672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1008
timestamp 1679585382
transform 1 0 97344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1015
timestamp 1679585382
transform 1 0 98016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1022
timestamp 1679585382
transform 1 0 98688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679585382
transform 1 0 576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679585382
transform 1 0 1248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679585382
transform 1 0 1920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679585382
transform 1 0 2592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679585382
transform 1 0 3264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679585382
transform 1 0 3936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679585382
transform 1 0 4608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679585382
transform 1 0 5280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679585382
transform 1 0 5952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679585382
transform 1 0 6624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679585382
transform 1 0 7296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679585382
transform 1 0 7968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679585382
transform 1 0 8640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1679585382
transform 1 0 9312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1679585382
transform 1 0 9984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679585382
transform 1 0 10656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679585382
transform 1 0 11328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1679585382
transform 1 0 12000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_126
timestamp 1679581501
transform 1 0 12672 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_130
timestamp 1677583704
transform 1 0 13056 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_136
timestamp 1679585382
transform 1 0 13632 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_143
timestamp 1679585382
transform 1 0 14304 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_150
timestamp 1679585382
transform 1 0 14976 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_157
timestamp 1679585382
transform 1 0 15648 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_164
timestamp 1679585382
transform 1 0 16320 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_171
timestamp 1679585382
transform 1 0 16992 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_178
timestamp 1679585382
transform 1 0 17664 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_185
timestamp 1679585382
transform 1 0 18336 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_192
timestamp 1679585382
transform 1 0 19008 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_199
timestamp 1679585382
transform 1 0 19680 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_206
timestamp 1679585382
transform 1 0 20352 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_213
timestamp 1679585382
transform 1 0 21024 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_220
timestamp 1679585382
transform 1 0 21696 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_227
timestamp 1679585382
transform 1 0 22368 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_234
timestamp 1679585382
transform 1 0 23040 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_241
timestamp 1679585382
transform 1 0 23712 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_248
timestamp 1679585382
transform 1 0 24384 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_255
timestamp 1679585382
transform 1 0 25056 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_262
timestamp 1679585382
transform 1 0 25728 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_269
timestamp 1679585382
transform 1 0 26400 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_276
timestamp 1679585382
transform 1 0 27072 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_283
timestamp 1679585382
transform 1 0 27744 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_290
timestamp 1679585382
transform 1 0 28416 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_297
timestamp 1679585382
transform 1 0 29088 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_304
timestamp 1679585382
transform 1 0 29760 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_311
timestamp 1679585382
transform 1 0 30432 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_318
timestamp 1679585382
transform 1 0 31104 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_325
timestamp 1679585382
transform 1 0 31776 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_332
timestamp 1679585382
transform 1 0 32448 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_339
timestamp 1679585382
transform 1 0 33120 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_346
timestamp 1679585382
transform 1 0 33792 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_353
timestamp 1679585382
transform 1 0 34464 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_360
timestamp 1679585382
transform 1 0 35136 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_367
timestamp 1679585382
transform 1 0 35808 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_374
timestamp 1679585382
transform 1 0 36480 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_381
timestamp 1679585382
transform 1 0 37152 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_388
timestamp 1679585382
transform 1 0 37824 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_395
timestamp 1679585382
transform 1 0 38496 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_402
timestamp 1679585382
transform 1 0 39168 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_409
timestamp 1679585382
transform 1 0 39840 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_416
timestamp 1679585382
transform 1 0 40512 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_423
timestamp 1679585382
transform 1 0 41184 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_430
timestamp 1679585382
transform 1 0 41856 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_437
timestamp 1679585382
transform 1 0 42528 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_444
timestamp 1679585382
transform 1 0 43200 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_451
timestamp 1679585382
transform 1 0 43872 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_458
timestamp 1679585382
transform 1 0 44544 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_465
timestamp 1679585382
transform 1 0 45216 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_472
timestamp 1679585382
transform 1 0 45888 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_479
timestamp 1679585382
transform 1 0 46560 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_486
timestamp 1679585382
transform 1 0 47232 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_493
timestamp 1679585382
transform 1 0 47904 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_500
timestamp 1679585382
transform 1 0 48576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_507
timestamp 1679585382
transform 1 0 49248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_514
timestamp 1679585382
transform 1 0 49920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_521
timestamp 1679585382
transform 1 0 50592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_528
timestamp 1679585382
transform 1 0 51264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_535
timestamp 1679585382
transform 1 0 51936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_542
timestamp 1679585382
transform 1 0 52608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_549
timestamp 1679585382
transform 1 0 53280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_556
timestamp 1679585382
transform 1 0 53952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_563
timestamp 1679585382
transform 1 0 54624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_570
timestamp 1679585382
transform 1 0 55296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_577
timestamp 1679585382
transform 1 0 55968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_584
timestamp 1679585382
transform 1 0 56640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_591
timestamp 1679585382
transform 1 0 57312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_598
timestamp 1679585382
transform 1 0 57984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_605
timestamp 1679585382
transform 1 0 58656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_612
timestamp 1679585382
transform 1 0 59328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_619
timestamp 1679585382
transform 1 0 60000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_626
timestamp 1679585382
transform 1 0 60672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_633
timestamp 1679585382
transform 1 0 61344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_640
timestamp 1679585382
transform 1 0 62016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_647
timestamp 1679585382
transform 1 0 62688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_654
timestamp 1679585382
transform 1 0 63360 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_661
timestamp 1679585382
transform 1 0 64032 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_668
timestamp 1679585382
transform 1 0 64704 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_675
timestamp 1679585382
transform 1 0 65376 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_682
timestamp 1679585382
transform 1 0 66048 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_689
timestamp 1679585382
transform 1 0 66720 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_696
timestamp 1679585382
transform 1 0 67392 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_703
timestamp 1679585382
transform 1 0 68064 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_710
timestamp 1679585382
transform 1 0 68736 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_717
timestamp 1679585382
transform 1 0 69408 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_724
timestamp 1679585382
transform 1 0 70080 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_731
timestamp 1679585382
transform 1 0 70752 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_738
timestamp 1679585382
transform 1 0 71424 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_745
timestamp 1679585382
transform 1 0 72096 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_752
timestamp 1679585382
transform 1 0 72768 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_759
timestamp 1679585382
transform 1 0 73440 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_766
timestamp 1679585382
transform 1 0 74112 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_773
timestamp 1679585382
transform 1 0 74784 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_780
timestamp 1679585382
transform 1 0 75456 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_787
timestamp 1679585382
transform 1 0 76128 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_794
timestamp 1679585382
transform 1 0 76800 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_801
timestamp 1679585382
transform 1 0 77472 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_808
timestamp 1679585382
transform 1 0 78144 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_815
timestamp 1679585382
transform 1 0 78816 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_822
timestamp 1679585382
transform 1 0 79488 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_829
timestamp 1679585382
transform 1 0 80160 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_836
timestamp 1679585382
transform 1 0 80832 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_843
timestamp 1679585382
transform 1 0 81504 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_850
timestamp 1679585382
transform 1 0 82176 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_857
timestamp 1679585382
transform 1 0 82848 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_864
timestamp 1679585382
transform 1 0 83520 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_871
timestamp 1679585382
transform 1 0 84192 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_878
timestamp 1679585382
transform 1 0 84864 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_885
timestamp 1679585382
transform 1 0 85536 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_892
timestamp 1679585382
transform 1 0 86208 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_899
timestamp 1679585382
transform 1 0 86880 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_906
timestamp 1679585382
transform 1 0 87552 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_913
timestamp 1679585382
transform 1 0 88224 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_920
timestamp 1679585382
transform 1 0 88896 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_927
timestamp 1679585382
transform 1 0 89568 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_934
timestamp 1679585382
transform 1 0 90240 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_941
timestamp 1679585382
transform 1 0 90912 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_948
timestamp 1679585382
transform 1 0 91584 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_955
timestamp 1679585382
transform 1 0 92256 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_962
timestamp 1679585382
transform 1 0 92928 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_969
timestamp 1679585382
transform 1 0 93600 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_976
timestamp 1679585382
transform 1 0 94272 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_983
timestamp 1679585382
transform 1 0 94944 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_990
timestamp 1679585382
transform 1 0 95616 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_997
timestamp 1679585382
transform 1 0 96288 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1004
timestamp 1679585382
transform 1 0 96960 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1011
timestamp 1679585382
transform 1 0 97632 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1018
timestamp 1679585382
transform 1 0 98304 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_1025
timestamp 1679581501
transform 1 0 98976 0 -1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_4
timestamp 1679585382
transform 1 0 960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_11
timestamp 1679585382
transform 1 0 1632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_18
timestamp 1679585382
transform 1 0 2304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_25
timestamp 1679585382
transform 1 0 2976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_32
timestamp 1679585382
transform 1 0 3648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_39
timestamp 1679585382
transform 1 0 4320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_46
timestamp 1679585382
transform 1 0 4992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_53
timestamp 1679585382
transform 1 0 5664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_60
timestamp 1679585382
transform 1 0 6336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_67
timestamp 1679585382
transform 1 0 7008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_74
timestamp 1679585382
transform 1 0 7680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_81
timestamp 1679585382
transform 1 0 8352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_88
timestamp 1679585382
transform 1 0 9024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_95
timestamp 1679585382
transform 1 0 9696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_102
timestamp 1679585382
transform 1 0 10368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_109
timestamp 1679585382
transform 1 0 11040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_116
timestamp 1679581501
transform 1 0 11712 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_120
timestamp 1677583258
transform 1 0 12096 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_157
timestamp 1679585382
transform 1 0 15648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_164
timestamp 1679581501
transform 1 0 16320 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_168
timestamp 1677583258
transform 1 0 16704 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_173
timestamp 1677583704
transform 1 0 17184 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_179
timestamp 1677583704
transform 1 0 17760 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_185
timestamp 1677583704
transform 1 0 18336 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_187
timestamp 1677583258
transform 1 0 18528 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_196
timestamp 1679585382
transform 1 0 19392 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_203
timestamp 1679585382
transform 1 0 20064 0 1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_210
timestamp 1677583258
transform 1 0 20736 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_238
timestamp 1677583704
transform 1 0 23424 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_240
timestamp 1677583258
transform 1 0 23616 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_277
timestamp 1677583258
transform 1 0 27168 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_314
timestamp 1679585382
transform 1 0 30720 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_321
timestamp 1679585382
transform 1 0 31392 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_328
timestamp 1679585382
transform 1 0 32064 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_335
timestamp 1679585382
transform 1 0 32736 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_342
timestamp 1679585382
transform 1 0 33408 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_349
timestamp 1679585382
transform 1 0 34080 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_356
timestamp 1679585382
transform 1 0 34752 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_363
timestamp 1679585382
transform 1 0 35424 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_370
timestamp 1679585382
transform 1 0 36096 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_377
timestamp 1679585382
transform 1 0 36768 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_384
timestamp 1679581501
transform 1 0 37440 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_388
timestamp 1677583704
transform 1 0 37824 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_444
timestamp 1679585382
transform 1 0 43200 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_451
timestamp 1679585382
transform 1 0 43872 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_458
timestamp 1679581501
transform 1 0 44544 0 1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_2_516
timestamp 1679585382
transform 1 0 50112 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_523
timestamp 1679585382
transform 1 0 50784 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_530
timestamp 1677583704
transform 1 0 51456 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_532
timestamp 1677583258
transform 1 0 51648 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_564
timestamp 1679585382
transform 1 0 54720 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_571
timestamp 1679585382
transform 1 0 55392 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_578
timestamp 1679585382
transform 1 0 56064 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_585
timestamp 1679585382
transform 1 0 56736 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_592
timestamp 1679585382
transform 1 0 57408 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_599
timestamp 1679585382
transform 1 0 58080 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_606
timestamp 1679585382
transform 1 0 58752 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_613
timestamp 1679585382
transform 1 0 59424 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_620
timestamp 1679585382
transform 1 0 60096 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_627
timestamp 1679585382
transform 1 0 60768 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_634
timestamp 1679585382
transform 1 0 61440 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_641
timestamp 1679585382
transform 1 0 62112 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_648
timestamp 1679585382
transform 1 0 62784 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_655
timestamp 1679585382
transform 1 0 63456 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_662
timestamp 1679585382
transform 1 0 64128 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_669
timestamp 1679585382
transform 1 0 64800 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_676
timestamp 1679585382
transform 1 0 65472 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_683
timestamp 1679585382
transform 1 0 66144 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_690
timestamp 1679585382
transform 1 0 66816 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_697
timestamp 1679585382
transform 1 0 67488 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_704
timestamp 1679585382
transform 1 0 68160 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_711
timestamp 1679585382
transform 1 0 68832 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_718
timestamp 1679585382
transform 1 0 69504 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_725
timestamp 1679585382
transform 1 0 70176 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_732
timestamp 1679585382
transform 1 0 70848 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_739
timestamp 1679585382
transform 1 0 71520 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_746
timestamp 1679585382
transform 1 0 72192 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_753
timestamp 1679585382
transform 1 0 72864 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_760
timestamp 1679585382
transform 1 0 73536 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_767
timestamp 1679585382
transform 1 0 74208 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_774
timestamp 1679585382
transform 1 0 74880 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_781
timestamp 1679585382
transform 1 0 75552 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_788
timestamp 1679585382
transform 1 0 76224 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_795
timestamp 1679585382
transform 1 0 76896 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_802
timestamp 1679585382
transform 1 0 77568 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_809
timestamp 1679585382
transform 1 0 78240 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_816
timestamp 1679585382
transform 1 0 78912 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_823
timestamp 1679585382
transform 1 0 79584 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_830
timestamp 1679585382
transform 1 0 80256 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_837
timestamp 1679585382
transform 1 0 80928 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_844
timestamp 1679585382
transform 1 0 81600 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_851
timestamp 1679585382
transform 1 0 82272 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_858
timestamp 1679585382
transform 1 0 82944 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_865
timestamp 1679585382
transform 1 0 83616 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_872
timestamp 1679585382
transform 1 0 84288 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_879
timestamp 1679585382
transform 1 0 84960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_886
timestamp 1679585382
transform 1 0 85632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_893
timestamp 1679585382
transform 1 0 86304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_900
timestamp 1679585382
transform 1 0 86976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_907
timestamp 1679585382
transform 1 0 87648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_914
timestamp 1679585382
transform 1 0 88320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_921
timestamp 1679585382
transform 1 0 88992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_928
timestamp 1679585382
transform 1 0 89664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_935
timestamp 1679585382
transform 1 0 90336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_942
timestamp 1679585382
transform 1 0 91008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_949
timestamp 1679585382
transform 1 0 91680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_956
timestamp 1679585382
transform 1 0 92352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_963
timestamp 1679585382
transform 1 0 93024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_970
timestamp 1679585382
transform 1 0 93696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_977
timestamp 1679585382
transform 1 0 94368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_984
timestamp 1679585382
transform 1 0 95040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_991
timestamp 1679585382
transform 1 0 95712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_998
timestamp 1679585382
transform 1 0 96384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1005
timestamp 1679585382
transform 1 0 97056 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1012
timestamp 1679585382
transform 1 0 97728 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1019
timestamp 1679585382
transform 1 0 98400 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_1026
timestamp 1677583704
transform 1 0 99072 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_1028
timestamp 1677583258
transform 1 0 99264 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_4
timestamp 1679585382
transform 1 0 960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_11
timestamp 1679585382
transform 1 0 1632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_18
timestamp 1679585382
transform 1 0 2304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_25
timestamp 1679585382
transform 1 0 2976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_32
timestamp 1679585382
transform 1 0 3648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_39
timestamp 1679585382
transform 1 0 4320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_46
timestamp 1679585382
transform 1 0 4992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_53
timestamp 1679585382
transform 1 0 5664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_60
timestamp 1679585382
transform 1 0 6336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_67
timestamp 1679585382
transform 1 0 7008 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_74
timestamp 1679585382
transform 1 0 7680 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_81
timestamp 1679585382
transform 1 0 8352 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_88
timestamp 1679585382
transform 1 0 9024 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_95
timestamp 1679585382
transform 1 0 9696 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_102
timestamp 1679585382
transform 1 0 10368 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_109
timestamp 1679585382
transform 1 0 11040 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_143
timestamp 1679585382
transform 1 0 14304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_150
timestamp 1679585382
transform 1 0 14976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_157
timestamp 1679581501
transform 1 0 15648 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_161
timestamp 1677583704
transform 1 0 16032 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_3_190
timestamp 1679581501
transform 1 0 18816 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_194
timestamp 1677583258
transform 1 0 19200 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_222
timestamp 1679585382
transform 1 0 21888 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_229
timestamp 1679585382
transform 1 0 22560 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_236
timestamp 1679585382
transform 1 0 23232 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_243
timestamp 1679585382
transform 1 0 23904 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_250
timestamp 1679585382
transform 1 0 24576 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_257
timestamp 1679585382
transform 1 0 25248 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_264
timestamp 1679585382
transform 1 0 25920 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_271
timestamp 1679585382
transform 1 0 26592 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_278
timestamp 1679585382
transform 1 0 27264 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_285
timestamp 1679585382
transform 1 0 27936 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_292
timestamp 1679585382
transform 1 0 28608 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_299
timestamp 1679585382
transform 1 0 29280 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_306
timestamp 1679585382
transform 1 0 29952 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_313
timestamp 1679581501
transform 1 0 30624 0 -1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_345
timestamp 1679585382
transform 1 0 33696 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_352
timestamp 1679585382
transform 1 0 34368 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_359
timestamp 1679585382
transform 1 0 35040 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_366
timestamp 1679585382
transform 1 0 35712 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_373
timestamp 1679585382
transform 1 0 36384 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_380
timestamp 1679585382
transform 1 0 37056 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_387
timestamp 1679585382
transform 1 0 37728 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_394
timestamp 1679585382
transform 1 0 38400 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_401
timestamp 1677583258
transform 1 0 39072 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_406
timestamp 1679581501
transform 1 0 39552 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_410
timestamp 1677583258
transform 1 0 39936 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_433
timestamp 1679585382
transform 1 0 42144 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_440
timestamp 1679585382
transform 1 0 42816 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_447
timestamp 1679585382
transform 1 0 43488 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_454
timestamp 1679585382
transform 1 0 44160 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_461
timestamp 1679585382
transform 1 0 44832 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_468
timestamp 1677583704
transform 1 0 45504 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_483
timestamp 1679585382
transform 1 0 46944 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_490
timestamp 1679585382
transform 1 0 47616 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_497
timestamp 1677583704
transform 1 0 48288 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_503
timestamp 1677583704
transform 1 0 48864 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_522
timestamp 1679585382
transform 1 0 50688 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_529
timestamp 1679585382
transform 1 0 51360 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_536
timestamp 1679585382
transform 1 0 52032 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_543
timestamp 1679581501
transform 1 0 52704 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_547
timestamp 1677583704
transform 1 0 53088 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_558
timestamp 1679585382
transform 1 0 54144 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_565
timestamp 1679585382
transform 1 0 54816 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_572
timestamp 1679585382
transform 1 0 55488 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_579
timestamp 1679585382
transform 1 0 56160 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_586
timestamp 1679585382
transform 1 0 56832 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_593
timestamp 1679585382
transform 1 0 57504 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_600
timestamp 1679585382
transform 1 0 58176 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_607
timestamp 1679585382
transform 1 0 58848 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_614
timestamp 1679585382
transform 1 0 59520 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_621
timestamp 1679585382
transform 1 0 60192 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_628
timestamp 1679585382
transform 1 0 60864 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_635
timestamp 1679585382
transform 1 0 61536 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_642
timestamp 1679585382
transform 1 0 62208 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_649
timestamp 1679585382
transform 1 0 62880 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_656
timestamp 1679585382
transform 1 0 63552 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_663
timestamp 1679585382
transform 1 0 64224 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_670
timestamp 1679585382
transform 1 0 64896 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_677
timestamp 1679585382
transform 1 0 65568 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_684
timestamp 1679585382
transform 1 0 66240 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_691
timestamp 1679585382
transform 1 0 66912 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_698
timestamp 1679585382
transform 1 0 67584 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_705
timestamp 1679585382
transform 1 0 68256 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_712
timestamp 1679585382
transform 1 0 68928 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_719
timestamp 1679585382
transform 1 0 69600 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_726
timestamp 1679585382
transform 1 0 70272 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_733
timestamp 1679585382
transform 1 0 70944 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_740
timestamp 1679585382
transform 1 0 71616 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_747
timestamp 1679585382
transform 1 0 72288 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_754
timestamp 1679585382
transform 1 0 72960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_761
timestamp 1679585382
transform 1 0 73632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_768
timestamp 1679585382
transform 1 0 74304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_775
timestamp 1679585382
transform 1 0 74976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_782
timestamp 1679585382
transform 1 0 75648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_789
timestamp 1679585382
transform 1 0 76320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_796
timestamp 1679585382
transform 1 0 76992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_803
timestamp 1679585382
transform 1 0 77664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_810
timestamp 1679585382
transform 1 0 78336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_817
timestamp 1679585382
transform 1 0 79008 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_824
timestamp 1679585382
transform 1 0 79680 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_831
timestamp 1679585382
transform 1 0 80352 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_838
timestamp 1679585382
transform 1 0 81024 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_845
timestamp 1679585382
transform 1 0 81696 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_852
timestamp 1679585382
transform 1 0 82368 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_859
timestamp 1679585382
transform 1 0 83040 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_866
timestamp 1679585382
transform 1 0 83712 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_873
timestamp 1679585382
transform 1 0 84384 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_880
timestamp 1679585382
transform 1 0 85056 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_887
timestamp 1679585382
transform 1 0 85728 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_894
timestamp 1679585382
transform 1 0 86400 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_901
timestamp 1679585382
transform 1 0 87072 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_908
timestamp 1679585382
transform 1 0 87744 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_915
timestamp 1679585382
transform 1 0 88416 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_922
timestamp 1679585382
transform 1 0 89088 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_929
timestamp 1679585382
transform 1 0 89760 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_936
timestamp 1679585382
transform 1 0 90432 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_943
timestamp 1679585382
transform 1 0 91104 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_950
timestamp 1679585382
transform 1 0 91776 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_957
timestamp 1679585382
transform 1 0 92448 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_964
timestamp 1679585382
transform 1 0 93120 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_971
timestamp 1679585382
transform 1 0 93792 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_978
timestamp 1679585382
transform 1 0 94464 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_985
timestamp 1679585382
transform 1 0 95136 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_992
timestamp 1679585382
transform 1 0 95808 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_999
timestamp 1679585382
transform 1 0 96480 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1006
timestamp 1679585382
transform 1 0 97152 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1013
timestamp 1679585382
transform 1 0 97824 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1020
timestamp 1679585382
transform 1 0 98496 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_1027
timestamp 1677583704
transform 1 0 99168 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_4
timestamp 1679585382
transform 1 0 960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_11
timestamp 1679585382
transform 1 0 1632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_18
timestamp 1679585382
transform 1 0 2304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_25
timestamp 1679585382
transform 1 0 2976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_32
timestamp 1679585382
transform 1 0 3648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_43
timestamp 1679585382
transform 1 0 4704 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_50
timestamp 1679585382
transform 1 0 5376 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_57
timestamp 1679585382
transform 1 0 6048 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_64
timestamp 1679585382
transform 1 0 6720 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_71
timestamp 1679585382
transform 1 0 7392 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_78
timestamp 1679585382
transform 1 0 8064 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_85
timestamp 1679585382
transform 1 0 8736 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_92
timestamp 1679585382
transform 1 0 9408 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_99
timestamp 1679585382
transform 1 0 10080 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_106
timestamp 1679585382
transform 1 0 10752 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_113
timestamp 1679585382
transform 1 0 11424 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_120
timestamp 1679581501
transform 1 0 12096 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_124
timestamp 1677583704
transform 1 0 12480 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_130
timestamp 1679585382
transform 1 0 13056 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_137
timestamp 1679585382
transform 1 0 13728 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_144
timestamp 1679585382
transform 1 0 14400 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_151
timestamp 1679585382
transform 1 0 15072 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_158
timestamp 1679581501
transform 1 0 15744 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_162
timestamp 1677583258
transform 1 0 16128 0 1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_172
timestamp 1679581501
transform 1 0 17088 0 1 3780
box -48 -56 432 834
use sg13g2_decap_8  FILLER_4_190
timestamp 1679585382
transform 1 0 18816 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_197
timestamp 1679585382
transform 1 0 19488 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_204
timestamp 1679585382
transform 1 0 20160 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_211
timestamp 1679585382
transform 1 0 20832 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_218
timestamp 1679585382
transform 1 0 21504 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_225
timestamp 1679585382
transform 1 0 22176 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_268
timestamp 1679585382
transform 1 0 26304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_275
timestamp 1679585382
transform 1 0 26976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_282
timestamp 1679585382
transform 1 0 27648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_289
timestamp 1679585382
transform 1 0 28320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_296
timestamp 1679585382
transform 1 0 28992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_303
timestamp 1679585382
transform 1 0 29664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_310
timestamp 1679581501
transform 1 0 30336 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_314
timestamp 1677583704
transform 1 0 30720 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_325
timestamp 1679585382
transform 1 0 31776 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_332
timestamp 1679585382
transform 1 0 32448 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_339
timestamp 1679585382
transform 1 0 33120 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_346
timestamp 1679585382
transform 1 0 33792 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_353
timestamp 1679585382
transform 1 0 34464 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_360
timestamp 1679585382
transform 1 0 35136 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_367
timestamp 1679585382
transform 1 0 35808 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_374
timestamp 1679585382
transform 1 0 36480 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_381
timestamp 1679585382
transform 1 0 37152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_388
timestamp 1679585382
transform 1 0 37824 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_395
timestamp 1679585382
transform 1 0 38496 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_402
timestamp 1679585382
transform 1 0 39168 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_409
timestamp 1679585382
transform 1 0 39840 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_416
timestamp 1679581501
transform 1 0 40512 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_420
timestamp 1677583258
transform 1 0 40896 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_425
timestamp 1679585382
transform 1 0 41376 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_432
timestamp 1679585382
transform 1 0 42048 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_439
timestamp 1679585382
transform 1 0 42720 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_446
timestamp 1679585382
transform 1 0 43392 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_453
timestamp 1679585382
transform 1 0 44064 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_460
timestamp 1679585382
transform 1 0 44736 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_467
timestamp 1679585382
transform 1 0 45408 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_474
timestamp 1679585382
transform 1 0 46080 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_481
timestamp 1679585382
transform 1 0 46752 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_488
timestamp 1679585382
transform 1 0 47424 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_495
timestamp 1679585382
transform 1 0 48096 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_502
timestamp 1677583704
transform 1 0 48768 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_512
timestamp 1679585382
transform 1 0 49728 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_519
timestamp 1679585382
transform 1 0 50400 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_526
timestamp 1679585382
transform 1 0 51072 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_533
timestamp 1677583258
transform 1 0 51744 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_538
timestamp 1679585382
transform 1 0 52224 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_545
timestamp 1679585382
transform 1 0 52896 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_552
timestamp 1679585382
transform 1 0 53568 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_559
timestamp 1679585382
transform 1 0 54240 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_566
timestamp 1679585382
transform 1 0 54912 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_573
timestamp 1679585382
transform 1 0 55584 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_580
timestamp 1679585382
transform 1 0 56256 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_587
timestamp 1679585382
transform 1 0 56928 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_594
timestamp 1679585382
transform 1 0 57600 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_601
timestamp 1679585382
transform 1 0 58272 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_608
timestamp 1679585382
transform 1 0 58944 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_615
timestamp 1679585382
transform 1 0 59616 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_622
timestamp 1679585382
transform 1 0 60288 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_629
timestamp 1679585382
transform 1 0 60960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_636
timestamp 1679585382
transform 1 0 61632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_643
timestamp 1679585382
transform 1 0 62304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_650
timestamp 1679585382
transform 1 0 62976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_657
timestamp 1679585382
transform 1 0 63648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_664
timestamp 1679585382
transform 1 0 64320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_671
timestamp 1679585382
transform 1 0 64992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_678
timestamp 1679585382
transform 1 0 65664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_685
timestamp 1679585382
transform 1 0 66336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_692
timestamp 1679585382
transform 1 0 67008 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_699
timestamp 1679585382
transform 1 0 67680 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_706
timestamp 1679585382
transform 1 0 68352 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_713
timestamp 1679585382
transform 1 0 69024 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_720
timestamp 1679585382
transform 1 0 69696 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_727
timestamp 1679585382
transform 1 0 70368 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_734
timestamp 1679585382
transform 1 0 71040 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_741
timestamp 1679585382
transform 1 0 71712 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_748
timestamp 1679585382
transform 1 0 72384 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_755
timestamp 1679585382
transform 1 0 73056 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_762
timestamp 1679585382
transform 1 0 73728 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_769
timestamp 1679585382
transform 1 0 74400 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_776
timestamp 1679585382
transform 1 0 75072 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_783
timestamp 1679585382
transform 1 0 75744 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_790
timestamp 1679585382
transform 1 0 76416 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_797
timestamp 1679585382
transform 1 0 77088 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_804
timestamp 1679585382
transform 1 0 77760 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_811
timestamp 1679585382
transform 1 0 78432 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_818
timestamp 1679585382
transform 1 0 79104 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_825
timestamp 1679585382
transform 1 0 79776 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_832
timestamp 1679585382
transform 1 0 80448 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_839
timestamp 1679585382
transform 1 0 81120 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_846
timestamp 1679585382
transform 1 0 81792 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_853
timestamp 1679585382
transform 1 0 82464 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_860
timestamp 1679585382
transform 1 0 83136 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_867
timestamp 1679585382
transform 1 0 83808 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_874
timestamp 1679585382
transform 1 0 84480 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_881
timestamp 1679585382
transform 1 0 85152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_888
timestamp 1679585382
transform 1 0 85824 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_895
timestamp 1679585382
transform 1 0 86496 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_902
timestamp 1679585382
transform 1 0 87168 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_909
timestamp 1679585382
transform 1 0 87840 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_916
timestamp 1679585382
transform 1 0 88512 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_923
timestamp 1679585382
transform 1 0 89184 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_930
timestamp 1679585382
transform 1 0 89856 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_937
timestamp 1679585382
transform 1 0 90528 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_944
timestamp 1679585382
transform 1 0 91200 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_951
timestamp 1679585382
transform 1 0 91872 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_958
timestamp 1679585382
transform 1 0 92544 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_965
timestamp 1679585382
transform 1 0 93216 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_972
timestamp 1679585382
transform 1 0 93888 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_979
timestamp 1679585382
transform 1 0 94560 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_986
timestamp 1679585382
transform 1 0 95232 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_993
timestamp 1679585382
transform 1 0 95904 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1000
timestamp 1679585382
transform 1 0 96576 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1007
timestamp 1679585382
transform 1 0 97248 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1014
timestamp 1679585382
transform 1 0 97920 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1021
timestamp 1679585382
transform 1 0 98592 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_1028
timestamp 1677583258
transform 1 0 99264 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_4
timestamp 1677583704
transform 1 0 960 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_6
timestamp 1677583258
transform 1 0 1152 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_61
timestamp 1679581501
transform 1 0 6432 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_65
timestamp 1677583258
transform 1 0 6816 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_93
timestamp 1679585382
transform 1 0 9504 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_100
timestamp 1679585382
transform 1 0 10176 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_107
timestamp 1679585382
transform 1 0 10848 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_114
timestamp 1679585382
transform 1 0 11520 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_121
timestamp 1679585382
transform 1 0 12192 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_128
timestamp 1679585382
transform 1 0 12864 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_135
timestamp 1679585382
transform 1 0 13536 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_142
timestamp 1679585382
transform 1 0 14208 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_149
timestamp 1679585382
transform 1 0 14880 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_156
timestamp 1679585382
transform 1 0 15552 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_163
timestamp 1679585382
transform 1 0 16224 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_170
timestamp 1679585382
transform 1 0 16896 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_177
timestamp 1679585382
transform 1 0 17568 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_184
timestamp 1679585382
transform 1 0 18240 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_191
timestamp 1679585382
transform 1 0 18912 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_198
timestamp 1679585382
transform 1 0 19584 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_205
timestamp 1679585382
transform 1 0 20256 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_212
timestamp 1679585382
transform 1 0 20928 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_219
timestamp 1679585382
transform 1 0 21600 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_226
timestamp 1679585382
transform 1 0 22272 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_233
timestamp 1679585382
transform 1 0 22944 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_240
timestamp 1679585382
transform 1 0 23616 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_247
timestamp 1679585382
transform 1 0 24288 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_254
timestamp 1679585382
transform 1 0 24960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_261
timestamp 1679585382
transform 1 0 25632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_268
timestamp 1679581501
transform 1 0 26304 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_272
timestamp 1677583258
transform 1 0 26688 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_309
timestamp 1679585382
transform 1 0 30240 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_316
timestamp 1679585382
transform 1 0 30912 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_323
timestamp 1679585382
transform 1 0 31584 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_330
timestamp 1679585382
transform 1 0 32256 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_337
timestamp 1679585382
transform 1 0 32928 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_344
timestamp 1679585382
transform 1 0 33600 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_351
timestamp 1679585382
transform 1 0 34272 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_358
timestamp 1679585382
transform 1 0 34944 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_365
timestamp 1677583704
transform 1 0 35616 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_367
timestamp 1677583258
transform 1 0 35808 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_395
timestamp 1679585382
transform 1 0 38496 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_402
timestamp 1677583704
transform 1 0 39168 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_429
timestamp 1679585382
transform 1 0 41760 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_436
timestamp 1679585382
transform 1 0 42432 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_443
timestamp 1679585382
transform 1 0 43104 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_450
timestamp 1679585382
transform 1 0 43776 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_457
timestamp 1679585382
transform 1 0 44448 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_464
timestamp 1679585382
transform 1 0 45120 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_471
timestamp 1679585382
transform 1 0 45792 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_478
timestamp 1679585382
transform 1 0 46464 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_485
timestamp 1679585382
transform 1 0 47136 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_492
timestamp 1679585382
transform 1 0 47808 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_499
timestamp 1679585382
transform 1 0 48480 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_506
timestamp 1679585382
transform 1 0 49152 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_513
timestamp 1677583704
transform 1 0 49824 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_520
timestamp 1679585382
transform 1 0 50496 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_527
timestamp 1679585382
transform 1 0 51168 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_561
timestamp 1679585382
transform 1 0 54432 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_568
timestamp 1679585382
transform 1 0 55104 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_575
timestamp 1679585382
transform 1 0 55776 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_582
timestamp 1679585382
transform 1 0 56448 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_589
timestamp 1679585382
transform 1 0 57120 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_596
timestamp 1679585382
transform 1 0 57792 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_603
timestamp 1679585382
transform 1 0 58464 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_610
timestamp 1679585382
transform 1 0 59136 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_617
timestamp 1679585382
transform 1 0 59808 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_624
timestamp 1679585382
transform 1 0 60480 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_631
timestamp 1679585382
transform 1 0 61152 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_638
timestamp 1679585382
transform 1 0 61824 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_645
timestamp 1679585382
transform 1 0 62496 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_652
timestamp 1679585382
transform 1 0 63168 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_659
timestamp 1679585382
transform 1 0 63840 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_666
timestamp 1679585382
transform 1 0 64512 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_673
timestamp 1679585382
transform 1 0 65184 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_680
timestamp 1679585382
transform 1 0 65856 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_687
timestamp 1679585382
transform 1 0 66528 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_694
timestamp 1679585382
transform 1 0 67200 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_701
timestamp 1679585382
transform 1 0 67872 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_708
timestamp 1679585382
transform 1 0 68544 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_715
timestamp 1679585382
transform 1 0 69216 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_722
timestamp 1679585382
transform 1 0 69888 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_729
timestamp 1679585382
transform 1 0 70560 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_736
timestamp 1679585382
transform 1 0 71232 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_743
timestamp 1679585382
transform 1 0 71904 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_750
timestamp 1679585382
transform 1 0 72576 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_757
timestamp 1679585382
transform 1 0 73248 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_764
timestamp 1679585382
transform 1 0 73920 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_771
timestamp 1679585382
transform 1 0 74592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_778
timestamp 1679585382
transform 1 0 75264 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_785
timestamp 1679585382
transform 1 0 75936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_792
timestamp 1679585382
transform 1 0 76608 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_799
timestamp 1679585382
transform 1 0 77280 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_806
timestamp 1679585382
transform 1 0 77952 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_813
timestamp 1679585382
transform 1 0 78624 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_820
timestamp 1679585382
transform 1 0 79296 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_827
timestamp 1679585382
transform 1 0 79968 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_834
timestamp 1679585382
transform 1 0 80640 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_841
timestamp 1679585382
transform 1 0 81312 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_848
timestamp 1679585382
transform 1 0 81984 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_855
timestamp 1679585382
transform 1 0 82656 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_862
timestamp 1679585382
transform 1 0 83328 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_869
timestamp 1679585382
transform 1 0 84000 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_876
timestamp 1679585382
transform 1 0 84672 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_883
timestamp 1679585382
transform 1 0 85344 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_890
timestamp 1679585382
transform 1 0 86016 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_897
timestamp 1679585382
transform 1 0 86688 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_904
timestamp 1679585382
transform 1 0 87360 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_911
timestamp 1679585382
transform 1 0 88032 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_918
timestamp 1679585382
transform 1 0 88704 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_925
timestamp 1679585382
transform 1 0 89376 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_932
timestamp 1679585382
transform 1 0 90048 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_939
timestamp 1679585382
transform 1 0 90720 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_946
timestamp 1679585382
transform 1 0 91392 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_953
timestamp 1679585382
transform 1 0 92064 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_960
timestamp 1679585382
transform 1 0 92736 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_967
timestamp 1679585382
transform 1 0 93408 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_974
timestamp 1679585382
transform 1 0 94080 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_981
timestamp 1679585382
transform 1 0 94752 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_988
timestamp 1679585382
transform 1 0 95424 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_995
timestamp 1679585382
transform 1 0 96096 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1002
timestamp 1679585382
transform 1 0 96768 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1009
timestamp 1679585382
transform 1 0 97440 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1016
timestamp 1679585382
transform 1 0 98112 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_1023
timestamp 1679581501
transform 1 0 98784 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_1027
timestamp 1677583704
transform 1 0 99168 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_4
timestamp 1679585382
transform 1 0 960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_11
timestamp 1679581501
transform 1 0 1632 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_28
timestamp 1679585382
transform 1 0 3264 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_35
timestamp 1679581501
transform 1 0 3936 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_39
timestamp 1677583258
transform 1 0 4320 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_44
timestamp 1677583704
transform 1 0 4800 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_60
timestamp 1679585382
transform 1 0 6336 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_67
timestamp 1679585382
transform 1 0 7008 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_74
timestamp 1679585382
transform 1 0 7680 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_81
timestamp 1679585382
transform 1 0 8352 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_88
timestamp 1679585382
transform 1 0 9024 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_131
timestamp 1679585382
transform 1 0 13152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_138
timestamp 1679585382
transform 1 0 13824 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_145
timestamp 1679585382
transform 1 0 14496 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_152
timestamp 1679585382
transform 1 0 15168 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_159
timestamp 1679585382
transform 1 0 15840 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_166
timestamp 1677583258
transform 1 0 16512 0 1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_194
timestamp 1679581501
transform 1 0 19200 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_211
timestamp 1679585382
transform 1 0 20832 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_218
timestamp 1679585382
transform 1 0 21504 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_225
timestamp 1679585382
transform 1 0 22176 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_232
timestamp 1679585382
transform 1 0 22848 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_239
timestamp 1679585382
transform 1 0 23520 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_246
timestamp 1679585382
transform 1 0 24192 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_253
timestamp 1679585382
transform 1 0 24864 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_260
timestamp 1679585382
transform 1 0 25536 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_267
timestamp 1679585382
transform 1 0 26208 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_274
timestamp 1679585382
transform 1 0 26880 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_281
timestamp 1679585382
transform 1 0 27552 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_288
timestamp 1679585382
transform 1 0 28224 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_295
timestamp 1679585382
transform 1 0 28896 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_302
timestamp 1679581501
transform 1 0 29568 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_306
timestamp 1677583704
transform 1 0 29952 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_344
timestamp 1679585382
transform 1 0 33600 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_351
timestamp 1679585382
transform 1 0 34272 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_358
timestamp 1679585382
transform 1 0 34944 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_365
timestamp 1679585382
transform 1 0 35616 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_372
timestamp 1677583704
transform 1 0 36288 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_387
timestamp 1679585382
transform 1 0 37728 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_394
timestamp 1679585382
transform 1 0 38400 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_401
timestamp 1677583704
transform 1 0 39072 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_407
timestamp 1679585382
transform 1 0 39648 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_414
timestamp 1679585382
transform 1 0 40320 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_421
timestamp 1679585382
transform 1 0 40992 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_428
timestamp 1679581501
transform 1 0 41664 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_432
timestamp 1677583258
transform 1 0 42048 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_460
timestamp 1679585382
transform 1 0 44736 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_467
timestamp 1679585382
transform 1 0 45408 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_474
timestamp 1677583704
transform 1 0 46080 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_503
timestamp 1679585382
transform 1 0 48864 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_510
timestamp 1679585382
transform 1 0 49536 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_517
timestamp 1679585382
transform 1 0 50208 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_524
timestamp 1679585382
transform 1 0 50880 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_531
timestamp 1679585382
transform 1 0 51552 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_538
timestamp 1679585382
transform 1 0 52224 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_545
timestamp 1679581501
transform 1 0 52896 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_558
timestamp 1679585382
transform 1 0 54144 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_565
timestamp 1679585382
transform 1 0 54816 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_572
timestamp 1679585382
transform 1 0 55488 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_579
timestamp 1679585382
transform 1 0 56160 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_586
timestamp 1679585382
transform 1 0 56832 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_593
timestamp 1679585382
transform 1 0 57504 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_600
timestamp 1679585382
transform 1 0 58176 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_607
timestamp 1679585382
transform 1 0 58848 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_614
timestamp 1679585382
transform 1 0 59520 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_621
timestamp 1679585382
transform 1 0 60192 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_628
timestamp 1679585382
transform 1 0 60864 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_635
timestamp 1679585382
transform 1 0 61536 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_642
timestamp 1679585382
transform 1 0 62208 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_649
timestamp 1679585382
transform 1 0 62880 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_656
timestamp 1679585382
transform 1 0 63552 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_663
timestamp 1679585382
transform 1 0 64224 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_670
timestamp 1679585382
transform 1 0 64896 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_677
timestamp 1679585382
transform 1 0 65568 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_684
timestamp 1679585382
transform 1 0 66240 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_691
timestamp 1679585382
transform 1 0 66912 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_698
timestamp 1679585382
transform 1 0 67584 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_705
timestamp 1679585382
transform 1 0 68256 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_712
timestamp 1679585382
transform 1 0 68928 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_719
timestamp 1679585382
transform 1 0 69600 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_726
timestamp 1679585382
transform 1 0 70272 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_733
timestamp 1679585382
transform 1 0 70944 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_740
timestamp 1679585382
transform 1 0 71616 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_747
timestamp 1679585382
transform 1 0 72288 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_754
timestamp 1679585382
transform 1 0 72960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_761
timestamp 1679585382
transform 1 0 73632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_768
timestamp 1679585382
transform 1 0 74304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_775
timestamp 1679585382
transform 1 0 74976 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_782
timestamp 1679585382
transform 1 0 75648 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_789
timestamp 1679585382
transform 1 0 76320 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_796
timestamp 1679585382
transform 1 0 76992 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_803
timestamp 1679585382
transform 1 0 77664 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_810
timestamp 1679585382
transform 1 0 78336 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_817
timestamp 1679585382
transform 1 0 79008 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_824
timestamp 1679585382
transform 1 0 79680 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_831
timestamp 1679585382
transform 1 0 80352 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_838
timestamp 1679585382
transform 1 0 81024 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_845
timestamp 1679585382
transform 1 0 81696 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_852
timestamp 1679585382
transform 1 0 82368 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_859
timestamp 1679585382
transform 1 0 83040 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_866
timestamp 1679585382
transform 1 0 83712 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_873
timestamp 1679585382
transform 1 0 84384 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_880
timestamp 1679585382
transform 1 0 85056 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_887
timestamp 1679585382
transform 1 0 85728 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_894
timestamp 1679585382
transform 1 0 86400 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_901
timestamp 1679585382
transform 1 0 87072 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_908
timestamp 1679585382
transform 1 0 87744 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_915
timestamp 1679585382
transform 1 0 88416 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_922
timestamp 1679585382
transform 1 0 89088 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_929
timestamp 1679585382
transform 1 0 89760 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_936
timestamp 1679585382
transform 1 0 90432 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_943
timestamp 1679585382
transform 1 0 91104 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_950
timestamp 1679585382
transform 1 0 91776 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_957
timestamp 1679585382
transform 1 0 92448 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_964
timestamp 1679585382
transform 1 0 93120 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_971
timestamp 1679585382
transform 1 0 93792 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_978
timestamp 1679585382
transform 1 0 94464 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_985
timestamp 1679585382
transform 1 0 95136 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_992
timestamp 1679585382
transform 1 0 95808 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_999
timestamp 1679585382
transform 1 0 96480 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1006
timestamp 1679585382
transform 1 0 97152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1013
timestamp 1679585382
transform 1 0 97824 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1020
timestamp 1679585382
transform 1 0 98496 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_1027
timestamp 1677583704
transform 1 0 99168 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679585382
transform 1 0 576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679585382
transform 1 0 1248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679585382
transform 1 0 1920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_21
timestamp 1679585382
transform 1 0 2592 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_28
timestamp 1679585382
transform 1 0 3264 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_35
timestamp 1679585382
transform 1 0 3936 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_42
timestamp 1679585382
transform 1 0 4608 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_49
timestamp 1679585382
transform 1 0 5280 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_56
timestamp 1679585382
transform 1 0 5952 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_63
timestamp 1679585382
transform 1 0 6624 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_70
timestamp 1679585382
transform 1 0 7296 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_77
timestamp 1679585382
transform 1 0 7968 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_84
timestamp 1679585382
transform 1 0 8640 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_91
timestamp 1677583704
transform 1 0 9312 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_93
timestamp 1677583258
transform 1 0 9504 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_103
timestamp 1679585382
transform 1 0 10464 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_110
timestamp 1679585382
transform 1 0 11136 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_117
timestamp 1677583704
transform 1 0 11808 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_119
timestamp 1677583258
transform 1 0 12000 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_133
timestamp 1679585382
transform 1 0 13344 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_140
timestamp 1679585382
transform 1 0 14016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_147
timestamp 1679585382
transform 1 0 14688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_154
timestamp 1679585382
transform 1 0 15360 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_161
timestamp 1679585382
transform 1 0 16032 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_168
timestamp 1679585382
transform 1 0 16704 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_179
timestamp 1679585382
transform 1 0 17760 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_195
timestamp 1679585382
transform 1 0 19296 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_202
timestamp 1679585382
transform 1 0 19968 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_209
timestamp 1679585382
transform 1 0 20640 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_216
timestamp 1679585382
transform 1 0 21312 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_223
timestamp 1679585382
transform 1 0 21984 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_230
timestamp 1679585382
transform 1 0 22656 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_237
timestamp 1679585382
transform 1 0 23328 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_244
timestamp 1679585382
transform 1 0 24000 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_251
timestamp 1679585382
transform 1 0 24672 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_258
timestamp 1679585382
transform 1 0 25344 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_265
timestamp 1679585382
transform 1 0 26016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_272
timestamp 1679585382
transform 1 0 26688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_279
timestamp 1679585382
transform 1 0 27360 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_286
timestamp 1679585382
transform 1 0 28032 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_293
timestamp 1679585382
transform 1 0 28704 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_300
timestamp 1679585382
transform 1 0 29376 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_307
timestamp 1679585382
transform 1 0 30048 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_314
timestamp 1679585382
transform 1 0 30720 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_321
timestamp 1679585382
transform 1 0 31392 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_328
timestamp 1679585382
transform 1 0 32064 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_335
timestamp 1679585382
transform 1 0 32736 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_364
timestamp 1679585382
transform 1 0 35520 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_371
timestamp 1679585382
transform 1 0 36192 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_378
timestamp 1679585382
transform 1 0 36864 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_385
timestamp 1677583704
transform 1 0 37536 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_387
timestamp 1677583258
transform 1 0 37728 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_415
timestamp 1677583704
transform 1 0 40416 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_422
timestamp 1679585382
transform 1 0 41088 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_429
timestamp 1679585382
transform 1 0 41760 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_436
timestamp 1679585382
transform 1 0 42432 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_443
timestamp 1679585382
transform 1 0 43104 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_450
timestamp 1679585382
transform 1 0 43776 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_457
timestamp 1679585382
transform 1 0 44448 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_464
timestamp 1679585382
transform 1 0 45120 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_471
timestamp 1679581501
transform 1 0 45792 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_475
timestamp 1677583704
transform 1 0 46176 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_485
timestamp 1679585382
transform 1 0 47136 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_492
timestamp 1679585382
transform 1 0 47808 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_499
timestamp 1679585382
transform 1 0 48480 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_506
timestamp 1679585382
transform 1 0 49152 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_513
timestamp 1679585382
transform 1 0 49824 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_520
timestamp 1679585382
transform 1 0 50496 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_527
timestamp 1679585382
transform 1 0 51168 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_534
timestamp 1679585382
transform 1 0 51840 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_541
timestamp 1679585382
transform 1 0 52512 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_548
timestamp 1679585382
transform 1 0 53184 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_555
timestamp 1679585382
transform 1 0 53856 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_562
timestamp 1679585382
transform 1 0 54528 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_569
timestamp 1679585382
transform 1 0 55200 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_576
timestamp 1679585382
transform 1 0 55872 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_583
timestamp 1679585382
transform 1 0 56544 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_590
timestamp 1679585382
transform 1 0 57216 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_597
timestamp 1679585382
transform 1 0 57888 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_604
timestamp 1679585382
transform 1 0 58560 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_611
timestamp 1679585382
transform 1 0 59232 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_618
timestamp 1679585382
transform 1 0 59904 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_625
timestamp 1679585382
transform 1 0 60576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_632
timestamp 1679585382
transform 1 0 61248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_639
timestamp 1679585382
transform 1 0 61920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_646
timestamp 1679585382
transform 1 0 62592 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_653
timestamp 1679585382
transform 1 0 63264 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_660
timestamp 1679585382
transform 1 0 63936 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_667
timestamp 1679585382
transform 1 0 64608 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_674
timestamp 1679585382
transform 1 0 65280 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_681
timestamp 1679585382
transform 1 0 65952 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_688
timestamp 1679585382
transform 1 0 66624 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_695
timestamp 1679585382
transform 1 0 67296 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_702
timestamp 1679585382
transform 1 0 67968 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_709
timestamp 1679585382
transform 1 0 68640 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_716
timestamp 1679585382
transform 1 0 69312 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_723
timestamp 1679585382
transform 1 0 69984 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_730
timestamp 1679585382
transform 1 0 70656 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_737
timestamp 1679585382
transform 1 0 71328 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_744
timestamp 1679585382
transform 1 0 72000 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_751
timestamp 1679585382
transform 1 0 72672 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_758
timestamp 1679585382
transform 1 0 73344 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_765
timestamp 1679585382
transform 1 0 74016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_772
timestamp 1679585382
transform 1 0 74688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_779
timestamp 1679585382
transform 1 0 75360 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_786
timestamp 1679585382
transform 1 0 76032 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_793
timestamp 1679585382
transform 1 0 76704 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_800
timestamp 1679585382
transform 1 0 77376 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_807
timestamp 1679585382
transform 1 0 78048 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_814
timestamp 1679585382
transform 1 0 78720 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_821
timestamp 1679585382
transform 1 0 79392 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_828
timestamp 1679585382
transform 1 0 80064 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_835
timestamp 1679585382
transform 1 0 80736 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_842
timestamp 1679585382
transform 1 0 81408 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_849
timestamp 1679585382
transform 1 0 82080 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_856
timestamp 1679585382
transform 1 0 82752 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_863
timestamp 1679585382
transform 1 0 83424 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_870
timestamp 1679585382
transform 1 0 84096 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_877
timestamp 1679585382
transform 1 0 84768 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_884
timestamp 1679585382
transform 1 0 85440 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_891
timestamp 1679585382
transform 1 0 86112 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_898
timestamp 1679585382
transform 1 0 86784 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_905
timestamp 1679585382
transform 1 0 87456 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_912
timestamp 1679585382
transform 1 0 88128 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_919
timestamp 1679585382
transform 1 0 88800 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_926
timestamp 1679585382
transform 1 0 89472 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_933
timestamp 1679585382
transform 1 0 90144 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_940
timestamp 1679585382
transform 1 0 90816 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_947
timestamp 1679585382
transform 1 0 91488 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_954
timestamp 1679585382
transform 1 0 92160 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_961
timestamp 1679585382
transform 1 0 92832 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_968
timestamp 1679585382
transform 1 0 93504 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_975
timestamp 1679585382
transform 1 0 94176 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_982
timestamp 1679585382
transform 1 0 94848 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_989
timestamp 1679585382
transform 1 0 95520 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_996
timestamp 1679585382
transform 1 0 96192 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1003
timestamp 1679585382
transform 1 0 96864 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1010
timestamp 1679585382
transform 1 0 97536 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_1017
timestamp 1679585382
transform 1 0 98208 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_1024
timestamp 1679581501
transform 1 0 98880 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_1028
timestamp 1677583258
transform 1 0 99264 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_4
timestamp 1679585382
transform 1 0 960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_11
timestamp 1679585382
transform 1 0 1632 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_18
timestamp 1679585382
transform 1 0 2304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_25
timestamp 1679585382
transform 1 0 2976 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_32
timestamp 1679585382
transform 1 0 3648 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_39
timestamp 1679585382
transform 1 0 4320 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_46
timestamp 1679585382
transform 1 0 4992 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_53
timestamp 1679585382
transform 1 0 5664 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_60
timestamp 1679585382
transform 1 0 6336 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_67
timestamp 1679585382
transform 1 0 7008 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_74
timestamp 1679585382
transform 1 0 7680 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_81
timestamp 1679585382
transform 1 0 8352 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_88
timestamp 1679585382
transform 1 0 9024 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_95
timestamp 1679585382
transform 1 0 9696 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_102
timestamp 1679585382
transform 1 0 10368 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_149
timestamp 1679585382
transform 1 0 14880 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_156
timestamp 1679585382
transform 1 0 15552 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_163
timestamp 1679585382
transform 1 0 16224 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_170
timestamp 1679585382
transform 1 0 16896 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_177
timestamp 1679585382
transform 1 0 17568 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_184
timestamp 1679585382
transform 1 0 18240 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_191
timestamp 1679585382
transform 1 0 18912 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_198
timestamp 1679585382
transform 1 0 19584 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_205
timestamp 1679585382
transform 1 0 20256 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_212
timestamp 1679585382
transform 1 0 20928 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_219
timestamp 1679585382
transform 1 0 21600 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_226
timestamp 1679585382
transform 1 0 22272 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_260
timestamp 1679585382
transform 1 0 25536 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_267
timestamp 1679585382
transform 1 0 26208 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_274
timestamp 1679585382
transform 1 0 26880 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_281
timestamp 1679585382
transform 1 0 27552 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_288
timestamp 1679585382
transform 1 0 28224 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_295
timestamp 1679585382
transform 1 0 28896 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_302
timestamp 1679585382
transform 1 0 29568 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_309
timestamp 1679585382
transform 1 0 30240 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_316
timestamp 1679585382
transform 1 0 30912 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_323
timestamp 1679585382
transform 1 0 31584 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_330
timestamp 1679585382
transform 1 0 32256 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_337
timestamp 1677583704
transform 1 0 32928 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_352
timestamp 1679585382
transform 1 0 34368 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_359
timestamp 1679585382
transform 1 0 35040 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_366
timestamp 1679585382
transform 1 0 35712 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_373
timestamp 1679585382
transform 1 0 36384 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_380
timestamp 1679585382
transform 1 0 37056 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_387
timestamp 1679585382
transform 1 0 37728 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_394
timestamp 1677583704
transform 1 0 38400 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_400
timestamp 1679585382
transform 1 0 38976 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_416
timestamp 1679585382
transform 1 0 40512 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_423
timestamp 1679585382
transform 1 0 41184 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_430
timestamp 1679585382
transform 1 0 41856 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_437
timestamp 1679585382
transform 1 0 42528 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_444
timestamp 1679585382
transform 1 0 43200 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_451
timestamp 1679585382
transform 1 0 43872 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_458
timestamp 1679585382
transform 1 0 44544 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_465
timestamp 1679585382
transform 1 0 45216 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_472
timestamp 1679585382
transform 1 0 45888 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_479
timestamp 1679585382
transform 1 0 46560 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_486
timestamp 1679585382
transform 1 0 47232 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_493
timestamp 1679585382
transform 1 0 47904 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_500
timestamp 1677583704
transform 1 0 48576 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_515
timestamp 1677583704
transform 1 0 50016 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_517
timestamp 1677583258
transform 1 0 50208 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_545
timestamp 1679585382
transform 1 0 52896 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_552
timestamp 1679585382
transform 1 0 53568 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_559
timestamp 1679585382
transform 1 0 54240 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_566
timestamp 1679585382
transform 1 0 54912 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_573
timestamp 1679585382
transform 1 0 55584 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_593
timestamp 1679585382
transform 1 0 57504 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_600
timestamp 1679585382
transform 1 0 58176 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_607
timestamp 1679585382
transform 1 0 58848 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_614
timestamp 1679585382
transform 1 0 59520 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_621
timestamp 1679585382
transform 1 0 60192 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_628
timestamp 1679585382
transform 1 0 60864 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_635
timestamp 1679585382
transform 1 0 61536 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_642
timestamp 1679585382
transform 1 0 62208 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_649
timestamp 1679585382
transform 1 0 62880 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_656
timestamp 1679585382
transform 1 0 63552 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_663
timestamp 1679585382
transform 1 0 64224 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_670
timestamp 1679585382
transform 1 0 64896 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_677
timestamp 1679585382
transform 1 0 65568 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_684
timestamp 1679585382
transform 1 0 66240 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_691
timestamp 1679585382
transform 1 0 66912 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_698
timestamp 1679585382
transform 1 0 67584 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_705
timestamp 1679585382
transform 1 0 68256 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_712
timestamp 1679585382
transform 1 0 68928 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_719
timestamp 1679585382
transform 1 0 69600 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_726
timestamp 1679585382
transform 1 0 70272 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_733
timestamp 1679585382
transform 1 0 70944 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_740
timestamp 1679585382
transform 1 0 71616 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_747
timestamp 1679585382
transform 1 0 72288 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_754
timestamp 1679585382
transform 1 0 72960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_761
timestamp 1679585382
transform 1 0 73632 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_768
timestamp 1679585382
transform 1 0 74304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_775
timestamp 1679585382
transform 1 0 74976 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_782
timestamp 1679585382
transform 1 0 75648 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_789
timestamp 1679585382
transform 1 0 76320 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_796
timestamp 1679585382
transform 1 0 76992 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_803
timestamp 1679585382
transform 1 0 77664 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_810
timestamp 1679585382
transform 1 0 78336 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_817
timestamp 1679585382
transform 1 0 79008 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_824
timestamp 1679585382
transform 1 0 79680 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_831
timestamp 1679585382
transform 1 0 80352 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_838
timestamp 1679585382
transform 1 0 81024 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_845
timestamp 1679585382
transform 1 0 81696 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_852
timestamp 1679585382
transform 1 0 82368 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_859
timestamp 1679585382
transform 1 0 83040 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_866
timestamp 1679585382
transform 1 0 83712 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_873
timestamp 1679585382
transform 1 0 84384 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_880
timestamp 1679585382
transform 1 0 85056 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_887
timestamp 1679585382
transform 1 0 85728 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_894
timestamp 1679585382
transform 1 0 86400 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_901
timestamp 1679585382
transform 1 0 87072 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_908
timestamp 1679585382
transform 1 0 87744 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_915
timestamp 1679585382
transform 1 0 88416 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_922
timestamp 1679585382
transform 1 0 89088 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_929
timestamp 1679585382
transform 1 0 89760 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_936
timestamp 1679585382
transform 1 0 90432 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_943
timestamp 1679585382
transform 1 0 91104 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_950
timestamp 1679585382
transform 1 0 91776 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_957
timestamp 1679585382
transform 1 0 92448 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_964
timestamp 1679585382
transform 1 0 93120 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_971
timestamp 1679585382
transform 1 0 93792 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_978
timestamp 1679585382
transform 1 0 94464 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_985
timestamp 1679585382
transform 1 0 95136 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_992
timestamp 1679585382
transform 1 0 95808 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_999
timestamp 1679585382
transform 1 0 96480 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1006
timestamp 1679585382
transform 1 0 97152 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1013
timestamp 1679585382
transform 1 0 97824 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_1020
timestamp 1679585382
transform 1 0 98496 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_1027
timestamp 1677583704
transform 1 0 99168 0 1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_4
timestamp 1679585382
transform 1 0 960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_11
timestamp 1679585382
transform 1 0 1632 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_18
timestamp 1679585382
transform 1 0 2304 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_25
timestamp 1679585382
transform 1 0 2976 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_36
timestamp 1677583704
transform 1 0 4032 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_38
timestamp 1677583258
transform 1 0 4224 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_60
timestamp 1677583704
transform 1 0 6336 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_75
timestamp 1679585382
transform 1 0 7776 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_82
timestamp 1679585382
transform 1 0 8448 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_89
timestamp 1679585382
transform 1 0 9120 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_96
timestamp 1679585382
transform 1 0 9792 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_103
timestamp 1679585382
transform 1 0 10464 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_110
timestamp 1679585382
transform 1 0 11136 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_117
timestamp 1679585382
transform 1 0 11808 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_124
timestamp 1679585382
transform 1 0 12480 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_131
timestamp 1679585382
transform 1 0 13152 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_138
timestamp 1679585382
transform 1 0 13824 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_145
timestamp 1679585382
transform 1 0 14496 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_152
timestamp 1679581501
transform 1 0 15168 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_156
timestamp 1677583704
transform 1 0 15552 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_167
timestamp 1679585382
transform 1 0 16608 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_174
timestamp 1679581501
transform 1 0 17280 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_178
timestamp 1677583704
transform 1 0 17664 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_193
timestamp 1679585382
transform 1 0 19104 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_200
timestamp 1679585382
transform 1 0 19776 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_207
timestamp 1679585382
transform 1 0 20448 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_214
timestamp 1679585382
transform 1 0 21120 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_221
timestamp 1677583258
transform 1 0 21792 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_249
timestamp 1679585382
transform 1 0 24480 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_264
timestamp 1679585382
transform 1 0 25920 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_271
timestamp 1679585382
transform 1 0 26592 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_278
timestamp 1677583704
transform 1 0 27264 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_280
timestamp 1677583258
transform 1 0 27456 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_308
timestamp 1679585382
transform 1 0 30144 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_315
timestamp 1679585382
transform 1 0 30816 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_322
timestamp 1679585382
transform 1 0 31488 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_329
timestamp 1679585382
transform 1 0 32160 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_336
timestamp 1677583704
transform 1 0 32832 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_354
timestamp 1679585382
transform 1 0 34560 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_361
timestamp 1679585382
transform 1 0 35232 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_368
timestamp 1679585382
transform 1 0 35904 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_375
timestamp 1679585382
transform 1 0 36576 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_382
timestamp 1679585382
transform 1 0 37248 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_389
timestamp 1679585382
transform 1 0 37920 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_396
timestamp 1679585382
transform 1 0 38592 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_403
timestamp 1679585382
transform 1 0 39264 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_410
timestamp 1679585382
transform 1 0 39936 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_417
timestamp 1679585382
transform 1 0 40608 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_424
timestamp 1679585382
transform 1 0 41280 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_431
timestamp 1679585382
transform 1 0 41952 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_438
timestamp 1679585382
transform 1 0 42624 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_445
timestamp 1679585382
transform 1 0 43296 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_452
timestamp 1679585382
transform 1 0 43968 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_459
timestamp 1679585382
transform 1 0 44640 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_466
timestamp 1679585382
transform 1 0 45312 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_473
timestamp 1679581501
transform 1 0 45984 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_477
timestamp 1677583258
transform 1 0 46368 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_490
timestamp 1679585382
transform 1 0 47616 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_497
timestamp 1677583704
transform 1 0 48288 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_508
timestamp 1679585382
transform 1 0 49344 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_515
timestamp 1679585382
transform 1 0 50016 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_522
timestamp 1679585382
transform 1 0 50688 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_529
timestamp 1679585382
transform 1 0 51360 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_536
timestamp 1679585382
transform 1 0 52032 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_543
timestamp 1679585382
transform 1 0 52704 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_550
timestamp 1679585382
transform 1 0 53376 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_557
timestamp 1679585382
transform 1 0 54048 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_564
timestamp 1679585382
transform 1 0 54720 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_571
timestamp 1677583258
transform 1 0 55392 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_576
timestamp 1679585382
transform 1 0 55872 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_583
timestamp 1679585382
transform 1 0 56544 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_590
timestamp 1679585382
transform 1 0 57216 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_597
timestamp 1679585382
transform 1 0 57888 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_604
timestamp 1679585382
transform 1 0 58560 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_611
timestamp 1679585382
transform 1 0 59232 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_618
timestamp 1679585382
transform 1 0 59904 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_625
timestamp 1679585382
transform 1 0 60576 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_632
timestamp 1679585382
transform 1 0 61248 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_639
timestamp 1679585382
transform 1 0 61920 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_646
timestamp 1679585382
transform 1 0 62592 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_653
timestamp 1679585382
transform 1 0 63264 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_660
timestamp 1679585382
transform 1 0 63936 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_667
timestamp 1679585382
transform 1 0 64608 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_674
timestamp 1679585382
transform 1 0 65280 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_681
timestamp 1679585382
transform 1 0 65952 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_688
timestamp 1679585382
transform 1 0 66624 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_695
timestamp 1679585382
transform 1 0 67296 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_702
timestamp 1679585382
transform 1 0 67968 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_709
timestamp 1679585382
transform 1 0 68640 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_716
timestamp 1679585382
transform 1 0 69312 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_723
timestamp 1679585382
transform 1 0 69984 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_730
timestamp 1679585382
transform 1 0 70656 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_737
timestamp 1679585382
transform 1 0 71328 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_744
timestamp 1679585382
transform 1 0 72000 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_751
timestamp 1679585382
transform 1 0 72672 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_758
timestamp 1679585382
transform 1 0 73344 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_765
timestamp 1679585382
transform 1 0 74016 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_772
timestamp 1679585382
transform 1 0 74688 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_779
timestamp 1679585382
transform 1 0 75360 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_786
timestamp 1679585382
transform 1 0 76032 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_793
timestamp 1679585382
transform 1 0 76704 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_800
timestamp 1679585382
transform 1 0 77376 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_807
timestamp 1679585382
transform 1 0 78048 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_814
timestamp 1679585382
transform 1 0 78720 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_821
timestamp 1679585382
transform 1 0 79392 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_828
timestamp 1679585382
transform 1 0 80064 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_835
timestamp 1679585382
transform 1 0 80736 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_842
timestamp 1679585382
transform 1 0 81408 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_849
timestamp 1679585382
transform 1 0 82080 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_856
timestamp 1679585382
transform 1 0 82752 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_863
timestamp 1679585382
transform 1 0 83424 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_870
timestamp 1679585382
transform 1 0 84096 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_877
timestamp 1679585382
transform 1 0 84768 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_884
timestamp 1679585382
transform 1 0 85440 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_891
timestamp 1679585382
transform 1 0 86112 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_898
timestamp 1679585382
transform 1 0 86784 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_905
timestamp 1679585382
transform 1 0 87456 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_912
timestamp 1679585382
transform 1 0 88128 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_919
timestamp 1679585382
transform 1 0 88800 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_926
timestamp 1679585382
transform 1 0 89472 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_933
timestamp 1679585382
transform 1 0 90144 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_940
timestamp 1679585382
transform 1 0 90816 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_947
timestamp 1679585382
transform 1 0 91488 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_954
timestamp 1679585382
transform 1 0 92160 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_961
timestamp 1679585382
transform 1 0 92832 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_968
timestamp 1679585382
transform 1 0 93504 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_975
timestamp 1679585382
transform 1 0 94176 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_982
timestamp 1679585382
transform 1 0 94848 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_989
timestamp 1679585382
transform 1 0 95520 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_996
timestamp 1679585382
transform 1 0 96192 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1003
timestamp 1679585382
transform 1 0 96864 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1010
timestamp 1679585382
transform 1 0 97536 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_1017
timestamp 1679585382
transform 1 0 98208 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_1024
timestamp 1679581501
transform 1 0 98880 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_1028
timestamp 1677583258
transform 1 0 99264 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_4
timestamp 1679585382
transform 1 0 960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_11
timestamp 1679585382
transform 1 0 1632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_18
timestamp 1679581501
transform 1 0 2304 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_22
timestamp 1677583704
transform 1 0 2688 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_51
timestamp 1679585382
transform 1 0 5472 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_58
timestamp 1679585382
transform 1 0 6144 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_65
timestamp 1679585382
transform 1 0 6816 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_72
timestamp 1679585382
transform 1 0 7488 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_79
timestamp 1679585382
transform 1 0 8160 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_86
timestamp 1679585382
transform 1 0 8832 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_93
timestamp 1679585382
transform 1 0 9504 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_100
timestamp 1679585382
transform 1 0 10176 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_107
timestamp 1679585382
transform 1 0 10848 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_114
timestamp 1679585382
transform 1 0 11520 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_121
timestamp 1679585382
transform 1 0 12192 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_128
timestamp 1679585382
transform 1 0 12864 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_135
timestamp 1679585382
transform 1 0 13536 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_142
timestamp 1679585382
transform 1 0 14208 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_149
timestamp 1679585382
transform 1 0 14880 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_156
timestamp 1679585382
transform 1 0 15552 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_163
timestamp 1679581501
transform 1 0 16224 0 1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_10_194
timestamp 1679585382
transform 1 0 19200 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_201
timestamp 1679585382
transform 1 0 19872 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_208
timestamp 1679585382
transform 1 0 20544 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_215
timestamp 1679585382
transform 1 0 21216 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_222
timestamp 1679585382
transform 1 0 21888 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_229
timestamp 1679585382
transform 1 0 22560 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_236
timestamp 1677583258
transform 1 0 23232 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_250
timestamp 1679585382
transform 1 0 24576 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_257
timestamp 1679581501
transform 1 0 25248 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_261
timestamp 1677583704
transform 1 0 25632 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_267
timestamp 1679585382
transform 1 0 26208 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_299
timestamp 1677583704
transform 1 0 29280 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_306
timestamp 1679585382
transform 1 0 29952 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_313
timestamp 1679585382
transform 1 0 30624 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_320
timestamp 1677583704
transform 1 0 31296 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_322
timestamp 1677583258
transform 1 0 31488 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_332
timestamp 1679585382
transform 1 0 32448 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_355
timestamp 1679585382
transform 1 0 34656 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_362
timestamp 1679585382
transform 1 0 35328 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_369
timestamp 1679585382
transform 1 0 36000 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_376
timestamp 1679585382
transform 1 0 36672 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_383
timestamp 1677583258
transform 1 0 37344 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_397
timestamp 1679585382
transform 1 0 38688 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_404
timestamp 1679585382
transform 1 0 39360 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_411
timestamp 1679585382
transform 1 0 40032 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_418
timestamp 1679585382
transform 1 0 40704 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_425
timestamp 1679585382
transform 1 0 41376 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_459
timestamp 1679585382
transform 1 0 44640 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_466
timestamp 1677583704
transform 1 0 45312 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_468
timestamp 1677583258
transform 1 0 45504 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_486
timestamp 1679585382
transform 1 0 47232 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_493
timestamp 1679585382
transform 1 0 47904 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_500
timestamp 1679585382
transform 1 0 48576 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_507
timestamp 1679585382
transform 1 0 49248 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_514
timestamp 1679585382
transform 1 0 49920 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_521
timestamp 1679585382
transform 1 0 50592 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_528
timestamp 1679585382
transform 1 0 51264 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_535
timestamp 1679585382
transform 1 0 51936 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_542
timestamp 1679585382
transform 1 0 52608 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_549
timestamp 1679585382
transform 1 0 53280 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_556
timestamp 1677583258
transform 1 0 53952 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_584
timestamp 1677583258
transform 1 0 56640 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_594
timestamp 1679585382
transform 1 0 57600 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_601
timestamp 1679585382
transform 1 0 58272 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_608
timestamp 1679585382
transform 1 0 58944 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_615
timestamp 1679585382
transform 1 0 59616 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_622
timestamp 1679585382
transform 1 0 60288 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_629
timestamp 1679585382
transform 1 0 60960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_636
timestamp 1679585382
transform 1 0 61632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_643
timestamp 1679585382
transform 1 0 62304 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_650
timestamp 1679585382
transform 1 0 62976 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_657
timestamp 1679585382
transform 1 0 63648 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_664
timestamp 1679585382
transform 1 0 64320 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_671
timestamp 1679585382
transform 1 0 64992 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_678
timestamp 1679585382
transform 1 0 65664 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_685
timestamp 1679585382
transform 1 0 66336 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_692
timestamp 1679585382
transform 1 0 67008 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_699
timestamp 1679585382
transform 1 0 67680 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_706
timestamp 1679585382
transform 1 0 68352 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_713
timestamp 1679585382
transform 1 0 69024 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_720
timestamp 1679585382
transform 1 0 69696 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_727
timestamp 1679585382
transform 1 0 70368 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_734
timestamp 1679585382
transform 1 0 71040 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_741
timestamp 1679585382
transform 1 0 71712 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_748
timestamp 1679585382
transform 1 0 72384 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_755
timestamp 1679585382
transform 1 0 73056 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_762
timestamp 1679585382
transform 1 0 73728 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_769
timestamp 1679585382
transform 1 0 74400 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_776
timestamp 1679585382
transform 1 0 75072 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_783
timestamp 1679585382
transform 1 0 75744 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_790
timestamp 1679585382
transform 1 0 76416 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_797
timestamp 1679585382
transform 1 0 77088 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_804
timestamp 1679585382
transform 1 0 77760 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_811
timestamp 1679585382
transform 1 0 78432 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_818
timestamp 1679585382
transform 1 0 79104 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_825
timestamp 1679585382
transform 1 0 79776 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_832
timestamp 1679585382
transform 1 0 80448 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_839
timestamp 1679585382
transform 1 0 81120 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_846
timestamp 1679585382
transform 1 0 81792 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_853
timestamp 1679585382
transform 1 0 82464 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_860
timestamp 1679585382
transform 1 0 83136 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_867
timestamp 1679585382
transform 1 0 83808 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_874
timestamp 1679585382
transform 1 0 84480 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_881
timestamp 1679585382
transform 1 0 85152 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_888
timestamp 1679585382
transform 1 0 85824 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_895
timestamp 1679585382
transform 1 0 86496 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_902
timestamp 1679585382
transform 1 0 87168 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_909
timestamp 1679585382
transform 1 0 87840 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_916
timestamp 1679585382
transform 1 0 88512 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_923
timestamp 1679585382
transform 1 0 89184 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_930
timestamp 1679585382
transform 1 0 89856 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_937
timestamp 1679585382
transform 1 0 90528 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_944
timestamp 1679585382
transform 1 0 91200 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_951
timestamp 1679585382
transform 1 0 91872 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_958
timestamp 1679585382
transform 1 0 92544 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_965
timestamp 1679585382
transform 1 0 93216 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_972
timestamp 1679585382
transform 1 0 93888 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_979
timestamp 1679585382
transform 1 0 94560 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_986
timestamp 1679585382
transform 1 0 95232 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_993
timestamp 1679585382
transform 1 0 95904 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1000
timestamp 1679585382
transform 1 0 96576 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1007
timestamp 1679585382
transform 1 0 97248 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1014
timestamp 1679585382
transform 1 0 97920 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_1021
timestamp 1679585382
transform 1 0 98592 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_1028
timestamp 1677583258
transform 1 0 99264 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_4
timestamp 1679585382
transform 1 0 960 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_11
timestamp 1679581501
transform 1 0 1632 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_15
timestamp 1677583704
transform 1 0 2016 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_44
timestamp 1679585382
transform 1 0 4800 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_51
timestamp 1679585382
transform 1 0 5472 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_58
timestamp 1679581501
transform 1 0 6144 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_62
timestamp 1677583704
transform 1 0 6528 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_91
timestamp 1679585382
transform 1 0 9312 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_98
timestamp 1677583704
transform 1 0 9984 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_100
timestamp 1677583258
transform 1 0 10176 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_128
timestamp 1679585382
transform 1 0 12864 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_135
timestamp 1679585382
transform 1 0 13536 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_142
timestamp 1679585382
transform 1 0 14208 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_149
timestamp 1679585382
transform 1 0 14880 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_156
timestamp 1679585382
transform 1 0 15552 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_163
timestamp 1679585382
transform 1 0 16224 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_170
timestamp 1679585382
transform 1 0 16896 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_177
timestamp 1679585382
transform 1 0 17568 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_184
timestamp 1679585382
transform 1 0 18240 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_191
timestamp 1679585382
transform 1 0 18912 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_198
timestamp 1679585382
transform 1 0 19584 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_214
timestamp 1679585382
transform 1 0 21120 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_230
timestamp 1679585382
transform 1 0 22656 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_237
timestamp 1679585382
transform 1 0 23328 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_244
timestamp 1679585382
transform 1 0 24000 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_251
timestamp 1679585382
transform 1 0 24672 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_258
timestamp 1679585382
transform 1 0 25344 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_265
timestamp 1679585382
transform 1 0 26016 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_272
timestamp 1679585382
transform 1 0 26688 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_279
timestamp 1679585382
transform 1 0 27360 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_286
timestamp 1679585382
transform 1 0 28032 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_293
timestamp 1679585382
transform 1 0 28704 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_300
timestamp 1679585382
transform 1 0 29376 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_307
timestamp 1679585382
transform 1 0 30048 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_314
timestamp 1679585382
transform 1 0 30720 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_321
timestamp 1679585382
transform 1 0 31392 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_328
timestamp 1679585382
transform 1 0 32064 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_335
timestamp 1677583704
transform 1 0 32736 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_351
timestamp 1679585382
transform 1 0 34272 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_358
timestamp 1679585382
transform 1 0 34944 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_374
timestamp 1679581501
transform 1 0 36480 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_378
timestamp 1677583704
transform 1 0 36864 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_407
timestamp 1679585382
transform 1 0 39648 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_414
timestamp 1679585382
transform 1 0 40320 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_421
timestamp 1679585382
transform 1 0 40992 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_428
timestamp 1679585382
transform 1 0 41664 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_435
timestamp 1679585382
transform 1 0 42336 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_442
timestamp 1679585382
transform 1 0 43008 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_449
timestamp 1679585382
transform 1 0 43680 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_456
timestamp 1679585382
transform 1 0 44352 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_463
timestamp 1679585382
transform 1 0 45024 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_470
timestamp 1679581501
transform 1 0 45696 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_474
timestamp 1677583704
transform 1 0 46080 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_521
timestamp 1679585382
transform 1 0 50592 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_528
timestamp 1679585382
transform 1 0 51264 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_535
timestamp 1679581501
transform 1 0 51936 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_539
timestamp 1677583704
transform 1 0 52320 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_554
timestamp 1679585382
transform 1 0 53760 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_561
timestamp 1677583704
transform 1 0 54432 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_567
timestamp 1677583704
transform 1 0 55008 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_596
timestamp 1679585382
transform 1 0 57792 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_603
timestamp 1679585382
transform 1 0 58464 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_641
timestamp 1679585382
transform 1 0 62112 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_648
timestamp 1679585382
transform 1 0 62784 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_655
timestamp 1679585382
transform 1 0 63456 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_662
timestamp 1679585382
transform 1 0 64128 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_669
timestamp 1679585382
transform 1 0 64800 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_676
timestamp 1679585382
transform 1 0 65472 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_683
timestamp 1679585382
transform 1 0 66144 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_690
timestamp 1679585382
transform 1 0 66816 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_697
timestamp 1679585382
transform 1 0 67488 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_704
timestamp 1679585382
transform 1 0 68160 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_711
timestamp 1679585382
transform 1 0 68832 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_718
timestamp 1679585382
transform 1 0 69504 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_725
timestamp 1679585382
transform 1 0 70176 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_732
timestamp 1679585382
transform 1 0 70848 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_739
timestamp 1679585382
transform 1 0 71520 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_746
timestamp 1679585382
transform 1 0 72192 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_753
timestamp 1679585382
transform 1 0 72864 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_760
timestamp 1679585382
transform 1 0 73536 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_767
timestamp 1679585382
transform 1 0 74208 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_774
timestamp 1679585382
transform 1 0 74880 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_781
timestamp 1679585382
transform 1 0 75552 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_788
timestamp 1679585382
transform 1 0 76224 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_795
timestamp 1679585382
transform 1 0 76896 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_802
timestamp 1679585382
transform 1 0 77568 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_809
timestamp 1679585382
transform 1 0 78240 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_816
timestamp 1679585382
transform 1 0 78912 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_823
timestamp 1679585382
transform 1 0 79584 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_830
timestamp 1679585382
transform 1 0 80256 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_837
timestamp 1679585382
transform 1 0 80928 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_844
timestamp 1679585382
transform 1 0 81600 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_851
timestamp 1679585382
transform 1 0 82272 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_858
timestamp 1679585382
transform 1 0 82944 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_865
timestamp 1679585382
transform 1 0 83616 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_872
timestamp 1679585382
transform 1 0 84288 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_879
timestamp 1679585382
transform 1 0 84960 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_886
timestamp 1679585382
transform 1 0 85632 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_893
timestamp 1679585382
transform 1 0 86304 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_900
timestamp 1679585382
transform 1 0 86976 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_907
timestamp 1679585382
transform 1 0 87648 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_914
timestamp 1679585382
transform 1 0 88320 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_921
timestamp 1679585382
transform 1 0 88992 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_928
timestamp 1679585382
transform 1 0 89664 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_935
timestamp 1679585382
transform 1 0 90336 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_942
timestamp 1679585382
transform 1 0 91008 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_949
timestamp 1679585382
transform 1 0 91680 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_956
timestamp 1679585382
transform 1 0 92352 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_963
timestamp 1679585382
transform 1 0 93024 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_970
timestamp 1679585382
transform 1 0 93696 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_977
timestamp 1679585382
transform 1 0 94368 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_984
timestamp 1679585382
transform 1 0 95040 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_991
timestamp 1679585382
transform 1 0 95712 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_998
timestamp 1679585382
transform 1 0 96384 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1005
timestamp 1679585382
transform 1 0 97056 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1012
timestamp 1679585382
transform 1 0 97728 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_1019
timestamp 1679585382
transform 1 0 98400 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_1026
timestamp 1677583704
transform 1 0 99072 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_1028
timestamp 1677583258
transform 1 0 99264 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_4
timestamp 1679585382
transform 1 0 960 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_11
timestamp 1679585382
transform 1 0 1632 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_18
timestamp 1679585382
transform 1 0 2304 0 1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_12_25
timestamp 1677583258
transform 1 0 2976 0 1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_12_30
timestamp 1679581501
transform 1 0 3456 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_34
timestamp 1677583704
transform 1 0 3840 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_45
timestamp 1679585382
transform 1 0 4896 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_52
timestamp 1679585382
transform 1 0 5568 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_59
timestamp 1679585382
transform 1 0 6240 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_66
timestamp 1679585382
transform 1 0 6912 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_73
timestamp 1679585382
transform 1 0 7584 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_80
timestamp 1679585382
transform 1 0 8256 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_87
timestamp 1679585382
transform 1 0 8928 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_94
timestamp 1677583704
transform 1 0 9600 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_105
timestamp 1679585382
transform 1 0 10656 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_112
timestamp 1679585382
transform 1 0 11328 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_119
timestamp 1679581501
transform 1 0 12000 0 1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_12_155
timestamp 1679585382
transform 1 0 15456 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_162
timestamp 1679585382
transform 1 0 16128 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_169
timestamp 1679585382
transform 1 0 16800 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_176
timestamp 1679585382
transform 1 0 17472 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_183
timestamp 1679585382
transform 1 0 18144 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_190
timestamp 1679585382
transform 1 0 18816 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_197
timestamp 1679585382
transform 1 0 19488 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_204
timestamp 1679585382
transform 1 0 20160 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_211
timestamp 1677583704
transform 1 0 20832 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_225
timestamp 1679585382
transform 1 0 22176 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_232
timestamp 1679585382
transform 1 0 22848 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_239
timestamp 1679585382
transform 1 0 23520 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_246
timestamp 1679585382
transform 1 0 24192 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_253
timestamp 1679585382
transform 1 0 24864 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_260
timestamp 1679585382
transform 1 0 25536 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_267
timestamp 1679585382
transform 1 0 26208 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_274
timestamp 1679585382
transform 1 0 26880 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_281
timestamp 1677583704
transform 1 0 27552 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_291
timestamp 1679585382
transform 1 0 28512 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_298
timestamp 1679585382
transform 1 0 29184 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_305
timestamp 1679585382
transform 1 0 29856 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_312
timestamp 1679585382
transform 1 0 30528 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_319
timestamp 1679585382
transform 1 0 31200 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_326
timestamp 1679585382
transform 1 0 31872 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_333
timestamp 1679585382
transform 1 0 32544 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_340
timestamp 1679585382
transform 1 0 33216 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_347
timestamp 1679585382
transform 1 0 33888 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_354
timestamp 1679585382
transform 1 0 34560 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_361
timestamp 1679585382
transform 1 0 35232 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_368
timestamp 1679585382
transform 1 0 35904 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_375
timestamp 1677583704
transform 1 0 36576 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_377
timestamp 1677583258
transform 1 0 36768 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_404
timestamp 1679585382
transform 1 0 39360 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_411
timestamp 1679585382
transform 1 0 40032 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_418
timestamp 1679581501
transform 1 0 40704 0 1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_12_430
timestamp 1679585382
transform 1 0 41856 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_437
timestamp 1679585382
transform 1 0 42528 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_444
timestamp 1679585382
transform 1 0 43200 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_451
timestamp 1679585382
transform 1 0 43872 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_458
timestamp 1679585382
transform 1 0 44544 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_465
timestamp 1679585382
transform 1 0 45216 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_472
timestamp 1679585382
transform 1 0 45888 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_479
timestamp 1677583704
transform 1 0 46560 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_508
timestamp 1679585382
transform 1 0 49344 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_515
timestamp 1679585382
transform 1 0 50016 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_522
timestamp 1679585382
transform 1 0 50688 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_529
timestamp 1679585382
transform 1 0 51360 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_536
timestamp 1679585382
transform 1 0 52032 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_543
timestamp 1679585382
transform 1 0 52704 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_550
timestamp 1679585382
transform 1 0 53376 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_557
timestamp 1679585382
transform 1 0 54048 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_564
timestamp 1679581501
transform 1 0 54720 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_573
timestamp 1677583704
transform 1 0 55584 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_584
timestamp 1679585382
transform 1 0 56640 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_591
timestamp 1679585382
transform 1 0 57312 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_598
timestamp 1679581501
transform 1 0 57984 0 1 9828
box -48 -56 432 834
use sg13g2_decap_4  FILLER_12_610
timestamp 1679581501
transform 1 0 59136 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_614
timestamp 1677583704
transform 1 0 59520 0 1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_12_620
timestamp 1679581501
transform 1 0 60096 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_624
timestamp 1677583704
transform 1 0 60480 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_635
timestamp 1679585382
transform 1 0 61536 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_642
timestamp 1679585382
transform 1 0 62208 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_649
timestamp 1679585382
transform 1 0 62880 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_656
timestamp 1679585382
transform 1 0 63552 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_663
timestamp 1679585382
transform 1 0 64224 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_670
timestamp 1679585382
transform 1 0 64896 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_677
timestamp 1679585382
transform 1 0 65568 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_684
timestamp 1679585382
transform 1 0 66240 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_691
timestamp 1679585382
transform 1 0 66912 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_698
timestamp 1679585382
transform 1 0 67584 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_705
timestamp 1679585382
transform 1 0 68256 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_712
timestamp 1679585382
transform 1 0 68928 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_719
timestamp 1679585382
transform 1 0 69600 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_726
timestamp 1679585382
transform 1 0 70272 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_733
timestamp 1679585382
transform 1 0 70944 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_740
timestamp 1679585382
transform 1 0 71616 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_747
timestamp 1679585382
transform 1 0 72288 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_754
timestamp 1679585382
transform 1 0 72960 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_761
timestamp 1679585382
transform 1 0 73632 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_768
timestamp 1679585382
transform 1 0 74304 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_775
timestamp 1679585382
transform 1 0 74976 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_782
timestamp 1679585382
transform 1 0 75648 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_789
timestamp 1679585382
transform 1 0 76320 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_796
timestamp 1679585382
transform 1 0 76992 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_803
timestamp 1679585382
transform 1 0 77664 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_810
timestamp 1679585382
transform 1 0 78336 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_817
timestamp 1679585382
transform 1 0 79008 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_824
timestamp 1679585382
transform 1 0 79680 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_831
timestamp 1679585382
transform 1 0 80352 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_838
timestamp 1679585382
transform 1 0 81024 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_845
timestamp 1679585382
transform 1 0 81696 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_852
timestamp 1679585382
transform 1 0 82368 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_859
timestamp 1679585382
transform 1 0 83040 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_866
timestamp 1679585382
transform 1 0 83712 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_873
timestamp 1679585382
transform 1 0 84384 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_880
timestamp 1679585382
transform 1 0 85056 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_887
timestamp 1679585382
transform 1 0 85728 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_894
timestamp 1679585382
transform 1 0 86400 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_901
timestamp 1679585382
transform 1 0 87072 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_908
timestamp 1679585382
transform 1 0 87744 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_915
timestamp 1679585382
transform 1 0 88416 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_922
timestamp 1679585382
transform 1 0 89088 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_929
timestamp 1679585382
transform 1 0 89760 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_936
timestamp 1679585382
transform 1 0 90432 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_943
timestamp 1679585382
transform 1 0 91104 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_950
timestamp 1679585382
transform 1 0 91776 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_957
timestamp 1679585382
transform 1 0 92448 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_964
timestamp 1679585382
transform 1 0 93120 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_971
timestamp 1679585382
transform 1 0 93792 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_978
timestamp 1679585382
transform 1 0 94464 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_985
timestamp 1679585382
transform 1 0 95136 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_992
timestamp 1679585382
transform 1 0 95808 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_999
timestamp 1679585382
transform 1 0 96480 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1006
timestamp 1679585382
transform 1 0 97152 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1013
timestamp 1679585382
transform 1 0 97824 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_1020
timestamp 1679585382
transform 1 0 98496 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_1027
timestamp 1677583704
transform 1 0 99168 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_4
timestamp 1679585382
transform 1 0 960 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_11
timestamp 1679585382
transform 1 0 1632 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_18
timestamp 1679585382
transform 1 0 2304 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_25
timestamp 1679585382
transform 1 0 2976 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_32
timestamp 1679585382
transform 1 0 3648 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_39
timestamp 1679585382
transform 1 0 4320 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_46
timestamp 1679585382
transform 1 0 4992 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_53
timestamp 1679585382
transform 1 0 5664 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_60
timestamp 1679585382
transform 1 0 6336 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_67
timestamp 1679585382
transform 1 0 7008 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_74
timestamp 1679585382
transform 1 0 7680 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_81
timestamp 1679585382
transform 1 0 8352 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_88
timestamp 1677583704
transform 1 0 9024 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_103
timestamp 1679585382
transform 1 0 10464 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_110
timestamp 1679585382
transform 1 0 11136 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_117
timestamp 1679585382
transform 1 0 11808 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_124
timestamp 1679581501
transform 1 0 12480 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_13_137
timestamp 1679585382
transform 1 0 13728 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_144
timestamp 1679585382
transform 1 0 14400 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_151
timestamp 1677583704
transform 1 0 15072 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_153
timestamp 1677583258
transform 1 0 15264 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_190
timestamp 1679585382
transform 1 0 18816 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_197
timestamp 1679585382
transform 1 0 19488 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_204
timestamp 1679581501
transform 1 0 20160 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_208
timestamp 1677583258
transform 1 0 20544 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_222
timestamp 1679585382
transform 1 0 21888 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_229
timestamp 1679585382
transform 1 0 22560 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_236
timestamp 1679585382
transform 1 0 23232 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_243
timestamp 1679581501
transform 1 0 23904 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_247
timestamp 1677583258
transform 1 0 24288 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_275
timestamp 1679585382
transform 1 0 26976 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_282
timestamp 1679585382
transform 1 0 27648 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_289
timestamp 1679585382
transform 1 0 28320 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_296
timestamp 1679585382
transform 1 0 28992 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_303
timestamp 1679585382
transform 1 0 29664 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_310
timestamp 1679581501
transform 1 0 30336 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_4  FILLER_13_322
timestamp 1679581501
transform 1 0 31488 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_13_331
timestamp 1679585382
transform 1 0 32352 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_347
timestamp 1679585382
transform 1 0 33888 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_354
timestamp 1679585382
transform 1 0 34560 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_361
timestamp 1679581501
transform 1 0 35232 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_365
timestamp 1677583258
transform 1 0 35616 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_394
timestamp 1679585382
transform 1 0 38400 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_401
timestamp 1679585382
transform 1 0 39072 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_408
timestamp 1679585382
transform 1 0 39744 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_424
timestamp 1679581501
transform 1 0 41280 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_13_428
timestamp 1677583704
transform 1 0 41664 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_457
timestamp 1679585382
transform 1 0 44448 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_464
timestamp 1679585382
transform 1 0 45120 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_471
timestamp 1679585382
transform 1 0 45792 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_478
timestamp 1679585382
transform 1 0 46464 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_485
timestamp 1679585382
transform 1 0 47136 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_492
timestamp 1679585382
transform 1 0 47808 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_499
timestamp 1679585382
transform 1 0 48480 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_506
timestamp 1679585382
transform 1 0 49152 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_513
timestamp 1679585382
transform 1 0 49824 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_520
timestamp 1679585382
transform 1 0 50496 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_527
timestamp 1679581501
transform 1 0 51168 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_13_544
timestamp 1679585382
transform 1 0 52800 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_551
timestamp 1679585382
transform 1 0 53472 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_558
timestamp 1679585382
transform 1 0 54144 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_565
timestamp 1679585382
transform 1 0 54816 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_572
timestamp 1679585382
transform 1 0 55488 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_579
timestamp 1679585382
transform 1 0 56160 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_586
timestamp 1679585382
transform 1 0 56832 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_593
timestamp 1679585382
transform 1 0 57504 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_600
timestamp 1679581501
transform 1 0 58176 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_604
timestamp 1677583258
transform 1 0 58560 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_613
timestamp 1677583258
transform 1 0 59424 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_641
timestamp 1679585382
transform 1 0 62112 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_648
timestamp 1679585382
transform 1 0 62784 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_655
timestamp 1679585382
transform 1 0 63456 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_662
timestamp 1679585382
transform 1 0 64128 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_669
timestamp 1679585382
transform 1 0 64800 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_676
timestamp 1679585382
transform 1 0 65472 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_683
timestamp 1679585382
transform 1 0 66144 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_690
timestamp 1679585382
transform 1 0 66816 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_697
timestamp 1679585382
transform 1 0 67488 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_704
timestamp 1679585382
transform 1 0 68160 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_711
timestamp 1679585382
transform 1 0 68832 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_718
timestamp 1679585382
transform 1 0 69504 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_725
timestamp 1679585382
transform 1 0 70176 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_732
timestamp 1679585382
transform 1 0 70848 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_739
timestamp 1679585382
transform 1 0 71520 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_746
timestamp 1679585382
transform 1 0 72192 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_753
timestamp 1679585382
transform 1 0 72864 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_760
timestamp 1679585382
transform 1 0 73536 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_767
timestamp 1679585382
transform 1 0 74208 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_774
timestamp 1679585382
transform 1 0 74880 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_781
timestamp 1679585382
transform 1 0 75552 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_788
timestamp 1679585382
transform 1 0 76224 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_795
timestamp 1679585382
transform 1 0 76896 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_802
timestamp 1679585382
transform 1 0 77568 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_809
timestamp 1679585382
transform 1 0 78240 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_816
timestamp 1679585382
transform 1 0 78912 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_823
timestamp 1679585382
transform 1 0 79584 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_830
timestamp 1679585382
transform 1 0 80256 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_837
timestamp 1679585382
transform 1 0 80928 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_844
timestamp 1679585382
transform 1 0 81600 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_851
timestamp 1679585382
transform 1 0 82272 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_858
timestamp 1679585382
transform 1 0 82944 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_865
timestamp 1679585382
transform 1 0 83616 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_872
timestamp 1679585382
transform 1 0 84288 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_879
timestamp 1679585382
transform 1 0 84960 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_886
timestamp 1679585382
transform 1 0 85632 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_893
timestamp 1679585382
transform 1 0 86304 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_900
timestamp 1679585382
transform 1 0 86976 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_907
timestamp 1679585382
transform 1 0 87648 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_914
timestamp 1679585382
transform 1 0 88320 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_921
timestamp 1679585382
transform 1 0 88992 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_928
timestamp 1679585382
transform 1 0 89664 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_935
timestamp 1679585382
transform 1 0 90336 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_942
timestamp 1679585382
transform 1 0 91008 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_949
timestamp 1679585382
transform 1 0 91680 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_956
timestamp 1679585382
transform 1 0 92352 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_963
timestamp 1679585382
transform 1 0 93024 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_970
timestamp 1679585382
transform 1 0 93696 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_977
timestamp 1679585382
transform 1 0 94368 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_984
timestamp 1679585382
transform 1 0 95040 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_991
timestamp 1679585382
transform 1 0 95712 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_998
timestamp 1679585382
transform 1 0 96384 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1005
timestamp 1679585382
transform 1 0 97056 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1012
timestamp 1679585382
transform 1 0 97728 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_1019
timestamp 1679585382
transform 1 0 98400 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_1026
timestamp 1677583704
transform 1 0 99072 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_1028
timestamp 1677583258
transform 1 0 99264 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_4
timestamp 1679585382
transform 1 0 960 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_11
timestamp 1679585382
transform 1 0 1632 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_18
timestamp 1679585382
transform 1 0 2304 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_25
timestamp 1679585382
transform 1 0 2976 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_32
timestamp 1679585382
transform 1 0 3648 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_39
timestamp 1679585382
transform 1 0 4320 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_46
timestamp 1679585382
transform 1 0 4992 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_53
timestamp 1679585382
transform 1 0 5664 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_60
timestamp 1679585382
transform 1 0 6336 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_67
timestamp 1679585382
transform 1 0 7008 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_74
timestamp 1679585382
transform 1 0 7680 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_81
timestamp 1679585382
transform 1 0 8352 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_88
timestamp 1679585382
transform 1 0 9024 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_95
timestamp 1679585382
transform 1 0 9696 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_102
timestamp 1679585382
transform 1 0 10368 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_109
timestamp 1679585382
transform 1 0 11040 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_116
timestamp 1679585382
transform 1 0 11712 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_123
timestamp 1679585382
transform 1 0 12384 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_130
timestamp 1679585382
transform 1 0 13056 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_137
timestamp 1679585382
transform 1 0 13728 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_144
timestamp 1679585382
transform 1 0 14400 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_151
timestamp 1679585382
transform 1 0 15072 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_158
timestamp 1679585382
transform 1 0 15744 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_165
timestamp 1679585382
transform 1 0 16416 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_172
timestamp 1679585382
transform 1 0 17088 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_179
timestamp 1677583704
transform 1 0 17760 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_181
timestamp 1677583258
transform 1 0 17952 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_195
timestamp 1679585382
transform 1 0 19296 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_202
timestamp 1679585382
transform 1 0 19968 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_209
timestamp 1679585382
transform 1 0 20640 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_216
timestamp 1679585382
transform 1 0 21312 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_223
timestamp 1679585382
transform 1 0 21984 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_230
timestamp 1679581501
transform 1 0 22656 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_242
timestamp 1677583704
transform 1 0 23808 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_244
timestamp 1677583258
transform 1 0 24000 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_254
timestamp 1679585382
transform 1 0 24960 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_261
timestamp 1679585382
transform 1 0 25632 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_268
timestamp 1679585382
transform 1 0 26304 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_275
timestamp 1679585382
transform 1 0 26976 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_282
timestamp 1679585382
transform 1 0 27648 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_289
timestamp 1679585382
transform 1 0 28320 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_296
timestamp 1679585382
transform 1 0 28992 0 1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_14_303
timestamp 1677583258
transform 1 0 29664 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_336
timestamp 1679585382
transform 1 0 32832 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_343
timestamp 1679585382
transform 1 0 33504 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_350
timestamp 1679585382
transform 1 0 34176 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_357
timestamp 1679585382
transform 1 0 34848 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_364
timestamp 1679585382
transform 1 0 35520 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_371
timestamp 1679585382
transform 1 0 36192 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_378
timestamp 1679585382
transform 1 0 36864 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_385
timestamp 1679585382
transform 1 0 37536 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_392
timestamp 1679585382
transform 1 0 38208 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_399
timestamp 1679585382
transform 1 0 38880 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_406
timestamp 1679585382
transform 1 0 39552 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_413
timestamp 1679581501
transform 1 0 40224 0 1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_14_447
timestamp 1679585382
transform 1 0 43488 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_454
timestamp 1679585382
transform 1 0 44160 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_461
timestamp 1679585382
transform 1 0 44832 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_468
timestamp 1679585382
transform 1 0 45504 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_475
timestamp 1679581501
transform 1 0 46176 0 1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_14_488
timestamp 1679585382
transform 1 0 47424 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_495
timestamp 1679581501
transform 1 0 48096 0 1 11340
box -48 -56 432 834
use sg13g2_fill_2  FILLER_14_499
timestamp 1677583704
transform 1 0 48480 0 1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_518
timestamp 1679585382
transform 1 0 50304 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_525
timestamp 1679585382
transform 1 0 50976 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_532
timestamp 1679585382
transform 1 0 51648 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_539
timestamp 1679585382
transform 1 0 52320 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_546
timestamp 1679581501
transform 1 0 52992 0 1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_14_563
timestamp 1679585382
transform 1 0 54624 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_570
timestamp 1679585382
transform 1 0 55296 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_577
timestamp 1679585382
transform 1 0 55968 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_584
timestamp 1679585382
transform 1 0 56640 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_591
timestamp 1679585382
transform 1 0 57312 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_598
timestamp 1679585382
transform 1 0 57984 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_605
timestamp 1679585382
transform 1 0 58656 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_612
timestamp 1679585382
transform 1 0 59328 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_619
timestamp 1679585382
transform 1 0 60000 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_626
timestamp 1679581501
transform 1 0 60672 0 1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_14_639
timestamp 1679585382
transform 1 0 61920 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_646
timestamp 1679585382
transform 1 0 62592 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_653
timestamp 1679585382
transform 1 0 63264 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_660
timestamp 1679585382
transform 1 0 63936 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_667
timestamp 1679585382
transform 1 0 64608 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_674
timestamp 1679585382
transform 1 0 65280 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_681
timestamp 1679585382
transform 1 0 65952 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_688
timestamp 1679585382
transform 1 0 66624 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_695
timestamp 1679585382
transform 1 0 67296 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_702
timestamp 1679585382
transform 1 0 67968 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_709
timestamp 1679585382
transform 1 0 68640 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_716
timestamp 1679585382
transform 1 0 69312 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_723
timestamp 1679585382
transform 1 0 69984 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_730
timestamp 1679585382
transform 1 0 70656 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_737
timestamp 1679585382
transform 1 0 71328 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_744
timestamp 1679585382
transform 1 0 72000 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_751
timestamp 1679585382
transform 1 0 72672 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_758
timestamp 1679585382
transform 1 0 73344 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_765
timestamp 1679585382
transform 1 0 74016 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_772
timestamp 1679585382
transform 1 0 74688 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_779
timestamp 1679585382
transform 1 0 75360 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_786
timestamp 1679585382
transform 1 0 76032 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_793
timestamp 1679585382
transform 1 0 76704 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_800
timestamp 1679585382
transform 1 0 77376 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_807
timestamp 1679585382
transform 1 0 78048 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_814
timestamp 1679585382
transform 1 0 78720 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_821
timestamp 1679585382
transform 1 0 79392 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_828
timestamp 1679585382
transform 1 0 80064 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_835
timestamp 1679585382
transform 1 0 80736 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_842
timestamp 1679585382
transform 1 0 81408 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_849
timestamp 1679585382
transform 1 0 82080 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_856
timestamp 1679585382
transform 1 0 82752 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_863
timestamp 1679585382
transform 1 0 83424 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_870
timestamp 1679585382
transform 1 0 84096 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_877
timestamp 1679585382
transform 1 0 84768 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_884
timestamp 1679585382
transform 1 0 85440 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_891
timestamp 1679585382
transform 1 0 86112 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_898
timestamp 1679585382
transform 1 0 86784 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_905
timestamp 1679585382
transform 1 0 87456 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_912
timestamp 1679585382
transform 1 0 88128 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_919
timestamp 1679585382
transform 1 0 88800 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_926
timestamp 1679585382
transform 1 0 89472 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_933
timestamp 1679585382
transform 1 0 90144 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_940
timestamp 1679585382
transform 1 0 90816 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_947
timestamp 1679585382
transform 1 0 91488 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_954
timestamp 1679585382
transform 1 0 92160 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_961
timestamp 1679585382
transform 1 0 92832 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_968
timestamp 1679585382
transform 1 0 93504 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_975
timestamp 1679585382
transform 1 0 94176 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_982
timestamp 1679585382
transform 1 0 94848 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_989
timestamp 1679585382
transform 1 0 95520 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_996
timestamp 1679585382
transform 1 0 96192 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1003
timestamp 1679585382
transform 1 0 96864 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1010
timestamp 1679585382
transform 1 0 97536 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_1017
timestamp 1679585382
transform 1 0 98208 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_1024
timestamp 1679581501
transform 1 0 98880 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_1028
timestamp 1677583258
transform 1 0 99264 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_4
timestamp 1679585382
transform 1 0 960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_11
timestamp 1679585382
transform 1 0 1632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_18
timestamp 1679585382
transform 1 0 2304 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_25
timestamp 1679585382
transform 1 0 2976 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_32
timestamp 1679585382
transform 1 0 3648 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_39
timestamp 1679585382
transform 1 0 4320 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_46
timestamp 1679585382
transform 1 0 4992 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_53
timestamp 1679585382
transform 1 0 5664 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_60
timestamp 1679585382
transform 1 0 6336 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_67
timestamp 1679585382
transform 1 0 7008 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_74
timestamp 1679585382
transform 1 0 7680 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_81
timestamp 1677583258
transform 1 0 8352 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_95
timestamp 1679585382
transform 1 0 9696 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_102
timestamp 1679585382
transform 1 0 10368 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_109
timestamp 1679585382
transform 1 0 11040 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_116
timestamp 1679585382
transform 1 0 11712 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_123
timestamp 1679585382
transform 1 0 12384 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_130
timestamp 1679585382
transform 1 0 13056 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_137
timestamp 1679585382
transform 1 0 13728 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_144
timestamp 1679585382
transform 1 0 14400 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_151
timestamp 1679585382
transform 1 0 15072 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_158
timestamp 1679585382
transform 1 0 15744 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_165
timestamp 1679585382
transform 1 0 16416 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_172
timestamp 1679585382
transform 1 0 17088 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_179
timestamp 1679585382
transform 1 0 17760 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_199
timestamp 1679585382
transform 1 0 19680 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_206
timestamp 1679585382
transform 1 0 20352 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_213
timestamp 1677583258
transform 1 0 21024 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_227
timestamp 1677583704
transform 1 0 22368 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_229
timestamp 1677583258
transform 1 0 22560 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_247
timestamp 1679585382
transform 1 0 24288 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_254
timestamp 1679585382
transform 1 0 24960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_261
timestamp 1679585382
transform 1 0 25632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_268
timestamp 1679585382
transform 1 0 26304 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_275
timestamp 1679585382
transform 1 0 26976 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_282
timestamp 1679581501
transform 1 0 27648 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_286
timestamp 1677583704
transform 1 0 28032 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_328
timestamp 1679585382
transform 1 0 32064 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_335
timestamp 1679585382
transform 1 0 32736 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_342
timestamp 1679585382
transform 1 0 33408 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_349
timestamp 1679585382
transform 1 0 34080 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_356
timestamp 1677583258
transform 1 0 34752 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_370
timestamp 1679585382
transform 1 0 36096 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_377
timestamp 1679585382
transform 1 0 36768 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_384
timestamp 1679585382
transform 1 0 37440 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_391
timestamp 1679585382
transform 1 0 38112 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_398
timestamp 1679585382
transform 1 0 38784 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_405
timestamp 1679585382
transform 1 0 39456 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_412
timestamp 1679585382
transform 1 0 40128 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_419
timestamp 1677583704
transform 1 0 40800 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_421
timestamp 1677583258
transform 1 0 40992 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_426
timestamp 1677583704
transform 1 0 41472 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_441
timestamp 1679585382
transform 1 0 42912 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_448
timestamp 1679585382
transform 1 0 43584 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_455
timestamp 1679585382
transform 1 0 44256 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_462
timestamp 1679585382
transform 1 0 44928 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_469
timestamp 1679585382
transform 1 0 45600 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_476
timestamp 1679585382
transform 1 0 46272 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_483
timestamp 1679585382
transform 1 0 46944 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_490
timestamp 1679585382
transform 1 0 47616 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_497
timestamp 1679585382
transform 1 0 48288 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_504
timestamp 1677583704
transform 1 0 48960 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_506
timestamp 1677583258
transform 1 0 49152 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_511
timestamp 1679585382
transform 1 0 49632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_526
timestamp 1679585382
transform 1 0 51072 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_533
timestamp 1679585382
transform 1 0 51744 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_540
timestamp 1679581501
transform 1 0 52416 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_544
timestamp 1677583704
transform 1 0 52800 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_559
timestamp 1677583258
transform 1 0 54240 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_587
timestamp 1679585382
transform 1 0 56928 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_594
timestamp 1679585382
transform 1 0 57600 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_601
timestamp 1679585382
transform 1 0 58272 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_608
timestamp 1679585382
transform 1 0 58944 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_615
timestamp 1679585382
transform 1 0 59616 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_622
timestamp 1679585382
transform 1 0 60288 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_629
timestamp 1679585382
transform 1 0 60960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_636
timestamp 1679585382
transform 1 0 61632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_643
timestamp 1679585382
transform 1 0 62304 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_650
timestamp 1679585382
transform 1 0 62976 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_657
timestamp 1679585382
transform 1 0 63648 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_664
timestamp 1679585382
transform 1 0 64320 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_671
timestamp 1679585382
transform 1 0 64992 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_678
timestamp 1679585382
transform 1 0 65664 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_685
timestamp 1679585382
transform 1 0 66336 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_692
timestamp 1679585382
transform 1 0 67008 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_699
timestamp 1679585382
transform 1 0 67680 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_706
timestamp 1679585382
transform 1 0 68352 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_713
timestamp 1679585382
transform 1 0 69024 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_720
timestamp 1679585382
transform 1 0 69696 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_727
timestamp 1679585382
transform 1 0 70368 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_734
timestamp 1679585382
transform 1 0 71040 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_741
timestamp 1679585382
transform 1 0 71712 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_748
timestamp 1679585382
transform 1 0 72384 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_755
timestamp 1679585382
transform 1 0 73056 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_762
timestamp 1679585382
transform 1 0 73728 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_769
timestamp 1679585382
transform 1 0 74400 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_776
timestamp 1679585382
transform 1 0 75072 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_783
timestamp 1679585382
transform 1 0 75744 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_790
timestamp 1679585382
transform 1 0 76416 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_797
timestamp 1679585382
transform 1 0 77088 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_804
timestamp 1679585382
transform 1 0 77760 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_811
timestamp 1679585382
transform 1 0 78432 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_818
timestamp 1679585382
transform 1 0 79104 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_825
timestamp 1679585382
transform 1 0 79776 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_832
timestamp 1679585382
transform 1 0 80448 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_839
timestamp 1679585382
transform 1 0 81120 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_846
timestamp 1679585382
transform 1 0 81792 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_853
timestamp 1679585382
transform 1 0 82464 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_860
timestamp 1679585382
transform 1 0 83136 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_867
timestamp 1679585382
transform 1 0 83808 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_874
timestamp 1679585382
transform 1 0 84480 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_881
timestamp 1679585382
transform 1 0 85152 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_888
timestamp 1679585382
transform 1 0 85824 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_895
timestamp 1679585382
transform 1 0 86496 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_902
timestamp 1679585382
transform 1 0 87168 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_909
timestamp 1679585382
transform 1 0 87840 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_916
timestamp 1679585382
transform 1 0 88512 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_923
timestamp 1679585382
transform 1 0 89184 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_930
timestamp 1679585382
transform 1 0 89856 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_937
timestamp 1679585382
transform 1 0 90528 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_944
timestamp 1679585382
transform 1 0 91200 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_951
timestamp 1679585382
transform 1 0 91872 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_958
timestamp 1679585382
transform 1 0 92544 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_965
timestamp 1679585382
transform 1 0 93216 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_972
timestamp 1679585382
transform 1 0 93888 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_979
timestamp 1679585382
transform 1 0 94560 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_986
timestamp 1679585382
transform 1 0 95232 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_993
timestamp 1679585382
transform 1 0 95904 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1000
timestamp 1679585382
transform 1 0 96576 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1007
timestamp 1679585382
transform 1 0 97248 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1014
timestamp 1679585382
transform 1 0 97920 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_1021
timestamp 1679585382
transform 1 0 98592 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_1028
timestamp 1677583258
transform 1 0 99264 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_4
timestamp 1679585382
transform 1 0 960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_11
timestamp 1679585382
transform 1 0 1632 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_18
timestamp 1679585382
transform 1 0 2304 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_25
timestamp 1679585382
transform 1 0 2976 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_32
timestamp 1677583704
transform 1 0 3648 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_34
timestamp 1677583258
transform 1 0 3840 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_62
timestamp 1679585382
transform 1 0 6528 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_69
timestamp 1679585382
transform 1 0 7200 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_76
timestamp 1679585382
transform 1 0 7872 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_83
timestamp 1679581501
transform 1 0 8544 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_87
timestamp 1677583258
transform 1 0 8928 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_123
timestamp 1679585382
transform 1 0 12384 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_130
timestamp 1679585382
transform 1 0 13056 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_137
timestamp 1679585382
transform 1 0 13728 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_144
timestamp 1679585382
transform 1 0 14400 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_151
timestamp 1679585382
transform 1 0 15072 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_158
timestamp 1679585382
transform 1 0 15744 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_165
timestamp 1679581501
transform 1 0 16416 0 1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_16_196
timestamp 1679585382
transform 1 0 19392 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_203
timestamp 1679585382
transform 1 0 20064 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_210
timestamp 1679585382
transform 1 0 20736 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_217
timestamp 1679585382
transform 1 0 21408 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_224
timestamp 1679585382
transform 1 0 22080 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_231
timestamp 1677583704
transform 1 0 22752 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_237
timestamp 1677583258
transform 1 0 23328 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_247
timestamp 1679585382
transform 1 0 24288 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_254
timestamp 1679585382
transform 1 0 24960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_261
timestamp 1679581501
transform 1 0 25632 0 1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_16_274
timestamp 1679585382
transform 1 0 26880 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_281
timestamp 1679585382
transform 1 0 27552 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_288
timestamp 1679585382
transform 1 0 28224 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_295
timestamp 1679585382
transform 1 0 28896 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_302
timestamp 1679585382
transform 1 0 29568 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_309
timestamp 1679585382
transform 1 0 30240 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_316
timestamp 1679585382
transform 1 0 30912 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_323
timestamp 1679585382
transform 1 0 31584 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_330
timestamp 1679585382
transform 1 0 32256 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_337
timestamp 1679585382
transform 1 0 32928 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_344
timestamp 1679585382
transform 1 0 33600 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_351
timestamp 1679585382
transform 1 0 34272 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_358
timestamp 1679585382
transform 1 0 34944 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_365
timestamp 1679585382
transform 1 0 35616 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_372
timestamp 1679585382
transform 1 0 36288 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_379
timestamp 1679585382
transform 1 0 36960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_386
timestamp 1679585382
transform 1 0 37632 0 1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_16_393
timestamp 1677583258
transform 1 0 38304 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_421
timestamp 1679581501
transform 1 0 40992 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_425
timestamp 1677583704
transform 1 0 41376 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_436
timestamp 1679585382
transform 1 0 42432 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_443
timestamp 1679585382
transform 1 0 43104 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_450
timestamp 1679585382
transform 1 0 43776 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_457
timestamp 1679585382
transform 1 0 44448 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_464
timestamp 1679585382
transform 1 0 45120 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_471
timestamp 1679585382
transform 1 0 45792 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_478
timestamp 1679585382
transform 1 0 46464 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_485
timestamp 1679585382
transform 1 0 47136 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_492
timestamp 1679585382
transform 1 0 47808 0 1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_16_499
timestamp 1677583258
transform 1 0 48480 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_517
timestamp 1679585382
transform 1 0 50208 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_524
timestamp 1679585382
transform 1 0 50880 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_531
timestamp 1679585382
transform 1 0 51552 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_538
timestamp 1679585382
transform 1 0 52224 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_545
timestamp 1679585382
transform 1 0 52896 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_579
timestamp 1679581501
transform 1 0 56160 0 1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_16_586
timestamp 1679585382
transform 1 0 56832 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_593
timestamp 1679585382
transform 1 0 57504 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_600
timestamp 1679585382
transform 1 0 58176 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_607
timestamp 1679585382
transform 1 0 58848 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_614
timestamp 1679585382
transform 1 0 59520 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_621
timestamp 1679585382
transform 1 0 60192 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_628
timestamp 1679585382
transform 1 0 60864 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_635
timestamp 1679585382
transform 1 0 61536 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_642
timestamp 1679585382
transform 1 0 62208 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_649
timestamp 1679585382
transform 1 0 62880 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_656
timestamp 1679585382
transform 1 0 63552 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_663
timestamp 1679585382
transform 1 0 64224 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_670
timestamp 1679585382
transform 1 0 64896 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_677
timestamp 1679585382
transform 1 0 65568 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_684
timestamp 1679585382
transform 1 0 66240 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_691
timestamp 1679585382
transform 1 0 66912 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_698
timestamp 1679585382
transform 1 0 67584 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_705
timestamp 1679585382
transform 1 0 68256 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_712
timestamp 1679585382
transform 1 0 68928 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_719
timestamp 1679585382
transform 1 0 69600 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_726
timestamp 1679585382
transform 1 0 70272 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_733
timestamp 1679585382
transform 1 0 70944 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_740
timestamp 1679585382
transform 1 0 71616 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_747
timestamp 1679585382
transform 1 0 72288 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_754
timestamp 1679585382
transform 1 0 72960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_761
timestamp 1679585382
transform 1 0 73632 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_768
timestamp 1679585382
transform 1 0 74304 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_775
timestamp 1679585382
transform 1 0 74976 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_782
timestamp 1679585382
transform 1 0 75648 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_789
timestamp 1679585382
transform 1 0 76320 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_796
timestamp 1679585382
transform 1 0 76992 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_803
timestamp 1679585382
transform 1 0 77664 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_810
timestamp 1679585382
transform 1 0 78336 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_817
timestamp 1679585382
transform 1 0 79008 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_824
timestamp 1679585382
transform 1 0 79680 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_831
timestamp 1679585382
transform 1 0 80352 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_838
timestamp 1679585382
transform 1 0 81024 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_845
timestamp 1679585382
transform 1 0 81696 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_852
timestamp 1679585382
transform 1 0 82368 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_859
timestamp 1679585382
transform 1 0 83040 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_866
timestamp 1679585382
transform 1 0 83712 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_873
timestamp 1679585382
transform 1 0 84384 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_880
timestamp 1679585382
transform 1 0 85056 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_887
timestamp 1679585382
transform 1 0 85728 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_894
timestamp 1679585382
transform 1 0 86400 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_901
timestamp 1679585382
transform 1 0 87072 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_908
timestamp 1679585382
transform 1 0 87744 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_915
timestamp 1679585382
transform 1 0 88416 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_922
timestamp 1679585382
transform 1 0 89088 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_929
timestamp 1679585382
transform 1 0 89760 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_936
timestamp 1679585382
transform 1 0 90432 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_943
timestamp 1679585382
transform 1 0 91104 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_950
timestamp 1679585382
transform 1 0 91776 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_957
timestamp 1679585382
transform 1 0 92448 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_964
timestamp 1679585382
transform 1 0 93120 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_971
timestamp 1679585382
transform 1 0 93792 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_978
timestamp 1679585382
transform 1 0 94464 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_985
timestamp 1679585382
transform 1 0 95136 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_992
timestamp 1679585382
transform 1 0 95808 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_999
timestamp 1679585382
transform 1 0 96480 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1006
timestamp 1679585382
transform 1 0 97152 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1013
timestamp 1679585382
transform 1 0 97824 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_1020
timestamp 1679585382
transform 1 0 98496 0 1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_16_1027
timestamp 1677583704
transform 1 0 99168 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_0
timestamp 1679585382
transform 1 0 576 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_7
timestamp 1679585382
transform 1 0 1248 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_14
timestamp 1679585382
transform 1 0 1920 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_21
timestamp 1677583704
transform 1 0 2592 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_23
timestamp 1677583258
transform 1 0 2784 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_55
timestamp 1677583704
transform 1 0 5856 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_57
timestamp 1677583258
transform 1 0 6048 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_71
timestamp 1679585382
transform 1 0 7392 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_78
timestamp 1679585382
transform 1 0 8064 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_85
timestamp 1677583704
transform 1 0 8736 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_87
timestamp 1677583258
transform 1 0 8928 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_128
timestamp 1679585382
transform 1 0 12864 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_135
timestamp 1679585382
transform 1 0 13536 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_142
timestamp 1679585382
transform 1 0 14208 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_149
timestamp 1679585382
transform 1 0 14880 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_156
timestamp 1679585382
transform 1 0 15552 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_163
timestamp 1679585382
transform 1 0 16224 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_170
timestamp 1679581501
transform 1 0 16896 0 -1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_17_178
timestamp 1679585382
transform 1 0 17664 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_185
timestamp 1677583258
transform 1 0 18336 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_195
timestamp 1679585382
transform 1 0 19296 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_202
timestamp 1679585382
transform 1 0 19968 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_209
timestamp 1679585382
transform 1 0 20640 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_216
timestamp 1679585382
transform 1 0 21312 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_223
timestamp 1679585382
transform 1 0 21984 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_230
timestamp 1679585382
transform 1 0 22656 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_237
timestamp 1679585382
transform 1 0 23328 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_244
timestamp 1679585382
transform 1 0 24000 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_251
timestamp 1679585382
transform 1 0 24672 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_258
timestamp 1679585382
transform 1 0 25344 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_265
timestamp 1679585382
transform 1 0 26016 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_272
timestamp 1677583258
transform 1 0 26688 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_286
timestamp 1679585382
transform 1 0 28032 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_293
timestamp 1679585382
transform 1 0 28704 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_300
timestamp 1679585382
transform 1 0 29376 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_307
timestamp 1679585382
transform 1 0 30048 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_314
timestamp 1679585382
transform 1 0 30720 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_321
timestamp 1679585382
transform 1 0 31392 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_328
timestamp 1679585382
transform 1 0 32064 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_335
timestamp 1679585382
transform 1 0 32736 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_342
timestamp 1679585382
transform 1 0 33408 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_349
timestamp 1679585382
transform 1 0 34080 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_356
timestamp 1679585382
transform 1 0 34752 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_363
timestamp 1679585382
transform 1 0 35424 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_370
timestamp 1679585382
transform 1 0 36096 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_377
timestamp 1679585382
transform 1 0 36768 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_384
timestamp 1679585382
transform 1 0 37440 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_391
timestamp 1677583704
transform 1 0 38112 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_393
timestamp 1677583258
transform 1 0 38304 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_403
timestamp 1679585382
transform 1 0 39264 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_410
timestamp 1679585382
transform 1 0 39936 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_417
timestamp 1679585382
transform 1 0 40608 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_424
timestamp 1679585382
transform 1 0 41280 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_431
timestamp 1679585382
transform 1 0 41952 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_438
timestamp 1679585382
transform 1 0 42624 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_445
timestamp 1677583258
transform 1 0 43296 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_17_481
timestamp 1679581501
transform 1 0 46752 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_17_485
timestamp 1677583258
transform 1 0 47136 0 -1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_522
timestamp 1679585382
transform 1 0 50688 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_529
timestamp 1679585382
transform 1 0 51360 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_536
timestamp 1679585382
transform 1 0 52032 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_543
timestamp 1679585382
transform 1 0 52704 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_550
timestamp 1679585382
transform 1 0 53376 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_557
timestamp 1679585382
transform 1 0 54048 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_564
timestamp 1677583704
transform 1 0 54720 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_566
timestamp 1677583258
transform 1 0 54912 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_575
timestamp 1677583704
transform 1 0 55776 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_599
timestamp 1679585382
transform 1 0 58080 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_606
timestamp 1677583704
transform 1 0 58752 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_635
timestamp 1679585382
transform 1 0 61536 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_642
timestamp 1679585382
transform 1 0 62208 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_649
timestamp 1679585382
transform 1 0 62880 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_656
timestamp 1679585382
transform 1 0 63552 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_663
timestamp 1679585382
transform 1 0 64224 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_670
timestamp 1679585382
transform 1 0 64896 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_677
timestamp 1679585382
transform 1 0 65568 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_684
timestamp 1679585382
transform 1 0 66240 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_691
timestamp 1679585382
transform 1 0 66912 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_698
timestamp 1679585382
transform 1 0 67584 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_705
timestamp 1679585382
transform 1 0 68256 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_712
timestamp 1679585382
transform 1 0 68928 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_719
timestamp 1679585382
transform 1 0 69600 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_726
timestamp 1679585382
transform 1 0 70272 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_733
timestamp 1679585382
transform 1 0 70944 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_740
timestamp 1679585382
transform 1 0 71616 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_747
timestamp 1679585382
transform 1 0 72288 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_754
timestamp 1679585382
transform 1 0 72960 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_761
timestamp 1679585382
transform 1 0 73632 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_768
timestamp 1679585382
transform 1 0 74304 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_775
timestamp 1679585382
transform 1 0 74976 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_782
timestamp 1679585382
transform 1 0 75648 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_789
timestamp 1679585382
transform 1 0 76320 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_796
timestamp 1679585382
transform 1 0 76992 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_803
timestamp 1679585382
transform 1 0 77664 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_810
timestamp 1679585382
transform 1 0 78336 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_817
timestamp 1679585382
transform 1 0 79008 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_824
timestamp 1679585382
transform 1 0 79680 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_831
timestamp 1679585382
transform 1 0 80352 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_838
timestamp 1679585382
transform 1 0 81024 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_845
timestamp 1679585382
transform 1 0 81696 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_852
timestamp 1679585382
transform 1 0 82368 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_859
timestamp 1679585382
transform 1 0 83040 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_866
timestamp 1679585382
transform 1 0 83712 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_873
timestamp 1679585382
transform 1 0 84384 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_880
timestamp 1679585382
transform 1 0 85056 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_887
timestamp 1679585382
transform 1 0 85728 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_894
timestamp 1679585382
transform 1 0 86400 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_901
timestamp 1679585382
transform 1 0 87072 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_908
timestamp 1679585382
transform 1 0 87744 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_915
timestamp 1679585382
transform 1 0 88416 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_922
timestamp 1679585382
transform 1 0 89088 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_929
timestamp 1679585382
transform 1 0 89760 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_936
timestamp 1679585382
transform 1 0 90432 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_943
timestamp 1679585382
transform 1 0 91104 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_950
timestamp 1679585382
transform 1 0 91776 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_957
timestamp 1679585382
transform 1 0 92448 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_964
timestamp 1679585382
transform 1 0 93120 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_971
timestamp 1679585382
transform 1 0 93792 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_978
timestamp 1679585382
transform 1 0 94464 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_985
timestamp 1679585382
transform 1 0 95136 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_992
timestamp 1679585382
transform 1 0 95808 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_999
timestamp 1679585382
transform 1 0 96480 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1006
timestamp 1679585382
transform 1 0 97152 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1013
timestamp 1679585382
transform 1 0 97824 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_1020
timestamp 1679585382
transform 1 0 98496 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_1027
timestamp 1677583704
transform 1 0 99168 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_4
timestamp 1679585382
transform 1 0 960 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_11
timestamp 1679585382
transform 1 0 1632 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_18
timestamp 1679585382
transform 1 0 2304 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_25
timestamp 1679585382
transform 1 0 2976 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_32
timestamp 1677583258
transform 1 0 3648 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_37
timestamp 1677583704
transform 1 0 4128 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_39
timestamp 1677583258
transform 1 0 4320 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_62
timestamp 1679585382
transform 1 0 6528 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_69
timestamp 1679585382
transform 1 0 7200 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_76
timestamp 1677583258
transform 1 0 7872 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_90
timestamp 1679585382
transform 1 0 9216 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_97
timestamp 1679585382
transform 1 0 9888 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_113
timestamp 1679585382
transform 1 0 11424 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_120
timestamp 1679585382
transform 1 0 12096 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_127
timestamp 1679585382
transform 1 0 12768 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_134
timestamp 1679585382
transform 1 0 13440 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_141
timestamp 1679585382
transform 1 0 14112 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_148
timestamp 1679585382
transform 1 0 14784 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_155
timestamp 1679585382
transform 1 0 15456 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_162
timestamp 1679585382
transform 1 0 16128 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_169
timestamp 1679585382
transform 1 0 16800 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_176
timestamp 1679585382
transform 1 0 17472 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_183
timestamp 1679585382
transform 1 0 18144 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_190
timestamp 1679585382
transform 1 0 18816 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_197
timestamp 1679585382
transform 1 0 19488 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_204
timestamp 1679585382
transform 1 0 20160 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_211
timestamp 1679581501
transform 1 0 20832 0 1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_18_242
timestamp 1679585382
transform 1 0 23808 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_249
timestamp 1679585382
transform 1 0 24480 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_256
timestamp 1679585382
transform 1 0 25152 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_263
timestamp 1679585382
transform 1 0 25824 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_270
timestamp 1679585382
transform 1 0 26496 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_277
timestamp 1679585382
transform 1 0 27168 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_284
timestamp 1679585382
transform 1 0 27840 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_291
timestamp 1679585382
transform 1 0 28512 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_298
timestamp 1679585382
transform 1 0 29184 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_305
timestamp 1679585382
transform 1 0 29856 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_312
timestamp 1679585382
transform 1 0 30528 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_319
timestamp 1679585382
transform 1 0 31200 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_326
timestamp 1679585382
transform 1 0 31872 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_333
timestamp 1679585382
transform 1 0 32544 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_340
timestamp 1679581501
transform 1 0 33216 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_352
timestamp 1677583258
transform 1 0 34368 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_389
timestamp 1677583704
transform 1 0 37920 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_391
timestamp 1677583258
transform 1 0 38112 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_400
timestamp 1679585382
transform 1 0 38976 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_407
timestamp 1679585382
transform 1 0 39648 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_414
timestamp 1679585382
transform 1 0 40320 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_421
timestamp 1679585382
transform 1 0 40992 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_428
timestamp 1679585382
transform 1 0 41664 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_435
timestamp 1679585382
transform 1 0 42336 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_442
timestamp 1679585382
transform 1 0 43008 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_449
timestamp 1679585382
transform 1 0 43680 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_456
timestamp 1679585382
transform 1 0 44352 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_463
timestamp 1679585382
transform 1 0 45024 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_470
timestamp 1679585382
transform 1 0 45696 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_477
timestamp 1679585382
transform 1 0 46368 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_484
timestamp 1679585382
transform 1 0 47040 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_491
timestamp 1679585382
transform 1 0 47712 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_498
timestamp 1679585382
transform 1 0 48384 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_505
timestamp 1679585382
transform 1 0 49056 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_512
timestamp 1679585382
transform 1 0 49728 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_519
timestamp 1679585382
transform 1 0 50400 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_526
timestamp 1677583258
transform 1 0 51072 0 1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_18_540
timestamp 1679581501
transform 1 0 52416 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_544
timestamp 1677583258
transform 1 0 52800 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_554
timestamp 1679585382
transform 1 0 53760 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_561
timestamp 1679585382
transform 1 0 54432 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_568
timestamp 1677583704
transform 1 0 55104 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_591
timestamp 1679585382
transform 1 0 57312 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_598
timestamp 1679585382
transform 1 0 57984 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_605
timestamp 1679581501
transform 1 0 58656 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_609
timestamp 1677583258
transform 1 0 59040 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_618
timestamp 1679585382
transform 1 0 59904 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_625
timestamp 1679585382
transform 1 0 60576 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_632
timestamp 1679585382
transform 1 0 61248 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_639
timestamp 1679585382
transform 1 0 61920 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_646
timestamp 1679585382
transform 1 0 62592 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_653
timestamp 1679585382
transform 1 0 63264 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_660
timestamp 1679585382
transform 1 0 63936 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_667
timestamp 1679585382
transform 1 0 64608 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_674
timestamp 1679585382
transform 1 0 65280 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_681
timestamp 1679585382
transform 1 0 65952 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_688
timestamp 1679585382
transform 1 0 66624 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_695
timestamp 1679585382
transform 1 0 67296 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_702
timestamp 1679585382
transform 1 0 67968 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_709
timestamp 1679585382
transform 1 0 68640 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_716
timestamp 1679585382
transform 1 0 69312 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_723
timestamp 1679585382
transform 1 0 69984 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_730
timestamp 1679585382
transform 1 0 70656 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_737
timestamp 1679585382
transform 1 0 71328 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_744
timestamp 1679585382
transform 1 0 72000 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_751
timestamp 1679585382
transform 1 0 72672 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_758
timestamp 1679585382
transform 1 0 73344 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_765
timestamp 1679585382
transform 1 0 74016 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_772
timestamp 1679585382
transform 1 0 74688 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_779
timestamp 1679585382
transform 1 0 75360 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_786
timestamp 1679585382
transform 1 0 76032 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_793
timestamp 1679585382
transform 1 0 76704 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_800
timestamp 1679585382
transform 1 0 77376 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_807
timestamp 1679585382
transform 1 0 78048 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_814
timestamp 1679585382
transform 1 0 78720 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_821
timestamp 1679585382
transform 1 0 79392 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_828
timestamp 1679585382
transform 1 0 80064 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_835
timestamp 1679585382
transform 1 0 80736 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_842
timestamp 1679585382
transform 1 0 81408 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_849
timestamp 1679585382
transform 1 0 82080 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_856
timestamp 1679585382
transform 1 0 82752 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_863
timestamp 1679585382
transform 1 0 83424 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_870
timestamp 1679585382
transform 1 0 84096 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_877
timestamp 1679585382
transform 1 0 84768 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_884
timestamp 1679585382
transform 1 0 85440 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_891
timestamp 1679585382
transform 1 0 86112 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_898
timestamp 1679585382
transform 1 0 86784 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_905
timestamp 1679585382
transform 1 0 87456 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_912
timestamp 1679585382
transform 1 0 88128 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_919
timestamp 1679585382
transform 1 0 88800 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_926
timestamp 1679585382
transform 1 0 89472 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_933
timestamp 1679585382
transform 1 0 90144 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_940
timestamp 1679585382
transform 1 0 90816 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_947
timestamp 1679585382
transform 1 0 91488 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_954
timestamp 1679585382
transform 1 0 92160 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_961
timestamp 1679585382
transform 1 0 92832 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_968
timestamp 1679585382
transform 1 0 93504 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_975
timestamp 1679585382
transform 1 0 94176 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_982
timestamp 1679585382
transform 1 0 94848 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_989
timestamp 1679585382
transform 1 0 95520 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_996
timestamp 1679585382
transform 1 0 96192 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1003
timestamp 1679585382
transform 1 0 96864 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1010
timestamp 1679585382
transform 1 0 97536 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_1017
timestamp 1679585382
transform 1 0 98208 0 1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_18_1024
timestamp 1679581501
transform 1 0 98880 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_1028
timestamp 1677583258
transform 1 0 99264 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_4
timestamp 1679585382
transform 1 0 960 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_11
timestamp 1679585382
transform 1 0 1632 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_18
timestamp 1679585382
transform 1 0 2304 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_25
timestamp 1679585382
transform 1 0 2976 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_32
timestamp 1679585382
transform 1 0 3648 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_39
timestamp 1679585382
transform 1 0 4320 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_46
timestamp 1679585382
transform 1 0 4992 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_53
timestamp 1679585382
transform 1 0 5664 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_60
timestamp 1679585382
transform 1 0 6336 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_67
timestamp 1679585382
transform 1 0 7008 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_74
timestamp 1679585382
transform 1 0 7680 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_81
timestamp 1679585382
transform 1 0 8352 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_88
timestamp 1679585382
transform 1 0 9024 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_95
timestamp 1679585382
transform 1 0 9696 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_102
timestamp 1679585382
transform 1 0 10368 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_109
timestamp 1679585382
transform 1 0 11040 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_116
timestamp 1679585382
transform 1 0 11712 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_123
timestamp 1679585382
transform 1 0 12384 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_130
timestamp 1679585382
transform 1 0 13056 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_137
timestamp 1679585382
transform 1 0 13728 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_144
timestamp 1679585382
transform 1 0 14400 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_151
timestamp 1679581501
transform 1 0 15072 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_155
timestamp 1677583258
transform 1 0 15456 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_173
timestamp 1677583704
transform 1 0 17184 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_191
timestamp 1679585382
transform 1 0 18912 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_198
timestamp 1677583704
transform 1 0 19584 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_200
timestamp 1677583258
transform 1 0 19776 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_209
timestamp 1679585382
transform 1 0 20640 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_216
timestamp 1679585382
transform 1 0 21312 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_223
timestamp 1677583704
transform 1 0 21984 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_234
timestamp 1679585382
transform 1 0 23040 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_241
timestamp 1679585382
transform 1 0 23712 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_248
timestamp 1679585382
transform 1 0 24384 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_255
timestamp 1677583704
transform 1 0 25056 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_284
timestamp 1679585382
transform 1 0 27840 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_291
timestamp 1679585382
transform 1 0 28512 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_298
timestamp 1679585382
transform 1 0 29184 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_305
timestamp 1679585382
transform 1 0 29856 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_312
timestamp 1679585382
transform 1 0 30528 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_319
timestamp 1679585382
transform 1 0 31200 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_326
timestamp 1679585382
transform 1 0 31872 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_333
timestamp 1679585382
transform 1 0 32544 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_340
timestamp 1677583704
transform 1 0 33216 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_355
timestamp 1679585382
transform 1 0 34656 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_362
timestamp 1679585382
transform 1 0 35328 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_369
timestamp 1679585382
transform 1 0 36000 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_376
timestamp 1679585382
transform 1 0 36672 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_383
timestamp 1679585382
transform 1 0 37344 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_390
timestamp 1679581501
transform 1 0 38016 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_394
timestamp 1677583704
transform 1 0 38400 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_4  FILLER_19_409
timestamp 1679581501
transform 1 0 39840 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_413
timestamp 1677583258
transform 1 0 40224 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_422
timestamp 1679581501
transform 1 0 41088 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_426
timestamp 1677583704
transform 1 0 41472 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_455
timestamp 1679585382
transform 1 0 44256 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_462
timestamp 1679585382
transform 1 0 44928 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_469
timestamp 1679585382
transform 1 0 45600 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_476
timestamp 1679585382
transform 1 0 46272 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_483
timestamp 1679585382
transform 1 0 46944 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_490
timestamp 1679585382
transform 1 0 47616 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_497
timestamp 1679585382
transform 1 0 48288 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_504
timestamp 1679585382
transform 1 0 48960 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_511
timestamp 1679585382
transform 1 0 49632 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_518
timestamp 1679585382
transform 1 0 50304 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_525
timestamp 1679585382
transform 1 0 50976 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_532
timestamp 1679585382
transform 1 0 51648 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_539
timestamp 1679585382
transform 1 0 52320 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_546
timestamp 1679585382
transform 1 0 52992 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_553
timestamp 1679585382
transform 1 0 53664 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_560
timestamp 1679585382
transform 1 0 54336 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_567
timestamp 1679585382
transform 1 0 55008 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_574
timestamp 1679585382
transform 1 0 55680 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_581
timestamp 1679585382
transform 1 0 56352 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_588
timestamp 1679585382
transform 1 0 57024 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_595
timestamp 1679585382
transform 1 0 57696 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_602
timestamp 1679585382
transform 1 0 58368 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_609
timestamp 1679585382
transform 1 0 59040 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_616
timestamp 1679585382
transform 1 0 59712 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_623
timestamp 1679585382
transform 1 0 60384 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_630
timestamp 1679585382
transform 1 0 61056 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_637
timestamp 1679585382
transform 1 0 61728 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_644
timestamp 1679585382
transform 1 0 62400 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_651
timestamp 1679585382
transform 1 0 63072 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_658
timestamp 1679585382
transform 1 0 63744 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_665
timestamp 1679585382
transform 1 0 64416 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_672
timestamp 1679585382
transform 1 0 65088 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_679
timestamp 1679585382
transform 1 0 65760 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_686
timestamp 1679585382
transform 1 0 66432 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_693
timestamp 1679585382
transform 1 0 67104 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_700
timestamp 1679585382
transform 1 0 67776 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_707
timestamp 1679585382
transform 1 0 68448 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_714
timestamp 1679585382
transform 1 0 69120 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_721
timestamp 1679585382
transform 1 0 69792 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_728
timestamp 1679585382
transform 1 0 70464 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_735
timestamp 1679585382
transform 1 0 71136 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_742
timestamp 1679585382
transform 1 0 71808 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_749
timestamp 1679585382
transform 1 0 72480 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_756
timestamp 1679585382
transform 1 0 73152 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_763
timestamp 1679585382
transform 1 0 73824 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_770
timestamp 1679585382
transform 1 0 74496 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_777
timestamp 1679585382
transform 1 0 75168 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_784
timestamp 1679585382
transform 1 0 75840 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_791
timestamp 1679585382
transform 1 0 76512 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_798
timestamp 1679585382
transform 1 0 77184 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_805
timestamp 1679585382
transform 1 0 77856 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_812
timestamp 1679585382
transform 1 0 78528 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_819
timestamp 1679585382
transform 1 0 79200 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_826
timestamp 1679585382
transform 1 0 79872 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_833
timestamp 1679585382
transform 1 0 80544 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_840
timestamp 1679585382
transform 1 0 81216 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_847
timestamp 1679585382
transform 1 0 81888 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_854
timestamp 1679585382
transform 1 0 82560 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_861
timestamp 1679585382
transform 1 0 83232 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_868
timestamp 1679585382
transform 1 0 83904 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_875
timestamp 1679585382
transform 1 0 84576 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_882
timestamp 1679585382
transform 1 0 85248 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_889
timestamp 1679585382
transform 1 0 85920 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_896
timestamp 1679585382
transform 1 0 86592 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_903
timestamp 1679585382
transform 1 0 87264 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_910
timestamp 1679585382
transform 1 0 87936 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_917
timestamp 1679585382
transform 1 0 88608 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_924
timestamp 1679585382
transform 1 0 89280 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_931
timestamp 1679585382
transform 1 0 89952 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_938
timestamp 1679585382
transform 1 0 90624 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_945
timestamp 1679585382
transform 1 0 91296 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_952
timestamp 1679585382
transform 1 0 91968 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_959
timestamp 1679585382
transform 1 0 92640 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_966
timestamp 1679585382
transform 1 0 93312 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_973
timestamp 1679585382
transform 1 0 93984 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_980
timestamp 1679585382
transform 1 0 94656 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_987
timestamp 1679585382
transform 1 0 95328 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_994
timestamp 1679585382
transform 1 0 96000 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1001
timestamp 1679585382
transform 1 0 96672 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1008
timestamp 1679585382
transform 1 0 97344 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1015
timestamp 1679585382
transform 1 0 98016 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_1022
timestamp 1679585382
transform 1 0 98688 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_4
timestamp 1679585382
transform 1 0 960 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_11
timestamp 1679585382
transform 1 0 1632 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_18
timestamp 1679585382
transform 1 0 2304 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_25
timestamp 1679585382
transform 1 0 2976 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_32
timestamp 1679585382
transform 1 0 3648 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_39
timestamp 1679585382
transform 1 0 4320 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_46
timestamp 1679585382
transform 1 0 4992 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_53
timestamp 1679585382
transform 1 0 5664 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_60
timestamp 1679585382
transform 1 0 6336 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_67
timestamp 1679585382
transform 1 0 7008 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_74
timestamp 1679585382
transform 1 0 7680 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_81
timestamp 1679585382
transform 1 0 8352 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_88
timestamp 1679585382
transform 1 0 9024 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_95
timestamp 1679581501
transform 1 0 9696 0 1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_20_112
timestamp 1679585382
transform 1 0 11328 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_119
timestamp 1679585382
transform 1 0 12000 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_126
timestamp 1679585382
transform 1 0 12672 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_133
timestamp 1679585382
transform 1 0 13344 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_140
timestamp 1679581501
transform 1 0 14016 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_144
timestamp 1677583258
transform 1 0 14400 0 1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_181
timestamp 1679581501
transform 1 0 17952 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_185
timestamp 1677583258
transform 1 0 18336 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_217
timestamp 1679585382
transform 1 0 21408 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_224
timestamp 1679585382
transform 1 0 22080 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_231
timestamp 1679585382
transform 1 0 22752 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_238
timestamp 1679585382
transform 1 0 23424 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_245
timestamp 1679585382
transform 1 0 24096 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_252
timestamp 1679585382
transform 1 0 24768 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_259
timestamp 1679585382
transform 1 0 25440 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_266
timestamp 1679585382
transform 1 0 26112 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_273
timestamp 1679585382
transform 1 0 26784 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_280
timestamp 1679585382
transform 1 0 27456 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_287
timestamp 1679585382
transform 1 0 28128 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_294
timestamp 1679585382
transform 1 0 28800 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_301
timestamp 1679585382
transform 1 0 29472 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_308
timestamp 1679585382
transform 1 0 30144 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_315
timestamp 1677583704
transform 1 0 30816 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_344
timestamp 1677583258
transform 1 0 33600 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_353
timestamp 1679585382
transform 1 0 34464 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_360
timestamp 1679585382
transform 1 0 35136 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_367
timestamp 1679585382
transform 1 0 35808 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_374
timestamp 1679585382
transform 1 0 36480 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_381
timestamp 1679585382
transform 1 0 37152 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_388
timestamp 1679585382
transform 1 0 37824 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_395
timestamp 1679585382
transform 1 0 38496 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_402
timestamp 1679585382
transform 1 0 39168 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_409
timestamp 1679585382
transform 1 0 39840 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_416
timestamp 1679585382
transform 1 0 40512 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_423
timestamp 1677583704
transform 1 0 41184 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_20_434
timestamp 1679585382
transform 1 0 42240 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_441
timestamp 1679585382
transform 1 0 42912 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_448
timestamp 1679585382
transform 1 0 43584 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_455
timestamp 1679585382
transform 1 0 44256 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_462
timestamp 1679585382
transform 1 0 44928 0 1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_469
timestamp 1677583258
transform 1 0 45600 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_483
timestamp 1679585382
transform 1 0 46944 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_490
timestamp 1679585382
transform 1 0 47616 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_497
timestamp 1679585382
transform 1 0 48288 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_504
timestamp 1679585382
transform 1 0 48960 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_511
timestamp 1679585382
transform 1 0 49632 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_518
timestamp 1679585382
transform 1 0 50304 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_525
timestamp 1679585382
transform 1 0 50976 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_532
timestamp 1679585382
transform 1 0 51648 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_539
timestamp 1679585382
transform 1 0 52320 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_546
timestamp 1679585382
transform 1 0 52992 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_553
timestamp 1679585382
transform 1 0 53664 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_560
timestamp 1679585382
transform 1 0 54336 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_567
timestamp 1677583704
transform 1 0 55008 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_569
timestamp 1677583258
transform 1 0 55200 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_579
timestamp 1679585382
transform 1 0 56160 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_586
timestamp 1679585382
transform 1 0 56832 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_593
timestamp 1679585382
transform 1 0 57504 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_600
timestamp 1679585382
transform 1 0 58176 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_607
timestamp 1679585382
transform 1 0 58848 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_614
timestamp 1679585382
transform 1 0 59520 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_621
timestamp 1679585382
transform 1 0 60192 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_628
timestamp 1679585382
transform 1 0 60864 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_635
timestamp 1679585382
transform 1 0 61536 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_642
timestamp 1679585382
transform 1 0 62208 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_649
timestamp 1679585382
transform 1 0 62880 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_656
timestamp 1679585382
transform 1 0 63552 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_663
timestamp 1679585382
transform 1 0 64224 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_670
timestamp 1679585382
transform 1 0 64896 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_677
timestamp 1679585382
transform 1 0 65568 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_684
timestamp 1679585382
transform 1 0 66240 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_691
timestamp 1679585382
transform 1 0 66912 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_698
timestamp 1679585382
transform 1 0 67584 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_705
timestamp 1679585382
transform 1 0 68256 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_712
timestamp 1679585382
transform 1 0 68928 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_719
timestamp 1679585382
transform 1 0 69600 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_726
timestamp 1679585382
transform 1 0 70272 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_733
timestamp 1679585382
transform 1 0 70944 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_740
timestamp 1679585382
transform 1 0 71616 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_747
timestamp 1679585382
transform 1 0 72288 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_754
timestamp 1679585382
transform 1 0 72960 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_761
timestamp 1679585382
transform 1 0 73632 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_768
timestamp 1679585382
transform 1 0 74304 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_775
timestamp 1679585382
transform 1 0 74976 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_782
timestamp 1679585382
transform 1 0 75648 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_789
timestamp 1679585382
transform 1 0 76320 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_796
timestamp 1679585382
transform 1 0 76992 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_803
timestamp 1679585382
transform 1 0 77664 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_810
timestamp 1679585382
transform 1 0 78336 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_817
timestamp 1679585382
transform 1 0 79008 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_824
timestamp 1679585382
transform 1 0 79680 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_831
timestamp 1679585382
transform 1 0 80352 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_838
timestamp 1679585382
transform 1 0 81024 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_845
timestamp 1679585382
transform 1 0 81696 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_852
timestamp 1679585382
transform 1 0 82368 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_859
timestamp 1679585382
transform 1 0 83040 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_866
timestamp 1679585382
transform 1 0 83712 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_873
timestamp 1679585382
transform 1 0 84384 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_880
timestamp 1679585382
transform 1 0 85056 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_887
timestamp 1679585382
transform 1 0 85728 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_894
timestamp 1679585382
transform 1 0 86400 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_901
timestamp 1679585382
transform 1 0 87072 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_908
timestamp 1679585382
transform 1 0 87744 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_915
timestamp 1679585382
transform 1 0 88416 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_922
timestamp 1679585382
transform 1 0 89088 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_929
timestamp 1679585382
transform 1 0 89760 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_936
timestamp 1679585382
transform 1 0 90432 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_943
timestamp 1679585382
transform 1 0 91104 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_950
timestamp 1679585382
transform 1 0 91776 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_957
timestamp 1679585382
transform 1 0 92448 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_964
timestamp 1679585382
transform 1 0 93120 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_971
timestamp 1679585382
transform 1 0 93792 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_978
timestamp 1679585382
transform 1 0 94464 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_985
timestamp 1679585382
transform 1 0 95136 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_992
timestamp 1679585382
transform 1 0 95808 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_999
timestamp 1679585382
transform 1 0 96480 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1006
timestamp 1679585382
transform 1 0 97152 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1013
timestamp 1679585382
transform 1 0 97824 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1020
timestamp 1679585382
transform 1 0 98496 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_1027
timestamp 1677583704
transform 1 0 99168 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_4
timestamp 1679585382
transform 1 0 960 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_11
timestamp 1679585382
transform 1 0 1632 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_18
timestamp 1679585382
transform 1 0 2304 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_29
timestamp 1679581501
transform 1 0 3360 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_21_33
timestamp 1677583704
transform 1 0 3744 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_44
timestamp 1679585382
transform 1 0 4800 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_51
timestamp 1679585382
transform 1 0 5472 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_58
timestamp 1679585382
transform 1 0 6144 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_65
timestamp 1679585382
transform 1 0 6816 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_72
timestamp 1679585382
transform 1 0 7488 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_79
timestamp 1679585382
transform 1 0 8160 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_86
timestamp 1679585382
transform 1 0 8832 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_120
timestamp 1679585382
transform 1 0 12096 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_127
timestamp 1679585382
transform 1 0 12768 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_134
timestamp 1679585382
transform 1 0 13440 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_141
timestamp 1679585382
transform 1 0 14112 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_175
timestamp 1679585382
transform 1 0 17376 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_182
timestamp 1679585382
transform 1 0 18048 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_189
timestamp 1679585382
transform 1 0 18720 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_218
timestamp 1679585382
transform 1 0 21504 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_225
timestamp 1679585382
transform 1 0 22176 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_232
timestamp 1679581501
transform 1 0 22848 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_236
timestamp 1677583258
transform 1 0 23232 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_246
timestamp 1679585382
transform 1 0 24192 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_253
timestamp 1679585382
transform 1 0 24864 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_260
timestamp 1679581501
transform 1 0 25536 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_21_264
timestamp 1677583704
transform 1 0 25920 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_293
timestamp 1679585382
transform 1 0 28704 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_300
timestamp 1679585382
transform 1 0 29376 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_307
timestamp 1679585382
transform 1 0 30048 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_314
timestamp 1679585382
transform 1 0 30720 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_321
timestamp 1679585382
transform 1 0 31392 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_328
timestamp 1679581501
transform 1 0 32064 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_21_332
timestamp 1677583704
transform 1 0 32448 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_21_342
timestamp 1677583704
transform 1 0 33408 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_344
timestamp 1677583258
transform 1 0 33600 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_354
timestamp 1679585382
transform 1 0 34560 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_21_361
timestamp 1677583258
transform 1 0 35232 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_398
timestamp 1679585382
transform 1 0 38784 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_405
timestamp 1679585382
transform 1 0 39456 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_412
timestamp 1677583704
transform 1 0 40128 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_422
timestamp 1679585382
transform 1 0 41088 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_429
timestamp 1679585382
transform 1 0 41760 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_436
timestamp 1679585382
transform 1 0 42432 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_443
timestamp 1679585382
transform 1 0 43104 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_450
timestamp 1679585382
transform 1 0 43776 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_457
timestamp 1679581501
transform 1 0 44448 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_461
timestamp 1677583258
transform 1 0 44832 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_475
timestamp 1679585382
transform 1 0 46176 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_482
timestamp 1679585382
transform 1 0 46848 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_489
timestamp 1677583704
transform 1 0 47520 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_518
timestamp 1679585382
transform 1 0 50304 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_525
timestamp 1679585382
transform 1 0 50976 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_532
timestamp 1679585382
transform 1 0 51648 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_539
timestamp 1679581501
transform 1 0 52320 0 -1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_21_570
timestamp 1679585382
transform 1 0 55296 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_577
timestamp 1679581501
transform 1 0 55968 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_21_581
timestamp 1677583704
transform 1 0 56352 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_610
timestamp 1679585382
transform 1 0 59136 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_617
timestamp 1679585382
transform 1 0 59808 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_624
timestamp 1679585382
transform 1 0 60480 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_631
timestamp 1679585382
transform 1 0 61152 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_638
timestamp 1679585382
transform 1 0 61824 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_645
timestamp 1679585382
transform 1 0 62496 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_652
timestamp 1679585382
transform 1 0 63168 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_659
timestamp 1679585382
transform 1 0 63840 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_666
timestamp 1679585382
transform 1 0 64512 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_673
timestamp 1679585382
transform 1 0 65184 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_680
timestamp 1679585382
transform 1 0 65856 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_687
timestamp 1679585382
transform 1 0 66528 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_694
timestamp 1679585382
transform 1 0 67200 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_701
timestamp 1679585382
transform 1 0 67872 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_708
timestamp 1679585382
transform 1 0 68544 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_715
timestamp 1679585382
transform 1 0 69216 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_722
timestamp 1679585382
transform 1 0 69888 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_729
timestamp 1679585382
transform 1 0 70560 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_736
timestamp 1679585382
transform 1 0 71232 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_743
timestamp 1679585382
transform 1 0 71904 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_750
timestamp 1679585382
transform 1 0 72576 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_757
timestamp 1679585382
transform 1 0 73248 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_764
timestamp 1679585382
transform 1 0 73920 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_771
timestamp 1679585382
transform 1 0 74592 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_778
timestamp 1679585382
transform 1 0 75264 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_785
timestamp 1679585382
transform 1 0 75936 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_792
timestamp 1679585382
transform 1 0 76608 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_799
timestamp 1679585382
transform 1 0 77280 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_806
timestamp 1679585382
transform 1 0 77952 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_813
timestamp 1679585382
transform 1 0 78624 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_820
timestamp 1679585382
transform 1 0 79296 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_827
timestamp 1679585382
transform 1 0 79968 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_834
timestamp 1679585382
transform 1 0 80640 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_841
timestamp 1679585382
transform 1 0 81312 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_848
timestamp 1679585382
transform 1 0 81984 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_855
timestamp 1679585382
transform 1 0 82656 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_862
timestamp 1679585382
transform 1 0 83328 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_869
timestamp 1679585382
transform 1 0 84000 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_876
timestamp 1679585382
transform 1 0 84672 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_883
timestamp 1679585382
transform 1 0 85344 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_890
timestamp 1679585382
transform 1 0 86016 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_897
timestamp 1679585382
transform 1 0 86688 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_904
timestamp 1679585382
transform 1 0 87360 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_911
timestamp 1679585382
transform 1 0 88032 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_918
timestamp 1679585382
transform 1 0 88704 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_925
timestamp 1679585382
transform 1 0 89376 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_932
timestamp 1679585382
transform 1 0 90048 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_939
timestamp 1679585382
transform 1 0 90720 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_946
timestamp 1679585382
transform 1 0 91392 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_953
timestamp 1679585382
transform 1 0 92064 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_960
timestamp 1679585382
transform 1 0 92736 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_967
timestamp 1679585382
transform 1 0 93408 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_974
timestamp 1679585382
transform 1 0 94080 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_981
timestamp 1679585382
transform 1 0 94752 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_988
timestamp 1679585382
transform 1 0 95424 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_995
timestamp 1679585382
transform 1 0 96096 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1002
timestamp 1679585382
transform 1 0 96768 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1009
timestamp 1679585382
transform 1 0 97440 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1016
timestamp 1679585382
transform 1 0 98112 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_1023
timestamp 1679581501
transform 1 0 98784 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_21_1027
timestamp 1677583704
transform 1 0 99168 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_4
timestamp 1679585382
transform 1 0 960 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_11
timestamp 1679581501
transform 1 0 1632 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_15
timestamp 1677583258
transform 1 0 2016 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_43
timestamp 1679585382
transform 1 0 4704 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_50
timestamp 1679585382
transform 1 0 5376 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_57
timestamp 1679585382
transform 1 0 6048 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_64
timestamp 1679585382
transform 1 0 6720 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_71
timestamp 1679585382
transform 1 0 7392 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_78
timestamp 1679581501
transform 1 0 8064 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_82
timestamp 1677583258
transform 1 0 8448 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_110
timestamp 1679585382
transform 1 0 11136 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_117
timestamp 1679585382
transform 1 0 11808 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_124
timestamp 1679585382
transform 1 0 12480 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_131
timestamp 1679585382
transform 1 0 13152 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_138
timestamp 1679585382
transform 1 0 13824 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_145
timestamp 1679585382
transform 1 0 14496 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_152
timestamp 1679581501
transform 1 0 15168 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_156
timestamp 1677583704
transform 1 0 15552 0 1 17388
box -48 -56 240 834
use sg13g2_decap_4  FILLER_22_162
timestamp 1679581501
transform 1 0 16128 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_166
timestamp 1677583704
transform 1 0 16512 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_177
timestamp 1679585382
transform 1 0 17568 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_184
timestamp 1679585382
transform 1 0 18240 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_191
timestamp 1679585382
transform 1 0 18912 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_198
timestamp 1679585382
transform 1 0 19584 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_205
timestamp 1679585382
transform 1 0 20256 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_212
timestamp 1679585382
transform 1 0 20928 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_219
timestamp 1679585382
transform 1 0 21600 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_226
timestamp 1679585382
transform 1 0 22272 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_233
timestamp 1679585382
transform 1 0 22944 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_240
timestamp 1679585382
transform 1 0 23616 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_247
timestamp 1679585382
transform 1 0 24288 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_254
timestamp 1679585382
transform 1 0 24960 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_302
timestamp 1679585382
transform 1 0 29568 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_309
timestamp 1679585382
transform 1 0 30240 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_316
timestamp 1679585382
transform 1 0 30912 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_323
timestamp 1679585382
transform 1 0 31584 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_330
timestamp 1679585382
transform 1 0 32256 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_337
timestamp 1679585382
transform 1 0 32928 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_344
timestamp 1679585382
transform 1 0 33600 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_351
timestamp 1679585382
transform 1 0 34272 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_358
timestamp 1679585382
transform 1 0 34944 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_365
timestamp 1679585382
transform 1 0 35616 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_372
timestamp 1679585382
transform 1 0 36288 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_379
timestamp 1679585382
transform 1 0 36960 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_386
timestamp 1677583704
transform 1 0 37632 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_397
timestamp 1679585382
transform 1 0 38688 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_404
timestamp 1679585382
transform 1 0 39360 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_411
timestamp 1679585382
transform 1 0 40032 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_418
timestamp 1679585382
transform 1 0 40704 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_425
timestamp 1679585382
transform 1 0 41376 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_432
timestamp 1679581501
transform 1 0 42048 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_436
timestamp 1677583704
transform 1 0 42432 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_451
timestamp 1679585382
transform 1 0 43872 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_458
timestamp 1679585382
transform 1 0 44544 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_465
timestamp 1679585382
transform 1 0 45216 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_472
timestamp 1679585382
transform 1 0 45888 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_479
timestamp 1679585382
transform 1 0 46560 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_486
timestamp 1679585382
transform 1 0 47232 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_493
timestamp 1679585382
transform 1 0 47904 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_500
timestamp 1677583704
transform 1 0 48576 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_506
timestamp 1677583258
transform 1 0 49152 0 1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_22_520
timestamp 1679581501
transform 1 0 50496 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_524
timestamp 1677583704
transform 1 0 50880 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_530
timestamp 1679585382
transform 1 0 51456 0 1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_22_537
timestamp 1677583258
transform 1 0 52128 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_543
timestamp 1679585382
transform 1 0 52704 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_550
timestamp 1679585382
transform 1 0 53376 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_557
timestamp 1679585382
transform 1 0 54048 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_564
timestamp 1679581501
transform 1 0 54720 0 1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_22_576
timestamp 1679585382
transform 1 0 55872 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_583
timestamp 1679585382
transform 1 0 56544 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_590
timestamp 1679585382
transform 1 0 57216 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_597
timestamp 1679585382
transform 1 0 57888 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_604
timestamp 1679585382
transform 1 0 58560 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_611
timestamp 1679585382
transform 1 0 59232 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_618
timestamp 1679585382
transform 1 0 59904 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_625
timestamp 1679585382
transform 1 0 60576 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_632
timestamp 1679585382
transform 1 0 61248 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_639
timestamp 1679585382
transform 1 0 61920 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_646
timestamp 1679585382
transform 1 0 62592 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_653
timestamp 1679585382
transform 1 0 63264 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_660
timestamp 1679585382
transform 1 0 63936 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_667
timestamp 1679585382
transform 1 0 64608 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_674
timestamp 1679585382
transform 1 0 65280 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_681
timestamp 1679585382
transform 1 0 65952 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_688
timestamp 1679585382
transform 1 0 66624 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_695
timestamp 1679585382
transform 1 0 67296 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_702
timestamp 1679585382
transform 1 0 67968 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_709
timestamp 1679585382
transform 1 0 68640 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_716
timestamp 1679585382
transform 1 0 69312 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_723
timestamp 1679585382
transform 1 0 69984 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_730
timestamp 1679585382
transform 1 0 70656 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_737
timestamp 1679585382
transform 1 0 71328 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_744
timestamp 1679585382
transform 1 0 72000 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_751
timestamp 1679585382
transform 1 0 72672 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_758
timestamp 1679585382
transform 1 0 73344 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_765
timestamp 1679585382
transform 1 0 74016 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_772
timestamp 1679585382
transform 1 0 74688 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_779
timestamp 1679585382
transform 1 0 75360 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_786
timestamp 1679585382
transform 1 0 76032 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_793
timestamp 1679585382
transform 1 0 76704 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_800
timestamp 1679585382
transform 1 0 77376 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_807
timestamp 1679585382
transform 1 0 78048 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_814
timestamp 1679585382
transform 1 0 78720 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_821
timestamp 1679585382
transform 1 0 79392 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_828
timestamp 1679585382
transform 1 0 80064 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_835
timestamp 1679585382
transform 1 0 80736 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_842
timestamp 1679585382
transform 1 0 81408 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_849
timestamp 1679585382
transform 1 0 82080 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_856
timestamp 1679585382
transform 1 0 82752 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_863
timestamp 1679585382
transform 1 0 83424 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_870
timestamp 1679585382
transform 1 0 84096 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_877
timestamp 1679585382
transform 1 0 84768 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_884
timestamp 1679585382
transform 1 0 85440 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_891
timestamp 1679585382
transform 1 0 86112 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_898
timestamp 1679585382
transform 1 0 86784 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_905
timestamp 1679585382
transform 1 0 87456 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_912
timestamp 1679585382
transform 1 0 88128 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_919
timestamp 1679585382
transform 1 0 88800 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_926
timestamp 1679585382
transform 1 0 89472 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_933
timestamp 1679585382
transform 1 0 90144 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_940
timestamp 1679585382
transform 1 0 90816 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_947
timestamp 1679585382
transform 1 0 91488 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_954
timestamp 1679585382
transform 1 0 92160 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_961
timestamp 1679585382
transform 1 0 92832 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_968
timestamp 1679585382
transform 1 0 93504 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_975
timestamp 1679585382
transform 1 0 94176 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_982
timestamp 1679585382
transform 1 0 94848 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_989
timestamp 1679585382
transform 1 0 95520 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_996
timestamp 1679585382
transform 1 0 96192 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1003
timestamp 1679585382
transform 1 0 96864 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1010
timestamp 1679585382
transform 1 0 97536 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1017
timestamp 1679585382
transform 1 0 98208 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_1024
timestamp 1679581501
transform 1 0 98880 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_1028
timestamp 1677583258
transform 1 0 99264 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_4
timestamp 1679585382
transform 1 0 960 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_11
timestamp 1679581501
transform 1 0 1632 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_15
timestamp 1677583704
transform 1 0 2016 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_44
timestamp 1679585382
transform 1 0 4800 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_51
timestamp 1679585382
transform 1 0 5472 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_58
timestamp 1679585382
transform 1 0 6144 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_65
timestamp 1679585382
transform 1 0 6816 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_72
timestamp 1679585382
transform 1 0 7488 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_79
timestamp 1679585382
transform 1 0 8160 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_86
timestamp 1679585382
transform 1 0 8832 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_93
timestamp 1679585382
transform 1 0 9504 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_100
timestamp 1679581501
transform 1 0 10176 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_104
timestamp 1677583258
transform 1 0 10560 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_113
timestamp 1679585382
transform 1 0 11424 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_120
timestamp 1679585382
transform 1 0 12096 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_127
timestamp 1679585382
transform 1 0 12768 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_134
timestamp 1679585382
transform 1 0 13440 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_141
timestamp 1679585382
transform 1 0 14112 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_148
timestamp 1679585382
transform 1 0 14784 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_155
timestamp 1679585382
transform 1 0 15456 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_162
timestamp 1679585382
transform 1 0 16128 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_169
timestamp 1679585382
transform 1 0 16800 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_176
timestamp 1679585382
transform 1 0 17472 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_183
timestamp 1679585382
transform 1 0 18144 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_190
timestamp 1679585382
transform 1 0 18816 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_197
timestamp 1679585382
transform 1 0 19488 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_204
timestamp 1679585382
transform 1 0 20160 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_211
timestamp 1679585382
transform 1 0 20832 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_218
timestamp 1679585382
transform 1 0 21504 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_225
timestamp 1679585382
transform 1 0 22176 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_232
timestamp 1679585382
transform 1 0 22848 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_239
timestamp 1679585382
transform 1 0 23520 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_246
timestamp 1679585382
transform 1 0 24192 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_253
timestamp 1679585382
transform 1 0 24864 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_260
timestamp 1679585382
transform 1 0 25536 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_267
timestamp 1679581501
transform 1 0 26208 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_279
timestamp 1677583704
transform 1 0 27360 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_290
timestamp 1679585382
transform 1 0 28416 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_297
timestamp 1679585382
transform 1 0 29088 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_304
timestamp 1679585382
transform 1 0 29760 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_311
timestamp 1679585382
transform 1 0 30432 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_318
timestamp 1679585382
transform 1 0 31104 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_325
timestamp 1679585382
transform 1 0 31776 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_332
timestamp 1679585382
transform 1 0 32448 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_339
timestamp 1677583704
transform 1 0 33120 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_350
timestamp 1679585382
transform 1 0 34176 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_357
timestamp 1679585382
transform 1 0 34848 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_364
timestamp 1679585382
transform 1 0 35520 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_371
timestamp 1679585382
transform 1 0 36192 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_23_378
timestamp 1677583258
transform 1 0 36864 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_406
timestamp 1679585382
transform 1 0 39552 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_413
timestamp 1679581501
transform 1 0 40224 0 -1 18900
box -48 -56 432 834
use sg13g2_decap_8  FILLER_23_444
timestamp 1679585382
transform 1 0 43200 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_451
timestamp 1679585382
transform 1 0 43872 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_458
timestamp 1679585382
transform 1 0 44544 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_465
timestamp 1679585382
transform 1 0 45216 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_472
timestamp 1679585382
transform 1 0 45888 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_479
timestamp 1679585382
transform 1 0 46560 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_486
timestamp 1679585382
transform 1 0 47232 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_493
timestamp 1679585382
transform 1 0 47904 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_23_500
timestamp 1677583258
transform 1 0 48576 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_537
timestamp 1679585382
transform 1 0 52128 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_544
timestamp 1679585382
transform 1 0 52800 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_551
timestamp 1679585382
transform 1 0 53472 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_558
timestamp 1679585382
transform 1 0 54144 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_565
timestamp 1677583704
transform 1 0 54816 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_567
timestamp 1677583258
transform 1 0 55008 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_572
timestamp 1679585382
transform 1 0 55488 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_579
timestamp 1679585382
transform 1 0 56160 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_586
timestamp 1679585382
transform 1 0 56832 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_593
timestamp 1679585382
transform 1 0 57504 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_600
timestamp 1679585382
transform 1 0 58176 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_607
timestamp 1679585382
transform 1 0 58848 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_614
timestamp 1679585382
transform 1 0 59520 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_621
timestamp 1679585382
transform 1 0 60192 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_628
timestamp 1679585382
transform 1 0 60864 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_635
timestamp 1679585382
transform 1 0 61536 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_642
timestamp 1679585382
transform 1 0 62208 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_649
timestamp 1679585382
transform 1 0 62880 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_656
timestamp 1679585382
transform 1 0 63552 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_663
timestamp 1679585382
transform 1 0 64224 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_670
timestamp 1679585382
transform 1 0 64896 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_677
timestamp 1679585382
transform 1 0 65568 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_684
timestamp 1679585382
transform 1 0 66240 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_691
timestamp 1679585382
transform 1 0 66912 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_698
timestamp 1679585382
transform 1 0 67584 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_705
timestamp 1679585382
transform 1 0 68256 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_712
timestamp 1679585382
transform 1 0 68928 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_719
timestamp 1679585382
transform 1 0 69600 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_726
timestamp 1679585382
transform 1 0 70272 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_733
timestamp 1679585382
transform 1 0 70944 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_740
timestamp 1679585382
transform 1 0 71616 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_747
timestamp 1679585382
transform 1 0 72288 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_754
timestamp 1679585382
transform 1 0 72960 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_761
timestamp 1679585382
transform 1 0 73632 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_768
timestamp 1679585382
transform 1 0 74304 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_775
timestamp 1679585382
transform 1 0 74976 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_782
timestamp 1679585382
transform 1 0 75648 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_789
timestamp 1679585382
transform 1 0 76320 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_796
timestamp 1679585382
transform 1 0 76992 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_803
timestamp 1679585382
transform 1 0 77664 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_810
timestamp 1679585382
transform 1 0 78336 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_817
timestamp 1679585382
transform 1 0 79008 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_824
timestamp 1679585382
transform 1 0 79680 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_831
timestamp 1679585382
transform 1 0 80352 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_838
timestamp 1679585382
transform 1 0 81024 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_845
timestamp 1679585382
transform 1 0 81696 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_852
timestamp 1679585382
transform 1 0 82368 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_859
timestamp 1679585382
transform 1 0 83040 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_866
timestamp 1679585382
transform 1 0 83712 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_873
timestamp 1679585382
transform 1 0 84384 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_880
timestamp 1679585382
transform 1 0 85056 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_887
timestamp 1679585382
transform 1 0 85728 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_894
timestamp 1679585382
transform 1 0 86400 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_901
timestamp 1679585382
transform 1 0 87072 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_908
timestamp 1679585382
transform 1 0 87744 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_915
timestamp 1679585382
transform 1 0 88416 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_922
timestamp 1679585382
transform 1 0 89088 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_929
timestamp 1679585382
transform 1 0 89760 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_936
timestamp 1679585382
transform 1 0 90432 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_943
timestamp 1679585382
transform 1 0 91104 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_950
timestamp 1679585382
transform 1 0 91776 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_957
timestamp 1679585382
transform 1 0 92448 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_964
timestamp 1679585382
transform 1 0 93120 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_971
timestamp 1679585382
transform 1 0 93792 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_978
timestamp 1679585382
transform 1 0 94464 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_985
timestamp 1679585382
transform 1 0 95136 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_992
timestamp 1679585382
transform 1 0 95808 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_999
timestamp 1679585382
transform 1 0 96480 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1006
timestamp 1679585382
transform 1 0 97152 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1013
timestamp 1679585382
transform 1 0 97824 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1020
timestamp 1679585382
transform 1 0 98496 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_1027
timestamp 1677583704
transform 1 0 99168 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_4
timestamp 1679585382
transform 1 0 960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_11
timestamp 1679585382
transform 1 0 1632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_18
timestamp 1679581501
transform 1 0 2304 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_22
timestamp 1677583704
transform 1 0 2688 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_50
timestamp 1679585382
transform 1 0 5376 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_57
timestamp 1679585382
transform 1 0 6048 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_64
timestamp 1679581501
transform 1 0 6720 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_68
timestamp 1677583704
transform 1 0 7104 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_97
timestamp 1679585382
transform 1 0 9888 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_104
timestamp 1679585382
transform 1 0 10560 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_111
timestamp 1679585382
transform 1 0 11232 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_118
timestamp 1677583704
transform 1 0 11904 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_129
timestamp 1679585382
transform 1 0 12960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_136
timestamp 1679585382
transform 1 0 13632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_143
timestamp 1679585382
transform 1 0 14304 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_150
timestamp 1679585382
transform 1 0 14976 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_157
timestamp 1679585382
transform 1 0 15648 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_164
timestamp 1679585382
transform 1 0 16320 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_171
timestamp 1679585382
transform 1 0 16992 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_178
timestamp 1679585382
transform 1 0 17664 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_185
timestamp 1679585382
transform 1 0 18336 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_192
timestamp 1679585382
transform 1 0 19008 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_199
timestamp 1677583704
transform 1 0 19680 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_229
timestamp 1679585382
transform 1 0 22560 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_236
timestamp 1679585382
transform 1 0 23232 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_243
timestamp 1679585382
transform 1 0 23904 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_250
timestamp 1679585382
transform 1 0 24576 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_257
timestamp 1679585382
transform 1 0 25248 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_264
timestamp 1679585382
transform 1 0 25920 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_271
timestamp 1679585382
transform 1 0 26592 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_278
timestamp 1679585382
transform 1 0 27264 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_285
timestamp 1679585382
transform 1 0 27936 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_292
timestamp 1677583704
transform 1 0 28608 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_302
timestamp 1679585382
transform 1 0 29568 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_309
timestamp 1679585382
transform 1 0 30240 0 1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_24_316
timestamp 1677583258
transform 1 0 30912 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_344
timestamp 1679585382
transform 1 0 33600 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_351
timestamp 1679581501
transform 1 0 34272 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_355
timestamp 1677583258
transform 1 0 34656 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_369
timestamp 1679585382
transform 1 0 36000 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_376
timestamp 1679585382
transform 1 0 36672 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_383
timestamp 1679585382
transform 1 0 37344 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_390
timestamp 1679585382
transform 1 0 38016 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_397
timestamp 1679585382
transform 1 0 38688 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_404
timestamp 1679585382
transform 1 0 39360 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_411
timestamp 1679585382
transform 1 0 40032 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_418
timestamp 1679585382
transform 1 0 40704 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_425
timestamp 1679585382
transform 1 0 41376 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_432
timestamp 1679585382
transform 1 0 42048 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_439
timestamp 1679585382
transform 1 0 42720 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_446
timestamp 1679585382
transform 1 0 43392 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_453
timestamp 1679585382
transform 1 0 44064 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_460
timestamp 1679585382
transform 1 0 44736 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_467
timestamp 1679585382
transform 1 0 45408 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_474
timestamp 1679585382
transform 1 0 46080 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_481
timestamp 1679585382
transform 1 0 46752 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_488
timestamp 1679585382
transform 1 0 47424 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_495
timestamp 1679585382
transform 1 0 48096 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_502
timestamp 1679585382
transform 1 0 48768 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_509
timestamp 1679585382
transform 1 0 49440 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_516
timestamp 1679585382
transform 1 0 50112 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_523
timestamp 1679585382
transform 1 0 50784 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_530
timestamp 1679585382
transform 1 0 51456 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_537
timestamp 1679585382
transform 1 0 52128 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_544
timestamp 1679585382
transform 1 0 52800 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_560
timestamp 1679585382
transform 1 0 54336 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_567
timestamp 1677583704
transform 1 0 55008 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_600
timestamp 1679585382
transform 1 0 58176 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_607
timestamp 1679585382
transform 1 0 58848 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_614
timestamp 1679585382
transform 1 0 59520 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_621
timestamp 1679585382
transform 1 0 60192 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_628
timestamp 1679585382
transform 1 0 60864 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_635
timestamp 1679585382
transform 1 0 61536 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_642
timestamp 1679585382
transform 1 0 62208 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_649
timestamp 1679585382
transform 1 0 62880 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_656
timestamp 1679585382
transform 1 0 63552 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_663
timestamp 1679585382
transform 1 0 64224 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_670
timestamp 1679585382
transform 1 0 64896 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_677
timestamp 1679585382
transform 1 0 65568 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_684
timestamp 1679585382
transform 1 0 66240 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_691
timestamp 1679585382
transform 1 0 66912 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_698
timestamp 1679585382
transform 1 0 67584 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_705
timestamp 1679585382
transform 1 0 68256 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_712
timestamp 1679585382
transform 1 0 68928 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_719
timestamp 1679585382
transform 1 0 69600 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_726
timestamp 1679585382
transform 1 0 70272 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_733
timestamp 1679585382
transform 1 0 70944 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_740
timestamp 1679585382
transform 1 0 71616 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_747
timestamp 1679585382
transform 1 0 72288 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_754
timestamp 1679585382
transform 1 0 72960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_761
timestamp 1679585382
transform 1 0 73632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_768
timestamp 1679585382
transform 1 0 74304 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_775
timestamp 1679585382
transform 1 0 74976 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_782
timestamp 1679585382
transform 1 0 75648 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_789
timestamp 1679585382
transform 1 0 76320 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_796
timestamp 1679585382
transform 1 0 76992 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_803
timestamp 1679585382
transform 1 0 77664 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_810
timestamp 1679585382
transform 1 0 78336 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_817
timestamp 1679585382
transform 1 0 79008 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_824
timestamp 1679585382
transform 1 0 79680 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_831
timestamp 1679585382
transform 1 0 80352 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_838
timestamp 1679585382
transform 1 0 81024 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_845
timestamp 1679585382
transform 1 0 81696 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_852
timestamp 1679585382
transform 1 0 82368 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_859
timestamp 1679585382
transform 1 0 83040 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_866
timestamp 1679585382
transform 1 0 83712 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_873
timestamp 1679585382
transform 1 0 84384 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_880
timestamp 1679585382
transform 1 0 85056 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_887
timestamp 1679585382
transform 1 0 85728 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_894
timestamp 1679585382
transform 1 0 86400 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_901
timestamp 1679585382
transform 1 0 87072 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_908
timestamp 1679585382
transform 1 0 87744 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_915
timestamp 1679585382
transform 1 0 88416 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_922
timestamp 1679585382
transform 1 0 89088 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_929
timestamp 1679585382
transform 1 0 89760 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_936
timestamp 1679585382
transform 1 0 90432 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_943
timestamp 1679585382
transform 1 0 91104 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_950
timestamp 1679585382
transform 1 0 91776 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_957
timestamp 1679585382
transform 1 0 92448 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_964
timestamp 1679585382
transform 1 0 93120 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_971
timestamp 1679585382
transform 1 0 93792 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_978
timestamp 1679585382
transform 1 0 94464 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_985
timestamp 1679585382
transform 1 0 95136 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_992
timestamp 1679585382
transform 1 0 95808 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_999
timestamp 1679585382
transform 1 0 96480 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1006
timestamp 1679585382
transform 1 0 97152 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1013
timestamp 1679585382
transform 1 0 97824 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1020
timestamp 1679585382
transform 1 0 98496 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_1027
timestamp 1677583704
transform 1 0 99168 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_4
timestamp 1679585382
transform 1 0 960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_11
timestamp 1679585382
transform 1 0 1632 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_18
timestamp 1679585382
transform 1 0 2304 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_25
timestamp 1679585382
transform 1 0 2976 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_32
timestamp 1679585382
transform 1 0 3648 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_25_39
timestamp 1677583258
transform 1 0 4320 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_52
timestamp 1679585382
transform 1 0 5568 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_59
timestamp 1679585382
transform 1 0 6240 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_66
timestamp 1679585382
transform 1 0 6912 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_73
timestamp 1679585382
transform 1 0 7584 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_80
timestamp 1679585382
transform 1 0 8256 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_87
timestamp 1679585382
transform 1 0 8928 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_94
timestamp 1679585382
transform 1 0 9600 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_101
timestamp 1679585382
transform 1 0 10272 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_108
timestamp 1679585382
transform 1 0 10944 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_115
timestamp 1677583704
transform 1 0 11616 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_125
timestamp 1679585382
transform 1 0 12576 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_132
timestamp 1679585382
transform 1 0 13248 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_139
timestamp 1679585382
transform 1 0 13920 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_146
timestamp 1679585382
transform 1 0 14592 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_153
timestamp 1679585382
transform 1 0 15264 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_160
timestamp 1679585382
transform 1 0 15936 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_167
timestamp 1679585382
transform 1 0 16608 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_174
timestamp 1679585382
transform 1 0 17280 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_181
timestamp 1679585382
transform 1 0 17952 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_188
timestamp 1679585382
transform 1 0 18624 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_195
timestamp 1679581501
transform 1 0 19296 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_25_240
timestamp 1679585382
transform 1 0 23616 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_247
timestamp 1679585382
transform 1 0 24288 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_254
timestamp 1679585382
transform 1 0 24960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_261
timestamp 1679585382
transform 1 0 25632 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_268
timestamp 1679585382
transform 1 0 26304 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_275
timestamp 1679585382
transform 1 0 26976 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_282
timestamp 1677583704
transform 1 0 27648 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_292
timestamp 1679585382
transform 1 0 28608 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_299
timestamp 1679585382
transform 1 0 29280 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_306
timestamp 1679585382
transform 1 0 29952 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_313
timestamp 1679581501
transform 1 0 30624 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_25_343
timestamp 1679585382
transform 1 0 33504 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_350
timestamp 1679585382
transform 1 0 34176 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_357
timestamp 1679585382
transform 1 0 34848 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_364
timestamp 1679585382
transform 1 0 35520 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_371
timestamp 1679585382
transform 1 0 36192 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_378
timestamp 1679585382
transform 1 0 36864 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_385
timestamp 1679585382
transform 1 0 37536 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_392
timestamp 1679581501
transform 1 0 38208 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_4  FILLER_25_413
timestamp 1679581501
transform 1 0 40224 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_25_417
timestamp 1677583258
transform 1 0 40608 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_427
timestamp 1679585382
transform 1 0 41568 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_434
timestamp 1679585382
transform 1 0 42240 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_441
timestamp 1679585382
transform 1 0 42912 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_448
timestamp 1679585382
transform 1 0 43584 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_455
timestamp 1679581501
transform 1 0 44256 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_25_459
timestamp 1677583258
transform 1 0 44640 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_464
timestamp 1679585382
transform 1 0 45120 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_471
timestamp 1677583704
transform 1 0 45792 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_482
timestamp 1679585382
transform 1 0 46848 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_489
timestamp 1679585382
transform 1 0 47520 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_496
timestamp 1679585382
transform 1 0 48192 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_503
timestamp 1679585382
transform 1 0 48864 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_510
timestamp 1679585382
transform 1 0 49536 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_517
timestamp 1679585382
transform 1 0 50208 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_524
timestamp 1679585382
transform 1 0 50880 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_531
timestamp 1679581501
transform 1 0 51552 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_25_535
timestamp 1677583258
transform 1 0 51936 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_563
timestamp 1679585382
transform 1 0 54624 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_570
timestamp 1679585382
transform 1 0 55296 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_577
timestamp 1679585382
transform 1 0 55968 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_25_584
timestamp 1677583258
transform 1 0 56640 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_594
timestamp 1679585382
transform 1 0 57600 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_601
timestamp 1679585382
transform 1 0 58272 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_608
timestamp 1679585382
transform 1 0 58944 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_615
timestamp 1679585382
transform 1 0 59616 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_622
timestamp 1679585382
transform 1 0 60288 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_629
timestamp 1679585382
transform 1 0 60960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_636
timestamp 1679585382
transform 1 0 61632 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_643
timestamp 1679585382
transform 1 0 62304 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_650
timestamp 1679585382
transform 1 0 62976 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_657
timestamp 1679585382
transform 1 0 63648 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_664
timestamp 1679585382
transform 1 0 64320 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_671
timestamp 1679585382
transform 1 0 64992 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_678
timestamp 1679585382
transform 1 0 65664 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_685
timestamp 1679585382
transform 1 0 66336 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_692
timestamp 1679585382
transform 1 0 67008 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_699
timestamp 1679585382
transform 1 0 67680 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_706
timestamp 1679585382
transform 1 0 68352 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_713
timestamp 1679585382
transform 1 0 69024 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_720
timestamp 1679585382
transform 1 0 69696 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_727
timestamp 1679585382
transform 1 0 70368 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_734
timestamp 1679585382
transform 1 0 71040 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_741
timestamp 1679585382
transform 1 0 71712 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_748
timestamp 1679585382
transform 1 0 72384 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_755
timestamp 1679585382
transform 1 0 73056 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_762
timestamp 1679585382
transform 1 0 73728 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_769
timestamp 1679585382
transform 1 0 74400 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_776
timestamp 1679585382
transform 1 0 75072 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_783
timestamp 1679585382
transform 1 0 75744 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_790
timestamp 1679585382
transform 1 0 76416 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_797
timestamp 1679585382
transform 1 0 77088 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_804
timestamp 1679585382
transform 1 0 77760 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_811
timestamp 1679585382
transform 1 0 78432 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_818
timestamp 1679585382
transform 1 0 79104 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_825
timestamp 1679585382
transform 1 0 79776 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_832
timestamp 1679585382
transform 1 0 80448 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_839
timestamp 1679585382
transform 1 0 81120 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_846
timestamp 1679585382
transform 1 0 81792 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_853
timestamp 1679585382
transform 1 0 82464 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_860
timestamp 1679585382
transform 1 0 83136 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_867
timestamp 1679585382
transform 1 0 83808 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_874
timestamp 1679585382
transform 1 0 84480 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_881
timestamp 1679585382
transform 1 0 85152 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_888
timestamp 1679585382
transform 1 0 85824 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_895
timestamp 1679585382
transform 1 0 86496 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_902
timestamp 1679585382
transform 1 0 87168 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_909
timestamp 1679585382
transform 1 0 87840 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_916
timestamp 1679585382
transform 1 0 88512 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_923
timestamp 1679585382
transform 1 0 89184 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_930
timestamp 1679585382
transform 1 0 89856 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_937
timestamp 1679585382
transform 1 0 90528 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_944
timestamp 1679585382
transform 1 0 91200 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_951
timestamp 1679585382
transform 1 0 91872 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_958
timestamp 1679585382
transform 1 0 92544 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_965
timestamp 1679585382
transform 1 0 93216 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_972
timestamp 1679585382
transform 1 0 93888 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_979
timestamp 1679585382
transform 1 0 94560 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_986
timestamp 1679585382
transform 1 0 95232 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_993
timestamp 1679585382
transform 1 0 95904 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1000
timestamp 1679585382
transform 1 0 96576 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1007
timestamp 1679585382
transform 1 0 97248 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1014
timestamp 1679585382
transform 1 0 97920 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1021
timestamp 1679585382
transform 1 0 98592 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_25_1028
timestamp 1677583258
transform 1 0 99264 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_4
timestamp 1679585382
transform 1 0 960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_11
timestamp 1679585382
transform 1 0 1632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_18
timestamp 1679585382
transform 1 0 2304 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_25
timestamp 1679585382
transform 1 0 2976 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_32
timestamp 1679585382
transform 1 0 3648 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_39
timestamp 1679585382
transform 1 0 4320 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_46
timestamp 1679581501
transform 1 0 4992 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_50
timestamp 1677583258
transform 1 0 5376 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_56
timestamp 1679585382
transform 1 0 5952 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_63
timestamp 1679585382
transform 1 0 6624 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_70
timestamp 1679585382
transform 1 0 7296 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_77
timestamp 1679585382
transform 1 0 7968 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_84
timestamp 1679585382
transform 1 0 8640 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_91
timestamp 1679585382
transform 1 0 9312 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_98
timestamp 1679585382
transform 1 0 9984 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_105
timestamp 1679585382
transform 1 0 10656 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_124
timestamp 1677583704
transform 1 0 12480 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_162
timestamp 1679585382
transform 1 0 16128 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_169
timestamp 1679585382
transform 1 0 16800 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_176
timestamp 1679585382
transform 1 0 17472 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_183
timestamp 1679585382
transform 1 0 18144 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_190
timestamp 1679585382
transform 1 0 18816 0 1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_210
timestamp 1677583258
transform 1 0 20736 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_224
timestamp 1679585382
transform 1 0 22080 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_231
timestamp 1679585382
transform 1 0 22752 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_238
timestamp 1679585382
transform 1 0 23424 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_245
timestamp 1679585382
transform 1 0 24096 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_252
timestamp 1679585382
transform 1 0 24768 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_259
timestamp 1679585382
transform 1 0 25440 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_266
timestamp 1677583704
transform 1 0 26112 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_268
timestamp 1677583258
transform 1 0 26304 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_277
timestamp 1679585382
transform 1 0 27168 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_284
timestamp 1679585382
transform 1 0 27840 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_291
timestamp 1679585382
transform 1 0 28512 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_298
timestamp 1679585382
transform 1 0 29184 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_305
timestamp 1679585382
transform 1 0 29856 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_312
timestamp 1679585382
transform 1 0 30528 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_319
timestamp 1679585382
transform 1 0 31200 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_326
timestamp 1679585382
transform 1 0 31872 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_333
timestamp 1679585382
transform 1 0 32544 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_340
timestamp 1679585382
transform 1 0 33216 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_347
timestamp 1679585382
transform 1 0 33888 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_354
timestamp 1679585382
transform 1 0 34560 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_361
timestamp 1679585382
transform 1 0 35232 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_368
timestamp 1679585382
transform 1 0 35904 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_375
timestamp 1679585382
transform 1 0 36576 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_382
timestamp 1679585382
transform 1 0 37248 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_389
timestamp 1679585382
transform 1 0 37920 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_396
timestamp 1679585382
transform 1 0 38592 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_403
timestamp 1679581501
transform 1 0 39264 0 1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_26_419
timestamp 1679585382
transform 1 0 40800 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_426
timestamp 1679585382
transform 1 0 41472 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_433
timestamp 1679585382
transform 1 0 42144 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_440
timestamp 1679585382
transform 1 0 42816 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_447
timestamp 1679585382
transform 1 0 43488 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_454
timestamp 1677583704
transform 1 0 44160 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_483
timestamp 1679585382
transform 1 0 46944 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_490
timestamp 1679585382
transform 1 0 47616 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_497
timestamp 1679585382
transform 1 0 48288 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_504
timestamp 1679585382
transform 1 0 48960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_511
timestamp 1679585382
transform 1 0 49632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_518
timestamp 1679585382
transform 1 0 50304 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_525
timestamp 1679585382
transform 1 0 50976 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_532
timestamp 1679585382
transform 1 0 51648 0 1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_539
timestamp 1677583258
transform 1 0 52320 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_544
timestamp 1679585382
transform 1 0 52800 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_551
timestamp 1679585382
transform 1 0 53472 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_558
timestamp 1679585382
transform 1 0 54144 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_565
timestamp 1679585382
transform 1 0 54816 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_572
timestamp 1679585382
transform 1 0 55488 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_579
timestamp 1679585382
transform 1 0 56160 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_586
timestamp 1679585382
transform 1 0 56832 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_593
timestamp 1679585382
transform 1 0 57504 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_600
timestamp 1679585382
transform 1 0 58176 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_607
timestamp 1679585382
transform 1 0 58848 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_614
timestamp 1679585382
transform 1 0 59520 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_621
timestamp 1679585382
transform 1 0 60192 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_628
timestamp 1679585382
transform 1 0 60864 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_635
timestamp 1679585382
transform 1 0 61536 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_642
timestamp 1679585382
transform 1 0 62208 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_649
timestamp 1679585382
transform 1 0 62880 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_656
timestamp 1679585382
transform 1 0 63552 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_663
timestamp 1679585382
transform 1 0 64224 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_670
timestamp 1679585382
transform 1 0 64896 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_677
timestamp 1679585382
transform 1 0 65568 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_684
timestamp 1679585382
transform 1 0 66240 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_691
timestamp 1679585382
transform 1 0 66912 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_698
timestamp 1679585382
transform 1 0 67584 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_705
timestamp 1679585382
transform 1 0 68256 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_712
timestamp 1679585382
transform 1 0 68928 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_719
timestamp 1679585382
transform 1 0 69600 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_726
timestamp 1679585382
transform 1 0 70272 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_733
timestamp 1679585382
transform 1 0 70944 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_740
timestamp 1679585382
transform 1 0 71616 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_747
timestamp 1679585382
transform 1 0 72288 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_754
timestamp 1679585382
transform 1 0 72960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_761
timestamp 1679585382
transform 1 0 73632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_768
timestamp 1679585382
transform 1 0 74304 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_775
timestamp 1679585382
transform 1 0 74976 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_782
timestamp 1679585382
transform 1 0 75648 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_789
timestamp 1679585382
transform 1 0 76320 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_796
timestamp 1679585382
transform 1 0 76992 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_803
timestamp 1679585382
transform 1 0 77664 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_810
timestamp 1679585382
transform 1 0 78336 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_817
timestamp 1679585382
transform 1 0 79008 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_824
timestamp 1679585382
transform 1 0 79680 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_831
timestamp 1679585382
transform 1 0 80352 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_838
timestamp 1679585382
transform 1 0 81024 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_845
timestamp 1679585382
transform 1 0 81696 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_852
timestamp 1679585382
transform 1 0 82368 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_859
timestamp 1679585382
transform 1 0 83040 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_866
timestamp 1679585382
transform 1 0 83712 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_873
timestamp 1679585382
transform 1 0 84384 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_880
timestamp 1679585382
transform 1 0 85056 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_887
timestamp 1679585382
transform 1 0 85728 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_894
timestamp 1679585382
transform 1 0 86400 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_901
timestamp 1679585382
transform 1 0 87072 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_908
timestamp 1679585382
transform 1 0 87744 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_915
timestamp 1679585382
transform 1 0 88416 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_922
timestamp 1679585382
transform 1 0 89088 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_929
timestamp 1679585382
transform 1 0 89760 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_936
timestamp 1679585382
transform 1 0 90432 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_943
timestamp 1679585382
transform 1 0 91104 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_950
timestamp 1679585382
transform 1 0 91776 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_957
timestamp 1679585382
transform 1 0 92448 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_964
timestamp 1679585382
transform 1 0 93120 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_971
timestamp 1679585382
transform 1 0 93792 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_978
timestamp 1679585382
transform 1 0 94464 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_985
timestamp 1679585382
transform 1 0 95136 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_992
timestamp 1679585382
transform 1 0 95808 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_999
timestamp 1679585382
transform 1 0 96480 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1006
timestamp 1679585382
transform 1 0 97152 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1013
timestamp 1679585382
transform 1 0 97824 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1020
timestamp 1679585382
transform 1 0 98496 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_1027
timestamp 1677583704
transform 1 0 99168 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1679585382
transform 1 0 576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_7
timestamp 1679585382
transform 1 0 1248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_14
timestamp 1679585382
transform 1 0 1920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_21
timestamp 1679585382
transform 1 0 2592 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_28
timestamp 1679585382
transform 1 0 3264 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_35
timestamp 1679581501
transform 1 0 3936 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_39
timestamp 1677583258
transform 1 0 4320 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_44
timestamp 1679585382
transform 1 0 4800 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_51
timestamp 1679585382
transform 1 0 5472 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_58
timestamp 1679585382
transform 1 0 6144 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_65
timestamp 1679585382
transform 1 0 6816 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_72
timestamp 1679581501
transform 1 0 7488 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_76
timestamp 1677583258
transform 1 0 7872 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_27_104
timestamp 1679581501
transform 1 0 10560 0 -1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_27_117
timestamp 1679585382
transform 1 0 11808 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_124
timestamp 1679581501
transform 1 0 12480 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_128
timestamp 1677583258
transform 1 0 12864 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_138
timestamp 1679585382
transform 1 0 13824 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_1  FILLER_27_145
timestamp 1677583258
transform 1 0 14496 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_159
timestamp 1679585382
transform 1 0 15840 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_166
timestamp 1679585382
transform 1 0 16512 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_173
timestamp 1679585382
transform 1 0 17184 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_180
timestamp 1679585382
transform 1 0 17856 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_187
timestamp 1679585382
transform 1 0 18528 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_194
timestamp 1679585382
transform 1 0 19200 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_201
timestamp 1679581501
transform 1 0 19872 0 -1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_27_214
timestamp 1679585382
transform 1 0 21120 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_221
timestamp 1679585382
transform 1 0 21792 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_228
timestamp 1679585382
transform 1 0 22464 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_235
timestamp 1679585382
transform 1 0 23136 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_242
timestamp 1679585382
transform 1 0 23808 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_249
timestamp 1679585382
transform 1 0 24480 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_256
timestamp 1679581501
transform 1 0 25152 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_260
timestamp 1677583704
transform 1 0 25536 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_298
timestamp 1679585382
transform 1 0 29184 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_305
timestamp 1679585382
transform 1 0 29856 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_312
timestamp 1679581501
transform 1 0 30528 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_316
timestamp 1677583704
transform 1 0 30912 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_358
timestamp 1679585382
transform 1 0 34944 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_365
timestamp 1679581501
transform 1 0 35616 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_369
timestamp 1677583704
transform 1 0 36000 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_398
timestamp 1677583258
transform 1 0 38784 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_408
timestamp 1679585382
transform 1 0 39744 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_415
timestamp 1679585382
transform 1 0 40416 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_422
timestamp 1679585382
transform 1 0 41088 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_429
timestamp 1679585382
transform 1 0 41760 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_436
timestamp 1679581501
transform 1 0 42432 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_440
timestamp 1677583704
transform 1 0 42816 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_455
timestamp 1677583258
transform 1 0 44256 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_483
timestamp 1679585382
transform 1 0 46944 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_490
timestamp 1679585382
transform 1 0 47616 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_497
timestamp 1679585382
transform 1 0 48288 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_504
timestamp 1679585382
transform 1 0 48960 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_511
timestamp 1679585382
transform 1 0 49632 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_518
timestamp 1679585382
transform 1 0 50304 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_525
timestamp 1679585382
transform 1 0 50976 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_532
timestamp 1679585382
transform 1 0 51648 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_539
timestamp 1679585382
transform 1 0 52320 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_546
timestamp 1679585382
transform 1 0 52992 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_553
timestamp 1679585382
transform 1 0 53664 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_560
timestamp 1679585382
transform 1 0 54336 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_567
timestamp 1679585382
transform 1 0 55008 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_574
timestamp 1679585382
transform 1 0 55680 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_581
timestamp 1679585382
transform 1 0 56352 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_588
timestamp 1679585382
transform 1 0 57024 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_595
timestamp 1679585382
transform 1 0 57696 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_602
timestamp 1679585382
transform 1 0 58368 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_609
timestamp 1679585382
transform 1 0 59040 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_616
timestamp 1679585382
transform 1 0 59712 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_623
timestamp 1679585382
transform 1 0 60384 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_630
timestamp 1679585382
transform 1 0 61056 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_637
timestamp 1679585382
transform 1 0 61728 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_644
timestamp 1679585382
transform 1 0 62400 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_651
timestamp 1679585382
transform 1 0 63072 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_658
timestamp 1679585382
transform 1 0 63744 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_665
timestamp 1679585382
transform 1 0 64416 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_672
timestamp 1679585382
transform 1 0 65088 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_679
timestamp 1679585382
transform 1 0 65760 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_686
timestamp 1679585382
transform 1 0 66432 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_693
timestamp 1679585382
transform 1 0 67104 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_700
timestamp 1679585382
transform 1 0 67776 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_707
timestamp 1679585382
transform 1 0 68448 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_714
timestamp 1679585382
transform 1 0 69120 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_721
timestamp 1679585382
transform 1 0 69792 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_728
timestamp 1679585382
transform 1 0 70464 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_735
timestamp 1679585382
transform 1 0 71136 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_742
timestamp 1679585382
transform 1 0 71808 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_749
timestamp 1679585382
transform 1 0 72480 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_756
timestamp 1679585382
transform 1 0 73152 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_763
timestamp 1679585382
transform 1 0 73824 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_770
timestamp 1679585382
transform 1 0 74496 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_777
timestamp 1679585382
transform 1 0 75168 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_784
timestamp 1679585382
transform 1 0 75840 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_791
timestamp 1679585382
transform 1 0 76512 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_798
timestamp 1679585382
transform 1 0 77184 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_805
timestamp 1679585382
transform 1 0 77856 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_812
timestamp 1679585382
transform 1 0 78528 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_819
timestamp 1679585382
transform 1 0 79200 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_826
timestamp 1679585382
transform 1 0 79872 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_833
timestamp 1679585382
transform 1 0 80544 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_840
timestamp 1679585382
transform 1 0 81216 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_847
timestamp 1679585382
transform 1 0 81888 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_854
timestamp 1679585382
transform 1 0 82560 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_861
timestamp 1679585382
transform 1 0 83232 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_868
timestamp 1679585382
transform 1 0 83904 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_875
timestamp 1679585382
transform 1 0 84576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_882
timestamp 1679585382
transform 1 0 85248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_889
timestamp 1679585382
transform 1 0 85920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_896
timestamp 1679585382
transform 1 0 86592 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_903
timestamp 1679585382
transform 1 0 87264 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_910
timestamp 1679585382
transform 1 0 87936 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_917
timestamp 1679585382
transform 1 0 88608 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_924
timestamp 1679585382
transform 1 0 89280 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_931
timestamp 1679585382
transform 1 0 89952 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_938
timestamp 1679585382
transform 1 0 90624 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_945
timestamp 1679585382
transform 1 0 91296 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_952
timestamp 1679585382
transform 1 0 91968 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_959
timestamp 1679585382
transform 1 0 92640 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_966
timestamp 1679585382
transform 1 0 93312 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_973
timestamp 1679585382
transform 1 0 93984 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_980
timestamp 1679585382
transform 1 0 94656 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_987
timestamp 1679585382
transform 1 0 95328 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_994
timestamp 1679585382
transform 1 0 96000 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1001
timestamp 1679585382
transform 1 0 96672 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1008
timestamp 1679585382
transform 1 0 97344 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1015
timestamp 1679585382
transform 1 0 98016 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1022
timestamp 1679585382
transform 1 0 98688 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_4
timestamp 1677583704
transform 1 0 960 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_60
timestamp 1679585382
transform 1 0 6336 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_67
timestamp 1679585382
transform 1 0 7008 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_74
timestamp 1679585382
transform 1 0 7680 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_81
timestamp 1679581501
transform 1 0 8352 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_85
timestamp 1677583704
transform 1 0 8736 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_100
timestamp 1679585382
transform 1 0 10176 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_107
timestamp 1679585382
transform 1 0 10848 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_114
timestamp 1679585382
transform 1 0 11520 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_121
timestamp 1679585382
transform 1 0 12192 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_128
timestamp 1679585382
transform 1 0 12864 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_162
timestamp 1679585382
transform 1 0 16128 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_169
timestamp 1679585382
transform 1 0 16800 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_176
timestamp 1679585382
transform 1 0 17472 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_183
timestamp 1679585382
transform 1 0 18144 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_190
timestamp 1679585382
transform 1 0 18816 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_197
timestamp 1679585382
transform 1 0 19488 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_204
timestamp 1679585382
transform 1 0 20160 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_211
timestamp 1679581501
transform 1 0 20832 0 1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_28_224
timestamp 1679585382
transform 1 0 22080 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_231
timestamp 1679585382
transform 1 0 22752 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_238
timestamp 1679585382
transform 1 0 23424 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_245
timestamp 1679585382
transform 1 0 24096 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_252
timestamp 1679585382
transform 1 0 24768 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_259
timestamp 1677583704
transform 1 0 25440 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_288
timestamp 1679585382
transform 1 0 28224 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_295
timestamp 1679585382
transform 1 0 28896 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_302
timestamp 1679585382
transform 1 0 29568 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_309
timestamp 1679585382
transform 1 0 30240 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_316
timestamp 1679585382
transform 1 0 30912 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_323
timestamp 1679585382
transform 1 0 31584 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_330
timestamp 1679585382
transform 1 0 32256 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_337
timestamp 1677583704
transform 1 0 32928 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_339
timestamp 1677583258
transform 1 0 33120 0 1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_28_344
timestamp 1679581501
transform 1 0 33600 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_348
timestamp 1677583704
transform 1 0 33984 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_364
timestamp 1679585382
transform 1 0 35520 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_371
timestamp 1679585382
transform 1 0 36192 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_378
timestamp 1679585382
transform 1 0 36864 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_385
timestamp 1679585382
transform 1 0 37536 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_392
timestamp 1679585382
transform 1 0 38208 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_399
timestamp 1679585382
transform 1 0 38880 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_406
timestamp 1679585382
transform 1 0 39552 0 1 21924
box -48 -56 720 834
use sg13g2_fill_1  FILLER_28_413
timestamp 1677583258
transform 1 0 40224 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_423
timestamp 1679585382
transform 1 0 41184 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_430
timestamp 1679585382
transform 1 0 41856 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_437
timestamp 1679585382
transform 1 0 42528 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_444
timestamp 1679585382
transform 1 0 43200 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_451
timestamp 1679585382
transform 1 0 43872 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_458
timestamp 1677583704
transform 1 0 44544 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_460
timestamp 1677583258
transform 1 0 44736 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_466
timestamp 1679585382
transform 1 0 45312 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_473
timestamp 1679585382
transform 1 0 45984 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_480
timestamp 1679585382
transform 1 0 46656 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_487
timestamp 1679585382
transform 1 0 47328 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_494
timestamp 1679585382
transform 1 0 48000 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_501
timestamp 1679581501
transform 1 0 48672 0 1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_505
timestamp 1677583258
transform 1 0 49056 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_519
timestamp 1679585382
transform 1 0 50400 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_526
timestamp 1679585382
transform 1 0 51072 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_533
timestamp 1679585382
transform 1 0 51744 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_540
timestamp 1679585382
transform 1 0 52416 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_547
timestamp 1679585382
transform 1 0 53088 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_554
timestamp 1679585382
transform 1 0 53760 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_561
timestamp 1679585382
transform 1 0 54432 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_568
timestamp 1679585382
transform 1 0 55104 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_575
timestamp 1679585382
transform 1 0 55776 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_582
timestamp 1679585382
transform 1 0 56448 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_589
timestamp 1679585382
transform 1 0 57120 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_596
timestamp 1679585382
transform 1 0 57792 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_603
timestamp 1679585382
transform 1 0 58464 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_610
timestamp 1679585382
transform 1 0 59136 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_617
timestamp 1679585382
transform 1 0 59808 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_624
timestamp 1679585382
transform 1 0 60480 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_631
timestamp 1679585382
transform 1 0 61152 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_638
timestamp 1679585382
transform 1 0 61824 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_645
timestamp 1679585382
transform 1 0 62496 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_652
timestamp 1679585382
transform 1 0 63168 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_659
timestamp 1679585382
transform 1 0 63840 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_666
timestamp 1679585382
transform 1 0 64512 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_673
timestamp 1679585382
transform 1 0 65184 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_680
timestamp 1679585382
transform 1 0 65856 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_687
timestamp 1679585382
transform 1 0 66528 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_694
timestamp 1679585382
transform 1 0 67200 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_701
timestamp 1679585382
transform 1 0 67872 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_708
timestamp 1679585382
transform 1 0 68544 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_715
timestamp 1679585382
transform 1 0 69216 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_722
timestamp 1679585382
transform 1 0 69888 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_729
timestamp 1679585382
transform 1 0 70560 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_736
timestamp 1679585382
transform 1 0 71232 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_743
timestamp 1679585382
transform 1 0 71904 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_750
timestamp 1679585382
transform 1 0 72576 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_757
timestamp 1679585382
transform 1 0 73248 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_764
timestamp 1679585382
transform 1 0 73920 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_771
timestamp 1679585382
transform 1 0 74592 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_778
timestamp 1679585382
transform 1 0 75264 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_785
timestamp 1679585382
transform 1 0 75936 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_792
timestamp 1679585382
transform 1 0 76608 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_799
timestamp 1679585382
transform 1 0 77280 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_806
timestamp 1679585382
transform 1 0 77952 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_813
timestamp 1679585382
transform 1 0 78624 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_820
timestamp 1679585382
transform 1 0 79296 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_827
timestamp 1679585382
transform 1 0 79968 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_834
timestamp 1679585382
transform 1 0 80640 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_841
timestamp 1679585382
transform 1 0 81312 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_848
timestamp 1679585382
transform 1 0 81984 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_855
timestamp 1679585382
transform 1 0 82656 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_862
timestamp 1679585382
transform 1 0 83328 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_869
timestamp 1679585382
transform 1 0 84000 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_876
timestamp 1679585382
transform 1 0 84672 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_883
timestamp 1679585382
transform 1 0 85344 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_890
timestamp 1679585382
transform 1 0 86016 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_897
timestamp 1679585382
transform 1 0 86688 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_904
timestamp 1679585382
transform 1 0 87360 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_911
timestamp 1679585382
transform 1 0 88032 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_918
timestamp 1679585382
transform 1 0 88704 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_925
timestamp 1679585382
transform 1 0 89376 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_932
timestamp 1679585382
transform 1 0 90048 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_939
timestamp 1679585382
transform 1 0 90720 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_946
timestamp 1679585382
transform 1 0 91392 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_953
timestamp 1679585382
transform 1 0 92064 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_960
timestamp 1679585382
transform 1 0 92736 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_967
timestamp 1679585382
transform 1 0 93408 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_974
timestamp 1679585382
transform 1 0 94080 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_981
timestamp 1679585382
transform 1 0 94752 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_988
timestamp 1679585382
transform 1 0 95424 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_995
timestamp 1679585382
transform 1 0 96096 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1002
timestamp 1679585382
transform 1 0 96768 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1009
timestamp 1679585382
transform 1 0 97440 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1016
timestamp 1679585382
transform 1 0 98112 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_1023
timestamp 1679581501
transform 1 0 98784 0 1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_28_1027
timestamp 1677583704
transform 1 0 99168 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_0
timestamp 1679585382
transform 1 0 576 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_7
timestamp 1679585382
transform 1 0 1248 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_29_14
timestamp 1677583258
transform 1 0 1920 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_28
timestamp 1679585382
transform 1 0 3264 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_35
timestamp 1677583704
transform 1 0 3936 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_37
timestamp 1677583258
transform 1 0 4128 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_42
timestamp 1679585382
transform 1 0 4608 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_29_49
timestamp 1677583258
transform 1 0 5280 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_59
timestamp 1679585382
transform 1 0 6240 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_66
timestamp 1679585382
transform 1 0 6912 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_73
timestamp 1679585382
transform 1 0 7584 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_80
timestamp 1679585382
transform 1 0 8256 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_87
timestamp 1679585382
transform 1 0 8928 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_94
timestamp 1679585382
transform 1 0 9600 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_101
timestamp 1679585382
transform 1 0 10272 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_108
timestamp 1679585382
transform 1 0 10944 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_115
timestamp 1679585382
transform 1 0 11616 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_122
timestamp 1679585382
transform 1 0 12288 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_129
timestamp 1679585382
transform 1 0 12960 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_136
timestamp 1679585382
transform 1 0 13632 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_143
timestamp 1679585382
transform 1 0 14304 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_150
timestamp 1679585382
transform 1 0 14976 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_157
timestamp 1679585382
transform 1 0 15648 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_164
timestamp 1679585382
transform 1 0 16320 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_171
timestamp 1679585382
transform 1 0 16992 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_178
timestamp 1679585382
transform 1 0 17664 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_185
timestamp 1679585382
transform 1 0 18336 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_192
timestamp 1679585382
transform 1 0 19008 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_199
timestamp 1679585382
transform 1 0 19680 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_206
timestamp 1677583704
transform 1 0 20352 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_216
timestamp 1679585382
transform 1 0 21312 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_223
timestamp 1679585382
transform 1 0 21984 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_230
timestamp 1679585382
transform 1 0 22656 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_237
timestamp 1679585382
transform 1 0 23328 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_244
timestamp 1679585382
transform 1 0 24000 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_251
timestamp 1679585382
transform 1 0 24672 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_258
timestamp 1679585382
transform 1 0 25344 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_265
timestamp 1679585382
transform 1 0 26016 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_272
timestamp 1679585382
transform 1 0 26688 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_29_279
timestamp 1677583258
transform 1 0 27360 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_289
timestamp 1679585382
transform 1 0 28320 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_296
timestamp 1679585382
transform 1 0 28992 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_303
timestamp 1679585382
transform 1 0 29664 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_310
timestamp 1679585382
transform 1 0 30336 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_317
timestamp 1679585382
transform 1 0 31008 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_324
timestamp 1679585382
transform 1 0 31680 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_331
timestamp 1679585382
transform 1 0 32352 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_338
timestamp 1679585382
transform 1 0 33024 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_354
timestamp 1679585382
transform 1 0 34560 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_361
timestamp 1679585382
transform 1 0 35232 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_368
timestamp 1679585382
transform 1 0 35904 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_375
timestamp 1677583704
transform 1 0 36576 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_404
timestamp 1679585382
transform 1 0 39360 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_29_411
timestamp 1677583258
transform 1 0 40032 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_420
timestamp 1679585382
transform 1 0 40896 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_427
timestamp 1679585382
transform 1 0 41568 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_434
timestamp 1679585382
transform 1 0 42240 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_441
timestamp 1679585382
transform 1 0 42912 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_448
timestamp 1679585382
transform 1 0 43584 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_455
timestamp 1679585382
transform 1 0 44256 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_462
timestamp 1679585382
transform 1 0 44928 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_469
timestamp 1679585382
transform 1 0 45600 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_476
timestamp 1679585382
transform 1 0 46272 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_483
timestamp 1679585382
transform 1 0 46944 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_490
timestamp 1679585382
transform 1 0 47616 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_497
timestamp 1679585382
transform 1 0 48288 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_504
timestamp 1679585382
transform 1 0 48960 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_511
timestamp 1679585382
transform 1 0 49632 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_518
timestamp 1679585382
transform 1 0 50304 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_525
timestamp 1679585382
transform 1 0 50976 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_532
timestamp 1679585382
transform 1 0 51648 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_539
timestamp 1679585382
transform 1 0 52320 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_546
timestamp 1679585382
transform 1 0 52992 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_553
timestamp 1679585382
transform 1 0 53664 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_560
timestamp 1679585382
transform 1 0 54336 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_567
timestamp 1679585382
transform 1 0 55008 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_574
timestamp 1679585382
transform 1 0 55680 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_581
timestamp 1679585382
transform 1 0 56352 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_588
timestamp 1679585382
transform 1 0 57024 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_595
timestamp 1679585382
transform 1 0 57696 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_602
timestamp 1679585382
transform 1 0 58368 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_609
timestamp 1679585382
transform 1 0 59040 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_616
timestamp 1679585382
transform 1 0 59712 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_623
timestamp 1679585382
transform 1 0 60384 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_630
timestamp 1679585382
transform 1 0 61056 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_637
timestamp 1679585382
transform 1 0 61728 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_644
timestamp 1679585382
transform 1 0 62400 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_651
timestamp 1679585382
transform 1 0 63072 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_658
timestamp 1679585382
transform 1 0 63744 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_665
timestamp 1679585382
transform 1 0 64416 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_672
timestamp 1679585382
transform 1 0 65088 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_679
timestamp 1679585382
transform 1 0 65760 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_686
timestamp 1679585382
transform 1 0 66432 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_693
timestamp 1679585382
transform 1 0 67104 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_700
timestamp 1679585382
transform 1 0 67776 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_707
timestamp 1679585382
transform 1 0 68448 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_714
timestamp 1679585382
transform 1 0 69120 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_721
timestamp 1679585382
transform 1 0 69792 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_728
timestamp 1679585382
transform 1 0 70464 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_735
timestamp 1679585382
transform 1 0 71136 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_742
timestamp 1679585382
transform 1 0 71808 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_749
timestamp 1679585382
transform 1 0 72480 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_756
timestamp 1679585382
transform 1 0 73152 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_763
timestamp 1679585382
transform 1 0 73824 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_770
timestamp 1679585382
transform 1 0 74496 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_777
timestamp 1679585382
transform 1 0 75168 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_784
timestamp 1679585382
transform 1 0 75840 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_791
timestamp 1679585382
transform 1 0 76512 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_798
timestamp 1679585382
transform 1 0 77184 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_805
timestamp 1679585382
transform 1 0 77856 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_812
timestamp 1679585382
transform 1 0 78528 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_819
timestamp 1679585382
transform 1 0 79200 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_826
timestamp 1679585382
transform 1 0 79872 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_833
timestamp 1679585382
transform 1 0 80544 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_840
timestamp 1679585382
transform 1 0 81216 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_847
timestamp 1679585382
transform 1 0 81888 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_854
timestamp 1679585382
transform 1 0 82560 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_861
timestamp 1679585382
transform 1 0 83232 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_868
timestamp 1679585382
transform 1 0 83904 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_875
timestamp 1679585382
transform 1 0 84576 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_882
timestamp 1679585382
transform 1 0 85248 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_889
timestamp 1679585382
transform 1 0 85920 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_896
timestamp 1679585382
transform 1 0 86592 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_903
timestamp 1679585382
transform 1 0 87264 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_910
timestamp 1679585382
transform 1 0 87936 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_917
timestamp 1679585382
transform 1 0 88608 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_924
timestamp 1679585382
transform 1 0 89280 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_931
timestamp 1679585382
transform 1 0 89952 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_938
timestamp 1679585382
transform 1 0 90624 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_945
timestamp 1679585382
transform 1 0 91296 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_952
timestamp 1679585382
transform 1 0 91968 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_959
timestamp 1679585382
transform 1 0 92640 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_966
timestamp 1679585382
transform 1 0 93312 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_973
timestamp 1679585382
transform 1 0 93984 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_980
timestamp 1679585382
transform 1 0 94656 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_987
timestamp 1679585382
transform 1 0 95328 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_994
timestamp 1679585382
transform 1 0 96000 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1001
timestamp 1679585382
transform 1 0 96672 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1008
timestamp 1679585382
transform 1 0 97344 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1015
timestamp 1679585382
transform 1 0 98016 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1022
timestamp 1679585382
transform 1 0 98688 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_0
timestamp 1679585382
transform 1 0 576 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_7
timestamp 1679585382
transform 1 0 1248 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_14
timestamp 1679585382
transform 1 0 1920 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_21
timestamp 1679585382
transform 1 0 2592 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_28
timestamp 1679585382
transform 1 0 3264 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_35
timestamp 1679585382
transform 1 0 3936 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_42
timestamp 1679585382
transform 1 0 4608 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_49
timestamp 1679585382
transform 1 0 5280 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_56
timestamp 1679585382
transform 1 0 5952 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_63
timestamp 1679585382
transform 1 0 6624 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_70
timestamp 1679585382
transform 1 0 7296 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_77
timestamp 1679585382
transform 1 0 7968 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_84
timestamp 1679585382
transform 1 0 8640 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_91
timestamp 1679585382
transform 1 0 9312 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_98
timestamp 1679585382
transform 1 0 9984 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_105
timestamp 1679585382
transform 1 0 10656 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_112
timestamp 1679585382
transform 1 0 11328 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_119
timestamp 1679585382
transform 1 0 12000 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_126
timestamp 1679585382
transform 1 0 12672 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_133
timestamp 1679585382
transform 1 0 13344 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_140
timestamp 1679585382
transform 1 0 14016 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_147
timestamp 1679585382
transform 1 0 14688 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_207
timestamp 1677583704
transform 1 0 20448 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_209
timestamp 1677583258
transform 1 0 20640 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_227
timestamp 1679585382
transform 1 0 22368 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_234
timestamp 1679585382
transform 1 0 23040 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_241
timestamp 1679585382
transform 1 0 23712 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_248
timestamp 1679585382
transform 1 0 24384 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_255
timestamp 1679585382
transform 1 0 25056 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_262
timestamp 1679585382
transform 1 0 25728 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_269
timestamp 1679585382
transform 1 0 26400 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_276
timestamp 1679585382
transform 1 0 27072 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_283
timestamp 1679585382
transform 1 0 27744 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_290
timestamp 1679585382
transform 1 0 28416 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_297
timestamp 1679585382
transform 1 0 29088 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_304
timestamp 1679581501
transform 1 0 29760 0 1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_30_335
timestamp 1679585382
transform 1 0 32736 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_342
timestamp 1679585382
transform 1 0 33408 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_349
timestamp 1679585382
transform 1 0 34080 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_368
timestamp 1679585382
transform 1 0 35904 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_375
timestamp 1679585382
transform 1 0 36576 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_382
timestamp 1679585382
transform 1 0 37248 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_389
timestamp 1679585382
transform 1 0 37920 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_396
timestamp 1679585382
transform 1 0 38592 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_403
timestamp 1679581501
transform 1 0 39264 0 1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_30_407
timestamp 1677583704
transform 1 0 39648 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_418
timestamp 1677583258
transform 1 0 40704 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_454
timestamp 1679585382
transform 1 0 44160 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_461
timestamp 1679581501
transform 1 0 44832 0 1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_30_465
timestamp 1677583704
transform 1 0 45216 0 1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_471
timestamp 1677583704
transform 1 0 45792 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_473
timestamp 1677583258
transform 1 0 45984 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_478
timestamp 1679585382
transform 1 0 46464 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_485
timestamp 1679581501
transform 1 0 47136 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_489
timestamp 1677583258
transform 1 0 47520 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_499
timestamp 1679585382
transform 1 0 48480 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_506
timestamp 1679585382
transform 1 0 49152 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_513
timestamp 1679585382
transform 1 0 49824 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_520
timestamp 1679585382
transform 1 0 50496 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_527
timestamp 1679585382
transform 1 0 51168 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_534
timestamp 1679585382
transform 1 0 51840 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_541
timestamp 1679585382
transform 1 0 52512 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_548
timestamp 1679585382
transform 1 0 53184 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_555
timestamp 1679585382
transform 1 0 53856 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_562
timestamp 1679585382
transform 1 0 54528 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_569
timestamp 1679585382
transform 1 0 55200 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_576
timestamp 1679585382
transform 1 0 55872 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_583
timestamp 1679585382
transform 1 0 56544 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_590
timestamp 1679585382
transform 1 0 57216 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_597
timestamp 1679585382
transform 1 0 57888 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_604
timestamp 1679585382
transform 1 0 58560 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_611
timestamp 1679585382
transform 1 0 59232 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_618
timestamp 1679585382
transform 1 0 59904 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_625
timestamp 1679585382
transform 1 0 60576 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_632
timestamp 1679585382
transform 1 0 61248 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_639
timestamp 1679585382
transform 1 0 61920 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_646
timestamp 1679585382
transform 1 0 62592 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_653
timestamp 1679585382
transform 1 0 63264 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_660
timestamp 1679585382
transform 1 0 63936 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_667
timestamp 1679585382
transform 1 0 64608 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_674
timestamp 1679585382
transform 1 0 65280 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_681
timestamp 1679585382
transform 1 0 65952 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_688
timestamp 1679585382
transform 1 0 66624 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_695
timestamp 1679585382
transform 1 0 67296 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_702
timestamp 1679585382
transform 1 0 67968 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_709
timestamp 1679585382
transform 1 0 68640 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_716
timestamp 1679585382
transform 1 0 69312 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_723
timestamp 1679585382
transform 1 0 69984 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_730
timestamp 1679585382
transform 1 0 70656 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_737
timestamp 1679585382
transform 1 0 71328 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_744
timestamp 1679585382
transform 1 0 72000 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_751
timestamp 1679585382
transform 1 0 72672 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_758
timestamp 1679585382
transform 1 0 73344 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_765
timestamp 1679585382
transform 1 0 74016 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_772
timestamp 1679585382
transform 1 0 74688 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_779
timestamp 1679585382
transform 1 0 75360 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_786
timestamp 1679585382
transform 1 0 76032 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_793
timestamp 1679585382
transform 1 0 76704 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_800
timestamp 1679585382
transform 1 0 77376 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_807
timestamp 1679585382
transform 1 0 78048 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_814
timestamp 1679585382
transform 1 0 78720 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_821
timestamp 1679585382
transform 1 0 79392 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_828
timestamp 1679585382
transform 1 0 80064 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_835
timestamp 1679585382
transform 1 0 80736 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_842
timestamp 1679585382
transform 1 0 81408 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_849
timestamp 1679585382
transform 1 0 82080 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_856
timestamp 1679585382
transform 1 0 82752 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_863
timestamp 1679585382
transform 1 0 83424 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_870
timestamp 1679585382
transform 1 0 84096 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_877
timestamp 1679585382
transform 1 0 84768 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_884
timestamp 1679585382
transform 1 0 85440 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_891
timestamp 1679585382
transform 1 0 86112 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_898
timestamp 1679585382
transform 1 0 86784 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_905
timestamp 1679585382
transform 1 0 87456 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_912
timestamp 1679585382
transform 1 0 88128 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_919
timestamp 1679585382
transform 1 0 88800 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_926
timestamp 1679585382
transform 1 0 89472 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_933
timestamp 1679585382
transform 1 0 90144 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_940
timestamp 1679585382
transform 1 0 90816 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_947
timestamp 1679585382
transform 1 0 91488 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_954
timestamp 1679585382
transform 1 0 92160 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_961
timestamp 1679585382
transform 1 0 92832 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_968
timestamp 1679585382
transform 1 0 93504 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_975
timestamp 1679585382
transform 1 0 94176 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_982
timestamp 1679585382
transform 1 0 94848 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_989
timestamp 1679585382
transform 1 0 95520 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_996
timestamp 1679585382
transform 1 0 96192 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1003
timestamp 1679585382
transform 1 0 96864 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1010
timestamp 1679585382
transform 1 0 97536 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1017
timestamp 1679585382
transform 1 0 98208 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_1024
timestamp 1679581501
transform 1 0 98880 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_1028
timestamp 1677583258
transform 1 0 99264 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_0
timestamp 1679585382
transform 1 0 576 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_7
timestamp 1679585382
transform 1 0 1248 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_14
timestamp 1679585382
transform 1 0 1920 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_21
timestamp 1679585382
transform 1 0 2592 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_28
timestamp 1679585382
transform 1 0 3264 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_35
timestamp 1679585382
transform 1 0 3936 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_42
timestamp 1679585382
transform 1 0 4608 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_49
timestamp 1679585382
transform 1 0 5280 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_56
timestamp 1679585382
transform 1 0 5952 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_63
timestamp 1679585382
transform 1 0 6624 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_70
timestamp 1679585382
transform 1 0 7296 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_77
timestamp 1679585382
transform 1 0 7968 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_84
timestamp 1679585382
transform 1 0 8640 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_91
timestamp 1679585382
transform 1 0 9312 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_98
timestamp 1679585382
transform 1 0 9984 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_105
timestamp 1679585382
transform 1 0 10656 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_112
timestamp 1679581501
transform 1 0 11328 0 -1 24948
box -48 -56 432 834
use sg13g2_decap_8  FILLER_31_129
timestamp 1679585382
transform 1 0 12960 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_136
timestamp 1679585382
transform 1 0 13632 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_143
timestamp 1679585382
transform 1 0 14304 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_150
timestamp 1677583704
transform 1 0 14976 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_173
timestamp 1679585382
transform 1 0 17184 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_180
timestamp 1679585382
transform 1 0 17856 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_187
timestamp 1679585382
transform 1 0 18528 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_194
timestamp 1679585382
transform 1 0 19200 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_201
timestamp 1679585382
transform 1 0 19872 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_208
timestamp 1677583704
transform 1 0 20544 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_210
timestamp 1677583258
transform 1 0 20736 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_215
timestamp 1679585382
transform 1 0 21216 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_222
timestamp 1679585382
transform 1 0 21888 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_229
timestamp 1677583704
transform 1 0 22560 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_231
timestamp 1677583258
transform 1 0 22752 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_241
timestamp 1679585382
transform 1 0 23712 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_248
timestamp 1677583704
transform 1 0 24384 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_250
timestamp 1677583258
transform 1 0 24576 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_278
timestamp 1679585382
transform 1 0 27264 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_285
timestamp 1679585382
transform 1 0 27936 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_292
timestamp 1679585382
transform 1 0 28608 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_299
timestamp 1679585382
transform 1 0 29280 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_306
timestamp 1679585382
transform 1 0 29952 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_313
timestamp 1679581501
transform 1 0 30624 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_317
timestamp 1677583704
transform 1 0 31008 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_323
timestamp 1679585382
transform 1 0 31584 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_330
timestamp 1679585382
transform 1 0 32256 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_337
timestamp 1679585382
transform 1 0 32928 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_344
timestamp 1677583704
transform 1 0 33600 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_31_363
timestamp 1679585382
transform 1 0 35424 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_370
timestamp 1679585382
transform 1 0 36096 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_377
timestamp 1679585382
transform 1 0 36768 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_384
timestamp 1679585382
transform 1 0 37440 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_391
timestamp 1679585382
transform 1 0 38112 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_398
timestamp 1679585382
transform 1 0 38784 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_405
timestamp 1679585382
transform 1 0 39456 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_412
timestamp 1679585382
transform 1 0 40128 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_419
timestamp 1679585382
transform 1 0 40800 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_426
timestamp 1679585382
transform 1 0 41472 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_433
timestamp 1679585382
transform 1 0 42144 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_440
timestamp 1679581501
transform 1 0 42816 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_31_444
timestamp 1677583258
transform 1 0 43200 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_449
timestamp 1679585382
transform 1 0 43680 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_456
timestamp 1679581501
transform 1 0 44352 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_31_460
timestamp 1677583258
transform 1 0 44736 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_505
timestamp 1679585382
transform 1 0 49056 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_512
timestamp 1679585382
transform 1 0 49728 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_519
timestamp 1679585382
transform 1 0 50400 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_526
timestamp 1679585382
transform 1 0 51072 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_533
timestamp 1679585382
transform 1 0 51744 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_540
timestamp 1679585382
transform 1 0 52416 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_547
timestamp 1679585382
transform 1 0 53088 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_554
timestamp 1679585382
transform 1 0 53760 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_561
timestamp 1679585382
transform 1 0 54432 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_568
timestamp 1679585382
transform 1 0 55104 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_575
timestamp 1679585382
transform 1 0 55776 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_582
timestamp 1679585382
transform 1 0 56448 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_589
timestamp 1679585382
transform 1 0 57120 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_596
timestamp 1679585382
transform 1 0 57792 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_603
timestamp 1679585382
transform 1 0 58464 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_610
timestamp 1679585382
transform 1 0 59136 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_617
timestamp 1679585382
transform 1 0 59808 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_624
timestamp 1679585382
transform 1 0 60480 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_631
timestamp 1679585382
transform 1 0 61152 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_638
timestamp 1679585382
transform 1 0 61824 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_645
timestamp 1679585382
transform 1 0 62496 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_652
timestamp 1679585382
transform 1 0 63168 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_659
timestamp 1679585382
transform 1 0 63840 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_666
timestamp 1679585382
transform 1 0 64512 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_673
timestamp 1679585382
transform 1 0 65184 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_680
timestamp 1679585382
transform 1 0 65856 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_687
timestamp 1679585382
transform 1 0 66528 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_694
timestamp 1679585382
transform 1 0 67200 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_701
timestamp 1679585382
transform 1 0 67872 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_708
timestamp 1679585382
transform 1 0 68544 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_715
timestamp 1679585382
transform 1 0 69216 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_722
timestamp 1679585382
transform 1 0 69888 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_729
timestamp 1679585382
transform 1 0 70560 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_736
timestamp 1679585382
transform 1 0 71232 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_743
timestamp 1679585382
transform 1 0 71904 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_750
timestamp 1679585382
transform 1 0 72576 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_757
timestamp 1679585382
transform 1 0 73248 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_764
timestamp 1679585382
transform 1 0 73920 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_771
timestamp 1679585382
transform 1 0 74592 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_778
timestamp 1679585382
transform 1 0 75264 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_785
timestamp 1679585382
transform 1 0 75936 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_792
timestamp 1679585382
transform 1 0 76608 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_799
timestamp 1679585382
transform 1 0 77280 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_806
timestamp 1679585382
transform 1 0 77952 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_813
timestamp 1679585382
transform 1 0 78624 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_820
timestamp 1679585382
transform 1 0 79296 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_827
timestamp 1679585382
transform 1 0 79968 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_834
timestamp 1679585382
transform 1 0 80640 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_841
timestamp 1679585382
transform 1 0 81312 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_848
timestamp 1679585382
transform 1 0 81984 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_855
timestamp 1679585382
transform 1 0 82656 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_862
timestamp 1679585382
transform 1 0 83328 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_869
timestamp 1679585382
transform 1 0 84000 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_876
timestamp 1679585382
transform 1 0 84672 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_883
timestamp 1679585382
transform 1 0 85344 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_890
timestamp 1679585382
transform 1 0 86016 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_897
timestamp 1679585382
transform 1 0 86688 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_904
timestamp 1679585382
transform 1 0 87360 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_911
timestamp 1679585382
transform 1 0 88032 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_918
timestamp 1679585382
transform 1 0 88704 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_925
timestamp 1679585382
transform 1 0 89376 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_932
timestamp 1679585382
transform 1 0 90048 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_939
timestamp 1679585382
transform 1 0 90720 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_946
timestamp 1679585382
transform 1 0 91392 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_953
timestamp 1679585382
transform 1 0 92064 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_960
timestamp 1679585382
transform 1 0 92736 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_967
timestamp 1679585382
transform 1 0 93408 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_974
timestamp 1679585382
transform 1 0 94080 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_981
timestamp 1679585382
transform 1 0 94752 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_988
timestamp 1679585382
transform 1 0 95424 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_995
timestamp 1679585382
transform 1 0 96096 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1002
timestamp 1679585382
transform 1 0 96768 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1009
timestamp 1679585382
transform 1 0 97440 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_1016
timestamp 1679585382
transform 1 0 98112 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_1023
timestamp 1679581501
transform 1 0 98784 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_1027
timestamp 1677583704
transform 1 0 99168 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_0
timestamp 1679585382
transform 1 0 576 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_7
timestamp 1679585382
transform 1 0 1248 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_14
timestamp 1679581501
transform 1 0 1920 0 1 24948
box -48 -56 432 834
use sg13g2_decap_8  FILLER_32_45
timestamp 1679585382
transform 1 0 4896 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_52
timestamp 1677583704
transform 1 0 5568 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_67
timestamp 1679585382
transform 1 0 7008 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_74
timestamp 1679585382
transform 1 0 7680 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_81
timestamp 1679585382
transform 1 0 8352 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_88
timestamp 1679585382
transform 1 0 9024 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_95
timestamp 1679585382
transform 1 0 9696 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_102
timestamp 1679585382
transform 1 0 10368 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_109
timestamp 1677583704
transform 1 0 11040 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_111
timestamp 1677583258
transform 1 0 11232 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_139
timestamp 1679585382
transform 1 0 13920 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_146
timestamp 1679585382
transform 1 0 14592 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_153
timestamp 1679585382
transform 1 0 15264 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_160
timestamp 1679581501
transform 1 0 15936 0 1 24948
box -48 -56 432 834
use sg13g2_decap_8  FILLER_32_172
timestamp 1679585382
transform 1 0 17088 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_179
timestamp 1679585382
transform 1 0 17760 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_186
timestamp 1679585382
transform 1 0 18432 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_193
timestamp 1679585382
transform 1 0 19104 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_200
timestamp 1679585382
transform 1 0 19776 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_207
timestamp 1679585382
transform 1 0 20448 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_214
timestamp 1679581501
transform 1 0 21120 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_218
timestamp 1677583704
transform 1 0 21504 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_228
timestamp 1679585382
transform 1 0 22464 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_235
timestamp 1679585382
transform 1 0 23136 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_242
timestamp 1677583704
transform 1 0 23808 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_244
timestamp 1677583258
transform 1 0 24000 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_258
timestamp 1679585382
transform 1 0 25344 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_265
timestamp 1679585382
transform 1 0 26016 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_272
timestamp 1679585382
transform 1 0 26688 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_279
timestamp 1679585382
transform 1 0 27360 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_286
timestamp 1679581501
transform 1 0 28032 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_290
timestamp 1677583258
transform 1 0 28416 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_304
timestamp 1679585382
transform 1 0 29760 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_311
timestamp 1679585382
transform 1 0 30432 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_318
timestamp 1679585382
transform 1 0 31104 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_325
timestamp 1679585382
transform 1 0 31776 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_332
timestamp 1679585382
transform 1 0 32448 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_339
timestamp 1679585382
transform 1 0 33120 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_346
timestamp 1679585382
transform 1 0 33792 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_353
timestamp 1679585382
transform 1 0 34464 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_360
timestamp 1679585382
transform 1 0 35136 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_367
timestamp 1679585382
transform 1 0 35808 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_374
timestamp 1679585382
transform 1 0 36480 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_381
timestamp 1679585382
transform 1 0 37152 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_388
timestamp 1679585382
transform 1 0 37824 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_395
timestamp 1679585382
transform 1 0 38496 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_402
timestamp 1679585382
transform 1 0 39168 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_409
timestamp 1679585382
transform 1 0 39840 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_416
timestamp 1679585382
transform 1 0 40512 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_423
timestamp 1679585382
transform 1 0 41184 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_430
timestamp 1679585382
transform 1 0 41856 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_437
timestamp 1679585382
transform 1 0 42528 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_444
timestamp 1679585382
transform 1 0 43200 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_451
timestamp 1679585382
transform 1 0 43872 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_458
timestamp 1679581501
transform 1 0 44544 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_462
timestamp 1677583704
transform 1 0 44928 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_32_491
timestamp 1679585382
transform 1 0 47712 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_498
timestamp 1679585382
transform 1 0 48384 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_505
timestamp 1679585382
transform 1 0 49056 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_512
timestamp 1679585382
transform 1 0 49728 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_519
timestamp 1679585382
transform 1 0 50400 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_526
timestamp 1679585382
transform 1 0 51072 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_533
timestamp 1679585382
transform 1 0 51744 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_540
timestamp 1679585382
transform 1 0 52416 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_547
timestamp 1679585382
transform 1 0 53088 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_554
timestamp 1679585382
transform 1 0 53760 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_561
timestamp 1679585382
transform 1 0 54432 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_568
timestamp 1679585382
transform 1 0 55104 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_575
timestamp 1679585382
transform 1 0 55776 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_582
timestamp 1679585382
transform 1 0 56448 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_589
timestamp 1679585382
transform 1 0 57120 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_596
timestamp 1679585382
transform 1 0 57792 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_603
timestamp 1679585382
transform 1 0 58464 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_610
timestamp 1679585382
transform 1 0 59136 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_617
timestamp 1679585382
transform 1 0 59808 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_624
timestamp 1679585382
transform 1 0 60480 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_631
timestamp 1679585382
transform 1 0 61152 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_638
timestamp 1679585382
transform 1 0 61824 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_645
timestamp 1679585382
transform 1 0 62496 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_652
timestamp 1679585382
transform 1 0 63168 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_659
timestamp 1679585382
transform 1 0 63840 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_666
timestamp 1679585382
transform 1 0 64512 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_673
timestamp 1679585382
transform 1 0 65184 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_680
timestamp 1679585382
transform 1 0 65856 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_687
timestamp 1679585382
transform 1 0 66528 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_694
timestamp 1679585382
transform 1 0 67200 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_701
timestamp 1679585382
transform 1 0 67872 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_708
timestamp 1679585382
transform 1 0 68544 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_715
timestamp 1679585382
transform 1 0 69216 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_722
timestamp 1679585382
transform 1 0 69888 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_729
timestamp 1679585382
transform 1 0 70560 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_736
timestamp 1679585382
transform 1 0 71232 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_743
timestamp 1679585382
transform 1 0 71904 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_750
timestamp 1679585382
transform 1 0 72576 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_757
timestamp 1679585382
transform 1 0 73248 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_764
timestamp 1679585382
transform 1 0 73920 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_771
timestamp 1679585382
transform 1 0 74592 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_778
timestamp 1679585382
transform 1 0 75264 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_785
timestamp 1679585382
transform 1 0 75936 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_792
timestamp 1679585382
transform 1 0 76608 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_799
timestamp 1679585382
transform 1 0 77280 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_806
timestamp 1679585382
transform 1 0 77952 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_813
timestamp 1679585382
transform 1 0 78624 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_820
timestamp 1679585382
transform 1 0 79296 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_827
timestamp 1679585382
transform 1 0 79968 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_834
timestamp 1679585382
transform 1 0 80640 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_841
timestamp 1679585382
transform 1 0 81312 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_848
timestamp 1679585382
transform 1 0 81984 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_855
timestamp 1679585382
transform 1 0 82656 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_862
timestamp 1679585382
transform 1 0 83328 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_869
timestamp 1679585382
transform 1 0 84000 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_876
timestamp 1679585382
transform 1 0 84672 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_883
timestamp 1679585382
transform 1 0 85344 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_890
timestamp 1679585382
transform 1 0 86016 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_897
timestamp 1679585382
transform 1 0 86688 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_904
timestamp 1679585382
transform 1 0 87360 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_911
timestamp 1679585382
transform 1 0 88032 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_918
timestamp 1679585382
transform 1 0 88704 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_925
timestamp 1679585382
transform 1 0 89376 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_932
timestamp 1679585382
transform 1 0 90048 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_939
timestamp 1679585382
transform 1 0 90720 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_946
timestamp 1679585382
transform 1 0 91392 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_953
timestamp 1679585382
transform 1 0 92064 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_960
timestamp 1679585382
transform 1 0 92736 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_967
timestamp 1679585382
transform 1 0 93408 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_974
timestamp 1679585382
transform 1 0 94080 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_981
timestamp 1679585382
transform 1 0 94752 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_988
timestamp 1679585382
transform 1 0 95424 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_995
timestamp 1679585382
transform 1 0 96096 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1002
timestamp 1679585382
transform 1 0 96768 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1009
timestamp 1679585382
transform 1 0 97440 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_1016
timestamp 1679585382
transform 1 0 98112 0 1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_32_1023
timestamp 1679581501
transform 1 0 98784 0 1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_32_1027
timestamp 1677583704
transform 1 0 99168 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_0
timestamp 1679585382
transform 1 0 576 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_7
timestamp 1679585382
transform 1 0 1248 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_14
timestamp 1679581501
transform 1 0 1920 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_33_18
timestamp 1677583258
transform 1 0 2304 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_46
timestamp 1679585382
transform 1 0 4992 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_53
timestamp 1679585382
transform 1 0 5664 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_60
timestamp 1679585382
transform 1 0 6336 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_94
timestamp 1679581501
transform 1 0 9600 0 -1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_33_142
timestamp 1679585382
transform 1 0 14208 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_149
timestamp 1679585382
transform 1 0 14880 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_156
timestamp 1679585382
transform 1 0 15552 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_163
timestamp 1679585382
transform 1 0 16224 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_170
timestamp 1679585382
transform 1 0 16896 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_177
timestamp 1677583704
transform 1 0 17568 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_33_215
timestamp 1677583704
transform 1 0 21216 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_217
timestamp 1677583258
transform 1 0 21408 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_245
timestamp 1679585382
transform 1 0 24096 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_252
timestamp 1679585382
transform 1 0 24768 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_259
timestamp 1679585382
transform 1 0 25440 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_266
timestamp 1679585382
transform 1 0 26112 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_273
timestamp 1679585382
transform 1 0 26784 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_280
timestamp 1677583704
transform 1 0 27456 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_299
timestamp 1679585382
transform 1 0 29280 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_306
timestamp 1679585382
transform 1 0 29952 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_313
timestamp 1679585382
transform 1 0 30624 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_320
timestamp 1679585382
transform 1 0 31296 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_327
timestamp 1679585382
transform 1 0 31968 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_334
timestamp 1679585382
transform 1 0 32640 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_345
timestamp 1677583704
transform 1 0 33696 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_347
timestamp 1677583258
transform 1 0 33888 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_361
timestamp 1677583704
transform 1 0 35232 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_363
timestamp 1677583258
transform 1 0 35424 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_377
timestamp 1679585382
transform 1 0 36768 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_384
timestamp 1679585382
transform 1 0 37440 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_391
timestamp 1679585382
transform 1 0 38112 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_398
timestamp 1679585382
transform 1 0 38784 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_405
timestamp 1679585382
transform 1 0 39456 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_412
timestamp 1679585382
transform 1 0 40128 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_419
timestamp 1679581501
transform 1 0 40800 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_33_423
timestamp 1677583704
transform 1 0 41184 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_429
timestamp 1679585382
transform 1 0 41760 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_436
timestamp 1679585382
transform 1 0 42432 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_443
timestamp 1677583704
transform 1 0 43104 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_445
timestamp 1677583258
transform 1 0 43296 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_459
timestamp 1679585382
transform 1 0 44640 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_466
timestamp 1679585382
transform 1 0 45312 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_473
timestamp 1677583704
transform 1 0 45984 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_475
timestamp 1677583258
transform 1 0 46176 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_485
timestamp 1679585382
transform 1 0 47136 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_492
timestamp 1679585382
transform 1 0 47808 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_499
timestamp 1679585382
transform 1 0 48480 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_506
timestamp 1679585382
transform 1 0 49152 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_513
timestamp 1679585382
transform 1 0 49824 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_520
timestamp 1679585382
transform 1 0 50496 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_527
timestamp 1679585382
transform 1 0 51168 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_534
timestamp 1679585382
transform 1 0 51840 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_541
timestamp 1679585382
transform 1 0 52512 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_548
timestamp 1679585382
transform 1 0 53184 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_555
timestamp 1679585382
transform 1 0 53856 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_562
timestamp 1679585382
transform 1 0 54528 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_569
timestamp 1679585382
transform 1 0 55200 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_576
timestamp 1679585382
transform 1 0 55872 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_583
timestamp 1679585382
transform 1 0 56544 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_590
timestamp 1679585382
transform 1 0 57216 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_597
timestamp 1679585382
transform 1 0 57888 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_604
timestamp 1679585382
transform 1 0 58560 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_611
timestamp 1679585382
transform 1 0 59232 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_618
timestamp 1679585382
transform 1 0 59904 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_625
timestamp 1679585382
transform 1 0 60576 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_632
timestamp 1679585382
transform 1 0 61248 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_639
timestamp 1679585382
transform 1 0 61920 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_646
timestamp 1679585382
transform 1 0 62592 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_653
timestamp 1679585382
transform 1 0 63264 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_660
timestamp 1679585382
transform 1 0 63936 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_667
timestamp 1679585382
transform 1 0 64608 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_674
timestamp 1679585382
transform 1 0 65280 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_681
timestamp 1679585382
transform 1 0 65952 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_688
timestamp 1679585382
transform 1 0 66624 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_695
timestamp 1679585382
transform 1 0 67296 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_702
timestamp 1679585382
transform 1 0 67968 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_709
timestamp 1679585382
transform 1 0 68640 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_716
timestamp 1679585382
transform 1 0 69312 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_723
timestamp 1679585382
transform 1 0 69984 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_730
timestamp 1679585382
transform 1 0 70656 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_737
timestamp 1679585382
transform 1 0 71328 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_744
timestamp 1679585382
transform 1 0 72000 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_751
timestamp 1679585382
transform 1 0 72672 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_758
timestamp 1679585382
transform 1 0 73344 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_765
timestamp 1679585382
transform 1 0 74016 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_772
timestamp 1679585382
transform 1 0 74688 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_779
timestamp 1679585382
transform 1 0 75360 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_786
timestamp 1679585382
transform 1 0 76032 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_793
timestamp 1679585382
transform 1 0 76704 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_800
timestamp 1679585382
transform 1 0 77376 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_807
timestamp 1679585382
transform 1 0 78048 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_814
timestamp 1679585382
transform 1 0 78720 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_821
timestamp 1679585382
transform 1 0 79392 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_828
timestamp 1679585382
transform 1 0 80064 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_835
timestamp 1679585382
transform 1 0 80736 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_842
timestamp 1679585382
transform 1 0 81408 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_849
timestamp 1679585382
transform 1 0 82080 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_856
timestamp 1679585382
transform 1 0 82752 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_863
timestamp 1679585382
transform 1 0 83424 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_870
timestamp 1679585382
transform 1 0 84096 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_877
timestamp 1679585382
transform 1 0 84768 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_884
timestamp 1679585382
transform 1 0 85440 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_891
timestamp 1679585382
transform 1 0 86112 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_898
timestamp 1679585382
transform 1 0 86784 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_905
timestamp 1679585382
transform 1 0 87456 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_912
timestamp 1679585382
transform 1 0 88128 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_919
timestamp 1679585382
transform 1 0 88800 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_926
timestamp 1679585382
transform 1 0 89472 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_933
timestamp 1679585382
transform 1 0 90144 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_940
timestamp 1679585382
transform 1 0 90816 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_947
timestamp 1679585382
transform 1 0 91488 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_954
timestamp 1679585382
transform 1 0 92160 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_961
timestamp 1679585382
transform 1 0 92832 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_968
timestamp 1679585382
transform 1 0 93504 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_975
timestamp 1679585382
transform 1 0 94176 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_982
timestamp 1679585382
transform 1 0 94848 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_989
timestamp 1679585382
transform 1 0 95520 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_996
timestamp 1679585382
transform 1 0 96192 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1003
timestamp 1679585382
transform 1 0 96864 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1010
timestamp 1679585382
transform 1 0 97536 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_1017
timestamp 1679585382
transform 1 0 98208 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_1024
timestamp 1679581501
transform 1 0 98880 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_33_1028
timestamp 1677583258
transform 1 0 99264 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_0
timestamp 1679585382
transform 1 0 576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_7
timestamp 1679585382
transform 1 0 1248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_14
timestamp 1679585382
transform 1 0 1920 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_21
timestamp 1679581501
transform 1 0 2592 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_25
timestamp 1677583704
transform 1 0 2976 0 1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_34_35
timestamp 1677583704
transform 1 0 3936 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_55
timestamp 1679585382
transform 1 0 5856 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_62
timestamp 1679585382
transform 1 0 6528 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_69
timestamp 1679585382
transform 1 0 7200 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_76
timestamp 1679585382
transform 1 0 7872 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_83
timestamp 1679585382
transform 1 0 8544 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_90
timestamp 1679585382
transform 1 0 9216 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_97
timestamp 1677583704
transform 1 0 9888 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_112
timestamp 1679585382
transform 1 0 11328 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_119
timestamp 1679585382
transform 1 0 12000 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_126
timestamp 1679585382
transform 1 0 12672 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_133
timestamp 1679585382
transform 1 0 13344 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_140
timestamp 1679585382
transform 1 0 14016 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_147
timestamp 1679585382
transform 1 0 14688 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_154
timestamp 1679585382
transform 1 0 15360 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_161
timestamp 1679585382
transform 1 0 16032 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_168
timestamp 1679585382
transform 1 0 16704 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_175
timestamp 1679585382
transform 1 0 17376 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_182
timestamp 1679585382
transform 1 0 18048 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_189
timestamp 1679585382
transform 1 0 18720 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_196
timestamp 1679585382
transform 1 0 19392 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_203
timestamp 1679585382
transform 1 0 20064 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_210
timestamp 1679585382
transform 1 0 20736 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_217
timestamp 1679585382
transform 1 0 21408 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_224
timestamp 1679585382
transform 1 0 22080 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_231
timestamp 1679585382
transform 1 0 22752 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_238
timestamp 1679585382
transform 1 0 23424 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_245
timestamp 1679585382
transform 1 0 24096 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_252
timestamp 1679585382
transform 1 0 24768 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_259
timestamp 1679585382
transform 1 0 25440 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_266
timestamp 1679585382
transform 1 0 26112 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_273
timestamp 1679585382
transform 1 0 26784 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_280
timestamp 1679585382
transform 1 0 27456 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_287
timestamp 1679581501
transform 1 0 28128 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_291
timestamp 1677583258
transform 1 0 28512 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_296
timestamp 1679585382
transform 1 0 28992 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_303
timestamp 1679585382
transform 1 0 29664 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_310
timestamp 1679585382
transform 1 0 30336 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_317
timestamp 1679585382
transform 1 0 31008 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_324
timestamp 1679585382
transform 1 0 31680 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_331
timestamp 1679585382
transform 1 0 32352 0 1 26460
box -48 -56 720 834
use sg13g2_fill_1  FILLER_34_338
timestamp 1677583258
transform 1 0 33024 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_375
timestamp 1679585382
transform 1 0 36576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_382
timestamp 1679585382
transform 1 0 37248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_389
timestamp 1679585382
transform 1 0 37920 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_396
timestamp 1679585382
transform 1 0 38592 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_403
timestamp 1679585382
transform 1 0 39264 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_410
timestamp 1677583704
transform 1 0 39936 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_412
timestamp 1677583258
transform 1 0 40128 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_449
timestamp 1679585382
transform 1 0 43680 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_456
timestamp 1679585382
transform 1 0 44352 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_463
timestamp 1679585382
transform 1 0 45024 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_470
timestamp 1679585382
transform 1 0 45696 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_477
timestamp 1679585382
transform 1 0 46368 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_484
timestamp 1679585382
transform 1 0 47040 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_491
timestamp 1679585382
transform 1 0 47712 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_498
timestamp 1679585382
transform 1 0 48384 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_505
timestamp 1679585382
transform 1 0 49056 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_512
timestamp 1679585382
transform 1 0 49728 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_519
timestamp 1679585382
transform 1 0 50400 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_526
timestamp 1679585382
transform 1 0 51072 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_533
timestamp 1679585382
transform 1 0 51744 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_540
timestamp 1679585382
transform 1 0 52416 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_547
timestamp 1679585382
transform 1 0 53088 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_554
timestamp 1679585382
transform 1 0 53760 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_561
timestamp 1679585382
transform 1 0 54432 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_568
timestamp 1679585382
transform 1 0 55104 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_575
timestamp 1679585382
transform 1 0 55776 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_582
timestamp 1679585382
transform 1 0 56448 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_589
timestamp 1679585382
transform 1 0 57120 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_596
timestamp 1679585382
transform 1 0 57792 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_603
timestamp 1679585382
transform 1 0 58464 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_610
timestamp 1679585382
transform 1 0 59136 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_617
timestamp 1679585382
transform 1 0 59808 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_624
timestamp 1679585382
transform 1 0 60480 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_631
timestamp 1679585382
transform 1 0 61152 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_638
timestamp 1679585382
transform 1 0 61824 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_645
timestamp 1679585382
transform 1 0 62496 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_652
timestamp 1679585382
transform 1 0 63168 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_659
timestamp 1679585382
transform 1 0 63840 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_666
timestamp 1679585382
transform 1 0 64512 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_673
timestamp 1679585382
transform 1 0 65184 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_680
timestamp 1679585382
transform 1 0 65856 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_687
timestamp 1679585382
transform 1 0 66528 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_694
timestamp 1679585382
transform 1 0 67200 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_701
timestamp 1679585382
transform 1 0 67872 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_708
timestamp 1679585382
transform 1 0 68544 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_715
timestamp 1679585382
transform 1 0 69216 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_722
timestamp 1679585382
transform 1 0 69888 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_729
timestamp 1679585382
transform 1 0 70560 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_736
timestamp 1679585382
transform 1 0 71232 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_743
timestamp 1679585382
transform 1 0 71904 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_750
timestamp 1679585382
transform 1 0 72576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_757
timestamp 1679585382
transform 1 0 73248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_764
timestamp 1679585382
transform 1 0 73920 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_771
timestamp 1679585382
transform 1 0 74592 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_778
timestamp 1679585382
transform 1 0 75264 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_785
timestamp 1679585382
transform 1 0 75936 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_792
timestamp 1679585382
transform 1 0 76608 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_799
timestamp 1679585382
transform 1 0 77280 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_806
timestamp 1679585382
transform 1 0 77952 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_813
timestamp 1679585382
transform 1 0 78624 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_820
timestamp 1679585382
transform 1 0 79296 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_827
timestamp 1679585382
transform 1 0 79968 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_834
timestamp 1679585382
transform 1 0 80640 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_841
timestamp 1679585382
transform 1 0 81312 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_848
timestamp 1679585382
transform 1 0 81984 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_855
timestamp 1679585382
transform 1 0 82656 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_862
timestamp 1679585382
transform 1 0 83328 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_869
timestamp 1679585382
transform 1 0 84000 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_876
timestamp 1679585382
transform 1 0 84672 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_883
timestamp 1679585382
transform 1 0 85344 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_890
timestamp 1679585382
transform 1 0 86016 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_897
timestamp 1679585382
transform 1 0 86688 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_904
timestamp 1679585382
transform 1 0 87360 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_911
timestamp 1679585382
transform 1 0 88032 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_918
timestamp 1679585382
transform 1 0 88704 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_925
timestamp 1679585382
transform 1 0 89376 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_932
timestamp 1679585382
transform 1 0 90048 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_939
timestamp 1679585382
transform 1 0 90720 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_946
timestamp 1679585382
transform 1 0 91392 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_953
timestamp 1679585382
transform 1 0 92064 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_960
timestamp 1679585382
transform 1 0 92736 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_967
timestamp 1679585382
transform 1 0 93408 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_974
timestamp 1679585382
transform 1 0 94080 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_981
timestamp 1679585382
transform 1 0 94752 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_988
timestamp 1679585382
transform 1 0 95424 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_995
timestamp 1679585382
transform 1 0 96096 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1002
timestamp 1679585382
transform 1 0 96768 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1009
timestamp 1679585382
transform 1 0 97440 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_1016
timestamp 1679585382
transform 1 0 98112 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_1023
timestamp 1679581501
transform 1 0 98784 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_1027
timestamp 1677583704
transform 1 0 99168 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_0
timestamp 1679585382
transform 1 0 576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_7
timestamp 1679585382
transform 1 0 1248 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_14
timestamp 1679585382
transform 1 0 1920 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_21
timestamp 1679585382
transform 1 0 2592 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_28
timestamp 1679585382
transform 1 0 3264 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_35
timestamp 1677583704
transform 1 0 3936 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_58
timestamp 1679585382
transform 1 0 6144 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_65
timestamp 1679585382
transform 1 0 6816 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_72
timestamp 1679585382
transform 1 0 7488 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_79
timestamp 1679581501
transform 1 0 8160 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_83
timestamp 1677583704
transform 1 0 8544 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_98
timestamp 1679585382
transform 1 0 9984 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_35_105
timestamp 1677583258
transform 1 0 10656 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_123
timestamp 1679585382
transform 1 0 12384 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_130
timestamp 1679585382
transform 1 0 13056 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_137
timestamp 1679585382
transform 1 0 13728 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_144
timestamp 1679585382
transform 1 0 14400 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_151
timestamp 1679585382
transform 1 0 15072 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_158
timestamp 1679585382
transform 1 0 15744 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_165
timestamp 1679585382
transform 1 0 16416 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_172
timestamp 1679585382
transform 1 0 17088 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_179
timestamp 1679585382
transform 1 0 17760 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_186
timestamp 1679585382
transform 1 0 18432 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_193
timestamp 1679585382
transform 1 0 19104 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_200
timestamp 1679585382
transform 1 0 19776 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_207
timestamp 1679585382
transform 1 0 20448 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_214
timestamp 1679585382
transform 1 0 21120 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_221
timestamp 1679585382
transform 1 0 21792 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_228
timestamp 1679585382
transform 1 0 22464 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_235
timestamp 1679585382
transform 1 0 23136 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_242
timestamp 1679585382
transform 1 0 23808 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_249
timestamp 1679585382
transform 1 0 24480 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_256
timestamp 1679585382
transform 1 0 25152 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_263
timestamp 1677583704
transform 1 0 25824 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_265
timestamp 1677583258
transform 1 0 26016 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_302
timestamp 1679585382
transform 1 0 29568 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_309
timestamp 1679585382
transform 1 0 30240 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_316
timestamp 1679585382
transform 1 0 30912 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_323
timestamp 1679585382
transform 1 0 31584 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_330
timestamp 1677583704
transform 1 0 32256 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_359
timestamp 1679585382
transform 1 0 35040 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_366
timestamp 1679585382
transform 1 0 35712 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_373
timestamp 1679585382
transform 1 0 36384 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_380
timestamp 1679585382
transform 1 0 37056 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_387
timestamp 1679581501
transform 1 0 37728 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_391
timestamp 1677583704
transform 1 0 38112 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_421
timestamp 1679585382
transform 1 0 40992 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_428
timestamp 1679585382
transform 1 0 41664 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_435
timestamp 1679585382
transform 1 0 42336 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_442
timestamp 1679585382
transform 1 0 43008 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_449
timestamp 1679585382
transform 1 0 43680 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_456
timestamp 1679585382
transform 1 0 44352 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_463
timestamp 1679585382
transform 1 0 45024 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_470
timestamp 1679585382
transform 1 0 45696 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_477
timestamp 1679585382
transform 1 0 46368 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_484
timestamp 1679585382
transform 1 0 47040 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_491
timestamp 1679585382
transform 1 0 47712 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_498
timestamp 1679585382
transform 1 0 48384 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_505
timestamp 1679585382
transform 1 0 49056 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_512
timestamp 1679585382
transform 1 0 49728 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_519
timestamp 1679585382
transform 1 0 50400 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_526
timestamp 1679585382
transform 1 0 51072 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_533
timestamp 1679585382
transform 1 0 51744 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_540
timestamp 1679585382
transform 1 0 52416 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_547
timestamp 1679585382
transform 1 0 53088 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_554
timestamp 1679585382
transform 1 0 53760 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_561
timestamp 1679585382
transform 1 0 54432 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_568
timestamp 1679585382
transform 1 0 55104 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_575
timestamp 1679585382
transform 1 0 55776 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_582
timestamp 1679585382
transform 1 0 56448 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_589
timestamp 1679585382
transform 1 0 57120 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_596
timestamp 1679585382
transform 1 0 57792 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_603
timestamp 1679585382
transform 1 0 58464 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_610
timestamp 1679585382
transform 1 0 59136 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_617
timestamp 1679585382
transform 1 0 59808 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_624
timestamp 1679585382
transform 1 0 60480 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_631
timestamp 1679585382
transform 1 0 61152 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_638
timestamp 1679585382
transform 1 0 61824 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_645
timestamp 1679585382
transform 1 0 62496 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_652
timestamp 1679585382
transform 1 0 63168 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_659
timestamp 1679585382
transform 1 0 63840 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_666
timestamp 1679585382
transform 1 0 64512 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_673
timestamp 1679585382
transform 1 0 65184 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_680
timestamp 1679585382
transform 1 0 65856 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_687
timestamp 1679585382
transform 1 0 66528 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_694
timestamp 1679585382
transform 1 0 67200 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_701
timestamp 1679585382
transform 1 0 67872 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_708
timestamp 1679585382
transform 1 0 68544 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_715
timestamp 1679585382
transform 1 0 69216 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_722
timestamp 1679585382
transform 1 0 69888 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_729
timestamp 1679585382
transform 1 0 70560 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_736
timestamp 1679585382
transform 1 0 71232 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_743
timestamp 1679585382
transform 1 0 71904 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_750
timestamp 1679585382
transform 1 0 72576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_757
timestamp 1679585382
transform 1 0 73248 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_764
timestamp 1679585382
transform 1 0 73920 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_771
timestamp 1679585382
transform 1 0 74592 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_778
timestamp 1679585382
transform 1 0 75264 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_785
timestamp 1679585382
transform 1 0 75936 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_792
timestamp 1679585382
transform 1 0 76608 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_799
timestamp 1679585382
transform 1 0 77280 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_806
timestamp 1679585382
transform 1 0 77952 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_813
timestamp 1679585382
transform 1 0 78624 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_820
timestamp 1679585382
transform 1 0 79296 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_827
timestamp 1679585382
transform 1 0 79968 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_834
timestamp 1679585382
transform 1 0 80640 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_841
timestamp 1679585382
transform 1 0 81312 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_848
timestamp 1679585382
transform 1 0 81984 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_855
timestamp 1679585382
transform 1 0 82656 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_862
timestamp 1679585382
transform 1 0 83328 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_869
timestamp 1679585382
transform 1 0 84000 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_876
timestamp 1679585382
transform 1 0 84672 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_883
timestamp 1679585382
transform 1 0 85344 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_890
timestamp 1679585382
transform 1 0 86016 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_897
timestamp 1679585382
transform 1 0 86688 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_904
timestamp 1679585382
transform 1 0 87360 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_911
timestamp 1679585382
transform 1 0 88032 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_918
timestamp 1679585382
transform 1 0 88704 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_925
timestamp 1679585382
transform 1 0 89376 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_932
timestamp 1679585382
transform 1 0 90048 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_939
timestamp 1679585382
transform 1 0 90720 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_946
timestamp 1679585382
transform 1 0 91392 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_953
timestamp 1679585382
transform 1 0 92064 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_960
timestamp 1679585382
transform 1 0 92736 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_967
timestamp 1679585382
transform 1 0 93408 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_974
timestamp 1679585382
transform 1 0 94080 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_981
timestamp 1679585382
transform 1 0 94752 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_988
timestamp 1679585382
transform 1 0 95424 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_995
timestamp 1679585382
transform 1 0 96096 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1002
timestamp 1679585382
transform 1 0 96768 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1009
timestamp 1679585382
transform 1 0 97440 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_1016
timestamp 1679585382
transform 1 0 98112 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_35_1023
timestamp 1679581501
transform 1 0 98784 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_1027
timestamp 1677583704
transform 1 0 99168 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_0
timestamp 1679585382
transform 1 0 576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_7
timestamp 1679585382
transform 1 0 1248 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_14
timestamp 1679585382
transform 1 0 1920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_21
timestamp 1679585382
transform 1 0 2592 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_28
timestamp 1679585382
transform 1 0 3264 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_35
timestamp 1679585382
transform 1 0 3936 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_42
timestamp 1679585382
transform 1 0 4608 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_49
timestamp 1679585382
transform 1 0 5280 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_56
timestamp 1679585382
transform 1 0 5952 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_63
timestamp 1679585382
transform 1 0 6624 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_70
timestamp 1679585382
transform 1 0 7296 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_77
timestamp 1679585382
transform 1 0 7968 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_84
timestamp 1679585382
transform 1 0 8640 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_91
timestamp 1679585382
transform 1 0 9312 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_98
timestamp 1679585382
transform 1 0 9984 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_105
timestamp 1679585382
transform 1 0 10656 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_112
timestamp 1679585382
transform 1 0 11328 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_119
timestamp 1679585382
transform 1 0 12000 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_126
timestamp 1679585382
transform 1 0 12672 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_133
timestamp 1679585382
transform 1 0 13344 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_140
timestamp 1679585382
transform 1 0 14016 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_147
timestamp 1679585382
transform 1 0 14688 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_154
timestamp 1679585382
transform 1 0 15360 0 1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_36_161
timestamp 1677583258
transform 1 0 16032 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_166
timestamp 1679585382
transform 1 0 16512 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_173
timestamp 1679585382
transform 1 0 17184 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_180
timestamp 1679585382
transform 1 0 17856 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_187
timestamp 1679585382
transform 1 0 18528 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_211
timestamp 1679585382
transform 1 0 20832 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_218
timestamp 1679585382
transform 1 0 21504 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_225
timestamp 1679585382
transform 1 0 22176 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_232
timestamp 1679585382
transform 1 0 22848 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_239
timestamp 1679585382
transform 1 0 23520 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_246
timestamp 1679585382
transform 1 0 24192 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_253
timestamp 1679585382
transform 1 0 24864 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_260
timestamp 1679585382
transform 1 0 25536 0 1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_36_267
timestamp 1677583704
transform 1 0 26208 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_278
timestamp 1679585382
transform 1 0 27264 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_285
timestamp 1679585382
transform 1 0 27936 0 1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_36_292
timestamp 1677583258
transform 1 0 28608 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_301
timestamp 1679585382
transform 1 0 29472 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_308
timestamp 1679585382
transform 1 0 30144 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_315
timestamp 1679585382
transform 1 0 30816 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_322
timestamp 1679585382
transform 1 0 31488 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_329
timestamp 1679581501
transform 1 0 32160 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_333
timestamp 1677583704
transform 1 0 32544 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_348
timestamp 1679585382
transform 1 0 33984 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_355
timestamp 1679585382
transform 1 0 34656 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_362
timestamp 1679585382
transform 1 0 35328 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_369
timestamp 1679585382
transform 1 0 36000 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_376
timestamp 1679585382
transform 1 0 36672 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_383
timestamp 1679585382
transform 1 0 37344 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_390
timestamp 1679585382
transform 1 0 38016 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_397
timestamp 1679585382
transform 1 0 38688 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_404
timestamp 1679581501
transform 1 0 39360 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_408
timestamp 1677583704
transform 1 0 39744 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_423
timestamp 1679585382
transform 1 0 41184 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_430
timestamp 1679585382
transform 1 0 41856 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_437
timestamp 1679585382
transform 1 0 42528 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_444
timestamp 1679585382
transform 1 0 43200 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_451
timestamp 1679581501
transform 1 0 43872 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_455
timestamp 1677583704
transform 1 0 44256 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_484
timestamp 1679585382
transform 1 0 47040 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_491
timestamp 1679585382
transform 1 0 47712 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_498
timestamp 1679585382
transform 1 0 48384 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_505
timestamp 1679585382
transform 1 0 49056 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_512
timestamp 1679585382
transform 1 0 49728 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_519
timestamp 1679585382
transform 1 0 50400 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_526
timestamp 1679585382
transform 1 0 51072 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_533
timestamp 1679585382
transform 1 0 51744 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_540
timestamp 1679585382
transform 1 0 52416 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_547
timestamp 1679585382
transform 1 0 53088 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_554
timestamp 1679585382
transform 1 0 53760 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_561
timestamp 1679585382
transform 1 0 54432 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_568
timestamp 1679585382
transform 1 0 55104 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_575
timestamp 1679585382
transform 1 0 55776 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_582
timestamp 1679585382
transform 1 0 56448 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_589
timestamp 1679585382
transform 1 0 57120 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_596
timestamp 1679585382
transform 1 0 57792 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_603
timestamp 1679585382
transform 1 0 58464 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_610
timestamp 1679585382
transform 1 0 59136 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_617
timestamp 1679585382
transform 1 0 59808 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_624
timestamp 1679585382
transform 1 0 60480 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_631
timestamp 1679585382
transform 1 0 61152 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_638
timestamp 1679585382
transform 1 0 61824 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_645
timestamp 1679585382
transform 1 0 62496 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_652
timestamp 1679585382
transform 1 0 63168 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_659
timestamp 1679585382
transform 1 0 63840 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_666
timestamp 1679585382
transform 1 0 64512 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_673
timestamp 1679585382
transform 1 0 65184 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_680
timestamp 1679585382
transform 1 0 65856 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_687
timestamp 1679585382
transform 1 0 66528 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_694
timestamp 1679585382
transform 1 0 67200 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_701
timestamp 1679585382
transform 1 0 67872 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_708
timestamp 1679585382
transform 1 0 68544 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_715
timestamp 1679585382
transform 1 0 69216 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_722
timestamp 1679585382
transform 1 0 69888 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_729
timestamp 1679585382
transform 1 0 70560 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_736
timestamp 1679585382
transform 1 0 71232 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_743
timestamp 1679585382
transform 1 0 71904 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_750
timestamp 1679585382
transform 1 0 72576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_757
timestamp 1679585382
transform 1 0 73248 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_764
timestamp 1679585382
transform 1 0 73920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_771
timestamp 1679585382
transform 1 0 74592 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_778
timestamp 1679585382
transform 1 0 75264 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_785
timestamp 1679585382
transform 1 0 75936 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_792
timestamp 1679585382
transform 1 0 76608 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_799
timestamp 1679585382
transform 1 0 77280 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_806
timestamp 1679585382
transform 1 0 77952 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_813
timestamp 1679585382
transform 1 0 78624 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_820
timestamp 1679585382
transform 1 0 79296 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_827
timestamp 1679585382
transform 1 0 79968 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_834
timestamp 1679585382
transform 1 0 80640 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_841
timestamp 1679585382
transform 1 0 81312 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_848
timestamp 1679585382
transform 1 0 81984 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_855
timestamp 1679585382
transform 1 0 82656 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_862
timestamp 1679585382
transform 1 0 83328 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_869
timestamp 1679585382
transform 1 0 84000 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_876
timestamp 1679585382
transform 1 0 84672 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_883
timestamp 1679585382
transform 1 0 85344 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_890
timestamp 1679585382
transform 1 0 86016 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_897
timestamp 1679585382
transform 1 0 86688 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_904
timestamp 1679585382
transform 1 0 87360 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_911
timestamp 1679585382
transform 1 0 88032 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_918
timestamp 1679585382
transform 1 0 88704 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_925
timestamp 1679585382
transform 1 0 89376 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_932
timestamp 1679585382
transform 1 0 90048 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_939
timestamp 1679585382
transform 1 0 90720 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_946
timestamp 1679585382
transform 1 0 91392 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_953
timestamp 1679585382
transform 1 0 92064 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_960
timestamp 1679585382
transform 1 0 92736 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_967
timestamp 1679585382
transform 1 0 93408 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_974
timestamp 1679585382
transform 1 0 94080 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_981
timestamp 1679585382
transform 1 0 94752 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_988
timestamp 1679585382
transform 1 0 95424 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_995
timestamp 1679585382
transform 1 0 96096 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1002
timestamp 1679585382
transform 1 0 96768 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1009
timestamp 1679585382
transform 1 0 97440 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_1016
timestamp 1679585382
transform 1 0 98112 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_1023
timestamp 1679581501
transform 1 0 98784 0 1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_36_1027
timestamp 1677583704
transform 1 0 99168 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_37_0
timestamp 1679585382
transform 1 0 576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_7
timestamp 1679585382
transform 1 0 1248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_14
timestamp 1679585382
transform 1 0 1920 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_21
timestamp 1677583258
transform 1 0 2592 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_49
timestamp 1679585382
transform 1 0 5280 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_56
timestamp 1679585382
transform 1 0 5952 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_63
timestamp 1679585382
transform 1 0 6624 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_70
timestamp 1679581501
transform 1 0 7296 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_37_74
timestamp 1677583258
transform 1 0 7680 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_102
timestamp 1679585382
transform 1 0 10368 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_109
timestamp 1677583258
transform 1 0 11040 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_119
timestamp 1679585382
transform 1 0 12000 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_126
timestamp 1679585382
transform 1 0 12672 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_133
timestamp 1679585382
transform 1 0 13344 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_140
timestamp 1679585382
transform 1 0 14016 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_147
timestamp 1677583704
transform 1 0 14688 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_149
timestamp 1677583258
transform 1 0 14880 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_181
timestamp 1679585382
transform 1 0 17952 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_188
timestamp 1679585382
transform 1 0 18624 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_195
timestamp 1679585382
transform 1 0 19296 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_202
timestamp 1679585382
transform 1 0 19968 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_209
timestamp 1679585382
transform 1 0 20640 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_216
timestamp 1679585382
transform 1 0 21312 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_223
timestamp 1677583258
transform 1 0 21984 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_237
timestamp 1679585382
transform 1 0 23328 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_244
timestamp 1679585382
transform 1 0 24000 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_251
timestamp 1679585382
transform 1 0 24672 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_258
timestamp 1679585382
transform 1 0 25344 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_274
timestamp 1679585382
transform 1 0 26880 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_281
timestamp 1679585382
transform 1 0 27552 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_288
timestamp 1679585382
transform 1 0 28224 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_295
timestamp 1679585382
transform 1 0 28896 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_302
timestamp 1677583704
transform 1 0 29568 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_304
timestamp 1677583258
transform 1 0 29760 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_314
timestamp 1679585382
transform 1 0 30720 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_321
timestamp 1679585382
transform 1 0 31392 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_328
timestamp 1679585382
transform 1 0 32064 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_335
timestamp 1679585382
transform 1 0 32736 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_342
timestamp 1679585382
transform 1 0 33408 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_349
timestamp 1679585382
transform 1 0 34080 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_356
timestamp 1679585382
transform 1 0 34752 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_363
timestamp 1679585382
transform 1 0 35424 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_370
timestamp 1679585382
transform 1 0 36096 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_377
timestamp 1679585382
transform 1 0 36768 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_384
timestamp 1679585382
transform 1 0 37440 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_391
timestamp 1679585382
transform 1 0 38112 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_398
timestamp 1679585382
transform 1 0 38784 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_405
timestamp 1677583704
transform 1 0 39456 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_407
timestamp 1677583258
transform 1 0 39648 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_421
timestamp 1679585382
transform 1 0 40992 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_428
timestamp 1679585382
transform 1 0 41664 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_435
timestamp 1679585382
transform 1 0 42336 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_442
timestamp 1679585382
transform 1 0 43008 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_449
timestamp 1679585382
transform 1 0 43680 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_469
timestamp 1679585382
transform 1 0 45600 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_476
timestamp 1679585382
transform 1 0 46272 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_483
timestamp 1679585382
transform 1 0 46944 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_490
timestamp 1679585382
transform 1 0 47616 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_497
timestamp 1679585382
transform 1 0 48288 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_504
timestamp 1679585382
transform 1 0 48960 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_511
timestamp 1679585382
transform 1 0 49632 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_518
timestamp 1679585382
transform 1 0 50304 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_525
timestamp 1679585382
transform 1 0 50976 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_532
timestamp 1679585382
transform 1 0 51648 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_539
timestamp 1679585382
transform 1 0 52320 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_546
timestamp 1679585382
transform 1 0 52992 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_553
timestamp 1679585382
transform 1 0 53664 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_560
timestamp 1679585382
transform 1 0 54336 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_567
timestamp 1679585382
transform 1 0 55008 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_574
timestamp 1679585382
transform 1 0 55680 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_581
timestamp 1679585382
transform 1 0 56352 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_588
timestamp 1679585382
transform 1 0 57024 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_595
timestamp 1679585382
transform 1 0 57696 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_602
timestamp 1679585382
transform 1 0 58368 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_609
timestamp 1679585382
transform 1 0 59040 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_616
timestamp 1679585382
transform 1 0 59712 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_623
timestamp 1679585382
transform 1 0 60384 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_630
timestamp 1679585382
transform 1 0 61056 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_637
timestamp 1679585382
transform 1 0 61728 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_644
timestamp 1679585382
transform 1 0 62400 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_651
timestamp 1679585382
transform 1 0 63072 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_658
timestamp 1679585382
transform 1 0 63744 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_665
timestamp 1679585382
transform 1 0 64416 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_672
timestamp 1679585382
transform 1 0 65088 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_679
timestamp 1679585382
transform 1 0 65760 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_686
timestamp 1679585382
transform 1 0 66432 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_693
timestamp 1679585382
transform 1 0 67104 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_700
timestamp 1679585382
transform 1 0 67776 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_707
timestamp 1679585382
transform 1 0 68448 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_714
timestamp 1679585382
transform 1 0 69120 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_721
timestamp 1679585382
transform 1 0 69792 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_728
timestamp 1679585382
transform 1 0 70464 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_735
timestamp 1679585382
transform 1 0 71136 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_742
timestamp 1679585382
transform 1 0 71808 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_749
timestamp 1679585382
transform 1 0 72480 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_756
timestamp 1679585382
transform 1 0 73152 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_763
timestamp 1679585382
transform 1 0 73824 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_770
timestamp 1679585382
transform 1 0 74496 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_777
timestamp 1679585382
transform 1 0 75168 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_784
timestamp 1679585382
transform 1 0 75840 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_791
timestamp 1679585382
transform 1 0 76512 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_798
timestamp 1679585382
transform 1 0 77184 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_805
timestamp 1679585382
transform 1 0 77856 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_812
timestamp 1679585382
transform 1 0 78528 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_819
timestamp 1679585382
transform 1 0 79200 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_826
timestamp 1679585382
transform 1 0 79872 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_833
timestamp 1679585382
transform 1 0 80544 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_840
timestamp 1679585382
transform 1 0 81216 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_847
timestamp 1679585382
transform 1 0 81888 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_854
timestamp 1679585382
transform 1 0 82560 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_861
timestamp 1679585382
transform 1 0 83232 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_868
timestamp 1679585382
transform 1 0 83904 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_875
timestamp 1679585382
transform 1 0 84576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_882
timestamp 1679585382
transform 1 0 85248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_889
timestamp 1679585382
transform 1 0 85920 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_896
timestamp 1679585382
transform 1 0 86592 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_903
timestamp 1679585382
transform 1 0 87264 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_910
timestamp 1679585382
transform 1 0 87936 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_917
timestamp 1679585382
transform 1 0 88608 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_924
timestamp 1679585382
transform 1 0 89280 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_931
timestamp 1679585382
transform 1 0 89952 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_938
timestamp 1679585382
transform 1 0 90624 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_945
timestamp 1679585382
transform 1 0 91296 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_952
timestamp 1679585382
transform 1 0 91968 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_959
timestamp 1679585382
transform 1 0 92640 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_966
timestamp 1679585382
transform 1 0 93312 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_973
timestamp 1679585382
transform 1 0 93984 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_980
timestamp 1679585382
transform 1 0 94656 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_987
timestamp 1679585382
transform 1 0 95328 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_994
timestamp 1679585382
transform 1 0 96000 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1001
timestamp 1679585382
transform 1 0 96672 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1008
timestamp 1679585382
transform 1 0 97344 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1015
timestamp 1679585382
transform 1 0 98016 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_1022
timestamp 1679585382
transform 1 0 98688 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_0
timestamp 1679585382
transform 1 0 576 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_7
timestamp 1679585382
transform 1 0 1248 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_14
timestamp 1679585382
transform 1 0 1920 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_21
timestamp 1679585382
transform 1 0 2592 0 1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_38_28
timestamp 1677583704
transform 1 0 3264 0 1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_38
timestamp 1677583704
transform 1 0 4224 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_40
timestamp 1677583258
transform 1 0 4416 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_50
timestamp 1679585382
transform 1 0 5376 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_57
timestamp 1679585382
transform 1 0 6048 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_64
timestamp 1679585382
transform 1 0 6720 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_71
timestamp 1679585382
transform 1 0 7392 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_78
timestamp 1679585382
transform 1 0 8064 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_85
timestamp 1679581501
transform 1 0 8736 0 1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_38_102
timestamp 1677583258
transform 1 0 10368 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_111
timestamp 1679585382
transform 1 0 11232 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_118
timestamp 1679585382
transform 1 0 11904 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_125
timestamp 1679585382
transform 1 0 12576 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_132
timestamp 1679585382
transform 1 0 13248 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_139
timestamp 1679581501
transform 1 0 13920 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_170
timestamp 1677583704
transform 1 0 16896 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_172
timestamp 1677583258
transform 1 0 17088 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_182
timestamp 1679585382
transform 1 0 18048 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_189
timestamp 1679585382
transform 1 0 18720 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_196
timestamp 1679585382
transform 1 0 19392 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_203
timestamp 1679585382
transform 1 0 20064 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_237
timestamp 1679585382
transform 1 0 23328 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_244
timestamp 1679585382
transform 1 0 24000 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_251
timestamp 1679581501
transform 1 0 24672 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_255
timestamp 1677583704
transform 1 0 25056 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_305
timestamp 1677583258
transform 1 0 29856 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_314
timestamp 1679585382
transform 1 0 30720 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_321
timestamp 1679585382
transform 1 0 31392 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_328
timestamp 1679585382
transform 1 0 32064 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_335
timestamp 1679585382
transform 1 0 32736 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_342
timestamp 1679585382
transform 1 0 33408 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_349
timestamp 1679585382
transform 1 0 34080 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_356
timestamp 1679585382
transform 1 0 34752 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_363
timestamp 1679585382
transform 1 0 35424 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_370
timestamp 1679585382
transform 1 0 36096 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_377
timestamp 1679585382
transform 1 0 36768 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_384
timestamp 1679585382
transform 1 0 37440 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_391
timestamp 1679585382
transform 1 0 38112 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_398
timestamp 1679585382
transform 1 0 38784 0 1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_38_405
timestamp 1677583258
transform 1 0 39456 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_415
timestamp 1679585382
transform 1 0 40416 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_422
timestamp 1679585382
transform 1 0 41088 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_429
timestamp 1679585382
transform 1 0 41760 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_436
timestamp 1679585382
transform 1 0 42432 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_443
timestamp 1679585382
transform 1 0 43104 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_450
timestamp 1679585382
transform 1 0 43776 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_477
timestamp 1679581501
transform 1 0 46368 0 1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_38_481
timestamp 1677583258
transform 1 0 46752 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_509
timestamp 1679585382
transform 1 0 49440 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_516
timestamp 1679585382
transform 1 0 50112 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_523
timestamp 1679585382
transform 1 0 50784 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_530
timestamp 1679585382
transform 1 0 51456 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_537
timestamp 1679585382
transform 1 0 52128 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_544
timestamp 1679585382
transform 1 0 52800 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_551
timestamp 1679585382
transform 1 0 53472 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_558
timestamp 1679585382
transform 1 0 54144 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_565
timestamp 1679585382
transform 1 0 54816 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_572
timestamp 1679585382
transform 1 0 55488 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_579
timestamp 1679585382
transform 1 0 56160 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_586
timestamp 1679585382
transform 1 0 56832 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_593
timestamp 1679585382
transform 1 0 57504 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_600
timestamp 1679585382
transform 1 0 58176 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_607
timestamp 1679585382
transform 1 0 58848 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_614
timestamp 1679585382
transform 1 0 59520 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_621
timestamp 1679585382
transform 1 0 60192 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_628
timestamp 1679585382
transform 1 0 60864 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_635
timestamp 1679585382
transform 1 0 61536 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_642
timestamp 1679585382
transform 1 0 62208 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_649
timestamp 1679585382
transform 1 0 62880 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_656
timestamp 1679585382
transform 1 0 63552 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_663
timestamp 1679585382
transform 1 0 64224 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_670
timestamp 1679585382
transform 1 0 64896 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_677
timestamp 1679585382
transform 1 0 65568 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_684
timestamp 1679585382
transform 1 0 66240 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_691
timestamp 1679585382
transform 1 0 66912 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_698
timestamp 1679585382
transform 1 0 67584 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_705
timestamp 1679585382
transform 1 0 68256 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_712
timestamp 1679585382
transform 1 0 68928 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_719
timestamp 1679585382
transform 1 0 69600 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_726
timestamp 1679585382
transform 1 0 70272 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_733
timestamp 1679585382
transform 1 0 70944 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_740
timestamp 1679585382
transform 1 0 71616 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_747
timestamp 1679585382
transform 1 0 72288 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_754
timestamp 1679585382
transform 1 0 72960 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_761
timestamp 1679585382
transform 1 0 73632 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_768
timestamp 1679585382
transform 1 0 74304 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_775
timestamp 1679585382
transform 1 0 74976 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_782
timestamp 1679585382
transform 1 0 75648 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_789
timestamp 1679585382
transform 1 0 76320 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_796
timestamp 1679585382
transform 1 0 76992 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_803
timestamp 1679585382
transform 1 0 77664 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_810
timestamp 1679585382
transform 1 0 78336 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_817
timestamp 1679585382
transform 1 0 79008 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_824
timestamp 1679585382
transform 1 0 79680 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_831
timestamp 1679585382
transform 1 0 80352 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_838
timestamp 1679585382
transform 1 0 81024 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_845
timestamp 1679585382
transform 1 0 81696 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_852
timestamp 1679585382
transform 1 0 82368 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_859
timestamp 1679585382
transform 1 0 83040 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_866
timestamp 1679585382
transform 1 0 83712 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_873
timestamp 1679585382
transform 1 0 84384 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_880
timestamp 1679585382
transform 1 0 85056 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_887
timestamp 1679585382
transform 1 0 85728 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_894
timestamp 1679585382
transform 1 0 86400 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_901
timestamp 1679585382
transform 1 0 87072 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_908
timestamp 1679585382
transform 1 0 87744 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_915
timestamp 1679585382
transform 1 0 88416 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_922
timestamp 1679585382
transform 1 0 89088 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_929
timestamp 1679585382
transform 1 0 89760 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_936
timestamp 1679585382
transform 1 0 90432 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_943
timestamp 1679585382
transform 1 0 91104 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_950
timestamp 1679585382
transform 1 0 91776 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_957
timestamp 1679585382
transform 1 0 92448 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_964
timestamp 1679585382
transform 1 0 93120 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_971
timestamp 1679585382
transform 1 0 93792 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_978
timestamp 1679585382
transform 1 0 94464 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_985
timestamp 1679585382
transform 1 0 95136 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_992
timestamp 1679585382
transform 1 0 95808 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_999
timestamp 1679585382
transform 1 0 96480 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1006
timestamp 1679585382
transform 1 0 97152 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1013
timestamp 1679585382
transform 1 0 97824 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_1020
timestamp 1679585382
transform 1 0 98496 0 1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_38_1027
timestamp 1677583704
transform 1 0 99168 0 1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_0
timestamp 1679585382
transform 1 0 576 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_7
timestamp 1679585382
transform 1 0 1248 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_14
timestamp 1679585382
transform 1 0 1920 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_21
timestamp 1677583704
transform 1 0 2592 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_59
timestamp 1679585382
transform 1 0 6240 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_66
timestamp 1679585382
transform 1 0 6912 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_73
timestamp 1679585382
transform 1 0 7584 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_80
timestamp 1679585382
transform 1 0 8256 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_87
timestamp 1679585382
transform 1 0 8928 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_94
timestamp 1679585382
transform 1 0 9600 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_101
timestamp 1679585382
transform 1 0 10272 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_108
timestamp 1679585382
transform 1 0 10944 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_115
timestamp 1679585382
transform 1 0 11616 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_122
timestamp 1679585382
transform 1 0 12288 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_129
timestamp 1679585382
transform 1 0 12960 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_136
timestamp 1679585382
transform 1 0 13632 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_143
timestamp 1679585382
transform 1 0 14304 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_150
timestamp 1677583704
transform 1 0 14976 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_4  FILLER_39_156
timestamp 1679581501
transform 1 0 15552 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_39_160
timestamp 1677583704
transform 1 0 15936 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_188
timestamp 1679585382
transform 1 0 18624 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_195
timestamp 1679585382
transform 1 0 19296 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_39_202
timestamp 1677583258
transform 1 0 19968 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_230
timestamp 1679585382
transform 1 0 22656 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_237
timestamp 1679585382
transform 1 0 23328 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_244
timestamp 1677583704
transform 1 0 24000 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_4  FILLER_39_267
timestamp 1679581501
transform 1 0 26208 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_39_271
timestamp 1677583258
transform 1 0 26592 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_281
timestamp 1679585382
transform 1 0 27552 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_288
timestamp 1679585382
transform 1 0 28224 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_295
timestamp 1679585382
transform 1 0 28896 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_302
timestamp 1679585382
transform 1 0 29568 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_39_309
timestamp 1677583258
transform 1 0 30240 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_337
timestamp 1679585382
transform 1 0 32928 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_344
timestamp 1679581501
transform 1 0 33600 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_39_348
timestamp 1677583258
transform 1 0 33984 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_362
timestamp 1677583704
transform 1 0 35328 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_364
timestamp 1677583258
transform 1 0 35520 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_395
timestamp 1679585382
transform 1 0 38496 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_402
timestamp 1677583704
transform 1 0 39168 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_431
timestamp 1679585382
transform 1 0 41952 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_438
timestamp 1679585382
transform 1 0 42624 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_445
timestamp 1679585382
transform 1 0 43296 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_452
timestamp 1679585382
transform 1 0 43968 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_459
timestamp 1677583704
transform 1 0 44640 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_461
timestamp 1677583258
transform 1 0 44832 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_470
timestamp 1679585382
transform 1 0 45696 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_481
timestamp 1679581501
transform 1 0 46752 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_39_485
timestamp 1677583258
transform 1 0 47136 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_490
timestamp 1679585382
transform 1 0 47616 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_497
timestamp 1677583704
transform 1 0 48288 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_508
timestamp 1679585382
transform 1 0 49344 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_515
timestamp 1679585382
transform 1 0 50016 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_522
timestamp 1679585382
transform 1 0 50688 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_529
timestamp 1679585382
transform 1 0 51360 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_536
timestamp 1679585382
transform 1 0 52032 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_543
timestamp 1679585382
transform 1 0 52704 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_550
timestamp 1679585382
transform 1 0 53376 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_557
timestamp 1679585382
transform 1 0 54048 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_564
timestamp 1679585382
transform 1 0 54720 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_571
timestamp 1679585382
transform 1 0 55392 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_578
timestamp 1679585382
transform 1 0 56064 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_585
timestamp 1679585382
transform 1 0 56736 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_592
timestamp 1679585382
transform 1 0 57408 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_599
timestamp 1679585382
transform 1 0 58080 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_606
timestamp 1679585382
transform 1 0 58752 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_613
timestamp 1679585382
transform 1 0 59424 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_620
timestamp 1679585382
transform 1 0 60096 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_627
timestamp 1679585382
transform 1 0 60768 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_634
timestamp 1679585382
transform 1 0 61440 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_641
timestamp 1679585382
transform 1 0 62112 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_648
timestamp 1679585382
transform 1 0 62784 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_655
timestamp 1679585382
transform 1 0 63456 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_662
timestamp 1679585382
transform 1 0 64128 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_669
timestamp 1679585382
transform 1 0 64800 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_676
timestamp 1679585382
transform 1 0 65472 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_683
timestamp 1679585382
transform 1 0 66144 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_690
timestamp 1679585382
transform 1 0 66816 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_697
timestamp 1679585382
transform 1 0 67488 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_704
timestamp 1679585382
transform 1 0 68160 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_711
timestamp 1679585382
transform 1 0 68832 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_718
timestamp 1679585382
transform 1 0 69504 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_725
timestamp 1679585382
transform 1 0 70176 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_732
timestamp 1679585382
transform 1 0 70848 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_739
timestamp 1679585382
transform 1 0 71520 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_746
timestamp 1679585382
transform 1 0 72192 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_753
timestamp 1679585382
transform 1 0 72864 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_760
timestamp 1679585382
transform 1 0 73536 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_767
timestamp 1679585382
transform 1 0 74208 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_774
timestamp 1679585382
transform 1 0 74880 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_781
timestamp 1679585382
transform 1 0 75552 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_788
timestamp 1679585382
transform 1 0 76224 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_795
timestamp 1679585382
transform 1 0 76896 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_802
timestamp 1679585382
transform 1 0 77568 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_809
timestamp 1679585382
transform 1 0 78240 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_816
timestamp 1679585382
transform 1 0 78912 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_823
timestamp 1679585382
transform 1 0 79584 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_830
timestamp 1679585382
transform 1 0 80256 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_837
timestamp 1679585382
transform 1 0 80928 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_844
timestamp 1679585382
transform 1 0 81600 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_851
timestamp 1679585382
transform 1 0 82272 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_858
timestamp 1679585382
transform 1 0 82944 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_865
timestamp 1679585382
transform 1 0 83616 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_872
timestamp 1679585382
transform 1 0 84288 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_879
timestamp 1679585382
transform 1 0 84960 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_886
timestamp 1679585382
transform 1 0 85632 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_893
timestamp 1679585382
transform 1 0 86304 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_900
timestamp 1679585382
transform 1 0 86976 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_907
timestamp 1679585382
transform 1 0 87648 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_914
timestamp 1679585382
transform 1 0 88320 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_921
timestamp 1679585382
transform 1 0 88992 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_928
timestamp 1679585382
transform 1 0 89664 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_935
timestamp 1679585382
transform 1 0 90336 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_942
timestamp 1679585382
transform 1 0 91008 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_949
timestamp 1679585382
transform 1 0 91680 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_956
timestamp 1679585382
transform 1 0 92352 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_963
timestamp 1679585382
transform 1 0 93024 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_970
timestamp 1679585382
transform 1 0 93696 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_977
timestamp 1679585382
transform 1 0 94368 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_984
timestamp 1679585382
transform 1 0 95040 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_991
timestamp 1679585382
transform 1 0 95712 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_998
timestamp 1679585382
transform 1 0 96384 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1005
timestamp 1679585382
transform 1 0 97056 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1012
timestamp 1679585382
transform 1 0 97728 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_1019
timestamp 1679585382
transform 1 0 98400 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_1026
timestamp 1677583704
transform 1 0 99072 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_1028
timestamp 1677583258
transform 1 0 99264 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_0
timestamp 1679585382
transform 1 0 576 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_7
timestamp 1679585382
transform 1 0 1248 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_14
timestamp 1679585382
transform 1 0 1920 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_21
timestamp 1679585382
transform 1 0 2592 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_28
timestamp 1679581501
transform 1 0 3264 0 1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_40_32
timestamp 1677583258
transform 1 0 3648 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_46
timestamp 1679585382
transform 1 0 4992 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_53
timestamp 1679585382
transform 1 0 5664 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_60
timestamp 1679585382
transform 1 0 6336 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_67
timestamp 1679585382
transform 1 0 7008 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_74
timestamp 1679585382
transform 1 0 7680 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_81
timestamp 1679585382
transform 1 0 8352 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_88
timestamp 1679585382
transform 1 0 9024 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_95
timestamp 1679585382
transform 1 0 9696 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_102
timestamp 1679585382
transform 1 0 10368 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_118
timestamp 1679585382
transform 1 0 11904 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_125
timestamp 1679585382
transform 1 0 12576 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_132
timestamp 1679585382
transform 1 0 13248 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_139
timestamp 1679585382
transform 1 0 13920 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_146
timestamp 1679585382
transform 1 0 14592 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_153
timestamp 1679585382
transform 1 0 15264 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_160
timestamp 1679585382
transform 1 0 15936 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_167
timestamp 1679585382
transform 1 0 16608 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_174
timestamp 1679585382
transform 1 0 17280 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_181
timestamp 1679585382
transform 1 0 17952 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_188
timestamp 1679585382
transform 1 0 18624 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_195
timestamp 1679585382
transform 1 0 19296 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_202
timestamp 1679585382
transform 1 0 19968 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_209
timestamp 1679585382
transform 1 0 20640 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_216
timestamp 1677583704
transform 1 0 21312 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_218
timestamp 1677583258
transform 1 0 21504 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_232
timestamp 1679585382
transform 1 0 22848 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_239
timestamp 1677583704
transform 1 0 23520 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_241
timestamp 1677583258
transform 1 0 23712 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_250
timestamp 1679585382
transform 1 0 24576 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_257
timestamp 1679585382
transform 1 0 25248 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_264
timestamp 1679585382
transform 1 0 25920 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_271
timestamp 1677583704
transform 1 0 26592 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_273
timestamp 1677583258
transform 1 0 26784 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_283
timestamp 1679585382
transform 1 0 27744 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_290
timestamp 1679585382
transform 1 0 28416 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_297
timestamp 1679585382
transform 1 0 29088 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_304
timestamp 1679585382
transform 1 0 29760 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_320
timestamp 1679585382
transform 1 0 31296 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_327
timestamp 1679585382
transform 1 0 31968 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_334
timestamp 1679581501
transform 1 0 32640 0 1 30996
box -48 -56 432 834
use sg13g2_decap_8  FILLER_40_351
timestamp 1679585382
transform 1 0 34272 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_358
timestamp 1679581501
transform 1 0 34944 0 1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_40_362
timestamp 1677583258
transform 1 0 35328 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_402
timestamp 1679585382
transform 1 0 39168 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_409
timestamp 1679585382
transform 1 0 39840 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_416
timestamp 1679585382
transform 1 0 40512 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_423
timestamp 1679585382
transform 1 0 41184 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_430
timestamp 1679585382
transform 1 0 41856 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_437
timestamp 1679585382
transform 1 0 42528 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_444
timestamp 1679585382
transform 1 0 43200 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_451
timestamp 1679581501
transform 1 0 43872 0 1 30996
box -48 -56 432 834
use sg13g2_decap_8  FILLER_40_460
timestamp 1679585382
transform 1 0 44736 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_467
timestamp 1679585382
transform 1 0 45408 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_474
timestamp 1679585382
transform 1 0 46080 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_481
timestamp 1679585382
transform 1 0 46752 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_488
timestamp 1679585382
transform 1 0 47424 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_495
timestamp 1679585382
transform 1 0 48096 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_502
timestamp 1679585382
transform 1 0 48768 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_509
timestamp 1679585382
transform 1 0 49440 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_516
timestamp 1679585382
transform 1 0 50112 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_523
timestamp 1679585382
transform 1 0 50784 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_530
timestamp 1679585382
transform 1 0 51456 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_537
timestamp 1679585382
transform 1 0 52128 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_544
timestamp 1679585382
transform 1 0 52800 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_551
timestamp 1679585382
transform 1 0 53472 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_558
timestamp 1679585382
transform 1 0 54144 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_565
timestamp 1679585382
transform 1 0 54816 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_572
timestamp 1679585382
transform 1 0 55488 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_579
timestamp 1679585382
transform 1 0 56160 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_586
timestamp 1679585382
transform 1 0 56832 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_593
timestamp 1679585382
transform 1 0 57504 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_600
timestamp 1679585382
transform 1 0 58176 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_607
timestamp 1679585382
transform 1 0 58848 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_614
timestamp 1679585382
transform 1 0 59520 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_621
timestamp 1679585382
transform 1 0 60192 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_628
timestamp 1679585382
transform 1 0 60864 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_635
timestamp 1679585382
transform 1 0 61536 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_642
timestamp 1679585382
transform 1 0 62208 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_649
timestamp 1679585382
transform 1 0 62880 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_656
timestamp 1679585382
transform 1 0 63552 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_663
timestamp 1679585382
transform 1 0 64224 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_670
timestamp 1679585382
transform 1 0 64896 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_677
timestamp 1679585382
transform 1 0 65568 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_684
timestamp 1679585382
transform 1 0 66240 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_691
timestamp 1679585382
transform 1 0 66912 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_698
timestamp 1679585382
transform 1 0 67584 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_705
timestamp 1679585382
transform 1 0 68256 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_712
timestamp 1679585382
transform 1 0 68928 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_719
timestamp 1679585382
transform 1 0 69600 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_726
timestamp 1679585382
transform 1 0 70272 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_733
timestamp 1679585382
transform 1 0 70944 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_740
timestamp 1679585382
transform 1 0 71616 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_747
timestamp 1679585382
transform 1 0 72288 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_754
timestamp 1679585382
transform 1 0 72960 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_761
timestamp 1679585382
transform 1 0 73632 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_768
timestamp 1679585382
transform 1 0 74304 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_775
timestamp 1679585382
transform 1 0 74976 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_782
timestamp 1679585382
transform 1 0 75648 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_789
timestamp 1679585382
transform 1 0 76320 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_796
timestamp 1679585382
transform 1 0 76992 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_803
timestamp 1679585382
transform 1 0 77664 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_810
timestamp 1679585382
transform 1 0 78336 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_817
timestamp 1679585382
transform 1 0 79008 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_824
timestamp 1679585382
transform 1 0 79680 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_831
timestamp 1679585382
transform 1 0 80352 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_838
timestamp 1679585382
transform 1 0 81024 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_845
timestamp 1679585382
transform 1 0 81696 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_852
timestamp 1679585382
transform 1 0 82368 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_859
timestamp 1679585382
transform 1 0 83040 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_866
timestamp 1679585382
transform 1 0 83712 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_873
timestamp 1679585382
transform 1 0 84384 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_880
timestamp 1679585382
transform 1 0 85056 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_887
timestamp 1679585382
transform 1 0 85728 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_894
timestamp 1679585382
transform 1 0 86400 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_901
timestamp 1679585382
transform 1 0 87072 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_908
timestamp 1679585382
transform 1 0 87744 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_915
timestamp 1679585382
transform 1 0 88416 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_922
timestamp 1679585382
transform 1 0 89088 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_929
timestamp 1679585382
transform 1 0 89760 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_936
timestamp 1679585382
transform 1 0 90432 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_943
timestamp 1679585382
transform 1 0 91104 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_950
timestamp 1679585382
transform 1 0 91776 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_957
timestamp 1679585382
transform 1 0 92448 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_964
timestamp 1679585382
transform 1 0 93120 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_971
timestamp 1679585382
transform 1 0 93792 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_978
timestamp 1679585382
transform 1 0 94464 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_985
timestamp 1679585382
transform 1 0 95136 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_992
timestamp 1679585382
transform 1 0 95808 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_999
timestamp 1679585382
transform 1 0 96480 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1006
timestamp 1679585382
transform 1 0 97152 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1013
timestamp 1679585382
transform 1 0 97824 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_1020
timestamp 1679585382
transform 1 0 98496 0 1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_40_1027
timestamp 1677583704
transform 1 0 99168 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_41_0
timestamp 1679585382
transform 1 0 576 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_7
timestamp 1679585382
transform 1 0 1248 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_14
timestamp 1679585382
transform 1 0 1920 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_21
timestamp 1679585382
transform 1 0 2592 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_28
timestamp 1679585382
transform 1 0 3264 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_35
timestamp 1679585382
transform 1 0 3936 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_42
timestamp 1679585382
transform 1 0 4608 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_49
timestamp 1679585382
transform 1 0 5280 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_56
timestamp 1679585382
transform 1 0 5952 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_63
timestamp 1679585382
transform 1 0 6624 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_70
timestamp 1679585382
transform 1 0 7296 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_77
timestamp 1679585382
transform 1 0 7968 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_41_84
timestamp 1677583258
transform 1 0 8640 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_112
timestamp 1679585382
transform 1 0 11328 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_119
timestamp 1679585382
transform 1 0 12000 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_126
timestamp 1679585382
transform 1 0 12672 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_133
timestamp 1679585382
transform 1 0 13344 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_140
timestamp 1679585382
transform 1 0 14016 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_147
timestamp 1679585382
transform 1 0 14688 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_154
timestamp 1679585382
transform 1 0 15360 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_161
timestamp 1679585382
transform 1 0 16032 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_41_168
timestamp 1677583704
transform 1 0 16704 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_41_174
timestamp 1679585382
transform 1 0 17280 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_181
timestamp 1679585382
transform 1 0 17952 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_188
timestamp 1679585382
transform 1 0 18624 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_195
timestamp 1679585382
transform 1 0 19296 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_202
timestamp 1679585382
transform 1 0 19968 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_209
timestamp 1679585382
transform 1 0 20640 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_216
timestamp 1679585382
transform 1 0 21312 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_223
timestamp 1679585382
transform 1 0 21984 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_230
timestamp 1679585382
transform 1 0 22656 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_237
timestamp 1679585382
transform 1 0 23328 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_244
timestamp 1679585382
transform 1 0 24000 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_251
timestamp 1679585382
transform 1 0 24672 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_258
timestamp 1679585382
transform 1 0 25344 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_265
timestamp 1679585382
transform 1 0 26016 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_272
timestamp 1679585382
transform 1 0 26688 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_279
timestamp 1679585382
transform 1 0 27360 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_286
timestamp 1679585382
transform 1 0 28032 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_293
timestamp 1679585382
transform 1 0 28704 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_300
timestamp 1679585382
transform 1 0 29376 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_307
timestamp 1679585382
transform 1 0 30048 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_314
timestamp 1679585382
transform 1 0 30720 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_321
timestamp 1679585382
transform 1 0 31392 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_328
timestamp 1679585382
transform 1 0 32064 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_335
timestamp 1679585382
transform 1 0 32736 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_342
timestamp 1679581501
transform 1 0 33408 0 -1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_41_373
timestamp 1679585382
transform 1 0 36384 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_41_380
timestamp 1677583258
transform 1 0 37056 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_393
timestamp 1679585382
transform 1 0 38304 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_400
timestamp 1679585382
transform 1 0 38976 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_41_407
timestamp 1677583258
transform 1 0 39648 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_416
timestamp 1679585382
transform 1 0 40512 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_423
timestamp 1679585382
transform 1 0 41184 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_430
timestamp 1679581501
transform 1 0 41856 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_41_434
timestamp 1677583704
transform 1 0 42240 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_4  FILLER_41_463
timestamp 1679581501
transform 1 0 45024 0 -1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_41_471
timestamp 1679585382
transform 1 0 45792 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_478
timestamp 1679585382
transform 1 0 46464 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_485
timestamp 1679585382
transform 1 0 47136 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_492
timestamp 1679585382
transform 1 0 47808 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_499
timestamp 1679585382
transform 1 0 48480 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_506
timestamp 1679585382
transform 1 0 49152 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_513
timestamp 1679585382
transform 1 0 49824 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_520
timestamp 1679585382
transform 1 0 50496 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_527
timestamp 1679585382
transform 1 0 51168 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_534
timestamp 1679585382
transform 1 0 51840 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_541
timestamp 1679585382
transform 1 0 52512 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_548
timestamp 1679585382
transform 1 0 53184 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_555
timestamp 1679585382
transform 1 0 53856 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_562
timestamp 1679585382
transform 1 0 54528 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_569
timestamp 1679585382
transform 1 0 55200 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_576
timestamp 1679585382
transform 1 0 55872 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_583
timestamp 1679585382
transform 1 0 56544 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_590
timestamp 1679585382
transform 1 0 57216 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_597
timestamp 1679585382
transform 1 0 57888 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_604
timestamp 1679585382
transform 1 0 58560 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_611
timestamp 1679585382
transform 1 0 59232 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_618
timestamp 1679585382
transform 1 0 59904 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_625
timestamp 1679585382
transform 1 0 60576 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_632
timestamp 1679585382
transform 1 0 61248 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_639
timestamp 1679585382
transform 1 0 61920 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_646
timestamp 1679585382
transform 1 0 62592 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_653
timestamp 1679585382
transform 1 0 63264 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_660
timestamp 1679585382
transform 1 0 63936 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_667
timestamp 1679585382
transform 1 0 64608 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_674
timestamp 1679585382
transform 1 0 65280 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_681
timestamp 1679585382
transform 1 0 65952 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_688
timestamp 1679585382
transform 1 0 66624 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_695
timestamp 1679585382
transform 1 0 67296 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_702
timestamp 1679585382
transform 1 0 67968 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_709
timestamp 1679585382
transform 1 0 68640 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_716
timestamp 1679585382
transform 1 0 69312 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_723
timestamp 1679585382
transform 1 0 69984 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_730
timestamp 1679585382
transform 1 0 70656 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_737
timestamp 1679585382
transform 1 0 71328 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_744
timestamp 1679585382
transform 1 0 72000 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_751
timestamp 1679585382
transform 1 0 72672 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_758
timestamp 1679585382
transform 1 0 73344 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_765
timestamp 1679585382
transform 1 0 74016 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_772
timestamp 1679585382
transform 1 0 74688 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_779
timestamp 1679585382
transform 1 0 75360 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_786
timestamp 1679585382
transform 1 0 76032 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_793
timestamp 1679585382
transform 1 0 76704 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_800
timestamp 1679585382
transform 1 0 77376 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_807
timestamp 1679585382
transform 1 0 78048 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_814
timestamp 1679585382
transform 1 0 78720 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_821
timestamp 1679585382
transform 1 0 79392 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_828
timestamp 1679585382
transform 1 0 80064 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_835
timestamp 1679585382
transform 1 0 80736 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_842
timestamp 1679585382
transform 1 0 81408 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_849
timestamp 1679585382
transform 1 0 82080 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_856
timestamp 1679585382
transform 1 0 82752 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_863
timestamp 1679585382
transform 1 0 83424 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_870
timestamp 1679585382
transform 1 0 84096 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_877
timestamp 1679585382
transform 1 0 84768 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_884
timestamp 1679585382
transform 1 0 85440 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_891
timestamp 1679585382
transform 1 0 86112 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_898
timestamp 1679585382
transform 1 0 86784 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_905
timestamp 1679585382
transform 1 0 87456 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_912
timestamp 1679585382
transform 1 0 88128 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_919
timestamp 1679585382
transform 1 0 88800 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_926
timestamp 1679585382
transform 1 0 89472 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_933
timestamp 1679585382
transform 1 0 90144 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_940
timestamp 1679585382
transform 1 0 90816 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_947
timestamp 1679585382
transform 1 0 91488 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_954
timestamp 1679585382
transform 1 0 92160 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_961
timestamp 1679585382
transform 1 0 92832 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_968
timestamp 1679585382
transform 1 0 93504 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_975
timestamp 1679585382
transform 1 0 94176 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_982
timestamp 1679585382
transform 1 0 94848 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_989
timestamp 1679585382
transform 1 0 95520 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_996
timestamp 1679585382
transform 1 0 96192 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1003
timestamp 1679585382
transform 1 0 96864 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1010
timestamp 1679585382
transform 1 0 97536 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_1017
timestamp 1679585382
transform 1 0 98208 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_1024
timestamp 1679581501
transform 1 0 98880 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_41_1028
timestamp 1677583258
transform 1 0 99264 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_0
timestamp 1679585382
transform 1 0 576 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_7
timestamp 1679585382
transform 1 0 1248 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_14
timestamp 1679585382
transform 1 0 1920 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_21
timestamp 1679585382
transform 1 0 2592 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_28
timestamp 1679585382
transform 1 0 3264 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_35
timestamp 1679585382
transform 1 0 3936 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_42
timestamp 1679585382
transform 1 0 4608 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_49
timestamp 1679585382
transform 1 0 5280 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_56
timestamp 1679581501
transform 1 0 5952 0 1 32508
box -48 -56 432 834
use sg13g2_fill_1  FILLER_42_60
timestamp 1677583258
transform 1 0 6336 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_74
timestamp 1679585382
transform 1 0 7680 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_81
timestamp 1679581501
transform 1 0 8352 0 1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_42_112
timestamp 1679585382
transform 1 0 11328 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_119
timestamp 1679585382
transform 1 0 12000 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_126
timestamp 1679585382
transform 1 0 12672 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_133
timestamp 1679585382
transform 1 0 13344 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_140
timestamp 1679585382
transform 1 0 14016 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_147
timestamp 1679585382
transform 1 0 14688 0 1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_42_158
timestamp 1677583258
transform 1 0 15744 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_163
timestamp 1679585382
transform 1 0 16224 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_170
timestamp 1679585382
transform 1 0 16896 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_177
timestamp 1679585382
transform 1 0 17568 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_184
timestamp 1679585382
transform 1 0 18240 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_191
timestamp 1679585382
transform 1 0 18912 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_198
timestamp 1679585382
transform 1 0 19584 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_205
timestamp 1679585382
transform 1 0 20256 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_212
timestamp 1679585382
transform 1 0 20928 0 1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_42_219
timestamp 1677583258
transform 1 0 21600 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_247
timestamp 1679585382
transform 1 0 24288 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_254
timestamp 1679581501
transform 1 0 24960 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_258
timestamp 1677583704
transform 1 0 25344 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_287
timestamp 1679585382
transform 1 0 28128 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_294
timestamp 1679585382
transform 1 0 28800 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_301
timestamp 1679585382
transform 1 0 29472 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_308
timestamp 1679585382
transform 1 0 30144 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_315
timestamp 1679585382
transform 1 0 30816 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_322
timestamp 1679585382
transform 1 0 31488 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_329
timestamp 1679585382
transform 1 0 32160 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_336
timestamp 1679585382
transform 1 0 32832 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_343
timestamp 1679585382
transform 1 0 33504 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_350
timestamp 1679585382
transform 1 0 34176 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_357
timestamp 1679585382
transform 1 0 34848 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_364
timestamp 1679585382
transform 1 0 35520 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_371
timestamp 1679585382
transform 1 0 36192 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_387
timestamp 1679585382
transform 1 0 37728 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_394
timestamp 1679585382
transform 1 0 38400 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_401
timestamp 1679585382
transform 1 0 39072 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_408
timestamp 1679585382
transform 1 0 39744 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_415
timestamp 1679585382
transform 1 0 40416 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_422
timestamp 1679585382
transform 1 0 41088 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_429
timestamp 1679585382
transform 1 0 41760 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_436
timestamp 1679585382
transform 1 0 42432 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_443
timestamp 1677583704
transform 1 0 43104 0 1 32508
box -48 -56 240 834
use sg13g2_decap_4  FILLER_42_449
timestamp 1679581501
transform 1 0 43680 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_453
timestamp 1677583704
transform 1 0 44064 0 1 32508
box -48 -56 240 834
use sg13g2_fill_2  FILLER_42_464
timestamp 1677583704
transform 1 0 45120 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_493
timestamp 1679585382
transform 1 0 47904 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_500
timestamp 1679585382
transform 1 0 48576 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_507
timestamp 1679585382
transform 1 0 49248 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_514
timestamp 1679585382
transform 1 0 49920 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_521
timestamp 1679585382
transform 1 0 50592 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_528
timestamp 1679585382
transform 1 0 51264 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_535
timestamp 1679585382
transform 1 0 51936 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_542
timestamp 1679585382
transform 1 0 52608 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_549
timestamp 1679585382
transform 1 0 53280 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_556
timestamp 1679585382
transform 1 0 53952 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_563
timestamp 1679585382
transform 1 0 54624 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_570
timestamp 1679585382
transform 1 0 55296 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_577
timestamp 1679585382
transform 1 0 55968 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_584
timestamp 1679585382
transform 1 0 56640 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_591
timestamp 1679585382
transform 1 0 57312 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_598
timestamp 1679585382
transform 1 0 57984 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_605
timestamp 1679585382
transform 1 0 58656 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_612
timestamp 1679585382
transform 1 0 59328 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_619
timestamp 1679585382
transform 1 0 60000 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_626
timestamp 1679585382
transform 1 0 60672 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_633
timestamp 1679585382
transform 1 0 61344 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_640
timestamp 1679585382
transform 1 0 62016 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_647
timestamp 1679585382
transform 1 0 62688 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_654
timestamp 1679585382
transform 1 0 63360 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_661
timestamp 1679585382
transform 1 0 64032 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_668
timestamp 1679585382
transform 1 0 64704 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_675
timestamp 1679585382
transform 1 0 65376 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_682
timestamp 1679585382
transform 1 0 66048 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_689
timestamp 1679585382
transform 1 0 66720 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_696
timestamp 1679585382
transform 1 0 67392 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_703
timestamp 1679585382
transform 1 0 68064 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_710
timestamp 1679585382
transform 1 0 68736 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_717
timestamp 1679585382
transform 1 0 69408 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_724
timestamp 1679585382
transform 1 0 70080 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_731
timestamp 1679585382
transform 1 0 70752 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_738
timestamp 1679585382
transform 1 0 71424 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_745
timestamp 1679585382
transform 1 0 72096 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_752
timestamp 1679585382
transform 1 0 72768 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_759
timestamp 1679585382
transform 1 0 73440 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_766
timestamp 1679585382
transform 1 0 74112 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_773
timestamp 1679585382
transform 1 0 74784 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_780
timestamp 1679585382
transform 1 0 75456 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_787
timestamp 1679585382
transform 1 0 76128 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_794
timestamp 1679585382
transform 1 0 76800 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_801
timestamp 1679585382
transform 1 0 77472 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_808
timestamp 1679585382
transform 1 0 78144 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_815
timestamp 1679585382
transform 1 0 78816 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_822
timestamp 1679585382
transform 1 0 79488 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_829
timestamp 1679585382
transform 1 0 80160 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_836
timestamp 1679585382
transform 1 0 80832 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_843
timestamp 1679585382
transform 1 0 81504 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_850
timestamp 1679585382
transform 1 0 82176 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_857
timestamp 1679585382
transform 1 0 82848 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_864
timestamp 1679585382
transform 1 0 83520 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_871
timestamp 1679585382
transform 1 0 84192 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_878
timestamp 1679585382
transform 1 0 84864 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_885
timestamp 1679585382
transform 1 0 85536 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_892
timestamp 1679585382
transform 1 0 86208 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_899
timestamp 1679585382
transform 1 0 86880 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_906
timestamp 1679585382
transform 1 0 87552 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_913
timestamp 1679585382
transform 1 0 88224 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_920
timestamp 1679585382
transform 1 0 88896 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_927
timestamp 1679585382
transform 1 0 89568 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_934
timestamp 1679585382
transform 1 0 90240 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_941
timestamp 1679585382
transform 1 0 90912 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_948
timestamp 1679585382
transform 1 0 91584 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_955
timestamp 1679585382
transform 1 0 92256 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_962
timestamp 1679585382
transform 1 0 92928 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_969
timestamp 1679585382
transform 1 0 93600 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_976
timestamp 1679585382
transform 1 0 94272 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_983
timestamp 1679585382
transform 1 0 94944 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_990
timestamp 1679585382
transform 1 0 95616 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_997
timestamp 1679585382
transform 1 0 96288 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1004
timestamp 1679585382
transform 1 0 96960 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1011
timestamp 1679585382
transform 1 0 97632 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_1018
timestamp 1679585382
transform 1 0 98304 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_1025
timestamp 1679581501
transform 1 0 98976 0 1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_43_0
timestamp 1679585382
transform 1 0 576 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_7
timestamp 1679585382
transform 1 0 1248 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_14
timestamp 1679585382
transform 1 0 1920 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_21
timestamp 1679585382
transform 1 0 2592 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_28
timestamp 1679585382
transform 1 0 3264 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_35
timestamp 1679585382
transform 1 0 3936 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_42
timestamp 1679585382
transform 1 0 4608 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_49
timestamp 1679585382
transform 1 0 5280 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_56
timestamp 1679585382
transform 1 0 5952 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_63
timestamp 1679585382
transform 1 0 6624 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_70
timestamp 1679585382
transform 1 0 7296 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_77
timestamp 1679585382
transform 1 0 7968 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_84
timestamp 1679585382
transform 1 0 8640 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_91
timestamp 1679585382
transform 1 0 9312 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_98
timestamp 1679585382
transform 1 0 9984 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_121
timestamp 1679585382
transform 1 0 12192 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_128
timestamp 1679585382
transform 1 0 12864 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_135
timestamp 1679585382
transform 1 0 13536 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_142
timestamp 1679585382
transform 1 0 14208 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_185
timestamp 1679585382
transform 1 0 18336 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_192
timestamp 1679585382
transform 1 0 19008 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_199
timestamp 1679585382
transform 1 0 19680 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_206
timestamp 1679585382
transform 1 0 20352 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_213
timestamp 1679585382
transform 1 0 21024 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_220
timestamp 1679585382
transform 1 0 21696 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_227
timestamp 1679585382
transform 1 0 22368 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_234
timestamp 1679585382
transform 1 0 23040 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_43_241
timestamp 1679581501
transform 1 0 23712 0 -1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_43_261
timestamp 1679585382
transform 1 0 25632 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_268
timestamp 1679585382
transform 1 0 26304 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_275
timestamp 1679585382
transform 1 0 26976 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_282
timestamp 1679585382
transform 1 0 27648 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_289
timestamp 1679585382
transform 1 0 28320 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_296
timestamp 1679585382
transform 1 0 28992 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_303
timestamp 1679585382
transform 1 0 29664 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_310
timestamp 1679585382
transform 1 0 30336 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_317
timestamp 1679585382
transform 1 0 31008 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_324
timestamp 1679585382
transform 1 0 31680 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_331
timestamp 1679585382
transform 1 0 32352 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_338
timestamp 1679585382
transform 1 0 33024 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_345
timestamp 1679585382
transform 1 0 33696 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_352
timestamp 1679585382
transform 1 0 34368 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_359
timestamp 1679585382
transform 1 0 35040 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_366
timestamp 1679585382
transform 1 0 35712 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_373
timestamp 1679585382
transform 1 0 36384 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_380
timestamp 1679585382
transform 1 0 37056 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_387
timestamp 1679585382
transform 1 0 37728 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_394
timestamp 1679585382
transform 1 0 38400 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_401
timestamp 1679585382
transform 1 0 39072 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_408
timestamp 1679585382
transform 1 0 39744 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_415
timestamp 1679585382
transform 1 0 40416 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_422
timestamp 1679585382
transform 1 0 41088 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_429
timestamp 1679585382
transform 1 0 41760 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_436
timestamp 1679585382
transform 1 0 42432 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_443
timestamp 1679585382
transform 1 0 43104 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_450
timestamp 1679585382
transform 1 0 43776 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_457
timestamp 1679585382
transform 1 0 44448 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_464
timestamp 1679585382
transform 1 0 45120 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_471
timestamp 1679585382
transform 1 0 45792 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_43_478
timestamp 1677583704
transform 1 0 46464 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_480
timestamp 1677583258
transform 1 0 46656 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_490
timestamp 1679585382
transform 1 0 47616 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_497
timestamp 1679585382
transform 1 0 48288 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_504
timestamp 1679585382
transform 1 0 48960 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_511
timestamp 1679585382
transform 1 0 49632 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_518
timestamp 1679585382
transform 1 0 50304 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_525
timestamp 1679585382
transform 1 0 50976 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_532
timestamp 1679585382
transform 1 0 51648 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_539
timestamp 1679585382
transform 1 0 52320 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_546
timestamp 1679585382
transform 1 0 52992 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_553
timestamp 1679585382
transform 1 0 53664 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_560
timestamp 1679585382
transform 1 0 54336 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_567
timestamp 1679585382
transform 1 0 55008 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_574
timestamp 1679585382
transform 1 0 55680 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_581
timestamp 1679585382
transform 1 0 56352 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_588
timestamp 1679585382
transform 1 0 57024 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_595
timestamp 1679585382
transform 1 0 57696 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_602
timestamp 1679585382
transform 1 0 58368 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_609
timestamp 1679585382
transform 1 0 59040 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_616
timestamp 1679585382
transform 1 0 59712 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_623
timestamp 1679585382
transform 1 0 60384 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_630
timestamp 1679585382
transform 1 0 61056 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_637
timestamp 1679585382
transform 1 0 61728 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_644
timestamp 1679585382
transform 1 0 62400 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_651
timestamp 1679585382
transform 1 0 63072 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_658
timestamp 1679585382
transform 1 0 63744 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_665
timestamp 1679585382
transform 1 0 64416 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_672
timestamp 1679585382
transform 1 0 65088 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_679
timestamp 1679585382
transform 1 0 65760 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_686
timestamp 1679585382
transform 1 0 66432 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_693
timestamp 1679585382
transform 1 0 67104 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_700
timestamp 1679585382
transform 1 0 67776 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_707
timestamp 1679585382
transform 1 0 68448 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_714
timestamp 1679585382
transform 1 0 69120 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_721
timestamp 1679585382
transform 1 0 69792 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_728
timestamp 1679585382
transform 1 0 70464 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_735
timestamp 1679585382
transform 1 0 71136 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_742
timestamp 1679585382
transform 1 0 71808 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_749
timestamp 1679585382
transform 1 0 72480 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_756
timestamp 1679585382
transform 1 0 73152 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_763
timestamp 1679585382
transform 1 0 73824 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_770
timestamp 1679585382
transform 1 0 74496 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_777
timestamp 1679585382
transform 1 0 75168 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_784
timestamp 1679585382
transform 1 0 75840 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_791
timestamp 1679585382
transform 1 0 76512 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_798
timestamp 1679585382
transform 1 0 77184 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_805
timestamp 1679585382
transform 1 0 77856 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_812
timestamp 1679585382
transform 1 0 78528 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_819
timestamp 1679585382
transform 1 0 79200 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_826
timestamp 1679585382
transform 1 0 79872 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_833
timestamp 1679585382
transform 1 0 80544 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_840
timestamp 1679585382
transform 1 0 81216 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_847
timestamp 1679585382
transform 1 0 81888 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_854
timestamp 1679585382
transform 1 0 82560 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_861
timestamp 1679585382
transform 1 0 83232 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_868
timestamp 1679585382
transform 1 0 83904 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_875
timestamp 1679585382
transform 1 0 84576 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_882
timestamp 1679585382
transform 1 0 85248 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_889
timestamp 1679585382
transform 1 0 85920 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_896
timestamp 1679585382
transform 1 0 86592 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_903
timestamp 1679585382
transform 1 0 87264 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_910
timestamp 1679585382
transform 1 0 87936 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_917
timestamp 1679585382
transform 1 0 88608 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_924
timestamp 1679585382
transform 1 0 89280 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_931
timestamp 1679585382
transform 1 0 89952 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_938
timestamp 1679585382
transform 1 0 90624 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_945
timestamp 1679585382
transform 1 0 91296 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_952
timestamp 1679585382
transform 1 0 91968 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_959
timestamp 1679585382
transform 1 0 92640 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_966
timestamp 1679585382
transform 1 0 93312 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_973
timestamp 1679585382
transform 1 0 93984 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_980
timestamp 1679585382
transform 1 0 94656 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_987
timestamp 1679585382
transform 1 0 95328 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_994
timestamp 1679585382
transform 1 0 96000 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1001
timestamp 1679585382
transform 1 0 96672 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1008
timestamp 1679585382
transform 1 0 97344 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1015
timestamp 1679585382
transform 1 0 98016 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_1022
timestamp 1679585382
transform 1 0 98688 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_0
timestamp 1679585382
transform 1 0 576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_7
timestamp 1679585382
transform 1 0 1248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_14
timestamp 1679585382
transform 1 0 1920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_21
timestamp 1679585382
transform 1 0 2592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_28
timestamp 1679581501
transform 1 0 3264 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_44_32
timestamp 1677583704
transform 1 0 3648 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_61
timestamp 1679585382
transform 1 0 6432 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_68
timestamp 1679585382
transform 1 0 7104 0 1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_44_75
timestamp 1677583258
transform 1 0 7776 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_89
timestamp 1679585382
transform 1 0 9120 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_96
timestamp 1679585382
transform 1 0 9792 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_103
timestamp 1679585382
transform 1 0 10464 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_110
timestamp 1679585382
transform 1 0 11136 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_117
timestamp 1679585382
transform 1 0 11808 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_124
timestamp 1679585382
transform 1 0 12480 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_131
timestamp 1679585382
transform 1 0 13152 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_138
timestamp 1679581501
transform 1 0 13824 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_44_142
timestamp 1677583704
transform 1 0 14208 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_180
timestamp 1679585382
transform 1 0 17856 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_187
timestamp 1679585382
transform 1 0 18528 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_194
timestamp 1679581501
transform 1 0 19200 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_44_198
timestamp 1677583704
transform 1 0 19584 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_213
timestamp 1679585382
transform 1 0 21024 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_220
timestamp 1679585382
transform 1 0 21696 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_227
timestamp 1679585382
transform 1 0 22368 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_234
timestamp 1679585382
transform 1 0 23040 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_241
timestamp 1679585382
transform 1 0 23712 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_248
timestamp 1679585382
transform 1 0 24384 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_255
timestamp 1679585382
transform 1 0 25056 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_262
timestamp 1679585382
transform 1 0 25728 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_269
timestamp 1679585382
transform 1 0 26400 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_276
timestamp 1679585382
transform 1 0 27072 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_283
timestamp 1679585382
transform 1 0 27744 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_290
timestamp 1679585382
transform 1 0 28416 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_297
timestamp 1679585382
transform 1 0 29088 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_304
timestamp 1679581501
transform 1 0 29760 0 1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_44_308
timestamp 1677583258
transform 1 0 30144 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_336
timestamp 1679585382
transform 1 0 32832 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_343
timestamp 1677583704
transform 1 0 33504 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_350
timestamp 1679585382
transform 1 0 34176 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_357
timestamp 1679585382
transform 1 0 34848 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_364
timestamp 1679585382
transform 1 0 35520 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_371
timestamp 1679585382
transform 1 0 36192 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_378
timestamp 1679581501
transform 1 0 36864 0 1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_44_409
timestamp 1679585382
transform 1 0 39840 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_416
timestamp 1679585382
transform 1 0 40512 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_423
timestamp 1679585382
transform 1 0 41184 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_430
timestamp 1679585382
transform 1 0 41856 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_437
timestamp 1679585382
transform 1 0 42528 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_444
timestamp 1679585382
transform 1 0 43200 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_451
timestamp 1679585382
transform 1 0 43872 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_458
timestamp 1679585382
transform 1 0 44544 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_465
timestamp 1679585382
transform 1 0 45216 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_472
timestamp 1679585382
transform 1 0 45888 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_479
timestamp 1679585382
transform 1 0 46560 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_486
timestamp 1679585382
transform 1 0 47232 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_493
timestamp 1679585382
transform 1 0 47904 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_500
timestamp 1679585382
transform 1 0 48576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_507
timestamp 1679585382
transform 1 0 49248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_514
timestamp 1679585382
transform 1 0 49920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_521
timestamp 1679585382
transform 1 0 50592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_528
timestamp 1679585382
transform 1 0 51264 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_535
timestamp 1679585382
transform 1 0 51936 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_542
timestamp 1679585382
transform 1 0 52608 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_549
timestamp 1679585382
transform 1 0 53280 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_556
timestamp 1679585382
transform 1 0 53952 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_563
timestamp 1679585382
transform 1 0 54624 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_570
timestamp 1679585382
transform 1 0 55296 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_577
timestamp 1679585382
transform 1 0 55968 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_584
timestamp 1679585382
transform 1 0 56640 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_591
timestamp 1679585382
transform 1 0 57312 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_598
timestamp 1679585382
transform 1 0 57984 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_605
timestamp 1679585382
transform 1 0 58656 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_612
timestamp 1679585382
transform 1 0 59328 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_619
timestamp 1679585382
transform 1 0 60000 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_626
timestamp 1679585382
transform 1 0 60672 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_633
timestamp 1679585382
transform 1 0 61344 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_640
timestamp 1679585382
transform 1 0 62016 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_647
timestamp 1679585382
transform 1 0 62688 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_654
timestamp 1679585382
transform 1 0 63360 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_661
timestamp 1679585382
transform 1 0 64032 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_668
timestamp 1679585382
transform 1 0 64704 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_675
timestamp 1679585382
transform 1 0 65376 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_682
timestamp 1679585382
transform 1 0 66048 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_689
timestamp 1679585382
transform 1 0 66720 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_696
timestamp 1679585382
transform 1 0 67392 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_703
timestamp 1679585382
transform 1 0 68064 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_710
timestamp 1679585382
transform 1 0 68736 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_717
timestamp 1679585382
transform 1 0 69408 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_724
timestamp 1679585382
transform 1 0 70080 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_731
timestamp 1679585382
transform 1 0 70752 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_738
timestamp 1679585382
transform 1 0 71424 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_745
timestamp 1679585382
transform 1 0 72096 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_752
timestamp 1679585382
transform 1 0 72768 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_759
timestamp 1679585382
transform 1 0 73440 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_766
timestamp 1679585382
transform 1 0 74112 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_773
timestamp 1679585382
transform 1 0 74784 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_780
timestamp 1679585382
transform 1 0 75456 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_787
timestamp 1679585382
transform 1 0 76128 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_794
timestamp 1679585382
transform 1 0 76800 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_801
timestamp 1679585382
transform 1 0 77472 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_808
timestamp 1679585382
transform 1 0 78144 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_815
timestamp 1679585382
transform 1 0 78816 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_822
timestamp 1679585382
transform 1 0 79488 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_829
timestamp 1679585382
transform 1 0 80160 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_836
timestamp 1679585382
transform 1 0 80832 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_843
timestamp 1679585382
transform 1 0 81504 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_850
timestamp 1679585382
transform 1 0 82176 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_857
timestamp 1679585382
transform 1 0 82848 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_864
timestamp 1679585382
transform 1 0 83520 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_871
timestamp 1679585382
transform 1 0 84192 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_878
timestamp 1679585382
transform 1 0 84864 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_885
timestamp 1679585382
transform 1 0 85536 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_892
timestamp 1679585382
transform 1 0 86208 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_899
timestamp 1679585382
transform 1 0 86880 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_906
timestamp 1679585382
transform 1 0 87552 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_913
timestamp 1679585382
transform 1 0 88224 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_920
timestamp 1679585382
transform 1 0 88896 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_927
timestamp 1679585382
transform 1 0 89568 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_934
timestamp 1679585382
transform 1 0 90240 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_941
timestamp 1679585382
transform 1 0 90912 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_948
timestamp 1679585382
transform 1 0 91584 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_955
timestamp 1679585382
transform 1 0 92256 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_962
timestamp 1679585382
transform 1 0 92928 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_969
timestamp 1679585382
transform 1 0 93600 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_976
timestamp 1679585382
transform 1 0 94272 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_983
timestamp 1679585382
transform 1 0 94944 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_990
timestamp 1679585382
transform 1 0 95616 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_997
timestamp 1679585382
transform 1 0 96288 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1004
timestamp 1679585382
transform 1 0 96960 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1011
timestamp 1679585382
transform 1 0 97632 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1018
timestamp 1679585382
transform 1 0 98304 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_1025
timestamp 1679581501
transform 1 0 98976 0 1 34020
box -48 -56 432 834
use sg13g2_decap_8  FILLER_45_0
timestamp 1679585382
transform 1 0 576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_7
timestamp 1679585382
transform 1 0 1248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_14
timestamp 1679585382
transform 1 0 1920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_21
timestamp 1679585382
transform 1 0 2592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_28
timestamp 1679585382
transform 1 0 3264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_35
timestamp 1679585382
transform 1 0 3936 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_42
timestamp 1677583704
transform 1 0 4608 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_4  FILLER_45_48
timestamp 1679581501
transform 1 0 5184 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_45_52
timestamp 1677583704
transform 1 0 5568 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_4  FILLER_45_63
timestamp 1679581501
transform 1 0 6624 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_45_67
timestamp 1677583704
transform 1 0 7008 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_73
timestamp 1679585382
transform 1 0 7584 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_80
timestamp 1679585382
transform 1 0 8256 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_87
timestamp 1677583704
transform 1 0 8928 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_89
timestamp 1677583258
transform 1 0 9120 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_103
timestamp 1679585382
transform 1 0 10464 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_110
timestamp 1679585382
transform 1 0 11136 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_117
timestamp 1679585382
transform 1 0 11808 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_124
timestamp 1679585382
transform 1 0 12480 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_131
timestamp 1679585382
transform 1 0 13152 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_138
timestamp 1679585382
transform 1 0 13824 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_145
timestamp 1679585382
transform 1 0 14496 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_152
timestamp 1679585382
transform 1 0 15168 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_159
timestamp 1679585382
transform 1 0 15840 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_166
timestamp 1679585382
transform 1 0 16512 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_173
timestamp 1679585382
transform 1 0 17184 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_180
timestamp 1679585382
transform 1 0 17856 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_187
timestamp 1679585382
transform 1 0 18528 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_194
timestamp 1679585382
transform 1 0 19200 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_201
timestamp 1679585382
transform 1 0 19872 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_208
timestamp 1679585382
transform 1 0 20544 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_227
timestamp 1679585382
transform 1 0 22368 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_234
timestamp 1679585382
transform 1 0 23040 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_241
timestamp 1679585382
transform 1 0 23712 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_248
timestamp 1677583704
transform 1 0 24384 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_45_254
timestamp 1677583704
transform 1 0 24960 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_261
timestamp 1679585382
transform 1 0 25632 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_268
timestamp 1679585382
transform 1 0 26304 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_275
timestamp 1679585382
transform 1 0 26976 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_282
timestamp 1679585382
transform 1 0 27648 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_289
timestamp 1679585382
transform 1 0 28320 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_296
timestamp 1679585382
transform 1 0 28992 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_303
timestamp 1679585382
transform 1 0 29664 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_310
timestamp 1679585382
transform 1 0 30336 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_317
timestamp 1677583704
transform 1 0 31008 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_4  FILLER_45_323
timestamp 1679581501
transform 1 0 31584 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_45_327
timestamp 1677583704
transform 1 0 31968 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_342
timestamp 1679585382
transform 1 0 33408 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_349
timestamp 1679585382
transform 1 0 34080 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_356
timestamp 1679585382
transform 1 0 34752 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_363
timestamp 1677583704
transform 1 0 35424 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_365
timestamp 1677583258
transform 1 0 35616 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_374
timestamp 1679585382
transform 1 0 36480 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_381
timestamp 1679585382
transform 1 0 37152 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_388
timestamp 1679585382
transform 1 0 37824 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_395
timestamp 1679585382
transform 1 0 38496 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_402
timestamp 1679585382
transform 1 0 39168 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_409
timestamp 1679585382
transform 1 0 39840 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_416
timestamp 1679585382
transform 1 0 40512 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_423
timestamp 1679585382
transform 1 0 41184 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_430
timestamp 1679585382
transform 1 0 41856 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_437
timestamp 1679585382
transform 1 0 42528 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_444
timestamp 1679585382
transform 1 0 43200 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_451
timestamp 1679585382
transform 1 0 43872 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_458
timestamp 1679585382
transform 1 0 44544 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_465
timestamp 1679585382
transform 1 0 45216 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_472
timestamp 1679585382
transform 1 0 45888 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_479
timestamp 1679585382
transform 1 0 46560 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_486
timestamp 1679585382
transform 1 0 47232 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_493
timestamp 1679585382
transform 1 0 47904 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_500
timestamp 1679585382
transform 1 0 48576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_507
timestamp 1679585382
transform 1 0 49248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_514
timestamp 1679585382
transform 1 0 49920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_521
timestamp 1679585382
transform 1 0 50592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_528
timestamp 1679585382
transform 1 0 51264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_535
timestamp 1679585382
transform 1 0 51936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_542
timestamp 1679585382
transform 1 0 52608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_549
timestamp 1679585382
transform 1 0 53280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_556
timestamp 1679585382
transform 1 0 53952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_563
timestamp 1679585382
transform 1 0 54624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_570
timestamp 1679585382
transform 1 0 55296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_577
timestamp 1679585382
transform 1 0 55968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_584
timestamp 1679585382
transform 1 0 56640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_591
timestamp 1679585382
transform 1 0 57312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_598
timestamp 1679585382
transform 1 0 57984 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_605
timestamp 1679585382
transform 1 0 58656 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_612
timestamp 1679585382
transform 1 0 59328 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_619
timestamp 1679585382
transform 1 0 60000 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_626
timestamp 1679585382
transform 1 0 60672 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_633
timestamp 1679585382
transform 1 0 61344 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_640
timestamp 1679585382
transform 1 0 62016 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_647
timestamp 1679585382
transform 1 0 62688 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_654
timestamp 1679585382
transform 1 0 63360 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_661
timestamp 1679585382
transform 1 0 64032 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_668
timestamp 1679585382
transform 1 0 64704 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_675
timestamp 1679585382
transform 1 0 65376 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_682
timestamp 1679585382
transform 1 0 66048 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_689
timestamp 1679585382
transform 1 0 66720 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_696
timestamp 1679585382
transform 1 0 67392 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_703
timestamp 1679585382
transform 1 0 68064 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_710
timestamp 1679585382
transform 1 0 68736 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_717
timestamp 1679585382
transform 1 0 69408 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_724
timestamp 1679585382
transform 1 0 70080 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_731
timestamp 1679585382
transform 1 0 70752 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_738
timestamp 1679585382
transform 1 0 71424 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_745
timestamp 1679585382
transform 1 0 72096 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_752
timestamp 1679585382
transform 1 0 72768 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_759
timestamp 1679585382
transform 1 0 73440 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_766
timestamp 1679585382
transform 1 0 74112 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_773
timestamp 1679585382
transform 1 0 74784 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_780
timestamp 1679585382
transform 1 0 75456 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_787
timestamp 1679585382
transform 1 0 76128 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_794
timestamp 1679585382
transform 1 0 76800 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_801
timestamp 1679585382
transform 1 0 77472 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_808
timestamp 1679585382
transform 1 0 78144 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_815
timestamp 1679585382
transform 1 0 78816 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_822
timestamp 1679585382
transform 1 0 79488 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_829
timestamp 1679585382
transform 1 0 80160 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_836
timestamp 1679585382
transform 1 0 80832 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_843
timestamp 1679585382
transform 1 0 81504 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_850
timestamp 1679585382
transform 1 0 82176 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_857
timestamp 1679585382
transform 1 0 82848 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_864
timestamp 1679585382
transform 1 0 83520 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_871
timestamp 1679585382
transform 1 0 84192 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_878
timestamp 1679585382
transform 1 0 84864 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_885
timestamp 1679585382
transform 1 0 85536 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_892
timestamp 1679585382
transform 1 0 86208 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_899
timestamp 1679585382
transform 1 0 86880 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_906
timestamp 1679585382
transform 1 0 87552 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_913
timestamp 1679585382
transform 1 0 88224 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_920
timestamp 1679585382
transform 1 0 88896 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_927
timestamp 1679585382
transform 1 0 89568 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_934
timestamp 1679585382
transform 1 0 90240 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_941
timestamp 1679585382
transform 1 0 90912 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_948
timestamp 1679585382
transform 1 0 91584 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_955
timestamp 1679585382
transform 1 0 92256 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_962
timestamp 1679585382
transform 1 0 92928 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_969
timestamp 1679585382
transform 1 0 93600 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_976
timestamp 1679585382
transform 1 0 94272 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_983
timestamp 1679585382
transform 1 0 94944 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_990
timestamp 1679585382
transform 1 0 95616 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_997
timestamp 1679585382
transform 1 0 96288 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1004
timestamp 1679585382
transform 1 0 96960 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1011
timestamp 1679585382
transform 1 0 97632 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1018
timestamp 1679585382
transform 1 0 98304 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_1025
timestamp 1679581501
transform 1 0 98976 0 -1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_46_0
timestamp 1679585382
transform 1 0 576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_7
timestamp 1679585382
transform 1 0 1248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_14
timestamp 1679585382
transform 1 0 1920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_21
timestamp 1679585382
transform 1 0 2592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_28
timestamp 1679585382
transform 1 0 3264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_35
timestamp 1679585382
transform 1 0 3936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_69
timestamp 1679585382
transform 1 0 7200 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_76
timestamp 1679585382
transform 1 0 7872 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_83
timestamp 1679581501
transform 1 0 8544 0 1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_87
timestamp 1677583704
transform 1 0 8928 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_120
timestamp 1679585382
transform 1 0 12096 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_127
timestamp 1679585382
transform 1 0 12768 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_134
timestamp 1679585382
transform 1 0 13440 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_141
timestamp 1679585382
transform 1 0 14112 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_148
timestamp 1679585382
transform 1 0 14784 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_155
timestamp 1679585382
transform 1 0 15456 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_162
timestamp 1679585382
transform 1 0 16128 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_169
timestamp 1679585382
transform 1 0 16800 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_176
timestamp 1679585382
transform 1 0 17472 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_183
timestamp 1679585382
transform 1 0 18144 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_190
timestamp 1679581501
transform 1 0 18816 0 1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_198
timestamp 1677583704
transform 1 0 19584 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_204
timestamp 1679585382
transform 1 0 20160 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_211
timestamp 1679585382
transform 1 0 20832 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_218
timestamp 1679581501
transform 1 0 21504 0 1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_222
timestamp 1677583704
transform 1 0 21888 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_228
timestamp 1679585382
transform 1 0 22464 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_275
timestamp 1679585382
transform 1 0 26976 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_282
timestamp 1679585382
transform 1 0 27648 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_289
timestamp 1679585382
transform 1 0 28320 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_296
timestamp 1679585382
transform 1 0 28992 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_303
timestamp 1679581501
transform 1 0 29664 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_307
timestamp 1677583258
transform 1 0 30048 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_335
timestamp 1679585382
transform 1 0 32736 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_342
timestamp 1679585382
transform 1 0 33408 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_349
timestamp 1679585382
transform 1 0 34080 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_356
timestamp 1679581501
transform 1 0 34752 0 1 35532
box -48 -56 432 834
use sg13g2_decap_4  FILLER_46_364
timestamp 1679581501
transform 1 0 35520 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_368
timestamp 1677583258
transform 1 0 35904 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_386
timestamp 1679585382
transform 1 0 37632 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_393
timestamp 1679585382
transform 1 0 38304 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_400
timestamp 1679585382
transform 1 0 38976 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_407
timestamp 1679585382
transform 1 0 39648 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_414
timestamp 1679585382
transform 1 0 40320 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_421
timestamp 1679585382
transform 1 0 40992 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_428
timestamp 1679585382
transform 1 0 41664 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_435
timestamp 1679585382
transform 1 0 42336 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_442
timestamp 1679585382
transform 1 0 43008 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_449
timestamp 1679585382
transform 1 0 43680 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_456
timestamp 1679585382
transform 1 0 44352 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_463
timestamp 1679585382
transform 1 0 45024 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_470
timestamp 1679585382
transform 1 0 45696 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_477
timestamp 1679585382
transform 1 0 46368 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_484
timestamp 1679585382
transform 1 0 47040 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_491
timestamp 1679585382
transform 1 0 47712 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_498
timestamp 1679585382
transform 1 0 48384 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_505
timestamp 1679585382
transform 1 0 49056 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_512
timestamp 1679585382
transform 1 0 49728 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_519
timestamp 1679585382
transform 1 0 50400 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_526
timestamp 1679585382
transform 1 0 51072 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_533
timestamp 1679585382
transform 1 0 51744 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_540
timestamp 1679585382
transform 1 0 52416 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_547
timestamp 1679585382
transform 1 0 53088 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_554
timestamp 1679585382
transform 1 0 53760 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_561
timestamp 1679585382
transform 1 0 54432 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_568
timestamp 1679585382
transform 1 0 55104 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_575
timestamp 1679585382
transform 1 0 55776 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_582
timestamp 1679585382
transform 1 0 56448 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_589
timestamp 1679585382
transform 1 0 57120 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_596
timestamp 1679585382
transform 1 0 57792 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_603
timestamp 1679585382
transform 1 0 58464 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_610
timestamp 1679585382
transform 1 0 59136 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_617
timestamp 1679585382
transform 1 0 59808 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_624
timestamp 1679585382
transform 1 0 60480 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_631
timestamp 1679585382
transform 1 0 61152 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_638
timestamp 1679585382
transform 1 0 61824 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_645
timestamp 1679585382
transform 1 0 62496 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_652
timestamp 1679585382
transform 1 0 63168 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_659
timestamp 1679585382
transform 1 0 63840 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_666
timestamp 1679585382
transform 1 0 64512 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_673
timestamp 1679585382
transform 1 0 65184 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_680
timestamp 1679585382
transform 1 0 65856 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_687
timestamp 1679585382
transform 1 0 66528 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_694
timestamp 1679585382
transform 1 0 67200 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_701
timestamp 1679585382
transform 1 0 67872 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_708
timestamp 1679585382
transform 1 0 68544 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_715
timestamp 1679585382
transform 1 0 69216 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_722
timestamp 1679585382
transform 1 0 69888 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_729
timestamp 1679585382
transform 1 0 70560 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_736
timestamp 1679585382
transform 1 0 71232 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_743
timestamp 1679585382
transform 1 0 71904 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_750
timestamp 1679585382
transform 1 0 72576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_757
timestamp 1679585382
transform 1 0 73248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_764
timestamp 1679585382
transform 1 0 73920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_771
timestamp 1679585382
transform 1 0 74592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_778
timestamp 1679585382
transform 1 0 75264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_785
timestamp 1679585382
transform 1 0 75936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_792
timestamp 1679585382
transform 1 0 76608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_799
timestamp 1679585382
transform 1 0 77280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_806
timestamp 1679585382
transform 1 0 77952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_813
timestamp 1679585382
transform 1 0 78624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_820
timestamp 1679585382
transform 1 0 79296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_827
timestamp 1679585382
transform 1 0 79968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_834
timestamp 1679585382
transform 1 0 80640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_841
timestamp 1679585382
transform 1 0 81312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_848
timestamp 1679585382
transform 1 0 81984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_855
timestamp 1679585382
transform 1 0 82656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_862
timestamp 1679585382
transform 1 0 83328 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_869
timestamp 1679585382
transform 1 0 84000 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_876
timestamp 1679585382
transform 1 0 84672 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_883
timestamp 1679585382
transform 1 0 85344 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_890
timestamp 1679585382
transform 1 0 86016 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_897
timestamp 1679585382
transform 1 0 86688 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_904
timestamp 1679585382
transform 1 0 87360 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_911
timestamp 1679585382
transform 1 0 88032 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_918
timestamp 1679585382
transform 1 0 88704 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_925
timestamp 1679585382
transform 1 0 89376 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_932
timestamp 1679585382
transform 1 0 90048 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_939
timestamp 1679585382
transform 1 0 90720 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_946
timestamp 1679585382
transform 1 0 91392 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_953
timestamp 1679585382
transform 1 0 92064 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_960
timestamp 1679585382
transform 1 0 92736 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_967
timestamp 1679585382
transform 1 0 93408 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_974
timestamp 1679585382
transform 1 0 94080 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_981
timestamp 1679585382
transform 1 0 94752 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_988
timestamp 1679585382
transform 1 0 95424 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_995
timestamp 1679585382
transform 1 0 96096 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1002
timestamp 1679585382
transform 1 0 96768 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1009
timestamp 1679585382
transform 1 0 97440 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1016
timestamp 1679585382
transform 1 0 98112 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_1023
timestamp 1679581501
transform 1 0 98784 0 1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_1027
timestamp 1677583704
transform 1 0 99168 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_0
timestamp 1679585382
transform 1 0 576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_7
timestamp 1679585382
transform 1 0 1248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_14
timestamp 1679585382
transform 1 0 1920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_21
timestamp 1679585382
transform 1 0 2592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_28
timestamp 1679585382
transform 1 0 3264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_35
timestamp 1679585382
transform 1 0 3936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_42
timestamp 1679585382
transform 1 0 4608 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_47_49
timestamp 1677583704
transform 1 0 5280 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_51
timestamp 1677583258
transform 1 0 5472 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_4  FILLER_47_56
timestamp 1679581501
transform 1 0 5952 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_47_60
timestamp 1677583704
transform 1 0 6336 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_71
timestamp 1679585382
transform 1 0 7392 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_78
timestamp 1679585382
transform 1 0 8064 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_85
timestamp 1679581501
transform 1 0 8736 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_47_89
timestamp 1677583704
transform 1 0 9120 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_118
timestamp 1679585382
transform 1 0 11904 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_125
timestamp 1679585382
transform 1 0 12576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_132
timestamp 1679585382
transform 1 0 13248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_139
timestamp 1679585382
transform 1 0 13920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_146
timestamp 1679585382
transform 1 0 14592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_153
timestamp 1679585382
transform 1 0 15264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_160
timestamp 1679585382
transform 1 0 15936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_167
timestamp 1679585382
transform 1 0 16608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_174
timestamp 1679585382
transform 1 0 17280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_181
timestamp 1679585382
transform 1 0 17952 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_1  FILLER_47_188
timestamp 1677583258
transform 1 0 18624 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_225
timestamp 1679585382
transform 1 0 22176 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_232
timestamp 1679585382
transform 1 0 22848 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_239
timestamp 1679585382
transform 1 0 23520 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_47_246
timestamp 1677583704
transform 1 0 24192 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_248
timestamp 1677583258
transform 1 0 24384 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_276
timestamp 1679585382
transform 1 0 27072 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_283
timestamp 1679585382
transform 1 0 27744 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_290
timestamp 1679585382
transform 1 0 28416 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_297
timestamp 1679585382
transform 1 0 29088 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_304
timestamp 1679585382
transform 1 0 29760 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_311
timestamp 1679585382
transform 1 0 30432 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_322
timestamp 1679581501
transform 1 0 31488 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_47_326
timestamp 1677583704
transform 1 0 31872 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_337
timestamp 1679585382
transform 1 0 32928 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_344
timestamp 1679585382
transform 1 0 33600 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_351
timestamp 1679585382
transform 1 0 34272 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_358
timestamp 1679585382
transform 1 0 34944 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_365
timestamp 1679585382
transform 1 0 35616 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_47_372
timestamp 1677583704
transform 1 0 36288 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_401
timestamp 1679585382
transform 1 0 39072 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_408
timestamp 1679585382
transform 1 0 39744 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_415
timestamp 1679585382
transform 1 0 40416 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_422
timestamp 1679585382
transform 1 0 41088 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_429
timestamp 1679585382
transform 1 0 41760 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_436
timestamp 1679585382
transform 1 0 42432 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_443
timestamp 1679585382
transform 1 0 43104 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_450
timestamp 1679585382
transform 1 0 43776 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_457
timestamp 1679585382
transform 1 0 44448 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_464
timestamp 1679585382
transform 1 0 45120 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_471
timestamp 1679585382
transform 1 0 45792 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_478
timestamp 1679585382
transform 1 0 46464 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_485
timestamp 1679585382
transform 1 0 47136 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_492
timestamp 1679585382
transform 1 0 47808 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_499
timestamp 1679585382
transform 1 0 48480 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_506
timestamp 1679585382
transform 1 0 49152 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_513
timestamp 1679585382
transform 1 0 49824 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_520
timestamp 1679585382
transform 1 0 50496 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_527
timestamp 1679585382
transform 1 0 51168 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_534
timestamp 1679585382
transform 1 0 51840 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_541
timestamp 1679585382
transform 1 0 52512 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_548
timestamp 1679585382
transform 1 0 53184 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_555
timestamp 1679585382
transform 1 0 53856 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_562
timestamp 1679585382
transform 1 0 54528 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_569
timestamp 1679585382
transform 1 0 55200 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_576
timestamp 1679585382
transform 1 0 55872 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_583
timestamp 1679585382
transform 1 0 56544 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_590
timestamp 1679585382
transform 1 0 57216 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_597
timestamp 1679585382
transform 1 0 57888 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_604
timestamp 1679585382
transform 1 0 58560 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_611
timestamp 1679585382
transform 1 0 59232 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_618
timestamp 1679585382
transform 1 0 59904 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_625
timestamp 1679585382
transform 1 0 60576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_632
timestamp 1679585382
transform 1 0 61248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_639
timestamp 1679585382
transform 1 0 61920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_646
timestamp 1679585382
transform 1 0 62592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_653
timestamp 1679585382
transform 1 0 63264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_660
timestamp 1679585382
transform 1 0 63936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_667
timestamp 1679585382
transform 1 0 64608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_674
timestamp 1679585382
transform 1 0 65280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_681
timestamp 1679585382
transform 1 0 65952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_688
timestamp 1679585382
transform 1 0 66624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_695
timestamp 1679585382
transform 1 0 67296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_702
timestamp 1679585382
transform 1 0 67968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_709
timestamp 1679585382
transform 1 0 68640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_716
timestamp 1679585382
transform 1 0 69312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_723
timestamp 1679585382
transform 1 0 69984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_730
timestamp 1679585382
transform 1 0 70656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_737
timestamp 1679585382
transform 1 0 71328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_744
timestamp 1679585382
transform 1 0 72000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_751
timestamp 1679585382
transform 1 0 72672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_758
timestamp 1679585382
transform 1 0 73344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_765
timestamp 1679585382
transform 1 0 74016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_772
timestamp 1679585382
transform 1 0 74688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_779
timestamp 1679585382
transform 1 0 75360 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_786
timestamp 1679585382
transform 1 0 76032 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_793
timestamp 1679585382
transform 1 0 76704 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_800
timestamp 1679585382
transform 1 0 77376 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_807
timestamp 1679585382
transform 1 0 78048 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_814
timestamp 1679585382
transform 1 0 78720 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_821
timestamp 1679585382
transform 1 0 79392 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_828
timestamp 1679585382
transform 1 0 80064 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_835
timestamp 1679585382
transform 1 0 80736 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_842
timestamp 1679585382
transform 1 0 81408 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_849
timestamp 1679585382
transform 1 0 82080 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_856
timestamp 1679585382
transform 1 0 82752 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_863
timestamp 1679585382
transform 1 0 83424 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_870
timestamp 1679585382
transform 1 0 84096 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_877
timestamp 1679585382
transform 1 0 84768 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_884
timestamp 1679585382
transform 1 0 85440 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_891
timestamp 1679585382
transform 1 0 86112 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_898
timestamp 1679585382
transform 1 0 86784 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_905
timestamp 1679585382
transform 1 0 87456 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_912
timestamp 1679585382
transform 1 0 88128 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_919
timestamp 1679585382
transform 1 0 88800 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_926
timestamp 1679585382
transform 1 0 89472 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_933
timestamp 1679585382
transform 1 0 90144 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_940
timestamp 1679585382
transform 1 0 90816 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_947
timestamp 1679585382
transform 1 0 91488 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_954
timestamp 1679585382
transform 1 0 92160 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_961
timestamp 1679585382
transform 1 0 92832 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_968
timestamp 1679585382
transform 1 0 93504 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_975
timestamp 1679585382
transform 1 0 94176 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_982
timestamp 1679585382
transform 1 0 94848 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_989
timestamp 1679585382
transform 1 0 95520 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_996
timestamp 1679585382
transform 1 0 96192 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1003
timestamp 1679585382
transform 1 0 96864 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1010
timestamp 1679585382
transform 1 0 97536 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1017
timestamp 1679585382
transform 1 0 98208 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_47_1024
timestamp 1679581501
transform 1 0 98880 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_47_1028
timestamp 1677583258
transform 1 0 99264 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_0
timestamp 1679585382
transform 1 0 576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_7
timestamp 1679585382
transform 1 0 1248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_14
timestamp 1679585382
transform 1 0 1920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_21
timestamp 1679585382
transform 1 0 2592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_28
timestamp 1679585382
transform 1 0 3264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_35
timestamp 1679585382
transform 1 0 3936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_42
timestamp 1679585382
transform 1 0 4608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_49
timestamp 1679585382
transform 1 0 5280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_56
timestamp 1679585382
transform 1 0 5952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_63
timestamp 1679585382
transform 1 0 6624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_70
timestamp 1679585382
transform 1 0 7296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_77
timestamp 1679585382
transform 1 0 7968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_48_84
timestamp 1679581501
transform 1 0 8640 0 1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_48_88
timestamp 1677583704
transform 1 0 9024 0 1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_48_103
timestamp 1679585382
transform 1 0 10464 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_110
timestamp 1679585382
transform 1 0 11136 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_117
timestamp 1679585382
transform 1 0 11808 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_124
timestamp 1679585382
transform 1 0 12480 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_131
timestamp 1679585382
transform 1 0 13152 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_138
timestamp 1679585382
transform 1 0 13824 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_145
timestamp 1679585382
transform 1 0 14496 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_152
timestamp 1679585382
transform 1 0 15168 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_159
timestamp 1679585382
transform 1 0 15840 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_166
timestamp 1679585382
transform 1 0 16512 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_173
timestamp 1679585382
transform 1 0 17184 0 1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_48_180
timestamp 1679581501
transform 1 0 17856 0 1 37044
box -48 -56 432 834
use sg13g2_decap_8  FILLER_48_220
timestamp 1679585382
transform 1 0 21696 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_227
timestamp 1679585382
transform 1 0 22368 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_234
timestamp 1679585382
transform 1 0 23040 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_241
timestamp 1679585382
transform 1 0 23712 0 1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_48_248
timestamp 1677583704
transform 1 0 24384 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_250
timestamp 1677583258
transform 1 0 24576 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_260
timestamp 1679585382
transform 1 0 25536 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_267
timestamp 1679585382
transform 1 0 26208 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_274
timestamp 1679585382
transform 1 0 26880 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_281
timestamp 1679585382
transform 1 0 27552 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_288
timestamp 1679585382
transform 1 0 28224 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_295
timestamp 1679585382
transform 1 0 28896 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_302
timestamp 1679585382
transform 1 0 29568 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_309
timestamp 1679585382
transform 1 0 30240 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_316
timestamp 1679585382
transform 1 0 30912 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_323
timestamp 1679585382
transform 1 0 31584 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_330
timestamp 1679585382
transform 1 0 32256 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_337
timestamp 1679585382
transform 1 0 32928 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_344
timestamp 1679585382
transform 1 0 33600 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_351
timestamp 1679585382
transform 1 0 34272 0 1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_48_358
timestamp 1677583704
transform 1 0 34944 0 1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_48_387
timestamp 1679585382
transform 1 0 37728 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_394
timestamp 1679585382
transform 1 0 38400 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_401
timestamp 1679585382
transform 1 0 39072 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_408
timestamp 1679585382
transform 1 0 39744 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_415
timestamp 1679585382
transform 1 0 40416 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_422
timestamp 1679585382
transform 1 0 41088 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_429
timestamp 1679585382
transform 1 0 41760 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_436
timestamp 1679585382
transform 1 0 42432 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_443
timestamp 1679585382
transform 1 0 43104 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_450
timestamp 1679585382
transform 1 0 43776 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_457
timestamp 1679585382
transform 1 0 44448 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_464
timestamp 1679585382
transform 1 0 45120 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_471
timestamp 1679585382
transform 1 0 45792 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_478
timestamp 1679585382
transform 1 0 46464 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_485
timestamp 1679585382
transform 1 0 47136 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_492
timestamp 1679585382
transform 1 0 47808 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_499
timestamp 1679585382
transform 1 0 48480 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_506
timestamp 1679585382
transform 1 0 49152 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_513
timestamp 1679585382
transform 1 0 49824 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_520
timestamp 1679585382
transform 1 0 50496 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_527
timestamp 1679585382
transform 1 0 51168 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_534
timestamp 1679585382
transform 1 0 51840 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_541
timestamp 1679585382
transform 1 0 52512 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_548
timestamp 1679585382
transform 1 0 53184 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_555
timestamp 1679585382
transform 1 0 53856 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_562
timestamp 1679585382
transform 1 0 54528 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_569
timestamp 1679585382
transform 1 0 55200 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_576
timestamp 1679585382
transform 1 0 55872 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_583
timestamp 1679585382
transform 1 0 56544 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_590
timestamp 1679585382
transform 1 0 57216 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_597
timestamp 1679585382
transform 1 0 57888 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_604
timestamp 1679585382
transform 1 0 58560 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_611
timestamp 1679585382
transform 1 0 59232 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_618
timestamp 1679585382
transform 1 0 59904 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_625
timestamp 1679585382
transform 1 0 60576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_632
timestamp 1679585382
transform 1 0 61248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_639
timestamp 1679585382
transform 1 0 61920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_646
timestamp 1679585382
transform 1 0 62592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_653
timestamp 1679585382
transform 1 0 63264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_660
timestamp 1679585382
transform 1 0 63936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_667
timestamp 1679585382
transform 1 0 64608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_674
timestamp 1679585382
transform 1 0 65280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_681
timestamp 1679585382
transform 1 0 65952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_688
timestamp 1679585382
transform 1 0 66624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_695
timestamp 1679585382
transform 1 0 67296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_702
timestamp 1679585382
transform 1 0 67968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_709
timestamp 1679585382
transform 1 0 68640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_716
timestamp 1679585382
transform 1 0 69312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_723
timestamp 1679585382
transform 1 0 69984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_730
timestamp 1679585382
transform 1 0 70656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_737
timestamp 1679585382
transform 1 0 71328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_744
timestamp 1679585382
transform 1 0 72000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_751
timestamp 1679585382
transform 1 0 72672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_758
timestamp 1679585382
transform 1 0 73344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_765
timestamp 1679585382
transform 1 0 74016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_772
timestamp 1679585382
transform 1 0 74688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_779
timestamp 1679585382
transform 1 0 75360 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_786
timestamp 1679585382
transform 1 0 76032 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_793
timestamp 1679585382
transform 1 0 76704 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_800
timestamp 1679585382
transform 1 0 77376 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_807
timestamp 1679585382
transform 1 0 78048 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_814
timestamp 1679585382
transform 1 0 78720 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_821
timestamp 1679585382
transform 1 0 79392 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_828
timestamp 1679585382
transform 1 0 80064 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_835
timestamp 1679585382
transform 1 0 80736 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_842
timestamp 1679585382
transform 1 0 81408 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_849
timestamp 1679585382
transform 1 0 82080 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_856
timestamp 1679585382
transform 1 0 82752 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_863
timestamp 1679585382
transform 1 0 83424 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_870
timestamp 1679585382
transform 1 0 84096 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_877
timestamp 1679585382
transform 1 0 84768 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_884
timestamp 1679585382
transform 1 0 85440 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_891
timestamp 1679585382
transform 1 0 86112 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_898
timestamp 1679585382
transform 1 0 86784 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_905
timestamp 1679585382
transform 1 0 87456 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_912
timestamp 1679585382
transform 1 0 88128 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_919
timestamp 1679585382
transform 1 0 88800 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_926
timestamp 1679585382
transform 1 0 89472 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_933
timestamp 1679585382
transform 1 0 90144 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_940
timestamp 1679585382
transform 1 0 90816 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_947
timestamp 1679585382
transform 1 0 91488 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_954
timestamp 1679585382
transform 1 0 92160 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_961
timestamp 1679585382
transform 1 0 92832 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_968
timestamp 1679585382
transform 1 0 93504 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_975
timestamp 1679585382
transform 1 0 94176 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_982
timestamp 1679585382
transform 1 0 94848 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_989
timestamp 1679585382
transform 1 0 95520 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_996
timestamp 1679585382
transform 1 0 96192 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1003
timestamp 1679585382
transform 1 0 96864 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1010
timestamp 1679585382
transform 1 0 97536 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1017
timestamp 1679585382
transform 1 0 98208 0 1 37044
box -48 -56 720 834
use sg13g2_decap_4  FILLER_48_1024
timestamp 1679581501
transform 1 0 98880 0 1 37044
box -48 -56 432 834
use sg13g2_fill_1  FILLER_48_1028
timestamp 1677583258
transform 1 0 99264 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_0
timestamp 1679585382
transform 1 0 576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_7
timestamp 1679585382
transform 1 0 1248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_14
timestamp 1679585382
transform 1 0 1920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_21
timestamp 1679585382
transform 1 0 2592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_28
timestamp 1679585382
transform 1 0 3264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_35
timestamp 1679585382
transform 1 0 3936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_42
timestamp 1679585382
transform 1 0 4608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_49
timestamp 1679585382
transform 1 0 5280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_56
timestamp 1679585382
transform 1 0 5952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_63
timestamp 1679585382
transform 1 0 6624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_70
timestamp 1679585382
transform 1 0 7296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_77
timestamp 1679585382
transform 1 0 7968 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_84
timestamp 1679585382
transform 1 0 8640 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_91
timestamp 1679585382
transform 1 0 9312 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_98
timestamp 1679585382
transform 1 0 9984 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_105
timestamp 1679585382
transform 1 0 10656 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_112
timestamp 1679585382
transform 1 0 11328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_119
timestamp 1679585382
transform 1 0 12000 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_126
timestamp 1679585382
transform 1 0 12672 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_133
timestamp 1679585382
transform 1 0 13344 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_140
timestamp 1679585382
transform 1 0 14016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_147
timestamp 1679585382
transform 1 0 14688 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_154
timestamp 1679585382
transform 1 0 15360 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_161
timestamp 1679585382
transform 1 0 16032 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_168
timestamp 1679585382
transform 1 0 16704 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_175
timestamp 1679585382
transform 1 0 17376 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_182
timestamp 1679585382
transform 1 0 18048 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_189
timestamp 1679585382
transform 1 0 18720 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_196
timestamp 1679585382
transform 1 0 19392 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_203
timestamp 1679585382
transform 1 0 20064 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_210
timestamp 1679585382
transform 1 0 20736 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_217
timestamp 1679585382
transform 1 0 21408 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_224
timestamp 1679585382
transform 1 0 22080 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_231
timestamp 1679585382
transform 1 0 22752 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_238
timestamp 1679585382
transform 1 0 23424 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_245
timestamp 1679585382
transform 1 0 24096 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_252
timestamp 1679585382
transform 1 0 24768 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_259
timestamp 1679585382
transform 1 0 25440 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_266
timestamp 1679585382
transform 1 0 26112 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_273
timestamp 1679585382
transform 1 0 26784 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_280
timestamp 1679585382
transform 1 0 27456 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_287
timestamp 1679585382
transform 1 0 28128 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_294
timestamp 1679585382
transform 1 0 28800 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_301
timestamp 1679585382
transform 1 0 29472 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_308
timestamp 1679585382
transform 1 0 30144 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_315
timestamp 1679585382
transform 1 0 30816 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_322
timestamp 1679585382
transform 1 0 31488 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_329
timestamp 1679585382
transform 1 0 32160 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_336
timestamp 1679585382
transform 1 0 32832 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_343
timestamp 1679585382
transform 1 0 33504 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_350
timestamp 1679585382
transform 1 0 34176 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_357
timestamp 1679585382
transform 1 0 34848 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_364
timestamp 1679585382
transform 1 0 35520 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_371
timestamp 1679581501
transform 1 0 36192 0 -1 38556
box -48 -56 432 834
use sg13g2_decap_8  FILLER_49_384
timestamp 1679585382
transform 1 0 37440 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_391
timestamp 1679585382
transform 1 0 38112 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_398
timestamp 1679585382
transform 1 0 38784 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_405
timestamp 1679585382
transform 1 0 39456 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_412
timestamp 1679585382
transform 1 0 40128 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_419
timestamp 1679585382
transform 1 0 40800 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_426
timestamp 1679585382
transform 1 0 41472 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_433
timestamp 1679585382
transform 1 0 42144 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_440
timestamp 1679585382
transform 1 0 42816 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_447
timestamp 1679585382
transform 1 0 43488 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_454
timestamp 1679585382
transform 1 0 44160 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_461
timestamp 1679585382
transform 1 0 44832 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_468
timestamp 1679585382
transform 1 0 45504 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_475
timestamp 1679585382
transform 1 0 46176 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_482
timestamp 1679585382
transform 1 0 46848 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_489
timestamp 1679585382
transform 1 0 47520 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_496
timestamp 1679585382
transform 1 0 48192 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_503
timestamp 1679585382
transform 1 0 48864 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_510
timestamp 1679585382
transform 1 0 49536 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_517
timestamp 1679585382
transform 1 0 50208 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_524
timestamp 1679585382
transform 1 0 50880 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_531
timestamp 1679585382
transform 1 0 51552 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_538
timestamp 1679585382
transform 1 0 52224 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_545
timestamp 1679585382
transform 1 0 52896 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_552
timestamp 1679585382
transform 1 0 53568 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_559
timestamp 1679585382
transform 1 0 54240 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_566
timestamp 1679585382
transform 1 0 54912 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_573
timestamp 1679585382
transform 1 0 55584 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_580
timestamp 1679585382
transform 1 0 56256 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_587
timestamp 1679585382
transform 1 0 56928 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_594
timestamp 1679585382
transform 1 0 57600 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_601
timestamp 1679585382
transform 1 0 58272 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_608
timestamp 1679585382
transform 1 0 58944 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_615
timestamp 1679585382
transform 1 0 59616 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_622
timestamp 1679585382
transform 1 0 60288 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_629
timestamp 1679585382
transform 1 0 60960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_636
timestamp 1679585382
transform 1 0 61632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_643
timestamp 1679585382
transform 1 0 62304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_650
timestamp 1679585382
transform 1 0 62976 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_657
timestamp 1679585382
transform 1 0 63648 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_664
timestamp 1679585382
transform 1 0 64320 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_671
timestamp 1679585382
transform 1 0 64992 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_678
timestamp 1679585382
transform 1 0 65664 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_685
timestamp 1679585382
transform 1 0 66336 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_692
timestamp 1679585382
transform 1 0 67008 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_699
timestamp 1679585382
transform 1 0 67680 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_706
timestamp 1679585382
transform 1 0 68352 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_713
timestamp 1679585382
transform 1 0 69024 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_720
timestamp 1679585382
transform 1 0 69696 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_727
timestamp 1679585382
transform 1 0 70368 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_734
timestamp 1679585382
transform 1 0 71040 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_741
timestamp 1679585382
transform 1 0 71712 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_748
timestamp 1679585382
transform 1 0 72384 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_755
timestamp 1679585382
transform 1 0 73056 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_762
timestamp 1679585382
transform 1 0 73728 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_769
timestamp 1679585382
transform 1 0 74400 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_776
timestamp 1679585382
transform 1 0 75072 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_783
timestamp 1679585382
transform 1 0 75744 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_790
timestamp 1679585382
transform 1 0 76416 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_797
timestamp 1679585382
transform 1 0 77088 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_804
timestamp 1679585382
transform 1 0 77760 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_811
timestamp 1679585382
transform 1 0 78432 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_818
timestamp 1679585382
transform 1 0 79104 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_825
timestamp 1679585382
transform 1 0 79776 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_832
timestamp 1679585382
transform 1 0 80448 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_839
timestamp 1679585382
transform 1 0 81120 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_846
timestamp 1679585382
transform 1 0 81792 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_853
timestamp 1679585382
transform 1 0 82464 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_860
timestamp 1679585382
transform 1 0 83136 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_867
timestamp 1679585382
transform 1 0 83808 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_874
timestamp 1679585382
transform 1 0 84480 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_881
timestamp 1679585382
transform 1 0 85152 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_888
timestamp 1679585382
transform 1 0 85824 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_895
timestamp 1679585382
transform 1 0 86496 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_902
timestamp 1679585382
transform 1 0 87168 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_909
timestamp 1679585382
transform 1 0 87840 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_916
timestamp 1679585382
transform 1 0 88512 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_923
timestamp 1679585382
transform 1 0 89184 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_930
timestamp 1679585382
transform 1 0 89856 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_937
timestamp 1679585382
transform 1 0 90528 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_944
timestamp 1679585382
transform 1 0 91200 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_951
timestamp 1679585382
transform 1 0 91872 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_958
timestamp 1679585382
transform 1 0 92544 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_965
timestamp 1679585382
transform 1 0 93216 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_972
timestamp 1679585382
transform 1 0 93888 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_979
timestamp 1679585382
transform 1 0 94560 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_986
timestamp 1679585382
transform 1 0 95232 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_993
timestamp 1679585382
transform 1 0 95904 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1000
timestamp 1679585382
transform 1 0 96576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1007
timestamp 1679585382
transform 1 0 97248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1014
timestamp 1679585382
transform 1 0 97920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1021
timestamp 1679585382
transform 1 0 98592 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_1  FILLER_49_1028
timestamp 1677583258
transform 1 0 99264 0 -1 38556
box -48 -56 144 834
use sg13g2_tielo  heichips25_template_5
timestamp 1680004237
transform -1 0 960 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_6
timestamp 1680004237
transform -1 0 960 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_7
timestamp 1680004237
transform -1 0 960 0 -1 11340
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_8
timestamp 1680004237
transform -1 0 960 0 1 11340
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_9
timestamp 1680004237
transform -1 0 960 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_10
timestamp 1680004237
transform -1 0 960 0 1 12852
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_11
timestamp 1680004237
transform -1 0 960 0 1 14364
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_12
timestamp 1680004237
transform -1 0 960 0 -1 15876
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_13
timestamp 1680004237
transform -1 0 960 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_14
timestamp 1680004237
transform -1 0 960 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_15
timestamp 1680004237
transform -1 0 960 0 -1 8316
box -48 -56 432 834
use sg13g2_tielo  heichips25_template_16
timestamp 1680004237
transform -1 0 960 0 1 8316
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_17
timestamp 1680004251
transform -1 0 960 0 1 15876
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_18
timestamp 1680004251
transform -1 0 960 0 -1 17388
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_19
timestamp 1680004251
transform -1 0 960 0 1 17388
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_20
timestamp 1680004251
transform -1 0 960 0 -1 18900
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_21
timestamp 1680004251
transform -1 0 960 0 1 18900
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_22
timestamp 1680004251
transform -1 0 960 0 -1 20412
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_23
timestamp 1680004251
transform -1 0 960 0 1 20412
box -48 -56 432 834
use sg13g2_tiehi  heichips25_template_24
timestamp 1680004251
transform -1 0 960 0 1 21924
box -48 -56 432 834
use sg13g2_dlygate4sd3_1  hold1
timestamp 1677675658
transform -1 0 13728 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold2
timestamp 1677675658
transform 1 0 27264 0 1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold3
timestamp 1677675658
transform 1 0 23712 0 1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold4
timestamp 1677675658
transform 1 0 9600 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold5
timestamp 1677675658
transform 1 0 30912 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold6
timestamp 1677675658
transform -1 0 13152 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold7
timestamp 1677675658
transform 1 0 30144 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold8
timestamp 1677675658
transform 1 0 9792 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold9
timestamp 1677675658
transform 1 0 15360 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold10
timestamp 1677675658
transform 1 0 26784 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold11
timestamp 1677675658
transform 1 0 22848 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold12
timestamp 1677675658
transform 1 0 15744 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold13
timestamp 1677675658
transform 1 0 33792 0 -1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold14
timestamp 1677675658
transform 1 0 34464 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold15
timestamp 1677675658
transform -1 0 37632 0 1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold16
timestamp 1677675658
transform -1 0 57600 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold17
timestamp 1677675658
transform -1 0 12864 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold18
timestamp 1677675658
transform -1 0 16992 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold19
timestamp 1677675658
transform 1 0 6144 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold20
timestamp 1677675658
transform -1 0 5856 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold21
timestamp 1677675658
transform -1 0 45600 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold22
timestamp 1677675658
transform -1 0 61536 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold23
timestamp 1677675658
transform 1 0 17088 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold24
timestamp 1677675658
transform -1 0 29184 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold25
timestamp 1677675658
transform -1 0 50496 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold26
timestamp 1677675658
transform -1 0 10464 0 1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold27
timestamp 1677675658
transform -1 0 49344 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold28
timestamp 1677675658
transform -1 0 7392 0 -1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold29
timestamp 1677675658
transform 1 0 40896 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold30
timestamp 1677675658
transform 1 0 21312 0 -1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold31
timestamp 1677675658
transform -1 0 61920 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold32
timestamp 1677675658
transform -1 0 32928 0 -1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold33
timestamp 1677675658
transform -1 0 4896 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold34
timestamp 1677675658
transform -1 0 48480 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold35
timestamp 1677675658
transform -1 0 4800 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold36
timestamp 1677675658
transform -1 0 54144 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold37
timestamp 1677675658
transform 1 0 2016 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold38
timestamp 1677675658
transform -1 0 17568 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold39
timestamp 1677675658
transform 1 0 42816 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold40
timestamp 1677675658
transform -1 0 17856 0 1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold41
timestamp 1677675658
transform -1 0 35232 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold42
timestamp 1677675658
transform 1 0 36480 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold43
timestamp 1677675658
transform -1 0 4992 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold44
timestamp 1677675658
transform 1 0 2016 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold45
timestamp 1677675658
transform -1 0 28320 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold46
timestamp 1677675658
transform 1 0 14784 0 1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold47
timestamp 1677675658
transform 1 0 38880 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold48
timestamp 1677675658
transform -1 0 40224 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold49
timestamp 1677675658
transform 1 0 20832 0 1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold50
timestamp 1677675658
transform 1 0 45696 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold51
timestamp 1677675658
transform 1 0 33120 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold52
timestamp 1677675658
transform 1 0 37824 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold53
timestamp 1677675658
transform -1 0 39264 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold54
timestamp 1677675658
transform -1 0 19296 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold55
timestamp 1677675658
transform 1 0 15168 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold56
timestamp 1677675658
transform 1 0 16992 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold57
timestamp 1677675658
transform 1 0 20256 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold58
timestamp 1677675658
transform 1 0 21792 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold59
timestamp 1677675658
transform -1 0 49344 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold60
timestamp 1677675658
transform 1 0 46272 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold61
timestamp 1677675658
transform 1 0 10080 0 1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold62
timestamp 1677675658
transform 1 0 10752 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold63
timestamp 1677675658
transform -1 0 12960 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold64
timestamp 1677675658
transform 1 0 12960 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold65
timestamp 1677675658
transform 1 0 41664 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold66
timestamp 1677675658
transform -1 0 41280 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold67
timestamp 1677675658
transform -1 0 27744 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold68
timestamp 1677675658
transform 1 0 26016 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold69
timestamp 1677675658
transform -1 0 18816 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold70
timestamp 1677675658
transform -1 0 20256 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold71
timestamp 1677675658
transform 1 0 28704 0 -1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold72
timestamp 1677675658
transform -1 0 28512 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold73
timestamp 1677675658
transform -1 0 40512 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold74
timestamp 1677675658
transform -1 0 6336 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold75
timestamp 1677675658
transform -1 0 11424 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold76
timestamp 1677675658
transform -1 0 56160 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold77
timestamp 1677675658
transform -1 0 53760 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold78
timestamp 1677675658
transform 1 0 51264 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold79
timestamp 1677675658
transform 1 0 48576 0 1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold80
timestamp 1677675658
transform -1 0 47424 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold81
timestamp 1677675658
transform -1 0 35040 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold82
timestamp 1677675658
transform -1 0 50304 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold83
timestamp 1677675658
transform -1 0 33024 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold84
timestamp 1677675658
transform -1 0 5376 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold85
timestamp 1677675658
transform -1 0 54336 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold86
timestamp 1677675658
transform 1 0 4512 0 1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold87
timestamp 1677675658
transform -1 0 6240 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold88
timestamp 1677675658
transform -1 0 10464 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold89
timestamp 1677675658
transform -1 0 25536 0 1 37044
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold90
timestamp 1677675658
transform -1 0 28416 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold91
timestamp 1677675658
transform -1 0 6240 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold92
timestamp 1677675658
transform -1 0 5568 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold93
timestamp 1677675658
transform -1 0 45120 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold94
timestamp 1677675658
transform -1 0 6624 0 -1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold95
timestamp 1677675658
transform -1 0 18048 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold96
timestamp 1677675658
transform -1 0 47616 0 -1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold97
timestamp 1677675658
transform 1 0 37536 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold98
timestamp 1677675658
transform 1 0 39552 0 1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold99
timestamp 1677675658
transform 1 0 17472 0 -1 34020
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold100
timestamp 1677675658
transform 1 0 16224 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold101
timestamp 1677675658
transform 1 0 28224 0 1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold102
timestamp 1677675658
transform -1 0 23712 0 -1 24948
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold103
timestamp 1677675658
transform -1 0 21120 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold104
timestamp 1677675658
transform -1 0 56640 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold105
timestamp 1677675658
transform -1 0 5280 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold106
timestamp 1677675658
transform -1 0 57600 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold107
timestamp 1677675658
transform 1 0 33696 0 -1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold108
timestamp 1677675658
transform -1 0 47136 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold109
timestamp 1677675658
transform -1 0 19296 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold110
timestamp 1677675658
transform -1 0 40896 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold111
timestamp 1677675658
transform -1 0 37440 0 -1 38556
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold112
timestamp 1677675658
transform -1 0 46848 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold113
timestamp 1677675658
transform -1 0 26976 0 1 35532
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold114
timestamp 1677675658
transform -1 0 54144 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold115
timestamp 1677675658
transform -1 0 36480 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold116
timestamp 1677675658
transform -1 0 29280 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold117
timestamp 1677675658
transform 1 0 33504 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold118
timestamp 1677675658
transform -1 0 34272 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold119
timestamp 1677675658
transform -1 0 33888 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold120
timestamp 1677675658
transform 1 0 23328 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold121
timestamp 1677675658
transform 1 0 23424 0 1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold122
timestamp 1677675658
transform 1 0 26016 0 1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold123
timestamp 1677675658
transform 1 0 38592 0 -1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold124
timestamp 1677675658
transform 1 0 41376 0 1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold125
timestamp 1677675658
transform -1 0 11904 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold126
timestamp 1677675658
transform -1 0 12000 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold127
timestamp 1677675658
transform 1 0 11520 0 -1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold128
timestamp 1677675658
transform -1 0 57312 0 1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold129
timestamp 1677675658
transform -1 0 56832 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold130
timestamp 1677675658
transform 1 0 10944 0 -1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold131
timestamp 1677675658
transform 1 0 12672 0 1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold132
timestamp 1677675658
transform 1 0 45600 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold133
timestamp 1677675658
transform 1 0 47136 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold134
timestamp 1677675658
transform 1 0 24192 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold135
timestamp 1677675658
transform 1 0 26688 0 -1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold136
timestamp 1677675658
transform 1 0 16128 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold137
timestamp 1677675658
transform 1 0 17760 0 -1 26460
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold138
timestamp 1677675658
transform 1 0 39840 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold139
timestamp 1677675658
transform -1 0 41184 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold140
timestamp 1677675658
transform 1 0 40704 0 -1 20412
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold141
timestamp 1677675658
transform -1 0 50304 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold142
timestamp 1677675658
transform -1 0 48096 0 -1 14364
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold143
timestamp 1677675658
transform -1 0 34176 0 -1 18900
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold144
timestamp 1677675658
transform 1 0 33696 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold145
timestamp 1677675658
transform 1 0 35328 0 -1 17388
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold146
timestamp 1677675658
transform 1 0 20736 0 1 23436
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold147
timestamp 1677675658
transform -1 0 22080 0 1 21924
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold148
timestamp 1677675658
transform -1 0 31296 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold149
timestamp 1677675658
transform -1 0 30720 0 -1 29484
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold150
timestamp 1677675658
transform -1 0 27264 0 1 27972
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold151
timestamp 1677675658
transform 1 0 36864 0 1 32508
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold152
timestamp 1677675658
transform -1 0 36288 0 1 30996
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold153
timestamp 1677675658
transform 1 0 41568 0 1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold154
timestamp 1677675658
transform -1 0 41472 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold155
timestamp 1677675658
transform -1 0 34272 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold156
timestamp 1677675658
transform -1 0 32448 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold157
timestamp 1677675658
transform -1 0 23040 0 -1 15876
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold158
timestamp 1677675658
transform 1 0 24096 0 1 11340
box -48 -56 912 834
use sg13g2_buf_1  output1
timestamp 1676385511
transform -1 0 960 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  output2
timestamp 1676385511
transform -1 0 960 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  output3
timestamp 1676385511
transform -1 0 960 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  output4
timestamp 1676385511
transform -1 0 960 0 -1 5292
box -48 -56 432 834
<< labels >>
flabel metal6 s 4316 630 4756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 19436 630 19876 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 34556 630 34996 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 49676 630 50116 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 64796 630 65236 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 79916 630 80356 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 95036 630 95476 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 3076 712 3516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 18196 712 18636 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 33316 712 33756 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 48436 712 48876 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 63556 712 63996 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 78676 712 79116 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 93796 712 94236 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 36668 80 36748 0 FreeSans 320 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 0 35828 80 35908 0 FreeSans 320 0 0 0 ena
port 3 nsew signal input
flabel metal3 s 0 37508 80 37588 0 FreeSans 320 0 0 0 rst_n
port 4 nsew signal input
flabel metal3 s 0 22388 80 22468 0 FreeSans 320 0 0 0 ui_in[0]
port 5 nsew signal input
flabel metal3 s 0 23228 80 23308 0 FreeSans 320 0 0 0 ui_in[1]
port 6 nsew signal input
flabel metal3 s 0 24068 80 24148 0 FreeSans 320 0 0 0 ui_in[2]
port 7 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 ui_in[3]
port 8 nsew signal input
flabel metal3 s 0 25748 80 25828 0 FreeSans 320 0 0 0 ui_in[4]
port 9 nsew signal input
flabel metal3 s 0 26588 80 26668 0 FreeSans 320 0 0 0 ui_in[5]
port 10 nsew signal input
flabel metal3 s 0 27428 80 27508 0 FreeSans 320 0 0 0 ui_in[6]
port 11 nsew signal input
flabel metal3 s 0 28268 80 28348 0 FreeSans 320 0 0 0 ui_in[7]
port 12 nsew signal input
flabel metal3 s 0 29108 80 29188 0 FreeSans 320 0 0 0 uio_in[0]
port 13 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 uio_in[1]
port 14 nsew signal input
flabel metal3 s 0 30788 80 30868 0 FreeSans 320 0 0 0 uio_in[2]
port 15 nsew signal input
flabel metal3 s 0 31628 80 31708 0 FreeSans 320 0 0 0 uio_in[3]
port 16 nsew signal input
flabel metal3 s 0 32468 80 32548 0 FreeSans 320 0 0 0 uio_in[4]
port 17 nsew signal input
flabel metal3 s 0 33308 80 33388 0 FreeSans 320 0 0 0 uio_in[5]
port 18 nsew signal input
flabel metal3 s 0 34148 80 34228 0 FreeSans 320 0 0 0 uio_in[6]
port 19 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 uio_in[7]
port 20 nsew signal input
flabel metal3 s 0 15668 80 15748 0 FreeSans 320 0 0 0 uio_oe[0]
port 21 nsew signal output
flabel metal3 s 0 16508 80 16588 0 FreeSans 320 0 0 0 uio_oe[1]
port 22 nsew signal output
flabel metal3 s 0 17348 80 17428 0 FreeSans 320 0 0 0 uio_oe[2]
port 23 nsew signal output
flabel metal3 s 0 18188 80 18268 0 FreeSans 320 0 0 0 uio_oe[3]
port 24 nsew signal output
flabel metal3 s 0 19028 80 19108 0 FreeSans 320 0 0 0 uio_oe[4]
port 25 nsew signal output
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 uio_oe[5]
port 26 nsew signal output
flabel metal3 s 0 20708 80 20788 0 FreeSans 320 0 0 0 uio_oe[6]
port 27 nsew signal output
flabel metal3 s 0 21548 80 21628 0 FreeSans 320 0 0 0 uio_oe[7]
port 28 nsew signal output
flabel metal3 s 0 8948 80 9028 0 FreeSans 320 0 0 0 uio_out[0]
port 29 nsew signal output
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 uio_out[1]
port 30 nsew signal output
flabel metal3 s 0 10628 80 10708 0 FreeSans 320 0 0 0 uio_out[2]
port 31 nsew signal output
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 uio_out[3]
port 32 nsew signal output
flabel metal3 s 0 12308 80 12388 0 FreeSans 320 0 0 0 uio_out[4]
port 33 nsew signal output
flabel metal3 s 0 13148 80 13228 0 FreeSans 320 0 0 0 uio_out[5]
port 34 nsew signal output
flabel metal3 s 0 13988 80 14068 0 FreeSans 320 0 0 0 uio_out[6]
port 35 nsew signal output
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 uio_out[7]
port 36 nsew signal output
flabel metal3 s 0 2228 80 2308 0 FreeSans 320 0 0 0 uo_out[0]
port 37 nsew signal output
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 uo_out[1]
port 38 nsew signal output
flabel metal3 s 0 3908 80 3988 0 FreeSans 320 0 0 0 uo_out[2]
port 39 nsew signal output
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 uo_out[3]
port 40 nsew signal output
flabel metal3 s 0 5588 80 5668 0 FreeSans 320 0 0 0 uo_out[4]
port 41 nsew signal output
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 uo_out[5]
port 42 nsew signal output
flabel metal3 s 0 7268 80 7348 0 FreeSans 320 0 0 0 uo_out[6]
port 43 nsew signal output
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 uo_out[7]
port 44 nsew signal output
rlabel via1 49968 38556 49968 38556 0 VGND
rlabel metal1 49968 37800 49968 37800 0 VPWR
rlabel metal2 56592 8484 56592 8484 0 DP_1.matrix\[0\]
rlabel metal2 19248 13440 19248 13440 0 DP_1.matrix\[112\]
rlabel metal2 17184 16254 17184 16254 0 DP_1.matrix\[113\]
rlabel metal2 18720 3864 18720 3864 0 DP_1.matrix\[128\]
rlabel metal2 19152 5880 19152 5880 0 DP_1.matrix\[129\]
rlabel metal2 51360 18522 51360 18522 0 DP_1.matrix\[16\]
rlabel metal3 57792 19488 57792 19488 0 DP_1.matrix\[17\]
rlabel metal2 62016 9912 62016 9912 0 DP_1.matrix\[1\]
rlabel metal2 40512 3150 40512 3150 0 DP_1.matrix\[32\]
rlabel metal2 36000 5250 36000 5250 0 DP_1.matrix\[33\]
rlabel metal2 54336 5250 54336 5250 0 DP_1.matrix\[48\]
rlabel metal3 54336 2856 54336 2856 0 DP_1.matrix\[49\]
rlabel metal2 34848 21714 34848 21714 0 DP_1.matrix\[64\]
rlabel metal3 32880 26796 32880 26796 0 DP_1.matrix\[65\]
rlabel metal2 46752 20706 46752 20706 0 DP_1.matrix\[80\]
rlabel metal2 42912 26838 42912 26838 0 DP_1.matrix\[81\]
rlabel metal2 28608 17472 28608 17472 0 DP_1.matrix\[96\]
rlabel metal2 29040 21504 29040 21504 0 DP_1.matrix\[97\]
rlabel metal2 57504 8946 57504 8946 0 DP_2.matrix\[0\]
rlabel metal3 20736 16380 20736 16380 0 DP_2.matrix\[112\]
rlabel metal2 17280 17472 17280 17472 0 DP_2.matrix\[113\]
rlabel metal2 14208 3864 14208 3864 0 DP_2.matrix\[128\]
rlabel metal2 14880 2646 14880 2646 0 DP_2.matrix\[129\]
rlabel metal2 54240 19530 54240 19530 0 DP_2.matrix\[16\]
rlabel metal2 50208 17262 50208 17262 0 DP_2.matrix\[17\]
rlabel metal2 62016 11424 62016 11424 0 DP_2.matrix\[1\]
rlabel metal2 40368 6636 40368 6636 0 DP_2.matrix\[32\]
rlabel metal2 40800 2856 40800 2856 0 DP_2.matrix\[33\]
rlabel metal2 50016 3150 50016 3150 0 DP_2.matrix\[48\]
rlabel metal3 45408 2856 45408 2856 0 DP_2.matrix\[49\]
rlabel metal3 33216 23100 33216 23100 0 DP_2.matrix\[64\]
rlabel metal2 35136 26376 35136 26376 0 DP_2.matrix\[65\]
rlabel metal2 47616 25830 47616 25830 0 DP_2.matrix\[80\]
rlabel metal2 48384 23856 48384 23856 0 DP_2.matrix\[81\]
rlabel metal2 28128 18270 28128 18270 0 DP_2.matrix\[96\]
rlabel metal2 28176 22512 28176 22512 0 DP_2.matrix\[97\]
rlabel metal2 47808 33390 47808 33390 0 DP_3.matrix\[0\]
rlabel metal3 11616 14196 11616 14196 0 DP_3.matrix\[112\]
rlabel metal2 6384 13440 6384 13440 0 DP_3.matrix\[113\]
rlabel metal2 5424 7980 5424 7980 0 DP_3.matrix\[128\]
rlabel metal2 1344 5376 1344 5376 0 DP_3.matrix\[129\]
rlabel metal2 37632 37926 37632 37926 0 DP_3.matrix\[16\]
rlabel metal2 32640 36414 32640 36414 0 DP_3.matrix\[17\]
rlabel metal2 46944 28854 46944 28854 0 DP_3.matrix\[1\]
rlabel metal2 26928 35868 26928 35868 0 DP_3.matrix\[32\]
rlabel metal2 20928 37422 20928 37422 0 DP_3.matrix\[33\]
rlabel metal2 17568 33642 17568 33642 0 DP_3.matrix\[48\]
rlabel metal2 16848 30072 16848 30072 0 DP_3.matrix\[49\]
rlabel metal2 6144 30618 6144 30618 0 DP_3.matrix\[64\]
rlabel metal2 4800 26166 4800 26166 0 DP_3.matrix\[65\]
rlabel metal2 10368 35448 10368 35448 0 DP_3.matrix\[80\]
rlabel metal2 7200 36120 7200 36120 0 DP_3.matrix\[81\]
rlabel metal2 6192 22512 6192 22512 0 DP_3.matrix\[96\]
rlabel metal2 4752 17052 4752 17052 0 DP_3.matrix\[97\]
rlabel metal2 44976 32340 44976 32340 0 DP_4.matrix\[0\]
rlabel metal2 5280 14196 5280 14196 0 DP_4.matrix\[112\]
rlabel metal2 12288 13734 12288 13734 0 DP_4.matrix\[113\]
rlabel metal2 6336 5250 6336 5250 0 DP_4.matrix\[128\]
rlabel metal2 4752 9660 4752 9660 0 DP_4.matrix\[129\]
rlabel metal2 32736 34902 32736 34902 0 DP_4.matrix\[16\]
rlabel metal2 37536 36204 37536 36204 0 DP_4.matrix\[17\]
rlabel metal2 49296 30072 49296 30072 0 DP_4.matrix\[1\]
rlabel metal2 26016 36750 26016 36750 0 DP_4.matrix\[32\]
rlabel metal2 21408 36666 21408 36666 0 DP_4.matrix\[33\]
rlabel metal2 17904 29316 17904 29316 0 DP_4.matrix\[48\]
rlabel metal2 17760 34398 17760 34398 0 DP_4.matrix\[49\]
rlabel metal2 5232 29316 5232 29316 0 DP_4.matrix\[64\]
rlabel metal2 4896 26376 4896 26376 0 DP_4.matrix\[65\]
rlabel metal2 6336 34902 6336 34902 0 DP_4.matrix\[80\]
rlabel metal3 11088 36876 11088 36876 0 DP_4.matrix\[81\]
rlabel metal2 4752 18732 4752 18732 0 DP_4.matrix\[96\]
rlabel metal2 1248 22806 1248 22806 0 DP_4.matrix\[97\]
rlabel metal3 54432 14196 54432 14196 0 _000_
rlabel metal2 56736 14280 56736 14280 0 _001_
rlabel metal2 46560 8568 46560 8568 0 _002_
rlabel metal2 47520 8820 47520 8820 0 _003_
rlabel metal2 40128 20118 40128 20118 0 _004_
rlabel metal2 40800 20328 40800 20328 0 _005_
rlabel metal2 34176 14658 34176 14658 0 _006_
rlabel metal2 34368 16338 34368 16338 0 _007_
rlabel metal2 48864 11634 48864 11634 0 _008_
rlabel metal2 49632 13650 49632 13650 0 _009_
rlabel metal3 38976 14028 38976 14028 0 _010_
rlabel metal2 40992 15960 40992 15960 0 _011_
rlabel metal2 41232 10080 41232 10080 0 _012_
rlabel metal2 41376 11760 41376 11760 0 _013_
rlabel metal2 33024 10332 33024 10332 0 _014_
rlabel metal2 33984 8190 33984 8190 0 _015_
rlabel metal2 32352 8400 32352 8400 0 _016_
rlabel metal3 38880 29820 38880 29820 0 _017_
rlabel metal2 36192 31374 36192 31374 0 _018_
rlabel metal2 26112 29400 26112 29400 0 _019_
rlabel metal2 26784 30618 26784 30618 0 _020_
rlabel metal2 10848 26166 10848 26166 0 _021_
rlabel metal2 11616 27594 11616 27594 0 _022_
rlabel metal2 12288 21126 12288 21126 0 _023_
rlabel metal2 12480 20370 12480 20370 0 _024_
rlabel metal2 28416 26166 28416 26166 0 _025_
rlabel metal2 27168 28350 27168 28350 0 _026_
rlabel metal2 15936 23730 15936 23730 0 _027_
rlabel metal3 17376 25536 17376 25536 0 _028_
rlabel metal2 20928 21588 20928 21588 0 _029_
rlabel metal2 21984 22932 21984 22932 0 _030_
rlabel metal2 26112 12894 26112 12894 0 _031_
rlabel metal3 21744 9492 21744 9492 0 _032_
rlabel metal3 23826 11760 23826 11760 0 _033_
rlabel metal2 9600 16086 9600 16086 0 _034_
rlabel metal2 8592 14616 8592 14616 0 _035_
rlabel metal2 5376 5250 5376 5250 0 _036_
rlabel metal2 6144 8820 6144 8820 0 _037_
rlabel metal2 8832 33516 8832 33516 0 _038_
rlabel metal2 8880 32256 8880 32256 0 _039_
rlabel metal2 8064 21294 8064 21294 0 _040_
rlabel metal2 5376 19698 5376 19698 0 _041_
rlabel metal2 54960 10416 54960 10416 0 _042_
rlabel metal2 59232 12600 59232 12600 0 _043_
rlabel metal2 44352 30912 44352 30912 0 _044_
rlabel metal3 43680 30744 43680 30744 0 _045_
rlabel metal3 30288 16212 30288 16212 0 _046_
rlabel metal3 30240 19152 30240 19152 0 _047_
rlabel metal3 46032 20748 46032 20748 0 _048_
rlabel metal2 43680 23604 43680 23604 0 _049_
rlabel metal2 36288 21882 36288 21882 0 _050_
rlabel metal3 36288 23184 36288 23184 0 _051_
rlabel metal2 52800 6048 52800 6048 0 _052_
rlabel metal2 49104 4032 49104 4032 0 _053_
rlabel metal2 40992 7602 40992 7602 0 _054_
rlabel metal2 41760 5334 41760 5334 0 _055_
rlabel metal2 52704 17136 52704 17136 0 _056_
rlabel metal2 56640 17346 56640 17346 0 _057_
rlabel metal2 19392 3738 19392 3738 0 _058_
rlabel metal3 20544 2520 20544 2520 0 _059_
rlabel metal2 7104 26796 7104 26796 0 _060_
rlabel metal2 5952 28434 5952 28434 0 _061_
rlabel metal3 20784 14700 20784 14700 0 _062_
rlabel metal3 22032 15624 22032 15624 0 _063_
rlabel metal2 18720 30156 18720 30156 0 _064_
rlabel metal3 19056 30744 19056 30744 0 _065_
rlabel metal2 25584 32844 25584 32844 0 _066_
rlabel metal2 21792 33432 21792 33432 0 _067_
rlabel metal2 34080 33474 34080 33474 0 _068_
rlabel metal3 36816 34356 36816 34356 0 _069_
rlabel metal2 54144 8946 54144 8946 0 _070_
rlabel metal2 59616 9618 59616 9618 0 _071_
rlabel metal2 49344 18270 49344 18270 0 _072_
rlabel metal2 55680 19110 55680 19110 0 _073_
rlabel metal2 38112 2898 38112 2898 0 _074_
rlabel metal3 38016 5040 38016 5040 0 _075_
rlabel metal2 51936 4662 51936 4662 0 _076_
rlabel metal2 52224 2688 52224 2688 0 _077_
rlabel metal3 32880 21672 32880 21672 0 _078_
rlabel metal2 33600 26376 33600 26376 0 _079_
rlabel metal2 44784 19908 44784 19908 0 _080_
rlabel metal2 41472 26502 41472 26502 0 _081_
rlabel metal2 26208 17724 26208 17724 0 _082_
rlabel metal2 26880 21294 26880 21294 0 _083_
rlabel metal2 16896 13482 16896 13482 0 _084_
rlabel metal2 14592 15918 14592 15918 0 _085_
rlabel metal3 16608 2856 16608 2856 0 _086_
rlabel metal2 16704 5922 16704 5922 0 _087_
rlabel metal2 55584 8820 55584 8820 0 _088_
rlabel metal2 59808 10710 59808 10710 0 _089_
rlabel metal2 52128 20370 52128 20370 0 _090_
rlabel metal2 47808 17514 47808 17514 0 _091_
rlabel metal2 37920 6762 37920 6762 0 _092_
rlabel metal2 43104 2898 43104 2898 0 _093_
rlabel metal2 47616 2898 47616 2898 0 _094_
rlabel metal2 47424 2898 47424 2898 0 _095_
rlabel metal2 30240 24066 30240 24066 0 _096_
rlabel metal2 34080 26502 34080 26502 0 _097_
rlabel metal2 45168 24780 45168 24780 0 _098_
rlabel metal2 46464 24024 46464 24024 0 _099_
rlabel metal3 26208 17724 26208 17724 0 _100_
rlabel metal2 26496 21588 26496 21588 0 _101_
rlabel metal2 18816 16128 18816 16128 0 _102_
rlabel metal2 14880 17514 14880 17514 0 _103_
rlabel metal2 11808 3738 11808 3738 0 _104_
rlabel metal3 12816 2100 12816 2100 0 _105_
rlabel metal2 45456 32340 45456 32340 0 _106_
rlabel metal2 44496 28308 44496 28308 0 _107_
rlabel metal2 35232 36708 35232 36708 0 _108_
rlabel metal2 30240 36204 30240 36204 0 _109_
rlabel metal2 24624 35028 24624 35028 0 _110_
rlabel metal2 19296 36708 19296 36708 0 _111_
rlabel metal2 14976 33390 14976 33390 0 _112_
rlabel metal2 14400 30114 14400 30114 0 _113_
rlabel metal2 3936 30366 3936 30366 0 _114_
rlabel metal2 2400 25872 2400 25872 0 _115_
rlabel metal2 9552 35364 9552 35364 0 _116_
rlabel metal2 4704 36204 4704 36204 0 _117_
rlabel metal2 3840 22554 3840 22554 0 _118_
rlabel metal3 2640 17220 2640 17220 0 _119_
rlabel metal2 9360 13440 9360 13440 0 _120_
rlabel metal2 4032 13524 4032 13524 0 _121_
rlabel metal2 3744 8190 3744 8190 0 _122_
rlabel metal2 3744 5250 3744 5250 0 _123_
rlabel metal3 42960 33012 42960 33012 0 _124_
rlabel metal2 46944 30114 46944 30114 0 _125_
rlabel metal2 30336 34650 30336 34650 0 _126_
rlabel metal2 36480 36330 36480 36330 0 _127_
rlabel metal2 23616 35742 23616 35742 0 _128_
rlabel metal2 19872 36414 19872 36414 0 _129_
rlabel metal2 16224 28602 16224 28602 0 _130_
rlabel metal2 15456 33684 15456 33684 0 _131_
rlabel metal2 2784 29442 2784 29442 0 _132_
rlabel metal2 2496 26418 2496 26418 0 _133_
rlabel metal2 3936 34650 3936 34650 0 _134_
rlabel metal2 9360 36792 9360 36792 0 _135_
rlabel metal2 2304 18858 2304 18858 0 _136_
rlabel metal2 3648 22554 3648 22554 0 _137_
rlabel metal3 3408 14112 3408 14112 0 _138_
rlabel metal2 9888 13062 9888 13062 0 _139_
rlabel metal2 4320 4368 4320 4368 0 _140_
rlabel metal2 2304 9954 2304 9954 0 _141_
rlabel metal2 27264 8610 27264 8610 0 _142_
rlabel metal2 29760 9366 29760 9366 0 _143_
rlabel metal2 29664 8736 29664 8736 0 _144_
rlabel metal2 27840 8610 27840 8610 0 _145_
rlabel metal2 31296 10482 31296 10482 0 _146_
rlabel metal2 31968 11634 31968 11634 0 _147_
rlabel metal2 31392 11088 31392 11088 0 _148_
rlabel metal2 31296 12474 31296 12474 0 _149_
rlabel metal2 56064 14784 56064 14784 0 _150_
rlabel metal3 56160 14658 56160 14658 0 _151_
rlabel metal2 43104 12138 43104 12138 0 _152_
rlabel metal2 43200 12894 43200 12894 0 _153_
rlabel metal3 40176 15540 40176 15540 0 _154_
rlabel metal2 40848 15540 40848 15540 0 _155_
rlabel metal2 49440 12894 49440 12894 0 _156_
rlabel metal2 50496 12936 50496 12936 0 _157_
rlabel metal3 33840 15540 33840 15540 0 _158_
rlabel metal2 33792 17094 33792 17094 0 _159_
rlabel metal3 40128 20748 40128 20748 0 _160_
rlabel metal2 41088 22722 41088 22722 0 _161_
rlabel metal3 46944 7980 46944 7980 0 _162_
rlabel metal2 46944 7308 46944 7308 0 _163_
rlabel metal2 38784 31626 38784 31626 0 _164_
rlabel metal2 38880 31794 38880 31794 0 _165_
rlabel metal2 33408 8148 33408 8148 0 _166_
rlabel metal3 33744 8820 33744 8820 0 _167_
rlabel metal2 34464 9114 34464 9114 0 _168_
rlabel metal2 33504 8232 33504 8232 0 _169_
rlabel metal3 21504 24360 21504 24360 0 _170_
rlabel metal2 22080 23856 22080 23856 0 _171_
rlabel metal2 16992 24990 16992 24990 0 _172_
rlabel metal2 16608 25032 16608 25032 0 _173_
rlabel metal2 28848 27048 28848 27048 0 _174_
rlabel metal2 30576 29148 30576 29148 0 _175_
rlabel metal2 12192 20244 12192 20244 0 _176_
rlabel metal2 11328 18732 11328 18732 0 _177_
rlabel metal2 11136 27342 11136 27342 0 _178_
rlabel metal3 11472 29148 11472 29148 0 _179_
rlabel metal3 25536 30660 25536 30660 0 _180_
rlabel metal3 25056 31164 25056 31164 0 _181_
rlabel metal2 23424 11046 23424 11046 0 _182_
rlabel metal2 23520 13272 23520 13272 0 _183_
rlabel metal2 23616 12432 23616 12432 0 _184_
rlabel metal2 23280 11676 23280 11676 0 _185_
rlabel metal3 7632 14112 7632 14112 0 _186_
rlabel metal3 8832 14112 8832 14112 0 _187_
rlabel metal3 5136 6636 5136 6636 0 _188_
rlabel metal3 5232 7980 5232 7980 0 _189_
rlabel metal2 8448 34818 8448 34818 0 _190_
rlabel metal2 8736 35070 8736 35070 0 _191_
rlabel metal2 4896 20034 4896 20034 0 _192_
rlabel metal2 5184 20118 5184 20118 0 _193_
rlabel metal2 58656 10416 58656 10416 0 _194_
rlabel metal2 58992 10416 58992 10416 0 _195_
rlabel metal2 44976 30072 44976 30072 0 _196_
rlabel metal3 45984 30660 45984 30660 0 _197_
rlabel metal3 28464 19236 28464 19236 0 _198_
rlabel metal3 28698 20160 28698 20160 0 _199_
rlabel metal2 43488 24066 43488 24066 0 _200_
rlabel metal3 44736 23772 44736 23772 0 _201_
rlabel metal2 35232 24066 35232 24066 0 _202_
rlabel metal3 35232 23772 35232 23772 0 _203_
rlabel metal2 50496 3822 50496 3822 0 _204_
rlabel metal2 49248 3822 49248 3822 0 _205_
rlabel metal2 41088 5250 41088 5250 0 _206_
rlabel metal2 41280 4368 41280 4368 0 _207_
rlabel metal2 55248 17724 55248 17724 0 _208_
rlabel metal2 55488 17682 55488 17682 0 _209_
rlabel metal2 18720 2730 18720 2730 0 _210_
rlabel metal2 19008 2688 19008 2688 0 _211_
rlabel metal2 5472 27678 5472 27678 0 _212_
rlabel metal2 4704 27762 4704 27762 0 _213_
rlabel metal2 18240 15456 18240 15456 0 _214_
rlabel metal3 18048 15372 18048 15372 0 _215_
rlabel metal2 17472 30576 17472 30576 0 _216_
rlabel metal2 17760 31290 17760 31290 0 _217_
rlabel metal2 21696 35112 21696 35112 0 _218_
rlabel metal2 22080 35322 22080 35322 0 _219_
rlabel metal3 34512 35196 34512 35196 0 _220_
rlabel metal2 36192 35490 36192 35490 0 _221_
rlabel via2 78 36708 78 36708 0 clk
rlabel metal2 21696 11760 21696 11760 0 clknet_0_clk
rlabel metal3 9408 7980 9408 7980 0 clknet_4_0_0_clk
rlabel metal2 53280 8190 53280 8190 0 clknet_4_10_0_clk
rlabel metal2 53856 13314 53856 13314 0 clknet_4_11_0_clk
rlabel metal2 35088 22260 35088 22260 0 clknet_4_12_0_clk
rlabel metal3 35376 30660 35376 30660 0 clknet_4_13_0_clk
rlabel metal3 45024 21588 45024 21588 0 clknet_4_14_0_clk
rlabel metal2 43968 27006 43968 27006 0 clknet_4_15_0_clk
rlabel metal2 9024 13104 9024 13104 0 clknet_4_1_0_clk
rlabel metal2 20688 11004 20688 11004 0 clknet_4_2_0_clk
rlabel metal3 19584 15960 19584 15960 0 clknet_4_3_0_clk
rlabel metal2 9504 26922 9504 26922 0 clknet_4_4_0_clk
rlabel metal3 10416 33684 10416 33684 0 clknet_4_5_0_clk
rlabel metal3 21408 28308 21408 28308 0 clknet_4_6_0_clk
rlabel metal2 22368 32760 22368 32760 0 clknet_4_7_0_clk
rlabel metal2 38016 8022 38016 8022 0 clknet_4_8_0_clk
rlabel metal2 38208 11340 38208 11340 0 clknet_4_9_0_clk
rlabel metal3 3840 4956 3840 4956 0 clknet_5_0__leaf_clk
rlabel metal2 5184 35112 5184 35112 0 clknet_5_10__leaf_clk
rlabel metal3 15648 32802 15648 32802 0 clknet_5_11__leaf_clk
rlabel metal2 19200 23856 19200 23856 0 clknet_5_12__leaf_clk
rlabel metal3 22512 20076 22512 20076 0 clknet_5_13__leaf_clk
rlabel metal2 19776 37380 19776 37380 0 clknet_5_14__leaf_clk
rlabel metal3 27744 32844 27744 32844 0 clknet_5_15__leaf_clk
rlabel metal2 32352 4536 32352 4536 0 clknet_5_16__leaf_clk
rlabel metal2 40224 3654 40224 3654 0 clknet_5_17__leaf_clk
rlabel metal2 37104 11004 37104 11004 0 clknet_5_18__leaf_clk
rlabel metal2 41184 12810 41184 12810 0 clknet_5_19__leaf_clk
rlabel metal2 11040 6510 11040 6510 0 clknet_5_1__leaf_clk
rlabel metal2 51552 7308 51552 7308 0 clknet_5_20__leaf_clk
rlabel metal3 54288 4956 54288 4956 0 clknet_5_21__leaf_clk
rlabel metal3 54432 14280 54432 14280 0 clknet_5_22__leaf_clk
rlabel metal2 56640 12852 56640 12852 0 clknet_5_23__leaf_clk
rlabel metal2 26976 19656 26976 19656 0 clknet_5_24__leaf_clk
rlabel metal3 34608 19488 34608 19488 0 clknet_5_25__leaf_clk
rlabel metal3 34896 30828 34896 30828 0 clknet_5_26__leaf_clk
rlabel metal3 37152 36708 37152 36708 0 clknet_5_27__leaf_clk
rlabel metal2 38112 22344 38112 22344 0 clknet_5_28__leaf_clk
rlabel metal3 55152 20076 55152 20076 0 clknet_5_29__leaf_clk
rlabel metal3 3840 17724 3840 17724 0 clknet_5_2__leaf_clk
rlabel metal2 39648 27216 39648 27216 0 clknet_5_30__leaf_clk
rlabel metal2 46656 32802 46656 32802 0 clknet_5_31__leaf_clk
rlabel metal2 9888 17766 9888 17766 0 clknet_5_3__leaf_clk
rlabel metal3 21408 3444 21408 3444 0 clknet_5_4__leaf_clk
rlabel metal3 24672 4116 24672 4116 0 clknet_5_5__leaf_clk
rlabel metal2 15888 16212 15888 16212 0 clknet_5_6__leaf_clk
rlabel metal2 21264 17136 21264 17136 0 clknet_5_7__leaf_clk
rlabel metal3 3744 22260 3744 22260 0 clknet_5_8__leaf_clk
rlabel metal2 9312 22764 9312 22764 0 clknet_5_9__leaf_clk
rlabel metal2 55680 14070 55680 14070 0 mac1.products_ff\[0\]
rlabel metal2 33648 15708 33648 15708 0 mac1.products_ff\[112\]
rlabel metal2 27744 16380 27744 16380 0 mac1.products_ff\[113\]
rlabel metal2 21792 3864 21792 3864 0 mac1.products_ff\[128\]
rlabel metal2 23808 2646 23808 2646 0 mac1.products_ff\[129\]
rlabel metal2 56064 16506 56064 16506 0 mac1.products_ff\[16\]
rlabel metal2 59040 15750 59040 15750 0 mac1.products_ff\[17\]
rlabel metal3 60624 14196 60624 14196 0 mac1.products_ff\[1\]
rlabel metal2 45696 8694 45696 8694 0 mac1.products_ff\[32\]
rlabel metal2 44640 6048 44640 6048 0 mac1.products_ff\[33\]
rlabel metal3 49824 7392 49824 7392 0 mac1.products_ff\[48\]
rlabel metal3 46560 6468 46560 6468 0 mac1.products_ff\[49\]
rlabel metal2 38976 21546 38976 21546 0 mac1.products_ff\[64\]
rlabel metal2 39264 23520 39264 23520 0 mac1.products_ff\[65\]
rlabel metal2 39936 20706 39936 20706 0 mac1.products_ff\[80\]
rlabel metal2 40848 23100 40848 23100 0 mac1.products_ff\[81\]
rlabel metal2 33888 15792 33888 15792 0 mac1.products_ff\[96\]
rlabel metal2 34080 18732 34080 18732 0 mac1.products_ff\[97\]
rlabel metal2 48528 13188 48528 13188 0 mac1.sum_lvl1_ff\[0\]
rlabel metal3 37488 17724 37488 17724 0 mac1.sum_lvl1_ff\[16\]
rlabel metal2 40704 17682 40704 17682 0 mac1.sum_lvl1_ff\[17\]
rlabel metal3 52128 12516 52128 12516 0 mac1.sum_lvl1_ff\[1\]
rlabel metal2 38688 15330 38688 15330 0 mac1.sum_lvl1_ff\[24\]
rlabel metal2 40416 17010 40416 17010 0 mac1.sum_lvl1_ff\[25\]
rlabel metal3 26544 4368 26544 4368 0 mac1.sum_lvl1_ff\[32\]
rlabel metal2 27360 2646 27360 2646 0 mac1.sum_lvl1_ff\[33\]
rlabel metal2 49296 11676 49296 11676 0 mac1.sum_lvl1_ff\[8\]
rlabel metal2 50496 10248 50496 10248 0 mac1.sum_lvl1_ff\[9\]
rlabel metal2 41904 11172 41904 11172 0 mac1.sum_lvl2_ff\[0\]
rlabel metal2 43776 13986 43776 13986 0 mac1.sum_lvl2_ff\[1\]
rlabel metal2 41664 12642 41664 12642 0 mac1.sum_lvl2_ff\[4\]
rlabel metal2 44160 15204 44160 15204 0 mac1.sum_lvl2_ff\[5\]
rlabel metal2 30192 4872 30192 4872 0 mac1.sum_lvl2_ff\[8\]
rlabel metal2 30624 3486 30624 3486 0 mac1.sum_lvl2_ff\[9\]
rlabel metal2 36384 9408 36384 9408 0 mac1.sum_lvl3_ff\[0\]
rlabel metal3 35232 8652 35232 8652 0 mac1.sum_lvl3_ff\[1\]
rlabel metal3 33744 5880 33744 5880 0 mac1.sum_lvl3_ff\[2\]
rlabel metal2 33696 3444 33696 3444 0 mac1.sum_lvl3_ff\[3\]
rlabel metal2 25824 7686 25824 7686 0 mac1.total_sum\[0\]
rlabel metal2 28320 8400 28320 8400 0 mac1.total_sum\[1\]
rlabel metal3 31008 11928 31008 11928 0 mac1.total_sum\[2\]
rlabel metal3 36816 30828 36816 30828 0 mac2.products_ff\[0\]
rlabel metal2 12000 17430 12000 17430 0 mac2.products_ff\[112\]
rlabel metal2 11040 18270 11040 18270 0 mac2.products_ff\[113\]
rlabel metal2 9408 5586 9408 5586 0 mac2.products_ff\[128\]
rlabel metal3 9552 9660 9552 9660 0 mac2.products_ff\[129\]
rlabel metal2 37632 32130 37632 32130 0 mac2.products_ff\[16\]
rlabel metal3 40080 32172 40080 32172 0 mac2.products_ff\[17\]
rlabel metal2 39744 30828 39744 30828 0 mac2.products_ff\[1\]
rlabel metal2 27648 32004 27648 32004 0 mac2.products_ff\[32\]
rlabel metal2 24192 32004 24192 32004 0 mac2.products_ff\[33\]
rlabel metal2 24288 30366 24288 30366 0 mac2.products_ff\[48\]
rlabel metal3 23232 30828 23232 30828 0 mac2.products_ff\[49\]
rlabel metal2 9552 26292 9552 26292 0 mac2.products_ff\[64\]
rlabel metal2 10272 29568 10272 29568 0 mac2.products_ff\[65\]
rlabel metal2 11280 26796 11280 26796 0 mac2.products_ff\[80\]
rlabel metal2 11808 31626 11808 31626 0 mac2.products_ff\[81\]
rlabel metal3 11424 21588 11424 21588 0 mac2.products_ff\[96\]
rlabel metal2 10752 18816 10752 18816 0 mac2.products_ff\[97\]
rlabel metal2 38496 27048 38496 27048 0 mac2.sum_lvl1_ff\[0\]
rlabel metal2 13824 24864 13824 24864 0 mac2.sum_lvl1_ff\[16\]
rlabel metal3 16416 24654 16416 24654 0 mac2.sum_lvl1_ff\[17\]
rlabel metal2 30432 31080 30432 31080 0 mac2.sum_lvl1_ff\[1\]
rlabel metal2 16224 23142 16224 23142 0 mac2.sum_lvl1_ff\[24\]
rlabel metal2 16080 21000 16080 21000 0 mac2.sum_lvl1_ff\[25\]
rlabel metal2 13056 5670 13056 5670 0 mac2.sum_lvl1_ff\[32\]
rlabel metal2 12816 9660 12816 9660 0 mac2.sum_lvl1_ff\[33\]
rlabel metal2 28800 27594 28800 27594 0 mac2.sum_lvl1_ff\[8\]
rlabel metal2 30048 29862 30048 29862 0 mac2.sum_lvl1_ff\[9\]
rlabel metal3 23778 24612 23778 24612 0 mac2.sum_lvl2_ff\[0\]
rlabel metal2 22080 25578 22080 25578 0 mac2.sum_lvl2_ff\[1\]
rlabel metal2 20832 23814 20832 23814 0 mac2.sum_lvl2_ff\[4\]
rlabel metal3 21456 25284 21456 25284 0 mac2.sum_lvl2_ff\[5\]
rlabel metal2 14784 7686 14784 7686 0 mac2.sum_lvl2_ff\[8\]
rlabel metal2 15408 10416 15408 10416 0 mac2.sum_lvl2_ff\[9\]
rlabel metal3 22704 15540 22704 15540 0 mac2.sum_lvl3_ff\[0\]
rlabel metal2 23424 18438 23424 18438 0 mac2.sum_lvl3_ff\[1\]
rlabel metal2 20352 9156 20352 9156 0 mac2.sum_lvl3_ff\[2\]
rlabel metal2 23040 12474 23040 12474 0 mac2.sum_lvl3_ff\[3\]
rlabel metal2 25440 7938 25440 7938 0 mac2.total_sum\[0\]
rlabel metal3 27456 10164 27456 10164 0 mac2.total_sum\[1\]
rlabel metal2 30720 12474 30720 12474 0 mac2.total_sum\[2\]
rlabel metal2 25344 5376 25344 5376 0 net1
rlabel metal3 366 13188 366 13188 0 net10
rlabel metal2 46656 3402 46656 3402 0 net100
rlabel metal2 33408 26334 33408 26334 0 net101
rlabel metal2 39552 15498 39552 15498 0 net102
rlabel metal2 38496 13482 38496 13482 0 net103
rlabel metal2 18528 6258 18528 6258 0 net104
rlabel metal2 15840 23856 15840 23856 0 net105
rlabel metal2 17856 23688 17856 23688 0 net106
rlabel metal3 21264 10164 21264 10164 0 net107
rlabel metal2 21984 8652 21984 8652 0 net108
rlabel metal2 46752 8022 46752 8022 0 net109
rlabel metal3 366 14028 366 14028 0 net11
rlabel metal2 47040 9870 47040 9870 0 net110
rlabel metal2 10560 26628 10560 26628 0 net111
rlabel metal2 11472 25284 11472 25284 0 net112
rlabel metal2 12192 20622 12192 20622 0 net113
rlabel metal2 13680 21756 13680 21756 0 net114
rlabel metal2 41472 11214 41472 11214 0 net115
rlabel metal2 39552 10164 39552 10164 0 net116
rlabel metal2 25344 30702 25344 30702 0 net117
rlabel metal3 26496 27720 26496 27720 0 net118
rlabel via2 17568 3945 17568 3945 0 net119
rlabel metal3 366 14868 366 14868 0 net12
rlabel metal3 19008 16296 19008 16296 0 net120
rlabel metal2 29184 26754 29184 26754 0 net121
rlabel metal2 27168 25284 27168 25284 0 net122
rlabel metal3 39312 7224 39312 7224 0 net123
rlabel metal2 4704 5544 4704 5544 0 net124
rlabel metal3 9792 14700 9792 14700 0 net125
rlabel metal2 55392 14364 55392 14364 0 net126
rlabel metal3 51792 14112 51792 14112 0 net127
rlabel metal2 51360 17808 51360 17808 0 net128
rlabel metal2 49344 12768 49344 12768 0 net129
rlabel metal3 366 5628 366 5628 0 net13
rlabel metal3 45504 11088 45504 11088 0 net130
rlabel metal3 35088 22092 35088 22092 0 net131
rlabel metal2 50399 3664 50399 3664 0 net132
rlabel metal2 33312 35154 33312 35154 0 net133
rlabel metal3 4176 29904 4176 29904 0 net134
rlabel metal2 53568 18984 53568 18984 0 net135
rlabel metal3 4224 19320 4224 19320 0 net136
rlabel metal2 4704 21546 4704 21546 0 net137
rlabel metal3 8688 35112 8688 35112 0 net138
rlabel metal2 23232 35910 23232 35910 0 net139
rlabel metal3 366 6468 366 6468 0 net14
rlabel metal2 27648 18018 27648 18018 0 net140
rlabel metal2 4128 29946 4128 29946 0 net141
rlabel metal3 4992 5628 4992 5628 0 net142
rlabel metal3 43968 32928 43968 32928 0 net143
rlabel metal2 5088 35154 5088 35154 0 net144
rlabel metal2 17280 30156 17280 30156 0 net145
rlabel metal3 46272 33432 46272 33432 0 net146
rlabel metal3 38160 32172 38160 32172 0 net147
rlabel metal2 40896 27678 40896 27678 0 net148
rlabel metal2 18192 33432 18192 33432 0 net149
rlabel metal3 366 7308 366 7308 0 net15
rlabel metal3 14976 4200 14976 4200 0 net150
rlabel metal3 28752 17976 28752 17976 0 net151
rlabel metal2 20928 24654 20928 24654 0 net152
rlabel metal2 19968 20286 19968 20286 0 net153
rlabel metal3 57360 10332 57360 10332 0 net154
rlabel metal2 4032 14658 4032 14658 0 net155
rlabel metal3 56640 8820 56640 8820 0 net156
rlabel metal2 34080 24570 34080 24570 0 net157
rlabel metal2 45024 23100 45024 23100 0 net158
rlabel metal3 19344 15372 19344 15372 0 net159
rlabel metal3 318 8148 318 8148 0 net16
rlabel metal3 40896 4116 40896 4116 0 net160
rlabel metal2 36096 36036 36096 36036 0 net161
rlabel metal2 45024 22092 45024 22092 0 net162
rlabel metal2 24864 35196 24864 35196 0 net163
rlabel metal2 52128 4830 52128 4830 0 net164
rlabel metal3 34896 7980 34896 7980 0 net165
rlabel metal2 28512 7770 28512 7770 0 net166
rlabel metal2 34224 8652 34224 8652 0 net167
rlabel metal2 33120 9618 33120 9618 0 net168
rlabel metal2 33120 11382 33120 11382 0 net169
rlabel metal3 318 15708 318 15708 0 net17
rlabel metal2 23280 13188 23280 13188 0 net170
rlabel metal2 23712 12768 23712 12768 0 net171
rlabel metal3 27552 12600 27552 12600 0 net172
rlabel metal2 39744 15624 39744 15624 0 net173
rlabel metal2 41760 15834 41760 15834 0 net174
rlabel metal2 10944 30492 10944 30492 0 net175
rlabel metal2 11232 28266 11232 28266 0 net176
rlabel metal3 12000 26208 12000 26208 0 net177
rlabel metal3 55584 14742 55584 14742 0 net178
rlabel metal2 56064 13482 56064 13482 0 net179
rlabel metal3 366 16548 366 16548 0 net18
rlabel metal2 11664 20748 11664 20748 0 net180
rlabel metal2 13536 20664 13536 20664 0 net181
rlabel metal2 46560 8232 46560 8232 0 net182
rlabel metal2 48000 9492 48000 9492 0 net183
rlabel metal2 25056 30660 25056 30660 0 net184
rlabel metal2 27408 29820 27408 29820 0 net185
rlabel metal2 16896 24318 16896 24318 0 net186
rlabel metal2 18624 26124 18624 26124 0 net187
rlabel metal2 40560 23100 40560 23100 0 net188
rlabel metal2 40512 21420 40512 21420 0 net189
rlabel metal3 366 17388 366 17388 0 net19
rlabel metal2 41472 19236 41472 19236 0 net190
rlabel metal2 49536 12222 49536 12222 0 net191
rlabel metal2 46992 14028 46992 14028 0 net192
rlabel metal2 33120 17682 33120 17682 0 net193
rlabel metal2 34176 16506 34176 16506 0 net194
rlabel metal2 36192 17052 36192 17052 0 net195
rlabel metal2 21504 24276 21504 24276 0 net196
rlabel metal2 21072 20076 21072 20076 0 net197
rlabel metal2 30480 29820 30480 29820 0 net198
rlabel metal2 29184 28602 29184 28602 0 net199
rlabel metal2 26976 5922 26976 5922 0 net2
rlabel metal3 366 18228 366 18228 0 net20
rlabel metal2 24000 27174 24000 27174 0 net200
rlabel metal2 37440 32424 37440 32424 0 net201
rlabel metal3 34176 30744 34176 30744 0 net202
rlabel metal2 42816 12768 42816 12768 0 net203
rlabel metal2 38304 11046 38304 11046 0 net204
rlabel metal2 33360 6636 33360 6636 0 net205
rlabel metal3 30864 8064 30864 8064 0 net206
rlabel metal2 22272 15204 22272 15204 0 net207
rlabel metal2 24480 11298 24480 11298 0 net208
rlabel metal3 366 19068 366 19068 0 net21
rlabel metal3 366 19908 366 19908 0 net22
rlabel metal3 366 20748 366 20748 0 net23
rlabel metal3 366 21588 366 21588 0 net24
rlabel metal2 12960 10458 12960 10458 0 net25
rlabel metal2 28128 2520 28128 2520 0 net26
rlabel metal2 24576 2520 24576 2520 0 net27
rlabel metal2 9792 5922 9792 5922 0 net28
rlabel metal2 31104 3696 31104 3696 0 net29
rlabel metal3 3582 4200 3582 4200 0 net3
rlabel metal2 12384 6468 12384 6468 0 net30
rlabel metal2 31008 5544 31008 5544 0 net31
rlabel metal2 10368 9786 10368 9786 0 net32
rlabel metal2 16224 11004 16224 11004 0 net33
rlabel metal2 27648 4956 27648 4956 0 net34
rlabel metal2 23712 4032 23712 4032 0 net35
rlabel metal2 16512 8358 16512 8358 0 net36
rlabel metal2 33696 15498 33696 15498 0 net37
rlabel metal2 35328 14616 35328 14616 0 net38
rlabel via2 36671 35952 36671 35952 0 net39
rlabel metal2 864 7770 864 7770 0 net4
rlabel metal3 56064 19320 56064 19320 0 net40
rlabel metal3 10704 14028 10704 14028 0 net41
rlabel metal3 16656 30660 16656 30660 0 net42
rlabel metal2 7104 13986 7104 13986 0 net43
rlabel metal3 4848 27636 4848 27636 0 net44
rlabel metal2 44832 29568 44832 29568 0 net45
rlabel metal3 58656 10122 58656 10122 0 net46
rlabel metal2 17856 15498 17856 15498 0 net47
rlabel metal2 28128 20328 28128 20328 0 net48
rlabel metal2 49056 17766 49056 17766 0 net49
rlabel metal3 366 8988 366 8988 0 net5
rlabel metal2 9504 36666 9504 36666 0 net50
rlabel metal3 48048 30576 48048 30576 0 net51
rlabel metal3 6078 36624 6078 36624 0 net52
rlabel metal2 41664 3864 41664 3864 0 net53
rlabel metal2 22176 35910 22176 35910 0 net54
rlabel metal3 60576 10248 60576 10248 0 net55
rlabel metal2 23424 7518 23424 7518 0 net56
rlabel metal2 4320 4914 4320 4914 0 net57
rlabel metal2 10752 9786 10752 9786 0 net58
rlabel metal2 12768 10206 12768 10206 0 net59
rlabel metal3 366 9828 366 9828 0 net6
rlabel metal2 21408 20034 21408 20034 0 net60
rlabel metal3 21504 2604 21504 2604 0 net61
rlabel metal3 20640 19824 20640 19824 0 net62
rlabel metal2 3264 22302 3264 22302 0 net63
rlabel metal3 3120 19236 3120 19236 0 net64
rlabel metal2 5088 35616 5088 35616 0 net65
rlabel metal2 15072 34020 15072 34020 0 net66
rlabel metal3 18720 23772 18720 23772 0 net67
rlabel metal2 20064 21504 20064 21504 0 net68
rlabel metal2 38496 2646 38496 2646 0 net69
rlabel metal3 366 10668 366 10668 0 net7
rlabel metal2 39072 18144 39072 18144 0 net70
rlabel metal2 52320 3780 52320 3780 0 net71
rlabel metal2 54528 9072 54528 9072 0 net72
rlabel metal3 56544 19236 56544 19236 0 net73
rlabel metal3 52896 11004 52896 11004 0 net74
rlabel metal2 31488 17724 31488 17724 0 net75
rlabel metal2 19200 36624 19200 36624 0 net76
rlabel metal2 30624 24528 30624 24528 0 net77
rlabel metal2 40512 27132 40512 27132 0 net78
rlabel metal2 36960 37044 36960 37044 0 net79
rlabel metal3 366 11508 366 11508 0 net8
rlabel metal2 39936 29694 39936 29694 0 net80
rlabel metal2 21984 20664 21984 20664 0 net81
rlabel metal2 33120 35868 33120 35868 0 net82
rlabel metal2 4128 9030 4128 9030 0 net83
rlabel metal3 46944 23856 46944 23856 0 net84
rlabel metal2 4032 18648 4032 18648 0 net85
rlabel metal3 52608 2688 52608 2688 0 net86
rlabel metal2 2976 5670 2976 5670 0 net87
rlabel metal3 17184 17640 17184 17640 0 net88
rlabel metal2 43392 25620 43392 25620 0 net89
rlabel metal3 366 12348 366 12348 0 net9
rlabel metal3 16368 32928 16368 32928 0 net90
rlabel metal2 34464 24822 34464 24822 0 net91
rlabel metal2 37440 5670 37440 5670 0 net92
rlabel metal2 4224 27342 4224 27342 0 net93
rlabel metal2 2976 22932 2976 22932 0 net94
rlabel metal2 26688 21294 26688 21294 0 net95
rlabel metal2 13584 1848 13584 1848 0 net96
rlabel metal2 39696 20748 39696 20748 0 net97
rlabel metal2 39456 19236 39456 19236 0 net98
rlabel metal2 19488 35910 19488 35910 0 net99
rlabel metal2 20784 20748 20784 20748 0 rst_n
rlabel metal3 366 2268 366 2268 0 uo_out[0]
rlabel metal3 366 3108 366 3108 0 uo_out[1]
rlabel metal3 366 3948 366 3948 0 uo_out[2]
rlabel metal3 366 4788 366 4788 0 uo_out[3]
<< properties >>
string FIXED_BBOX 0 0 100000 40000
<< end >>
