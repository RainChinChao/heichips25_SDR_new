module heichips25_template (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \DP_1.matrix[0] ;
 wire \DP_1.matrix[10] ;
 wire \DP_1.matrix[18] ;
 wire \DP_1.matrix[19] ;
 wire \DP_1.matrix[1] ;
 wire \DP_1.matrix[27] ;
 wire \DP_1.matrix[28] ;
 wire \DP_1.matrix[36] ;
 wire \DP_1.matrix[37] ;
 wire \DP_1.matrix[45] ;
 wire \DP_1.matrix[46] ;
 wire \DP_1.matrix[54] ;
 wire \DP_1.matrix[55] ;
 wire \DP_1.matrix[63] ;
 wire \DP_1.matrix[64] ;
 wire \DP_1.matrix[72] ;
 wire \DP_1.matrix[73] ;
 wire \DP_1.matrix[9] ;
 wire \DP_2.matrix[0] ;
 wire \DP_2.matrix[10] ;
 wire \DP_2.matrix[18] ;
 wire \DP_2.matrix[19] ;
 wire \DP_2.matrix[1] ;
 wire \DP_2.matrix[27] ;
 wire \DP_2.matrix[28] ;
 wire \DP_2.matrix[36] ;
 wire \DP_2.matrix[37] ;
 wire \DP_2.matrix[45] ;
 wire \DP_2.matrix[46] ;
 wire \DP_2.matrix[54] ;
 wire \DP_2.matrix[55] ;
 wire \DP_2.matrix[63] ;
 wire \DP_2.matrix[64] ;
 wire \DP_2.matrix[72] ;
 wire \DP_2.matrix[73] ;
 wire \DP_2.matrix[9] ;
 wire \DP_3.matrix[0] ;
 wire \DP_3.matrix[10] ;
 wire \DP_3.matrix[18] ;
 wire \DP_3.matrix[19] ;
 wire \DP_3.matrix[1] ;
 wire \DP_3.matrix[27] ;
 wire \DP_3.matrix[28] ;
 wire \DP_3.matrix[36] ;
 wire \DP_3.matrix[37] ;
 wire \DP_3.matrix[45] ;
 wire \DP_3.matrix[46] ;
 wire \DP_3.matrix[54] ;
 wire \DP_3.matrix[55] ;
 wire \DP_3.matrix[63] ;
 wire \DP_3.matrix[64] ;
 wire \DP_3.matrix[72] ;
 wire \DP_3.matrix[73] ;
 wire \DP_3.matrix[9] ;
 wire \DP_4.matrix[0] ;
 wire \DP_4.matrix[10] ;
 wire \DP_4.matrix[18] ;
 wire \DP_4.matrix[19] ;
 wire \DP_4.matrix[1] ;
 wire \DP_4.matrix[27] ;
 wire \DP_4.matrix[28] ;
 wire \DP_4.matrix[36] ;
 wire \DP_4.matrix[37] ;
 wire \DP_4.matrix[45] ;
 wire \DP_4.matrix[46] ;
 wire \DP_4.matrix[54] ;
 wire \DP_4.matrix[55] ;
 wire \DP_4.matrix[63] ;
 wire \DP_4.matrix[64] ;
 wire \DP_4.matrix[72] ;
 wire \DP_4.matrix[73] ;
 wire \DP_4.matrix[9] ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire \mac1.products_ff[0] ;
 wire \mac1.products_ff[102] ;
 wire \mac1.products_ff[103] ;
 wire \mac1.products_ff[119] ;
 wire \mac1.products_ff[120] ;
 wire \mac1.products_ff[136] ;
 wire \mac1.products_ff[137] ;
 wire \mac1.products_ff[17] ;
 wire \mac1.products_ff[18] ;
 wire \mac1.products_ff[1] ;
 wire \mac1.products_ff[34] ;
 wire \mac1.products_ff[35] ;
 wire \mac1.products_ff[51] ;
 wire \mac1.products_ff[52] ;
 wire \mac1.products_ff[68] ;
 wire \mac1.products_ff[69] ;
 wire \mac1.products_ff[85] ;
 wire \mac1.products_ff[86] ;
 wire \mac1.sum_lvl1_ff[0] ;
 wire \mac1.sum_lvl1_ff[16] ;
 wire \mac1.sum_lvl1_ff[17] ;
 wire \mac1.sum_lvl1_ff[1] ;
 wire \mac1.sum_lvl1_ff[24] ;
 wire \mac1.sum_lvl1_ff[25] ;
 wire \mac1.sum_lvl1_ff[32] ;
 wire \mac1.sum_lvl1_ff[33] ;
 wire \mac1.sum_lvl1_ff[8] ;
 wire \mac1.sum_lvl1_ff[9] ;
 wire \mac1.sum_lvl2_ff[0] ;
 wire \mac1.sum_lvl2_ff[1] ;
 wire \mac1.sum_lvl2_ff[4] ;
 wire \mac1.sum_lvl2_ff[5] ;
 wire \mac1.sum_lvl2_ff[8] ;
 wire \mac1.sum_lvl2_ff[9] ;
 wire \mac1.sum_lvl3_ff[0] ;
 wire \mac1.sum_lvl3_ff[1] ;
 wire \mac1.sum_lvl3_ff[2] ;
 wire \mac1.sum_lvl3_ff[3] ;
 wire \mac1.total_sum[0] ;
 wire \mac1.total_sum[1] ;
 wire \mac1.total_sum[2] ;
 wire \mac2.products_ff[0] ;
 wire \mac2.products_ff[102] ;
 wire \mac2.products_ff[103] ;
 wire \mac2.products_ff[119] ;
 wire \mac2.products_ff[120] ;
 wire \mac2.products_ff[136] ;
 wire \mac2.products_ff[137] ;
 wire \mac2.products_ff[17] ;
 wire \mac2.products_ff[18] ;
 wire \mac2.products_ff[1] ;
 wire \mac2.products_ff[34] ;
 wire \mac2.products_ff[35] ;
 wire \mac2.products_ff[51] ;
 wire \mac2.products_ff[52] ;
 wire \mac2.products_ff[68] ;
 wire \mac2.products_ff[69] ;
 wire \mac2.products_ff[85] ;
 wire \mac2.products_ff[86] ;
 wire \mac2.sum_lvl1_ff[0] ;
 wire \mac2.sum_lvl1_ff[16] ;
 wire \mac2.sum_lvl1_ff[17] ;
 wire \mac2.sum_lvl1_ff[1] ;
 wire \mac2.sum_lvl1_ff[24] ;
 wire \mac2.sum_lvl1_ff[25] ;
 wire \mac2.sum_lvl1_ff[32] ;
 wire \mac2.sum_lvl1_ff[33] ;
 wire \mac2.sum_lvl1_ff[8] ;
 wire \mac2.sum_lvl1_ff[9] ;
 wire \mac2.sum_lvl2_ff[0] ;
 wire \mac2.sum_lvl2_ff[1] ;
 wire \mac2.sum_lvl2_ff[4] ;
 wire \mac2.sum_lvl2_ff[5] ;
 wire \mac2.sum_lvl2_ff[8] ;
 wire \mac2.sum_lvl2_ff[9] ;
 wire \mac2.sum_lvl3_ff[0] ;
 wire \mac2.sum_lvl3_ff[1] ;
 wire \mac2.sum_lvl3_ff[2] ;
 wire \mac2.sum_lvl3_ff[3] ;
 wire \mac2.total_sum[0] ;
 wire \mac2.total_sum[1] ;
 wire \mac2.total_sum[2] ;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire clknet_0_clk;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net5;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;

 sg13g2_and2_1 _222_ (.A(net148),
    .B(net130),
    .X(_066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _223_ (.A(net118),
    .B(net133),
    .X(_068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _224_ (.Y(_142_),
    .A(net203),
    .B(net165),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _225_ (.B(net165),
    .A(\mac1.sum_lvl3_ff[0] ),
    .X(_017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _226_ (.A(net141),
    .B(net121),
    .X(_034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _227_ (.A(net156),
    .B(net131),
    .X(_036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _228_ (.A(net127),
    .B(net140),
    .X(_038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _229_ (.Y(_143_),
    .A(net167),
    .B(\mac1.sum_lvl3_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _230_ (.A(net167),
    .B(\mac1.sum_lvl3_ff[3] ),
    .Y(_144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _231_ (.B(\mac1.sum_lvl3_ff[3] ),
    .A(net167),
    .X(_145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _232_ (.Y(_018_),
    .A(_142_),
    .B(_145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _233_ (.A(net157),
    .B(net152),
    .X(_040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _234_ (.A(net159),
    .B(net142),
    .X(_042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _235_ (.A(net128),
    .B(net147),
    .X(_044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _236_ (.A(net129),
    .B(net134),
    .X(_046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _237_ (.A(net160),
    .B(net117),
    .X(_048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _238_ (.A(net122),
    .B(net139),
    .X(_050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _239_ (.A(net150),
    .B(net138),
    .X(_052_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _240_ (.A(net120),
    .B(net151),
    .X(_054_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _241_ (.A(net135),
    .B(net126),
    .X(_056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _242_ (.A(net149),
    .B(net155),
    .X(_058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _243_ (.A(net125),
    .B(net158),
    .X(_060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _244_ (.A(net144),
    .B(net143),
    .X(_062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _245_ (.A(net132),
    .B(net119),
    .X(_064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _246_ (.Y(_146_),
    .A(net197),
    .B(net153),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _247_ (.B(net153),
    .A(\mac1.sum_lvl2_ff[0] ),
    .X(_014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _248_ (.B(\mac1.sum_lvl2_ff[5] ),
    .A(\mac1.sum_lvl2_ff[1] ),
    .X(_147_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _249_ (.Y(_015_),
    .A(_146_),
    .B(_147_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _250_ (.Y(_148_),
    .A(net185),
    .B(net107),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _251_ (.B(\mac2.sum_lvl1_ff[9] ),
    .A(\mac2.sum_lvl1_ff[1] ),
    .X(_149_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _252_ (.Y(_031_),
    .A(_148_),
    .B(_149_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _253_ (.B(net107),
    .A(\mac2.sum_lvl1_ff[0] ),
    .X(_030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _254_ (.Y(_150_),
    .A(net163),
    .B(net199),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _255_ (.B(\mac2.sum_lvl2_ff[5] ),
    .A(\mac2.sum_lvl2_ff[1] ),
    .X(_151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _256_ (.Y(_001_),
    .A(_150_),
    .B(_151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _257_ (.B(\mac2.sum_lvl2_ff[4] ),
    .A(net163),
    .X(_000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _258_ (.Y(_152_),
    .A(\mac1.total_sum[0] ),
    .B(\mac2.total_sum[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _259_ (.Y(_153_),
    .A(\mac1.total_sum[1] ),
    .B(\mac2.total_sum[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _260_ (.A(\mac1.total_sum[1] ),
    .B(\mac2.total_sum[1] ),
    .Y(_154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _261_ (.B(\mac2.total_sum[1] ),
    .A(\mac1.total_sum[1] ),
    .X(_155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _262_ (.Y(net2),
    .A(_152_),
    .B(_155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _263_ (.B1(_153_),
    .VDD(VPWR),
    .Y(_156_),
    .VSS(VGND),
    .A1(_152_),
    .A2(_154_));
 sg13g2_and2_1 _264_ (.A(\mac1.total_sum[2] ),
    .B(\mac2.total_sum[2] ),
    .X(_157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _265_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_158_),
    .B(\mac2.total_sum[2] ),
    .A(\mac1.total_sum[2] ));
 sg13g2_nand2b_1 _266_ (.Y(_159_),
    .B(_158_),
    .A_N(_157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _267_ (.Y(net3),
    .A(_156_),
    .B(_159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _268_ (.B(\mac2.total_sum[0] ),
    .A(\mac1.total_sum[0] ),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _269_ (.Y(_160_),
    .A(net177),
    .B(net93),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _270_ (.B(\mac1.products_ff[1] ),
    .A(\mac1.products_ff[18] ),
    .X(_161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _271_ (.Y(_003_),
    .A(_160_),
    .B(_161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _272_ (.B(net93),
    .A(\mac1.products_ff[17] ),
    .X(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _273_ (.Y(_162_),
    .A(net183),
    .B(net111),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _274_ (.B(\mac1.products_ff[52] ),
    .A(\mac1.products_ff[35] ),
    .X(_163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _275_ (.Y(_005_),
    .A(_162_),
    .B(_163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _276_ (.B(net111),
    .A(\mac1.products_ff[34] ),
    .X(_004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _277_ (.Y(_164_),
    .A(net187),
    .B(net113),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _278_ (.B(\mac1.products_ff[69] ),
    .A(\mac1.products_ff[86] ),
    .X(_165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _279_ (.Y(_007_),
    .A(_164_),
    .B(_165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _280_ (.B(net113),
    .A(\mac1.products_ff[85] ),
    .X(_006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _281_ (.Y(_166_),
    .A(net193),
    .B(net99),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _282_ (.B(\mac1.products_ff[120] ),
    .A(\mac1.products_ff[103] ),
    .X(_167_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _283_ (.Y(_009_),
    .A(_166_),
    .B(_167_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _284_ (.B(net99),
    .A(\mac1.products_ff[102] ),
    .X(_008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _285_ (.Y(_168_),
    .A(net175),
    .B(net145),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _286_ (.B(\mac1.sum_lvl1_ff[1] ),
    .A(\mac1.sum_lvl1_ff[9] ),
    .X(_169_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _287_ (.Y(_011_),
    .A(_168_),
    .B(_169_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _288_ (.B(net145),
    .A(\mac1.sum_lvl1_ff[8] ),
    .X(_010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _289_ (.Y(_170_),
    .A(net173),
    .B(net161),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _290_ (.B(\mac1.sum_lvl1_ff[17] ),
    .A(\mac1.sum_lvl1_ff[25] ),
    .X(_171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _291_ (.Y(_013_),
    .A(_170_),
    .B(_171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _292_ (.B(net161),
    .A(\mac1.sum_lvl1_ff[24] ),
    .X(_012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _293_ (.Y(_172_),
    .A(net201),
    .B(net115),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _294_ (.Y(_173_),
    .A(net170),
    .B(\mac2.sum_lvl3_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _295_ (.A(net170),
    .B(\mac2.sum_lvl3_ff[1] ),
    .Y(_174_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _296_ (.B(\mac2.sum_lvl3_ff[1] ),
    .A(net170),
    .X(_175_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _297_ (.Y(_021_),
    .A(_172_),
    .B(_175_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _298_ (.B(net115),
    .A(\mac2.sum_lvl3_ff[2] ),
    .X(_020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _299_ (.Y(_176_),
    .A(net179),
    .B(net109),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _300_ (.B(\mac2.products_ff[35] ),
    .A(\mac2.products_ff[52] ),
    .X(_177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _301_ (.Y(_025_),
    .A(_176_),
    .B(_177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _302_ (.B(net109),
    .A(\mac2.products_ff[51] ),
    .X(_024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _303_ (.Y(_178_),
    .A(net181),
    .B(net103),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _304_ (.B(\mac2.products_ff[86] ),
    .A(\mac2.products_ff[69] ),
    .X(_179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _305_ (.Y(_027_),
    .A(_178_),
    .B(_179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _306_ (.B(net103),
    .A(\mac2.products_ff[68] ),
    .X(_026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _307_ (.Y(_180_),
    .A(net195),
    .B(net123),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _308_ (.B(\mac2.products_ff[103] ),
    .A(\mac2.products_ff[120] ),
    .X(_181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _309_ (.Y(_029_),
    .A(_180_),
    .B(_181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _310_ (.B(net123),
    .A(\mac2.products_ff[119] ),
    .X(_028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _311_ (.Y(_182_),
    .A(net189),
    .B(net136),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _312_ (.B(\mac2.sum_lvl1_ff[25] ),
    .A(\mac2.sum_lvl1_ff[17] ),
    .X(_183_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _313_ (.Y(_033_),
    .A(_182_),
    .B(_183_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _314_ (.B(net136),
    .A(\mac2.sum_lvl1_ff[16] ),
    .X(_032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _315_ (.Y(_184_),
    .A(net191),
    .B(net95),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _316_ (.B(\mac2.products_ff[18] ),
    .A(\mac2.products_ff[1] ),
    .X(_185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _317_ (.Y(_023_),
    .A(_184_),
    .B(_185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _318_ (.B(net95),
    .A(\mac2.products_ff[0] ),
    .X(_022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _319_ (.B1(net168),
    .VDD(VPWR),
    .Y(_016_),
    .VSS(VGND),
    .A1(_142_),
    .A2(_144_));
 sg13g2_nand2_1 _320_ (.Y(_186_),
    .A(net148),
    .B(net45),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _321_ (.Y(_187_),
    .A(net130),
    .B(net56),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _322_ (.B(_187_),
    .A(_186_),
    .X(_067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _323_ (.Y(_188_),
    .A(net118),
    .B(net91),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _324_ (.Y(_189_),
    .A(net133),
    .B(net106),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _325_ (.B(_189_),
    .A(_188_),
    .X(_069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _326_ (.Y(_190_),
    .A(net121),
    .B(net86),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _327_ (.Y(_191_),
    .A(net141),
    .B(net51),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _328_ (.B(_191_),
    .A(_190_),
    .X(_035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _329_ (.Y(_192_),
    .A(net131),
    .B(net58),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _330_ (.Y(_193_),
    .A(net156),
    .B(net52),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _331_ (.B(_193_),
    .A(_192_),
    .X(_037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _332_ (.A2(_158_),
    .A1(_156_),
    .B1(_157_),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _333_ (.Y(_194_),
    .A(net140),
    .B(net41),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _334_ (.Y(_195_),
    .A(net127),
    .B(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _335_ (.B(_195_),
    .A(_194_),
    .X(_039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _336_ (.Y(_196_),
    .A(net152),
    .B(net57),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _337_ (.Y(_197_),
    .A(net157),
    .B(net42),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _338_ (.B(_197_),
    .A(_196_),
    .X(_041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _339_ (.Y(_198_),
    .A(net142),
    .B(net46),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _340_ (.Y(_199_),
    .A(net159),
    .B(net38),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _341_ (.B(_199_),
    .A(_198_),
    .X(_043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _342_ (.Y(_200_),
    .A(net128),
    .B(net97),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _343_ (.Y(_201_),
    .A(net147),
    .B(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _344_ (.B(_201_),
    .A(_200_),
    .X(_045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _345_ (.Y(_202_),
    .A(net129),
    .B(net55),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _346_ (.Y(_203_),
    .A(net134),
    .B(net98),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _347_ (.B(_203_),
    .A(_202_),
    .X(_047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _348_ (.Y(_204_),
    .A(net160),
    .B(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _349_ (.Y(_205_),
    .A(net117),
    .B(net53),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _350_ (.B(_205_),
    .A(_204_),
    .X(_049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _351_ (.Y(_206_),
    .A(net122),
    .B(net87),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _352_ (.Y(_207_),
    .A(net139),
    .B(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _353_ (.B(_207_),
    .A(_206_),
    .X(_051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _354_ (.Y(_208_),
    .A(net150),
    .B(net105),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _355_ (.Y(_209_),
    .A(net138),
    .B(net59),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _356_ (.B(_209_),
    .A(_208_),
    .X(_053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _357_ (.Y(_210_),
    .A(net120),
    .B(net54),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _358_ (.Y(_211_),
    .A(net151),
    .B(net90),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _359_ (.B(_211_),
    .A(_210_),
    .X(_055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _360_ (.Y(_212_),
    .A(net135),
    .B(net92),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _361_ (.Y(_213_),
    .A(net126),
    .B(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _362_ (.B(_213_),
    .A(_212_),
    .X(_057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _363_ (.B1(net171),
    .VDD(VPWR),
    .Y(_019_),
    .VSS(VGND),
    .A1(_172_),
    .A2(_174_));
 sg13g2_nand2_1 _364_ (.Y(_214_),
    .A(net155),
    .B(net50),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _365_ (.Y(_215_),
    .A(net149),
    .B(net49),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _366_ (.B(_215_),
    .A(_214_),
    .X(_059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _367_ (.Y(_216_),
    .A(net158),
    .B(net102),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _368_ (.Y(_217_),
    .A(net125),
    .B(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _369_ (.B(_217_),
    .A(_216_),
    .X(_061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _370_ (.Y(_218_),
    .A(net143),
    .B(net89),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _371_ (.Y(_219_),
    .A(net144),
    .B(net37),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _372_ (.B(_219_),
    .A(_218_),
    .X(_063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _373_ (.Y(_220_),
    .A(net119),
    .B(net88),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _374_ (.Y(_221_),
    .A(net132),
    .B(net101),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _375_ (.B(_221_),
    .A(_220_),
    .X(_065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _376_ (.A(net159),
    .X(_070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _377_ (.A(net46),
    .X(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _378_ (.A(net147),
    .X(_072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _379_ (.A(net97),
    .X(_073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _380_ (.A(net134),
    .X(_074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _381_ (.A(net55),
    .X(_075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _382_ (.A(net117),
    .X(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _383_ (.A(net47),
    .X(_077_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _384_ (.A(net139),
    .X(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _385_ (.A(net87),
    .X(_079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _386_ (.A(net138),
    .X(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _387_ (.A(net105),
    .X(_081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _388_ (.A(net151),
    .X(_082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _389_ (.A(net54),
    .X(_083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _390_ (.A(net126),
    .X(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _391_ (.A(net92),
    .X(_085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _392_ (.A(net133),
    .X(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _393_ (.A(net91),
    .X(_087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _394_ (.A(net142),
    .X(_088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _395_ (.A(net38),
    .X(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _396_ (.A(net128),
    .X(_090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _397_ (.A(net48),
    .X(_091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _398_ (.A(net129),
    .X(_092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _399_ (.A(net98),
    .X(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _400_ (.A(net160),
    .X(_094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _401_ (.A(net53),
    .X(_095_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _402_ (.A(net122),
    .X(_096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _403_ (.A(net44),
    .X(_097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _404_ (.A(net150),
    .X(_098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _405_ (.A(net59),
    .X(_099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _406_ (.A(net120),
    .X(_100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _407_ (.A(net90),
    .X(_101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _408_ (.A(net135),
    .X(_102_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _409_ (.A(net40),
    .X(_103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _410_ (.A(net118),
    .X(_104_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _411_ (.A(net106),
    .X(_105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _412_ (.A(net132),
    .X(_106_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _413_ (.A(net88),
    .X(_107_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _414_ (.A(net157),
    .X(_108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _415_ (.A(net57),
    .X(_109_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _416_ (.A(net148),
    .X(_110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _417_ (.A(net56),
    .X(_111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _418_ (.A(net149),
    .X(_112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _419_ (.A(net50),
    .X(_113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _420_ (.A(net156),
    .X(_114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _421_ (.A(net58),
    .X(_115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _422_ (.A(net125),
    .X(_116_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _423_ (.A(net102),
    .X(_117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _424_ (.A(net144),
    .X(_118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _425_ (.A(net89),
    .X(_119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _426_ (.A(net141),
    .X(_120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _427_ (.A(net86),
    .X(_121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _428_ (.A(net127),
    .X(_122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _429_ (.A(net41),
    .X(_123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _430_ (.A(net119),
    .X(_124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _431_ (.A(net101),
    .X(_125_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _432_ (.A(net152),
    .X(_126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _433_ (.A(net42),
    .X(_127_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _434_ (.A(net130),
    .X(_128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _435_ (.A(net45),
    .X(_129_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _436_ (.A(net155),
    .X(_130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _437_ (.A(net49),
    .X(_131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _438_ (.A(net131),
    .X(_132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _439_ (.A(net52),
    .X(_133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _440_ (.A(net158),
    .X(_134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _441_ (.A(net39),
    .X(_135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _442_ (.A(net143),
    .X(_136_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _443_ (.A(net37),
    .X(_137_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _444_ (.A(net121),
    .X(_138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _445_ (.A(net51),
    .X(_139_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _446_ (.A(net140),
    .X(_140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _447_ (.A(net43),
    .X(_141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbpq_1 _448_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_042_),
    .Q(\mac1.products_ff[0] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _449_ (.RESET_B(net81),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_043_),
    .Q(\mac1.products_ff[1] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _450_ (.RESET_B(net74),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_044_),
    .Q(\mac1.products_ff[17] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _451_ (.RESET_B(net81),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_045_),
    .Q(\mac1.products_ff[18] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _452_ (.RESET_B(net85),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_046_),
    .Q(\mac1.products_ff[34] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _453_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_047_),
    .Q(\mac1.products_ff[35] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _454_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_048_),
    .Q(\mac1.products_ff[51] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _455_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_049_),
    .Q(\mac1.products_ff[52] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _456_ (.RESET_B(net78),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_050_),
    .Q(\mac1.products_ff[68] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _457_ (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_051_),
    .Q(\mac1.products_ff[69] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _458_ (.RESET_B(net78),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_052_),
    .Q(\mac1.products_ff[85] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _459_ (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_053_),
    .Q(\mac1.products_ff[86] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _460_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_054_),
    .Q(\mac1.products_ff[102] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _461_ (.RESET_B(net75),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_055_),
    .Q(\mac1.products_ff[103] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _462_ (.RESET_B(net75),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_056_),
    .Q(\mac1.products_ff[119] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _463_ (.RESET_B(net75),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_057_),
    .Q(\mac1.products_ff[120] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _464_ (.RESET_B(net61),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_068_),
    .Q(\mac1.products_ff[136] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _465_ (.RESET_B(net61),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_069_),
    .Q(\mac1.products_ff[137] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _466_ (.RESET_B(net74),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net94),
    .Q(\mac1.sum_lvl1_ff[0] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _467_ (.RESET_B(net74),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net178),
    .Q(\mac1.sum_lvl1_ff[1] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _468_ (.RESET_B(net74),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net112),
    .Q(\mac1.sum_lvl1_ff[8] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _469_ (.RESET_B(net74),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net184),
    .Q(\mac1.sum_lvl1_ff[9] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _470_ (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net114),
    .Q(\mac1.sum_lvl1_ff[16] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _471_ (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net188),
    .Q(\mac1.sum_lvl1_ff[17] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _472_ (.RESET_B(net75),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net100),
    .Q(\mac1.sum_lvl1_ff[24] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _473_ (.RESET_B(net75),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net194),
    .Q(\mac1.sum_lvl1_ff[25] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _474_ (.RESET_B(net61),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net27),
    .Q(\mac1.sum_lvl1_ff[32] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _475_ (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net33),
    .Q(\mac1.sum_lvl1_ff[33] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _476_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net146),
    .Q(\mac1.sum_lvl2_ff[0] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _477_ (.RESET_B(net74),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net176),
    .Q(\mac1.sum_lvl2_ff[1] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _478_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net162),
    .Q(\mac1.sum_lvl2_ff[4] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _479_ (.RESET_B(net75),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net174),
    .Q(\mac1.sum_lvl2_ff[5] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _480_ (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net35),
    .Q(\mac1.sum_lvl2_ff[8] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _481_ (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net31),
    .Q(\mac1.sum_lvl2_ff[9] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _482_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net154),
    .Q(\mac1.sum_lvl3_ff[0] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _483_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net198),
    .Q(\mac1.sum_lvl3_ff[1] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _484_ (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net36),
    .Q(\mac1.sum_lvl3_ff[2] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _485_ (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net30),
    .Q(\mac1.sum_lvl3_ff[3] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _486_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net166),
    .Q(\mac1.total_sum[0] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _487_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net204),
    .Q(\mac1.total_sum[1] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _488_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net169),
    .Q(\mac1.total_sum[2] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _489_ (.RESET_B(net69),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_064_),
    .Q(\mac2.products_ff[0] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _490_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_065_),
    .Q(\mac2.products_ff[1] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _491_ (.RESET_B(net69),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_040_),
    .Q(\mac2.products_ff[17] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _492_ (.RESET_B(net69),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_041_),
    .Q(\mac2.products_ff[18] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _493_ (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_066_),
    .Q(\mac2.products_ff[34] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _494_ (.RESET_B(net68),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_067_),
    .Q(\mac2.products_ff[35] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _495_ (.RESET_B(net68),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_058_),
    .Q(\mac2.products_ff[51] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _496_ (.RESET_B(net68),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_059_),
    .Q(\mac2.products_ff[52] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _497_ (.RESET_B(net80),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_036_),
    .Q(\mac2.products_ff[68] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _498_ (.RESET_B(net80),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_037_),
    .Q(\mac2.products_ff[69] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _499_ (.RESET_B(net80),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_060_),
    .Q(\mac2.products_ff[85] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _500_ (.RESET_B(net80),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_061_),
    .Q(\mac2.products_ff[86] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _501_ (.RESET_B(net82),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_062_),
    .Q(\mac2.products_ff[102] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _502_ (.RESET_B(net84),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_063_),
    .Q(\mac2.products_ff[103] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _503_ (.RESET_B(net82),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_034_),
    .Q(\mac2.products_ff[119] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _504_ (.RESET_B(net82),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_035_),
    .Q(\mac2.products_ff[120] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _505_ (.RESET_B(net62),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_038_),
    .Q(\mac2.products_ff[136] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _506_ (.RESET_B(net62),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_039_),
    .Q(\mac2.products_ff[137] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _507_ (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net96),
    .Q(\mac2.sum_lvl1_ff[0] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _508_ (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net192),
    .Q(\mac2.sum_lvl1_ff[1] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _509_ (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net110),
    .Q(\mac2.sum_lvl1_ff[8] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _510_ (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net180),
    .Q(\mac2.sum_lvl1_ff[9] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _511_ (.RESET_B(net80),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net104),
    .Q(\mac2.sum_lvl1_ff[16] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _512_ (.RESET_B(net80),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net182),
    .Q(\mac2.sum_lvl1_ff[17] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _513_ (.RESET_B(net81),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net124),
    .Q(\mac2.sum_lvl1_ff[24] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _514_ (.RESET_B(net82),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net196),
    .Q(\mac2.sum_lvl1_ff[25] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _515_ (.RESET_B(net62),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net25),
    .Q(\mac2.sum_lvl1_ff[32] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _516_ (.RESET_B(net63),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net29),
    .Q(\mac2.sum_lvl1_ff[33] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _517_ (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net108),
    .Q(\mac2.sum_lvl2_ff[0] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _518_ (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net186),
    .Q(\mac2.sum_lvl2_ff[1] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _519_ (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net137),
    .Q(\mac2.sum_lvl2_ff[4] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _520_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net190),
    .Q(\mac2.sum_lvl2_ff[5] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _521_ (.RESET_B(net63),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net26),
    .Q(\mac2.sum_lvl2_ff[8] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _522_ (.RESET_B(net63),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net28),
    .Q(\mac2.sum_lvl2_ff[9] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _523_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net164),
    .Q(\mac2.sum_lvl3_ff[0] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _524_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net200),
    .Q(\mac2.sum_lvl3_ff[1] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _525_ (.RESET_B(net62),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net32),
    .Q(\mac2.sum_lvl3_ff[2] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _526_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net34),
    .Q(\mac2.sum_lvl3_ff[3] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _527_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net116),
    .Q(\mac2.total_sum[0] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _528_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net202),
    .Q(\mac2.total_sum[1] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _529_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net172),
    .Q(\mac2.total_sum[2] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _530_ (.RESET_B(net83),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_070_),
    .Q(\DP_1.matrix[0] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _531_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_071_),
    .Q(\DP_1.matrix[1] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _532_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_072_),
    .Q(\DP_1.matrix[9] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _533_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_073_),
    .Q(\DP_1.matrix[10] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _534_ (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_074_),
    .Q(\DP_1.matrix[18] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _535_ (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_075_),
    .Q(\DP_1.matrix[19] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _536_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_076_),
    .Q(\DP_1.matrix[27] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _537_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_077_),
    .Q(\DP_1.matrix[28] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _538_ (.RESET_B(net75),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_078_),
    .Q(\DP_1.matrix[36] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _539_ (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_079_),
    .Q(\DP_1.matrix[37] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _540_ (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_080_),
    .Q(\DP_1.matrix[45] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _541_ (.RESET_B(net83),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_081_),
    .Q(\DP_1.matrix[46] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _542_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_082_),
    .Q(\DP_1.matrix[54] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _543_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_083_),
    .Q(\DP_1.matrix[55] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _544_ (.RESET_B(net76),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_084_),
    .Q(\DP_1.matrix[63] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _545_ (.RESET_B(net76),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_085_),
    .Q(\DP_1.matrix[64] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _546_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_086_),
    .Q(\DP_1.matrix[72] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _547_ (.RESET_B(net61),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_087_),
    .Q(\DP_1.matrix[73] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _548_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_088_),
    .Q(\DP_2.matrix[0] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _549_ (.RESET_B(net83),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_089_),
    .Q(\DP_2.matrix[1] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _550_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_090_),
    .Q(\DP_2.matrix[9] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _551_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_091_),
    .Q(\DP_2.matrix[10] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _552_ (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_092_),
    .Q(\DP_2.matrix[18] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _553_ (.RESET_B(net66),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_093_),
    .Q(\DP_2.matrix[19] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _554_ (.RESET_B(net66),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_094_),
    .Q(\DP_2.matrix[27] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _555_ (.RESET_B(net66),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_095_),
    .Q(\DP_2.matrix[28] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _556_ (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_096_),
    .Q(\DP_2.matrix[36] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _557_ (.RESET_B(net76),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_097_),
    .Q(\DP_2.matrix[37] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _558_ (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_098_),
    .Q(\DP_2.matrix[45] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _559_ (.RESET_B(net83),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_099_),
    .Q(\DP_2.matrix[46] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _560_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_100_),
    .Q(\DP_2.matrix[54] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _561_ (.RESET_B(net74),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_101_),
    .Q(\DP_2.matrix[55] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _562_ (.RESET_B(net75),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_102_),
    .Q(\DP_2.matrix[63] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _563_ (.RESET_B(net76),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_103_),
    .Q(\DP_2.matrix[64] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _564_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_104_),
    .Q(\DP_2.matrix[72] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _565_ (.RESET_B(net61),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_105_),
    .Q(\DP_2.matrix[73] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _566_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_106_),
    .Q(\DP_3.matrix[0] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _567_ (.RESET_B(net68),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_107_),
    .Q(\DP_3.matrix[1] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _568_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_108_),
    .Q(\DP_3.matrix[9] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _569_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_109_),
    .Q(\DP_3.matrix[10] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _570_ (.RESET_B(net69),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_110_),
    .Q(\DP_3.matrix[18] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _571_ (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_111_),
    .Q(\DP_3.matrix[19] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _572_ (.RESET_B(net68),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_112_),
    .Q(\DP_3.matrix[27] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _573_ (.RESET_B(net68),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_113_),
    .Q(\DP_3.matrix[28] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _574_ (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_114_),
    .Q(\DP_3.matrix[36] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _575_ (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_115_),
    .Q(\DP_3.matrix[37] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _576_ (.RESET_B(net80),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_116_),
    .Q(\DP_3.matrix[45] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _577_ (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_117_),
    .Q(\DP_3.matrix[46] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _578_ (.RESET_B(net83),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_118_),
    .Q(\DP_3.matrix[54] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _579_ (.RESET_B(net83),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_119_),
    .Q(\DP_3.matrix[55] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _580_ (.RESET_B(net82),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_120_),
    .Q(\DP_3.matrix[63] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _581_ (.RESET_B(net82),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_121_),
    .Q(\DP_3.matrix[64] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _582_ (.RESET_B(net62),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_122_),
    .Q(\DP_3.matrix[72] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _583_ (.RESET_B(net62),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_123_),
    .Q(\DP_3.matrix[73] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _584_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_124_),
    .Q(\DP_4.matrix[0] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _585_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_125_),
    .Q(\DP_4.matrix[1] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _586_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_126_),
    .Q(\DP_4.matrix[9] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _587_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_127_),
    .Q(\DP_4.matrix[10] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _588_ (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_128_),
    .Q(\DP_4.matrix[18] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _589_ (.RESET_B(net69),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_129_),
    .Q(\DP_4.matrix[19] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _590_ (.RESET_B(net68),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_130_),
    .Q(\DP_4.matrix[27] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _591_ (.RESET_B(net68),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_131_),
    .Q(\DP_4.matrix[28] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _592_ (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_132_),
    .Q(\DP_4.matrix[36] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _593_ (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_133_),
    .Q(\DP_4.matrix[37] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_2 _594_ (.RESET_B(net72),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_134_),
    .Q(\DP_4.matrix[45] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _595_ (.RESET_B(net80),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_135_),
    .Q(\DP_4.matrix[46] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _596_ (.RESET_B(net84),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_136_),
    .Q(\DP_4.matrix[54] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _597_ (.RESET_B(net83),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_137_),
    .Q(\DP_4.matrix[55] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _598_ (.RESET_B(net82),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_138_),
    .Q(\DP_4.matrix[63] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _599_ (.RESET_B(net82),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_139_),
    .Q(\DP_4.matrix[64] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _600_ (.RESET_B(net62),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_140_),
    .Q(\DP_4.matrix[72] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _601_ (.RESET_B(net62),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_141_),
    .Q(\DP_4.matrix[73] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_tiehi heichips25_template_18 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net18));
 sg13g2_tiehi heichips25_template_19 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net19));
 sg13g2_tiehi heichips25_template_20 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net20));
 sg13g2_tiehi heichips25_template_21 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net21));
 sg13g2_tiehi heichips25_template_22 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net22));
 sg13g2_tiehi heichips25_template_23 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net23));
 sg13g2_tiehi heichips25_template_24 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net24));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_template_6 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net6));
 sg13g2_tielo heichips25_template_7 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net7));
 sg13g2_tielo heichips25_template_8 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net8));
 sg13g2_tielo heichips25_template_9 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net9));
 sg13g2_tielo heichips25_template_10 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net10));
 sg13g2_tielo heichips25_template_11 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net11));
 sg13g2_tielo heichips25_template_12 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net12));
 sg13g2_tielo heichips25_template_13 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net13));
 sg13g2_tielo heichips25_template_14 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net14));
 sg13g2_tielo heichips25_template_15 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net15));
 sg13g2_tielo heichips25_template_16 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net16));
 sg13g2_tiehi heichips25_template_17 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net17));
 sg13g2_buf_8 fanout60 (.A(net61),
    .X(net60),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout61 (.A(net63),
    .X(net61),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout62 (.A(net63),
    .X(net62),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout63 (.A(net72),
    .X(net63),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout64 (.A(net66),
    .X(net64),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout65 (.A(net66),
    .X(net65),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout66 (.A(net72),
    .X(net66),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout67 (.A(net69),
    .X(net67),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout68 (.A(net69),
    .X(net68),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout69 (.A(net72),
    .X(net69),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout70 (.A(net71),
    .X(net70),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout71 (.A(net72),
    .X(net71),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout72 (.A(rst_n),
    .X(net72),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout73 (.A(net74),
    .X(net73),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout74 (.A(net85),
    .X(net74),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout75 (.A(net78),
    .X(net75),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout76 (.A(net78),
    .X(net76),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout77 (.A(net78),
    .X(net77),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout78 (.A(net85),
    .X(net78),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout79 (.A(net81),
    .X(net79),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout80 (.A(net81),
    .X(net80),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout81 (.A(net84),
    .X(net81),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout82 (.A(net83),
    .X(net82),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout83 (.A(net84),
    .X(net83),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout84 (.A(net85),
    .X(net84),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout85 (.A(rst_n),
    .X(net85),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output1 (.A(net1),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uo_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_template_5 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net5));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload0 (.VDD(VPWR),
    .A(clknet_5_7__leaf_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload1 (.VDD(VPWR),
    .A(clknet_5_11__leaf_clk),
    .VSS(VGND));
 sg13g2_buf_1 clkload2 (.A(clknet_5_12__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload3 (.VDD(VPWR),
    .A(clknet_5_15__leaf_clk),
    .VSS(VGND));
 sg13g2_buf_1 clkload4 (.A(clknet_5_17__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload5 (.VDD(VPWR),
    .A(clknet_5_23__leaf_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload6 (.VDD(VPWR),
    .A(clknet_5_27__leaf_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload7 (.VDD(VPWR),
    .A(clknet_5_31__leaf_clk),
    .VSS(VGND));
 sg13g2_dlygate4sd3_1 hold1 (.A(\mac2.products_ff[136] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold2 (.A(\mac2.sum_lvl1_ff[32] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold3 (.A(\mac1.products_ff[136] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold4 (.A(\mac2.sum_lvl1_ff[33] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold5 (.A(\mac2.products_ff[137] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold6 (.A(\mac1.sum_lvl2_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold7 (.A(\mac1.sum_lvl1_ff[33] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold8 (.A(\mac2.sum_lvl2_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold9 (.A(\mac1.products_ff[137] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold10 (.A(\mac2.sum_lvl2_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold11 (.A(\mac1.sum_lvl1_ff[32] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold12 (.A(\mac1.sum_lvl2_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold13 (.A(\DP_4.matrix[55] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold14 (.A(\DP_2.matrix[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold15 (.A(\DP_4.matrix[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold16 (.A(\DP_2.matrix[64] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold17 (.A(\DP_3.matrix[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold18 (.A(\DP_4.matrix[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold19 (.A(\DP_4.matrix[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold20 (.A(\DP_2.matrix[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold21 (.A(\DP_4.matrix[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold22 (.A(\DP_1.matrix[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold23 (.A(\DP_1.matrix[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold24 (.A(\DP_2.matrix[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold25 (.A(\DP_4.matrix[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold26 (.A(\DP_3.matrix[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold27 (.A(\DP_4.matrix[64] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold28 (.A(\DP_4.matrix[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold29 (.A(\DP_2.matrix[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold30 (.A(\DP_1.matrix[55] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold31 (.A(\DP_1.matrix[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold32 (.A(\DP_3.matrix[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold33 (.A(\DP_3.matrix[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold34 (.A(\DP_3.matrix[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold35 (.A(\DP_2.matrix[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold36 (.A(\DP_3.matrix[64] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold37 (.A(\DP_1.matrix[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold38 (.A(\DP_3.matrix[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold39 (.A(\DP_3.matrix[55] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold40 (.A(\DP_2.matrix[55] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold41 (.A(\DP_1.matrix[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold42 (.A(\DP_1.matrix[64] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold43 (.A(\mac1.products_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold44 (.A(_002_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold45 (.A(\mac2.products_ff[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold46 (.A(_022_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold47 (.A(\DP_1.matrix[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold48 (.A(\DP_2.matrix[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold49 (.A(\mac1.products_ff[119] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold50 (.A(_008_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold51 (.A(\DP_4.matrix[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold52 (.A(\DP_3.matrix[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold53 (.A(\mac2.products_ff[85] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold54 (.A(_026_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold55 (.A(\DP_1.matrix[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold56 (.A(\DP_2.matrix[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold57 (.A(\mac2.sum_lvl1_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold58 (.A(_030_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold59 (.A(\mac2.products_ff[34] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold60 (.A(_024_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold61 (.A(\mac1.products_ff[51] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold62 (.A(_004_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold63 (.A(\mac1.products_ff[68] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold64 (.A(_006_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold65 (.A(\mac2.sum_lvl3_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold66 (.A(_020_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold67 (.A(\DP_1.matrix[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold68 (.A(\DP_2.matrix[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold69 (.A(\DP_4.matrix[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold70 (.A(\DP_2.matrix[54] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold71 (.A(\DP_4.matrix[63] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold72 (.A(\DP_2.matrix[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold73 (.A(\mac2.products_ff[102] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold74 (.A(_028_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold75 (.A(\DP_3.matrix[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold76 (.A(\DP_1.matrix[63] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold77 (.A(\DP_3.matrix[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold78 (.A(\DP_2.matrix[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold79 (.A(\DP_2.matrix[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold80 (.A(\DP_4.matrix[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold81 (.A(\DP_4.matrix[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold82 (.A(\DP_3.matrix[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold83 (.A(\DP_1.matrix[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold84 (.A(\DP_1.matrix[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold85 (.A(\DP_2.matrix[63] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold86 (.A(\mac2.sum_lvl1_ff[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold87 (.A(_032_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold88 (.A(\DP_1.matrix[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold89 (.A(\DP_1.matrix[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold90 (.A(\DP_4.matrix[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold91 (.A(\DP_3.matrix[63] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold92 (.A(\DP_2.matrix[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold93 (.A(\DP_4.matrix[54] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold94 (.A(\DP_3.matrix[54] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold95 (.A(\mac1.sum_lvl1_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold96 (.A(_010_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold97 (.A(\DP_1.matrix[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold98 (.A(\DP_3.matrix[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold99 (.A(\DP_3.matrix[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold100 (.A(\DP_2.matrix[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold101 (.A(\DP_1.matrix[54] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold102 (.A(\DP_4.matrix[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold103 (.A(\mac1.sum_lvl2_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold104 (.A(_014_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold105 (.A(\DP_4.matrix[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold106 (.A(\DP_3.matrix[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold107 (.A(\DP_3.matrix[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold108 (.A(\DP_4.matrix[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold109 (.A(\DP_1.matrix[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold110 (.A(\DP_2.matrix[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold111 (.A(\mac1.sum_lvl1_ff[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold112 (.A(_012_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold113 (.A(\mac2.sum_lvl2_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold114 (.A(_000_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold115 (.A(\mac1.sum_lvl3_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold116 (.A(_017_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold117 (.A(\mac1.sum_lvl3_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold118 (.A(_143_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold119 (.A(_016_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold120 (.A(\mac2.sum_lvl3_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold121 (.A(_173_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold122 (.A(_019_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold123 (.A(\mac1.sum_lvl1_ff[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold124 (.A(_013_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold125 (.A(\mac1.sum_lvl1_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold126 (.A(_011_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold127 (.A(\mac1.products_ff[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold128 (.A(_003_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold129 (.A(\mac2.products_ff[51] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold130 (.A(_025_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold131 (.A(\mac2.products_ff[68] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold132 (.A(_027_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold133 (.A(\mac1.products_ff[34] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold134 (.A(_005_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold135 (.A(\mac2.sum_lvl1_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold136 (.A(_031_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold137 (.A(\mac1.products_ff[85] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold138 (.A(_007_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold139 (.A(\mac2.sum_lvl1_ff[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold140 (.A(_033_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold141 (.A(\mac2.products_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold142 (.A(_023_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold143 (.A(\mac1.products_ff[102] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold144 (.A(_009_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold145 (.A(\mac2.products_ff[119] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold146 (.A(_029_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold147 (.A(\mac1.sum_lvl2_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold148 (.A(_015_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold149 (.A(\mac2.sum_lvl2_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold150 (.A(_001_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold151 (.A(\mac2.sum_lvl3_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold152 (.A(_021_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold153 (.A(\mac1.sum_lvl3_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold154 (.A(_018_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net204));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_1028 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net17;
 assign uio_oe[1] = net18;
 assign uio_oe[2] = net19;
 assign uio_oe[3] = net20;
 assign uio_oe[4] = net21;
 assign uio_oe[5] = net22;
 assign uio_oe[6] = net23;
 assign uio_oe[7] = net24;
 assign uio_out[0] = net5;
 assign uio_out[1] = net6;
 assign uio_out[2] = net7;
 assign uio_out[3] = net8;
 assign uio_out[4] = net9;
 assign uio_out[5] = net10;
 assign uio_out[6] = net11;
 assign uio_out[7] = net12;
 assign uo_out[4] = net13;
 assign uo_out[5] = net14;
 assign uo_out[6] = net15;
 assign uo_out[7] = net16;
endmodule
