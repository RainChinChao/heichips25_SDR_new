module heichips25_template (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \DP_1.I_range.data_plus_4[6] ;
 wire \DP_1.I_range.out_data[2] ;
 wire \DP_1.I_range.out_data[3] ;
 wire \DP_1.I_range.out_data[4] ;
 wire \DP_1.I_range.out_data[5] ;
 wire \DP_1.I_range.out_data[6] ;
 wire \DP_1.Q_range.data_plus_4[6] ;
 wire \DP_1.Q_range.out_data[2] ;
 wire \DP_1.Q_range.out_data[3] ;
 wire \DP_1.Q_range.out_data[4] ;
 wire \DP_1.Q_range.out_data[5] ;
 wire \DP_1.Q_range.out_data[6] ;
 wire \DP_1.matrix[0] ;
 wire \DP_1.matrix[1] ;
 wire \DP_1.matrix[2] ;
 wire \DP_1.matrix[36] ;
 wire \DP_1.matrix[37] ;
 wire \DP_1.matrix[38] ;
 wire \DP_1.matrix[39] ;
 wire \DP_1.matrix[3] ;
 wire \DP_1.matrix[40] ;
 wire \DP_1.matrix[41] ;
 wire \DP_1.matrix[42] ;
 wire \DP_1.matrix[43] ;
 wire \DP_1.matrix[44] ;
 wire \DP_1.matrix[4] ;
 wire \DP_1.matrix[5] ;
 wire \DP_1.matrix[6] ;
 wire \DP_1.matrix[72] ;
 wire \DP_1.matrix[73] ;
 wire \DP_1.matrix[74] ;
 wire \DP_1.matrix[75] ;
 wire \DP_1.matrix[76] ;
 wire \DP_1.matrix[77] ;
 wire \DP_1.matrix[78] ;
 wire \DP_1.matrix[79] ;
 wire \DP_1.matrix[7] ;
 wire \DP_1.matrix[80] ;
 wire \DP_1.matrix[8] ;
 wire \DP_2.I_range.data_plus_4[6] ;
 wire \DP_2.I_range.out_data[2] ;
 wire \DP_2.I_range.out_data[3] ;
 wire \DP_2.I_range.out_data[4] ;
 wire \DP_2.I_range.out_data[5] ;
 wire \DP_2.I_range.out_data[6] ;
 wire \DP_2.Q_range.data_plus_4[6] ;
 wire \DP_2.Q_range.out_data[2] ;
 wire \DP_2.Q_range.out_data[3] ;
 wire \DP_2.Q_range.out_data[4] ;
 wire \DP_2.Q_range.out_data[5] ;
 wire \DP_2.Q_range.out_data[6] ;
 wire \DP_2.matrix[0] ;
 wire \DP_2.matrix[1] ;
 wire \DP_2.matrix[2] ;
 wire \DP_2.matrix[36] ;
 wire \DP_2.matrix[37] ;
 wire \DP_2.matrix[38] ;
 wire \DP_2.matrix[39] ;
 wire \DP_2.matrix[3] ;
 wire \DP_2.matrix[40] ;
 wire \DP_2.matrix[41] ;
 wire \DP_2.matrix[42] ;
 wire \DP_2.matrix[43] ;
 wire \DP_2.matrix[44] ;
 wire \DP_2.matrix[4] ;
 wire \DP_2.matrix[5] ;
 wire \DP_2.matrix[6] ;
 wire \DP_2.matrix[72] ;
 wire \DP_2.matrix[73] ;
 wire \DP_2.matrix[74] ;
 wire \DP_2.matrix[75] ;
 wire \DP_2.matrix[76] ;
 wire \DP_2.matrix[77] ;
 wire \DP_2.matrix[78] ;
 wire \DP_2.matrix[79] ;
 wire \DP_2.matrix[7] ;
 wire \DP_2.matrix[80] ;
 wire \DP_2.matrix[8] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire \mac1.products_ff[0] ;
 wire \mac1.products_ff[10] ;
 wire \mac1.products_ff[11] ;
 wire \mac1.products_ff[12] ;
 wire \mac1.products_ff[136] ;
 wire \mac1.products_ff[137] ;
 wire \mac1.products_ff[138] ;
 wire \mac1.products_ff[139] ;
 wire \mac1.products_ff[13] ;
 wire \mac1.products_ff[140] ;
 wire \mac1.products_ff[141] ;
 wire \mac1.products_ff[142] ;
 wire \mac1.products_ff[143] ;
 wire \mac1.products_ff[144] ;
 wire \mac1.products_ff[145] ;
 wire \mac1.products_ff[146] ;
 wire \mac1.products_ff[147] ;
 wire \mac1.products_ff[148] ;
 wire \mac1.products_ff[149] ;
 wire \mac1.products_ff[14] ;
 wire \mac1.products_ff[150] ;
 wire \mac1.products_ff[151] ;
 wire \mac1.products_ff[15] ;
 wire \mac1.products_ff[1] ;
 wire \mac1.products_ff[2] ;
 wire \mac1.products_ff[3] ;
 wire \mac1.products_ff[4] ;
 wire \mac1.products_ff[5] ;
 wire \mac1.products_ff[68] ;
 wire \mac1.products_ff[69] ;
 wire \mac1.products_ff[6] ;
 wire \mac1.products_ff[70] ;
 wire \mac1.products_ff[71] ;
 wire \mac1.products_ff[72] ;
 wire \mac1.products_ff[73] ;
 wire \mac1.products_ff[74] ;
 wire \mac1.products_ff[75] ;
 wire \mac1.products_ff[76] ;
 wire \mac1.products_ff[77] ;
 wire \mac1.products_ff[78] ;
 wire \mac1.products_ff[79] ;
 wire \mac1.products_ff[7] ;
 wire \mac1.products_ff[80] ;
 wire \mac1.products_ff[81] ;
 wire \mac1.products_ff[82] ;
 wire \mac1.products_ff[83] ;
 wire \mac1.products_ff[8] ;
 wire \mac1.products_ff[9] ;
 wire \mac1.sum_lvl1_ff[0] ;
 wire \mac1.sum_lvl1_ff[10] ;
 wire \mac1.sum_lvl1_ff[11] ;
 wire \mac1.sum_lvl1_ff[12] ;
 wire \mac1.sum_lvl1_ff[13] ;
 wire \mac1.sum_lvl1_ff[14] ;
 wire \mac1.sum_lvl1_ff[15] ;
 wire \mac1.sum_lvl1_ff[1] ;
 wire \mac1.sum_lvl1_ff[2] ;
 wire \mac1.sum_lvl1_ff[36] ;
 wire \mac1.sum_lvl1_ff[37] ;
 wire \mac1.sum_lvl1_ff[38] ;
 wire \mac1.sum_lvl1_ff[39] ;
 wire \mac1.sum_lvl1_ff[3] ;
 wire \mac1.sum_lvl1_ff[40] ;
 wire \mac1.sum_lvl1_ff[41] ;
 wire \mac1.sum_lvl1_ff[42] ;
 wire \mac1.sum_lvl1_ff[43] ;
 wire \mac1.sum_lvl1_ff[44] ;
 wire \mac1.sum_lvl1_ff[45] ;
 wire \mac1.sum_lvl1_ff[46] ;
 wire \mac1.sum_lvl1_ff[47] ;
 wire \mac1.sum_lvl1_ff[48] ;
 wire \mac1.sum_lvl1_ff[49] ;
 wire \mac1.sum_lvl1_ff[4] ;
 wire \mac1.sum_lvl1_ff[50] ;
 wire \mac1.sum_lvl1_ff[51] ;
 wire \mac1.sum_lvl1_ff[5] ;
 wire \mac1.sum_lvl1_ff[6] ;
 wire \mac1.sum_lvl1_ff[72] ;
 wire \mac1.sum_lvl1_ff[73] ;
 wire \mac1.sum_lvl1_ff[74] ;
 wire \mac1.sum_lvl1_ff[75] ;
 wire \mac1.sum_lvl1_ff[76] ;
 wire \mac1.sum_lvl1_ff[77] ;
 wire \mac1.sum_lvl1_ff[78] ;
 wire \mac1.sum_lvl1_ff[79] ;
 wire \mac1.sum_lvl1_ff[7] ;
 wire \mac1.sum_lvl1_ff[80] ;
 wire \mac1.sum_lvl1_ff[81] ;
 wire \mac1.sum_lvl1_ff[82] ;
 wire \mac1.sum_lvl1_ff[83] ;
 wire \mac1.sum_lvl1_ff[84] ;
 wire \mac1.sum_lvl1_ff[85] ;
 wire \mac1.sum_lvl1_ff[86] ;
 wire \mac1.sum_lvl1_ff[87] ;
 wire \mac1.sum_lvl1_ff[8] ;
 wire \mac1.sum_lvl1_ff[9] ;
 wire \mac1.sum_lvl2_ff[0] ;
 wire \mac1.sum_lvl2_ff[10] ;
 wire \mac1.sum_lvl2_ff[11] ;
 wire \mac1.sum_lvl2_ff[12] ;
 wire \mac1.sum_lvl2_ff[13] ;
 wire \mac1.sum_lvl2_ff[14] ;
 wire \mac1.sum_lvl2_ff[15] ;
 wire \mac1.sum_lvl2_ff[19] ;
 wire \mac1.sum_lvl2_ff[1] ;
 wire \mac1.sum_lvl2_ff[20] ;
 wire \mac1.sum_lvl2_ff[21] ;
 wire \mac1.sum_lvl2_ff[22] ;
 wire \mac1.sum_lvl2_ff[23] ;
 wire \mac1.sum_lvl2_ff[24] ;
 wire \mac1.sum_lvl2_ff[25] ;
 wire \mac1.sum_lvl2_ff[26] ;
 wire \mac1.sum_lvl2_ff[27] ;
 wire \mac1.sum_lvl2_ff[28] ;
 wire \mac1.sum_lvl2_ff[29] ;
 wire \mac1.sum_lvl2_ff[2] ;
 wire \mac1.sum_lvl2_ff[30] ;
 wire \mac1.sum_lvl2_ff[31] ;
 wire \mac1.sum_lvl2_ff[32] ;
 wire \mac1.sum_lvl2_ff[33] ;
 wire \mac1.sum_lvl2_ff[34] ;
 wire \mac1.sum_lvl2_ff[38] ;
 wire \mac1.sum_lvl2_ff[39] ;
 wire \mac1.sum_lvl2_ff[3] ;
 wire \mac1.sum_lvl2_ff[40] ;
 wire \mac1.sum_lvl2_ff[41] ;
 wire \mac1.sum_lvl2_ff[42] ;
 wire \mac1.sum_lvl2_ff[43] ;
 wire \mac1.sum_lvl2_ff[44] ;
 wire \mac1.sum_lvl2_ff[45] ;
 wire \mac1.sum_lvl2_ff[46] ;
 wire \mac1.sum_lvl2_ff[47] ;
 wire \mac1.sum_lvl2_ff[48] ;
 wire \mac1.sum_lvl2_ff[49] ;
 wire \mac1.sum_lvl2_ff[4] ;
 wire \mac1.sum_lvl2_ff[50] ;
 wire \mac1.sum_lvl2_ff[51] ;
 wire \mac1.sum_lvl2_ff[52] ;
 wire \mac1.sum_lvl2_ff[53] ;
 wire \mac1.sum_lvl2_ff[5] ;
 wire \mac1.sum_lvl2_ff[6] ;
 wire \mac1.sum_lvl2_ff[7] ;
 wire \mac1.sum_lvl2_ff[8] ;
 wire \mac1.sum_lvl2_ff[9] ;
 wire \mac1.sum_lvl3_ff[0] ;
 wire \mac1.sum_lvl3_ff[10] ;
 wire \mac1.sum_lvl3_ff[11] ;
 wire \mac1.sum_lvl3_ff[12] ;
 wire \mac1.sum_lvl3_ff[13] ;
 wire \mac1.sum_lvl3_ff[14] ;
 wire \mac1.sum_lvl3_ff[15] ;
 wire \mac1.sum_lvl3_ff[1] ;
 wire \mac1.sum_lvl3_ff[20] ;
 wire \mac1.sum_lvl3_ff[21] ;
 wire \mac1.sum_lvl3_ff[22] ;
 wire \mac1.sum_lvl3_ff[23] ;
 wire \mac1.sum_lvl3_ff[24] ;
 wire \mac1.sum_lvl3_ff[25] ;
 wire \mac1.sum_lvl3_ff[26] ;
 wire \mac1.sum_lvl3_ff[27] ;
 wire \mac1.sum_lvl3_ff[28] ;
 wire \mac1.sum_lvl3_ff[29] ;
 wire \mac1.sum_lvl3_ff[2] ;
 wire \mac1.sum_lvl3_ff[30] ;
 wire \mac1.sum_lvl3_ff[31] ;
 wire \mac1.sum_lvl3_ff[32] ;
 wire \mac1.sum_lvl3_ff[33] ;
 wire \mac1.sum_lvl3_ff[34] ;
 wire \mac1.sum_lvl3_ff[35] ;
 wire \mac1.sum_lvl3_ff[3] ;
 wire \mac1.sum_lvl3_ff[4] ;
 wire \mac1.sum_lvl3_ff[5] ;
 wire \mac1.sum_lvl3_ff[6] ;
 wire \mac1.sum_lvl3_ff[7] ;
 wire \mac1.sum_lvl3_ff[8] ;
 wire \mac1.sum_lvl3_ff[9] ;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire clknet_leaf_0_clk;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net33;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;

 sg13g2_inv_1 _1501_ (.VDD(VPWR),
    .Y(_0842_),
    .A(\DP_2.Q_range.out_data[5] ),
    .VSS(VGND));
 sg13g2_inv_1 _1502_ (.VDD(VPWR),
    .Y(\DP_1.I_range.data_plus_4[6] ),
    .A(net4),
    .VSS(VGND));
 sg13g2_inv_1 _1503_ (.VDD(VPWR),
    .Y(\DP_2.I_range.data_plus_4[6] ),
    .A(net16),
    .VSS(VGND));
 sg13g2_inv_1 _1504_ (.VDD(VPWR),
    .Y(\DP_2.Q_range.data_plus_4[6] ),
    .A(net12),
    .VSS(VGND));
 sg13g2_inv_1 _1505_ (.VDD(VPWR),
    .Y(\DP_1.Q_range.data_plus_4[6] ),
    .A(net8),
    .VSS(VGND));
 sg13g2_nand2_1 _1506_ (.Y(_0843_),
    .A(net474),
    .B(net410),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1507_ (.Y(_0844_),
    .A(net417),
    .B(net472),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1508_ (.A(net472),
    .B(net412),
    .X(_0845_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _1509_ (.A(net417),
    .B(net470),
    .C(net472),
    .D(net412),
    .X(_0846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1510_ (.Y(_0847_),
    .B1(net472),
    .B2(net412),
    .A2(net470),
    .A1(net417),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1511_ (.A(_0843_),
    .B(_0846_),
    .C(_0847_),
    .Y(_0848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1512_ (.B1(_0843_),
    .VDD(VPWR),
    .Y(_0849_),
    .VSS(VGND),
    .A1(_0846_),
    .A2(_0847_));
 sg13g2_nor2b_1 _1513_ (.A(_0848_),
    .B_N(_0849_),
    .Y(_0850_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1514_ (.A(net474),
    .B(net417),
    .X(_0042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1515_ (.Y(_0851_),
    .A(_0845_),
    .B(_0042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1516_ (.B(_0850_),
    .C(_0042_),
    .A(_0845_),
    .Y(_0852_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1517_ (.Y(_0044_),
    .A(_0850_),
    .B(_0851_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1518_ (.Y(_0853_),
    .A(net474),
    .B(net408),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1519_ (.A(_0846_),
    .B(_0848_),
    .Y(_0854_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1520_ (.Y(_0855_),
    .A(net472),
    .B(net410),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _1521_ (.A(net417),
    .B(net470),
    .C(net412),
    .D(net468),
    .X(_0856_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1522_ (.Y(_0857_),
    .B1(net468),
    .B2(net417),
    .A2(net413),
    .A1(net470),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1523_ (.A(_0855_),
    .B(_0856_),
    .C(_0857_),
    .Y(_0858_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1524_ (.B1(_0855_),
    .VDD(VPWR),
    .Y(_0859_),
    .VSS(VGND),
    .A1(_0856_),
    .A2(_0857_));
 sg13g2_nor2b_1 _1525_ (.A(_0858_),
    .B_N(_0859_),
    .Y(_0860_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1526_ (.Y(_0861_),
    .B(_0860_),
    .A_N(_0854_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1527_ (.Y(_0862_),
    .A(_0854_),
    .B(_0860_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1528_ (.Y(_0863_),
    .B(_0862_),
    .A_N(_0853_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1529_ (.Y(_0864_),
    .A(_0853_),
    .B(_0862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _1530_ (.Y(_0865_),
    .B(_0864_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0852_));
 sg13g2_xnor2_1 _1531_ (.Y(_0045_),
    .A(_0852_),
    .B(_0864_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1532_ (.Y(_0866_),
    .B1(net406),
    .B2(net474),
    .A2(net408),
    .A1(net472),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _1533_ (.Y(_0867_),
    .A(net473),
    .B(net406),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1534_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0868_),
    .B(_0867_),
    .A(_0853_));
 sg13g2_nor2b_1 _1535_ (.A(_0866_),
    .B_N(_0868_),
    .Y(_0869_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1536_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0870_),
    .B(_0858_),
    .A(_0856_));
 sg13g2_nand2_1 _1537_ (.Y(_0871_),
    .A(net470),
    .B(net410),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _1538_ (.A(net417),
    .B(net412),
    .C(net468),
    .D(net466),
    .X(_0872_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _1539_ (.B(net413),
    .C(net468),
    .A(net418),
    .Y(_0873_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net466));
 sg13g2_a22oi_1 _1540_ (.Y(_0874_),
    .B1(net466),
    .B2(net418),
    .A2(net468),
    .A1(net412),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _1541_ (.A(_0871_),
    .B(_0872_),
    .C(_0874_),
    .X(_0875_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1542_ (.B1(_0871_),
    .VDD(VPWR),
    .Y(_0876_),
    .VSS(VGND),
    .A1(_0872_),
    .A2(_0874_));
 sg13g2_and3_1 _1543_ (.X(_0877_),
    .A(_0870_),
    .B(_0875_),
    .C(_0876_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _1544_ (.A2(_0876_),
    .A1(_0875_),
    .B1(_0870_),
    .X(_0878_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1545_ (.Y(_0879_),
    .B(_0878_),
    .A_N(_0877_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1546_ (.B(_0879_),
    .A(_0869_),
    .X(_0880_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1547_ (.Y(_0881_),
    .A(_0861_),
    .B(_0863_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1548_ (.A(_0880_),
    .B_N(_0881_),
    .Y(_0882_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1549_ (.Y(_0883_),
    .B(_0881_),
    .A_N(_0880_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1550_ (.A(_0881_),
    .B_N(_0880_),
    .Y(_0884_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1551_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0885_),
    .B(_0884_),
    .A(_0882_));
 sg13g2_nor2_1 _1552_ (.A(_0865_),
    .B(_0885_),
    .Y(_0886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1553_ (.B(_0885_),
    .A(_0865_),
    .X(_0046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _1554_ (.A2(_0878_),
    .A1(_0869_),
    .B1(_0877_),
    .X(_0887_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1555_ (.Y(_0888_),
    .A(net475),
    .B(net405),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1556_ (.Y(_0889_),
    .A(net471),
    .B(net406),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1557_ (.Y(_0890_),
    .A(net470),
    .B(net408),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1558_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0891_),
    .B(_0890_),
    .A(_0867_));
 sg13g2_and2_1 _1559_ (.A(_0867_),
    .B(_0890_),
    .X(_0892_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1560_ (.Y(_0893_),
    .A(_0867_),
    .B(_0890_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1561_ (.Y(_0894_),
    .A(_0888_),
    .B(_0893_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1562_ (.B1(_0873_),
    .VDD(VPWR),
    .Y(_0895_),
    .VSS(VGND),
    .A1(_0871_),
    .A2(_0874_));
 sg13g2_nand2_1 _1563_ (.Y(_0896_),
    .A(net410),
    .B(net468),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _1564_ (.A(net419),
    .B(net413),
    .C(net466),
    .D(net464),
    .X(_0897_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _1565_ (.B(net414),
    .C(net466),
    .A(net419),
    .Y(_0898_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net464));
 sg13g2_a22oi_1 _1566_ (.Y(_0899_),
    .B1(net464),
    .B2(net419),
    .A2(net466),
    .A1(net413),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _1567_ (.A(_0896_),
    .B(_0897_),
    .C(_0899_),
    .X(_0900_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1568_ (.B1(_0896_),
    .VDD(VPWR),
    .Y(_0901_),
    .VSS(VGND),
    .A1(_0897_),
    .A2(_0899_));
 sg13g2_and3_1 _1569_ (.X(_0902_),
    .A(_0895_),
    .B(_0900_),
    .C(_0901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1570_ (.B(_0900_),
    .C(_0901_),
    .A(_0895_),
    .Y(_0903_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1571_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0900_),
    .A2(_0901_),
    .Y(_0904_),
    .B1(_0895_));
 sg13g2_or3_1 _1572_ (.A(_0894_),
    .B(_0902_),
    .C(_0904_),
    .X(_0905_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1573_ (.B1(_0894_),
    .VDD(VPWR),
    .Y(_0906_),
    .VSS(VGND),
    .A1(_0902_),
    .A2(_0904_));
 sg13g2_nand2_1 _1574_ (.Y(_0907_),
    .A(_0905_),
    .B(_0906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1575_ (.B(_0905_),
    .C(_0906_),
    .A(_0887_),
    .Y(_0908_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1576_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0905_),
    .A2(_0906_),
    .Y(_0909_),
    .B1(_0887_));
 sg13g2_xnor2_1 _1577_ (.Y(_0910_),
    .A(_0887_),
    .B(_0907_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1578_ (.B(_0910_),
    .A(_0868_),
    .X(_0911_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1579_ (.A(_0883_),
    .B(_0911_),
    .Y(_0912_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1580_ (.Y(_0913_),
    .A(_0883_),
    .B(_0911_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _1581_ (.A(_0865_),
    .B(_0882_),
    .C(_0884_),
    .D(_0911_),
    .Y(_0914_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1582_ (.Y(_0069_),
    .A(_0886_),
    .B(_0913_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1583_ (.B1(_0908_),
    .VDD(VPWR),
    .Y(_0915_),
    .VSS(VGND),
    .A1(_0868_),
    .A2(_0909_));
 sg13g2_o21ai_1 _1584_ (.B1(_0891_),
    .VDD(VPWR),
    .Y(_0916_),
    .VSS(VGND),
    .A1(_0888_),
    .A2(_0892_));
 sg13g2_nand2_1 _1585_ (.Y(_0917_),
    .A(net475),
    .B(net403),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1586_ (.Y(_0918_),
    .B(_0916_),
    .A_N(_0917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1587_ (.Y(_0919_),
    .A(_0916_),
    .B(_0917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1588_ (.VDD(VPWR),
    .Y(_0920_),
    .A(_0919_),
    .VSS(VGND));
 sg13g2_o21ai_1 _1589_ (.B1(_0903_),
    .VDD(VPWR),
    .Y(_0921_),
    .VSS(VGND),
    .A1(_0894_),
    .A2(_0904_));
 sg13g2_nand2_1 _1590_ (.Y(_0922_),
    .A(net473),
    .B(net405),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1591_ (.Y(_0923_),
    .A(net469),
    .B(net406),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1592_ (.Y(_0924_),
    .A(net469),
    .B(net408),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1593_ (.B(_0924_),
    .A(_0889_),
    .X(_0925_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1594_ (.Y(_0926_),
    .B(_0925_),
    .A_N(_0922_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1595_ (.Y(_0927_),
    .A(_0922_),
    .B(_0925_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1596_ (.B1(_0898_),
    .VDD(VPWR),
    .Y(_0928_),
    .VSS(VGND),
    .A1(_0896_),
    .A2(_0899_));
 sg13g2_nand2_1 _1597_ (.Y(_0929_),
    .A(net411),
    .B(net466),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _1598_ (.A(net419),
    .B(net414),
    .C(net464),
    .D(net463),
    .X(_0930_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _1599_ (.B(net414),
    .C(net464),
    .A(net419),
    .Y(_0931_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net463));
 sg13g2_a22oi_1 _1600_ (.Y(_0932_),
    .B1(net463),
    .B2(net419),
    .A2(net464),
    .A1(net414),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _1601_ (.A(_0929_),
    .B(_0930_),
    .C(_0932_),
    .X(_0933_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1602_ (.B1(_0929_),
    .VDD(VPWR),
    .Y(_0934_),
    .VSS(VGND),
    .A1(_0930_),
    .A2(_0932_));
 sg13g2_and3_1 _1603_ (.X(_0935_),
    .A(_0928_),
    .B(_0933_),
    .C(_0934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1604_ (.B(_0933_),
    .C(_0934_),
    .A(_0928_),
    .Y(_0936_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _1605_ (.A2(_0934_),
    .A1(_0933_),
    .B1(_0928_),
    .X(_0937_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1606_ (.B(_0936_),
    .C(_0937_),
    .A(_0927_),
    .Y(_0938_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _1607_ (.A2(_0937_),
    .A1(_0936_),
    .B1(_0927_),
    .X(_0939_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _1608_ (.X(_0940_),
    .A(_0921_),
    .B(_0938_),
    .C(_0939_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1609_ (.B(_0938_),
    .C(_0939_),
    .A(_0921_),
    .Y(_0941_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1610_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0938_),
    .A2(_0939_),
    .Y(_0942_),
    .B1(_0921_));
 sg13g2_nor2_1 _1611_ (.A(_0940_),
    .B(_0942_),
    .Y(_0943_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1612_ (.Y(_0944_),
    .A(_0919_),
    .B(_0943_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1613_ (.A(_0944_),
    .B_N(_0915_),
    .Y(_0945_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1614_ (.Y(_0946_),
    .A(_0915_),
    .B(_0944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1615_ (.Y(_0947_),
    .A(_0912_),
    .B(_0946_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1616_ (.Y(_0076_),
    .A(_0914_),
    .B(_0947_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1617_ (.B1(_0946_),
    .VDD(VPWR),
    .Y(_0948_),
    .VSS(VGND),
    .A1(_0912_),
    .A2(_0914_));
 sg13g2_o21ai_1 _1618_ (.B1(_0941_),
    .VDD(VPWR),
    .Y(_0949_),
    .VSS(VGND),
    .A1(_0920_),
    .A2(_0942_));
 sg13g2_o21ai_1 _1619_ (.B1(_0926_),
    .VDD(VPWR),
    .Y(_0950_),
    .VSS(VGND),
    .A1(_0889_),
    .A2(_0924_));
 sg13g2_a22oi_1 _1620_ (.Y(_0951_),
    .B1(net402),
    .B2(net475),
    .A2(net403),
    .A1(net473),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _1621_ (.B(net473),
    .C(net403),
    .A(net474),
    .Y(_0952_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net402));
 sg13g2_nor2b_1 _1622_ (.A(_0951_),
    .B_N(_0952_),
    .Y(_0953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1623_ (.Y(_0954_),
    .A(_0950_),
    .B(_0953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1624_ (.Y(_0955_),
    .A(_0950_),
    .B(_0953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _1625_ (.A2(_0937_),
    .A1(_0927_),
    .B1(_0935_),
    .X(_0956_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1626_ (.Y(_0957_),
    .A(net471),
    .B(net405),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1627_ (.Y(_0958_),
    .A(net467),
    .B(net406),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1628_ (.Y(_0959_),
    .A(net409),
    .B(net467),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1629_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0960_),
    .B(_0958_),
    .A(_0924_));
 sg13g2_and2_1 _1630_ (.A(_0923_),
    .B(_0959_),
    .X(_0961_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1631_ (.Y(_0962_),
    .A(_0923_),
    .B(_0959_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1632_ (.Y(_0963_),
    .A(_0957_),
    .B(_0962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1633_ (.B1(_0931_),
    .VDD(VPWR),
    .Y(_0964_),
    .VSS(VGND),
    .A1(_0929_),
    .A2(_0932_));
 sg13g2_nand2_1 _1634_ (.Y(_0965_),
    .A(net411),
    .B(net465),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _1635_ (.A(net420),
    .B(net414),
    .C(net463),
    .D(net461),
    .X(_0966_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _1636_ (.B(net415),
    .C(net462),
    .A(net419),
    .Y(_0967_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net461));
 sg13g2_a22oi_1 _1637_ (.Y(_0968_),
    .B1(net461),
    .B2(net419),
    .A2(net462),
    .A1(net415),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _1638_ (.A(_0965_),
    .B(_0966_),
    .C(_0968_),
    .X(_0969_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1639_ (.B1(_0965_),
    .VDD(VPWR),
    .Y(_0970_),
    .VSS(VGND),
    .A1(_0966_),
    .A2(_0968_));
 sg13g2_and3_1 _1640_ (.X(_0971_),
    .A(_0964_),
    .B(_0969_),
    .C(_0970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1641_ (.B(_0969_),
    .C(_0970_),
    .A(_0964_),
    .Y(_0972_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1642_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0969_),
    .A2(_0970_),
    .Y(_0973_),
    .B1(_0964_));
 sg13g2_or3_1 _1643_ (.A(_0963_),
    .B(_0971_),
    .C(_0973_),
    .X(_0974_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1644_ (.B1(_0963_),
    .VDD(VPWR),
    .Y(_0975_),
    .VSS(VGND),
    .A1(_0971_),
    .A2(_0973_));
 sg13g2_and3_1 _1645_ (.X(_0976_),
    .A(_0956_),
    .B(_0974_),
    .C(_0975_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1646_ (.B(_0974_),
    .C(_0975_),
    .A(_0956_),
    .Y(_0977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1647_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0974_),
    .A2(_0975_),
    .Y(_0978_),
    .B1(_0956_));
 sg13g2_or3_1 _1648_ (.A(_0955_),
    .B(_0976_),
    .C(_0978_),
    .X(_0979_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1649_ (.B1(_0955_),
    .VDD(VPWR),
    .Y(_0980_),
    .VSS(VGND),
    .A1(_0976_),
    .A2(_0978_));
 sg13g2_and3_1 _1650_ (.X(_0981_),
    .A(_0949_),
    .B(_0979_),
    .C(_0980_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1651_ (.B(_0979_),
    .C(_0980_),
    .A(_0949_),
    .Y(_0982_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1652_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0979_),
    .A2(_0980_),
    .Y(_0983_),
    .B1(_0949_));
 sg13g2_or3_1 _1653_ (.A(_0918_),
    .B(_0981_),
    .C(_0983_),
    .X(_0984_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1654_ (.B1(_0918_),
    .VDD(VPWR),
    .Y(_0985_),
    .VSS(VGND),
    .A1(_0981_),
    .A2(_0983_));
 sg13g2_and3_1 _1655_ (.X(_0986_),
    .A(_0945_),
    .B(_0984_),
    .C(_0985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1656_ (.B(_0984_),
    .C(_0985_),
    .A(_0945_),
    .Y(_0987_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1657_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0984_),
    .A2(_0985_),
    .Y(_0988_),
    .B1(_0945_));
 sg13g2_nor2_1 _1658_ (.A(_0986_),
    .B(_0988_),
    .Y(_0989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1659_ (.Y(_0077_),
    .A(_0948_),
    .B(_0989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1660_ (.B1(_0977_),
    .VDD(VPWR),
    .Y(_0990_),
    .VSS(VGND),
    .A1(_0955_),
    .A2(_0978_));
 sg13g2_o21ai_1 _1661_ (.B1(_0960_),
    .VDD(VPWR),
    .Y(_0991_),
    .VSS(VGND),
    .A1(_0957_),
    .A2(_0961_));
 sg13g2_nand2_1 _1662_ (.Y(_0992_),
    .A(net475),
    .B(net494),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1663_ (.Y(_0993_),
    .A(net471),
    .B(net401),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _1664_ (.A(net471),
    .B(net473),
    .C(net403),
    .D(net401),
    .X(_0994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1665_ (.Y(_0995_),
    .B1(net401),
    .B2(net473),
    .A2(net404),
    .A1(net471),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1666_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0996_),
    .B(_0995_),
    .A(_0994_));
 sg13g2_nor2_1 _1667_ (.A(_0992_),
    .B(_0996_),
    .Y(_0997_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1668_ (.B(_0996_),
    .A(_0992_),
    .X(_0998_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1669_ (.Y(_0999_),
    .A(_0991_),
    .B(_0998_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1670_ (.Y(_1000_),
    .A(_0991_),
    .B(_0998_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1671_ (.Y(_1001_),
    .A(_0952_),
    .B(_1000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1672_ (.B1(_0972_),
    .VDD(VPWR),
    .Y(_1002_),
    .VSS(VGND),
    .A1(_0963_),
    .A2(_0973_));
 sg13g2_nand2_1 _1673_ (.Y(_1003_),
    .A(net469),
    .B(net405),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _1674_ (.Y(_1004_),
    .A(net407),
    .B(net465),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1675_ (.Y(_1005_),
    .A(net409),
    .B(net465),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1676_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1006_),
    .B(_1004_),
    .A(_0959_));
 sg13g2_xnor2_1 _1677_ (.Y(_1007_),
    .A(_0958_),
    .B(_1005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1678_ (.Y(_1008_),
    .A(_1003_),
    .B(_1007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1679_ (.B1(_0967_),
    .VDD(VPWR),
    .Y(_1009_),
    .VSS(VGND),
    .A1(_0965_),
    .A2(_0968_));
 sg13g2_nand2_1 _1680_ (.Y(_1010_),
    .A(net411),
    .B(net462),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _1681_ (.A(net420),
    .B(net414),
    .C(net459),
    .D(net498),
    .X(_1011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _1682_ (.B(net415),
    .C(net459),
    .A(net420),
    .Y(_1012_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net498));
 sg13g2_a22oi_1 _1683_ (.Y(_1013_),
    .B1(net498),
    .B2(net420),
    .A2(net459),
    .A1(net414),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _1684_ (.A(_1010_),
    .B(_1011_),
    .C(_1013_),
    .X(_1014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1685_ (.B1(_1010_),
    .VDD(VPWR),
    .Y(_1015_),
    .VSS(VGND),
    .A1(_1011_),
    .A2(_1013_));
 sg13g2_and3_1 _1686_ (.X(_1016_),
    .A(_1009_),
    .B(_1014_),
    .C(_1015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1687_ (.B(_1014_),
    .C(_1015_),
    .A(_1009_),
    .Y(_1017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1688_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1014_),
    .A2(_1015_),
    .Y(_1018_),
    .B1(_1009_));
 sg13g2_or3_1 _1689_ (.A(_1008_),
    .B(_1016_),
    .C(_1018_),
    .X(_1019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1690_ (.B1(_1008_),
    .VDD(VPWR),
    .Y(_1020_),
    .VSS(VGND),
    .A1(_1016_),
    .A2(_1018_));
 sg13g2_and3_1 _1691_ (.X(_1021_),
    .A(_1002_),
    .B(_1019_),
    .C(_1020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1692_ (.B(_1019_),
    .C(_1020_),
    .A(_1002_),
    .Y(_1022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1693_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1019_),
    .A2(_1020_),
    .Y(_1023_),
    .B1(_1002_));
 sg13g2_or3_1 _1694_ (.A(_1001_),
    .B(_1021_),
    .C(_1023_),
    .X(_1024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1695_ (.B1(_1001_),
    .VDD(VPWR),
    .Y(_1025_),
    .VSS(VGND),
    .A1(_1021_),
    .A2(_1023_));
 sg13g2_and3_1 _1696_ (.X(_1026_),
    .A(_0990_),
    .B(_1024_),
    .C(_1025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1697_ (.B(_1024_),
    .C(_1025_),
    .A(_0990_),
    .Y(_1027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1698_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1024_),
    .A2(_1025_),
    .Y(_1028_),
    .B1(_0990_));
 sg13g2_or3_1 _1699_ (.A(_0954_),
    .B(_1026_),
    .C(_1028_),
    .X(_1029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1700_ (.B1(_0954_),
    .VDD(VPWR),
    .Y(_1030_),
    .VSS(VGND),
    .A1(_1026_),
    .A2(_1028_));
 sg13g2_o21ai_1 _1701_ (.B1(_0982_),
    .VDD(VPWR),
    .Y(_1031_),
    .VSS(VGND),
    .A1(_0918_),
    .A2(_0983_));
 sg13g2_nand3_1 _1702_ (.B(_1030_),
    .C(_1031_),
    .A(_1029_),
    .Y(_1032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _1703_ (.A2(_1030_),
    .A1(_1029_),
    .B1(_1031_),
    .X(_1033_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1704_ (.A(_1032_),
    .B(_1033_),
    .X(_1034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1705_ (.B1(_0987_),
    .VDD(VPWR),
    .Y(_1035_),
    .VSS(VGND),
    .A1(_0948_),
    .A2(_0988_));
 sg13g2_nand2_1 _1706_ (.Y(_1036_),
    .A(_1034_),
    .B(_1035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1707_ (.B(_1035_),
    .A(_1034_),
    .X(_0078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1708_ (.Y(_1037_),
    .A(_1032_),
    .B(_1036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1709_ (.B1(_1027_),
    .VDD(VPWR),
    .Y(_1038_),
    .VSS(VGND),
    .A1(_0954_),
    .A2(_1028_));
 sg13g2_o21ai_1 _1710_ (.B1(_0999_),
    .VDD(VPWR),
    .Y(_1039_),
    .VSS(VGND),
    .A1(_0952_),
    .A2(_1000_));
 sg13g2_o21ai_1 _1711_ (.B1(_1022_),
    .VDD(VPWR),
    .Y(_1040_),
    .VSS(VGND),
    .A1(_1001_),
    .A2(_1023_));
 sg13g2_nor2_1 _1712_ (.A(_0994_),
    .B(_0997_),
    .Y(_1041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1713_ (.B1(_1006_),
    .VDD(VPWR),
    .Y(_1042_),
    .VSS(VGND),
    .A1(_1003_),
    .A2(_1007_));
 sg13g2_nand2_1 _1714_ (.Y(_1043_),
    .A(net473),
    .B(net494),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1715_ (.Y(_1044_),
    .A(net469),
    .B(net401),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1716_ (.Y(_1045_),
    .A(net469),
    .B(net404),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1717_ (.B(_1045_),
    .A(_0993_),
    .X(_1046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1718_ (.Y(_1047_),
    .B(_1046_),
    .A_N(_1043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1719_ (.Y(_1048_),
    .A(_1043_),
    .B(_1046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1720_ (.Y(_1049_),
    .A(_1042_),
    .B(_1048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1721_ (.A(_1041_),
    .B(_1049_),
    .Y(_1050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1722_ (.Y(_1051_),
    .A(_1041_),
    .B(_1049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1723_ (.B1(_1017_),
    .VDD(VPWR),
    .Y(_1052_),
    .VSS(VGND),
    .A1(_1008_),
    .A2(_1018_));
 sg13g2_nand2_1 _1724_ (.Y(_1053_),
    .A(net467),
    .B(\DP_2.matrix[41] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1725_ (.Y(_1054_),
    .A(net409),
    .B(\DP_1.matrix[42] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1726_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1055_),
    .B(_1054_),
    .A(_1004_));
 sg13g2_and2_1 _1727_ (.A(_1004_),
    .B(_1054_),
    .X(_1056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1728_ (.Y(_1057_),
    .A(_1004_),
    .B(_1054_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1729_ (.Y(_1058_),
    .A(_1053_),
    .B(_1057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1730_ (.B1(_1012_),
    .VDD(VPWR),
    .Y(_1059_),
    .VSS(VGND),
    .A1(_1010_),
    .A2(_1013_));
 sg13g2_nand2_1 _1731_ (.Y(_1060_),
    .A(net410),
    .B(net498),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _1732_ (.A(net414),
    .B(net410),
    .C(net459),
    .D(net498),
    .X(_1061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1733_ (.Y(_1062_),
    .B1(net498),
    .B2(net415),
    .A2(net459),
    .A1(net411),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1734_ (.A(_1061_),
    .B(_1062_),
    .Y(_1063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1735_ (.Y(_1064_),
    .A(_1059_),
    .B(_1063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1736_ (.Y(_1065_),
    .A(_1059_),
    .B(_1063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1737_ (.B(_1065_),
    .A(_1058_),
    .X(_1066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1738_ (.Y(_1067_),
    .A(_1052_),
    .B(_1066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1739_ (.Y(_1068_),
    .A(_1052_),
    .B(_1066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1740_ (.B(_1068_),
    .A(_1051_),
    .X(_1069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1741_ (.Y(_1070_),
    .A(_1040_),
    .B(_1069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1742_ (.Y(_1071_),
    .A(_1040_),
    .B(_1069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1743_ (.Y(_1072_),
    .B(_1039_),
    .A_N(_1071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1744_ (.Y(_1073_),
    .A(_1039_),
    .B(_1071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1745_ (.A(_1038_),
    .B(_1073_),
    .Y(_1074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1746_ (.Y(_1075_),
    .A(_1038_),
    .B(_1073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1747_ (.Y(_1076_),
    .A(_1038_),
    .B(_1073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _1748_ (.VDD(VPWR),
    .Y(_1077_),
    .A(_1076_),
    .VSS(VGND));
 sg13g2_xnor2_1 _1749_ (.Y(_0079_),
    .A(_1037_),
    .B(_1076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1750_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1042_),
    .A2(_1048_),
    .Y(_1078_),
    .B1(_1050_));
 sg13g2_o21ai_1 _1751_ (.B1(_1067_),
    .VDD(VPWR),
    .Y(_1079_),
    .VSS(VGND),
    .A1(_1051_),
    .A2(_1068_));
 sg13g2_o21ai_1 _1752_ (.B1(_1047_),
    .VDD(VPWR),
    .Y(_1080_),
    .VSS(VGND),
    .A1(_0993_),
    .A2(_1045_));
 sg13g2_o21ai_1 _1753_ (.B1(_1055_),
    .VDD(VPWR),
    .Y(_1081_),
    .VSS(VGND),
    .A1(_1053_),
    .A2(_1056_));
 sg13g2_nand2_1 _1754_ (.Y(_1082_),
    .A(net471),
    .B(net494),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1755_ (.Y(_1083_),
    .A(net467),
    .B(net401),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1756_ (.Y(_1084_),
    .A(net467),
    .B(net404),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1757_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1085_),
    .B(_1083_),
    .A(_1045_));
 sg13g2_xnor2_1 _1758_ (.Y(_1086_),
    .A(_1044_),
    .B(_1084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1759_ (.B(_1086_),
    .A(_1082_),
    .X(_1087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1760_ (.Y(_1088_),
    .A(_1081_),
    .B(_1087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1761_ (.A(_1088_),
    .B_N(_1080_),
    .Y(_1089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1762_ (.B(_1088_),
    .A(_1080_),
    .X(_1090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1763_ (.B1(_1064_),
    .VDD(VPWR),
    .Y(_1091_),
    .VSS(VGND),
    .A1(_1058_),
    .A2(_1065_));
 sg13g2_a21oi_1 _1764_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net415),
    .A2(net459),
    .Y(_1092_),
    .B1(_1060_));
 sg13g2_nand2_1 _1765_ (.Y(_1093_),
    .A(net465),
    .B(\DP_2.matrix[41] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1766_ (.Y(_1094_),
    .A(net406),
    .B(net460),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _1767_ (.A(net408),
    .B(net407),
    .C(net463),
    .D(net460),
    .X(_1095_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1768_ (.Y(_1096_),
    .B1(net460),
    .B2(net409),
    .A2(\DP_1.matrix[42] ),
    .A1(net407),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _1769_ (.A(_1093_),
    .B(_1095_),
    .C(_1096_),
    .Y(_1097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1770_ (.B1(_1093_),
    .VDD(VPWR),
    .Y(_1098_),
    .VSS(VGND),
    .A1(_1095_),
    .A2(_1096_));
 sg13g2_nor2b_1 _1771_ (.A(_1097_),
    .B_N(_1098_),
    .Y(_1099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1772_ (.Y(_1100_),
    .A(_1092_),
    .B(_1099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1773_ (.Y(_1101_),
    .B(_1091_),
    .A_N(_1100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1774_ (.B(_1100_),
    .A(_1091_),
    .X(_1102_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1775_ (.B(_1102_),
    .A(_1090_),
    .X(_1103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1776_ (.Y(_1104_),
    .A(_1079_),
    .B(_1103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1777_ (.B(_1103_),
    .A(_1079_),
    .X(_1105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1778_ (.Y(_1106_),
    .B(_1105_),
    .A_N(_1078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1779_ (.B(_1105_),
    .A(_1078_),
    .X(_1107_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1780_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1070_),
    .A2(_1072_),
    .Y(_1108_),
    .B1(_1107_));
 sg13g2_nand3_1 _1781_ (.B(_1072_),
    .C(_1107_),
    .A(_1070_),
    .Y(_1109_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1782_ (.Y(_1110_),
    .B(_1109_),
    .A_N(_1108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1783_ (.B(_1035_),
    .C(_1077_),
    .A(_1034_),
    .Y(_1111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1784_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1032_),
    .A2(_1075_),
    .Y(_1112_),
    .B1(_1074_));
 sg13g2_nor2b_1 _1785_ (.A(_1112_),
    .B_N(_1111_),
    .Y(_1113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1786_ (.A(_1110_),
    .B(_1113_),
    .Y(_1114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1787_ (.B(_1113_),
    .A(_1110_),
    .X(_0070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _1788_ (.A2(_1087_),
    .A1(_1081_),
    .B1(_1089_),
    .X(_1115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1789_ (.B1(_1101_),
    .VDD(VPWR),
    .Y(_1116_),
    .VSS(VGND),
    .A1(_1090_),
    .A2(_1102_));
 sg13g2_a21o_2 _1790_ (.A2(_1099_),
    .A1(_1092_),
    .B1(_1061_),
    .X(_1117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1791_ (.Y(_1118_),
    .A(net405),
    .B(net462),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1792_ (.Y(_1119_),
    .A(net408),
    .B(net499),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1793_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1120_),
    .B(_1119_),
    .A(_1094_));
 sg13g2_xnor2_1 _1794_ (.Y(_1121_),
    .A(_1094_),
    .B(_1119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1795_ (.B(_1121_),
    .A(_1118_),
    .X(_1122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1796_ (.A(_1117_),
    .B(_1122_),
    .X(_1123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1797_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1124_),
    .B(_1122_),
    .A(_1117_));
 sg13g2_xnor2_1 _1798_ (.Y(_1125_),
    .A(_1117_),
    .B(_1122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1799_ (.B1(_1085_),
    .VDD(VPWR),
    .Y(_1126_),
    .VSS(VGND),
    .A1(_1082_),
    .A2(_1086_));
 sg13g2_or2_1 _1800_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1127_),
    .B(_1097_),
    .A(_1095_));
 sg13g2_nand2_1 _1801_ (.Y(_1128_),
    .A(net469),
    .B(net494),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1802_ (.Y(_1129_),
    .A(net465),
    .B(net403),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1803_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1130_),
    .B(_1129_),
    .A(_1083_));
 sg13g2_xnor2_1 _1804_ (.Y(_1131_),
    .A(_1083_),
    .B(_1129_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1805_ (.B(_1131_),
    .A(_1128_),
    .X(_1132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1806_ (.Y(_1133_),
    .A(_1127_),
    .B(_1132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1807_ (.A(_1133_),
    .B_N(_1126_),
    .Y(_1134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1808_ (.Y(_1135_),
    .A(_1126_),
    .B(_1133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1809_ (.Y(_1136_),
    .A(_1125_),
    .B(_1135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1810_ (.Y(_1137_),
    .A(_1116_),
    .B(_1136_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1811_ (.A(_1137_),
    .B_N(_1115_),
    .Y(_1138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1812_ (.B(_1137_),
    .A(_1115_),
    .X(_1139_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _1813_ (.B(_1106_),
    .C(_1139_),
    .A(_1104_),
    .Y(_1140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1814_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1104_),
    .A2(_1106_),
    .Y(_1141_),
    .B1(_1139_));
 sg13g2_inv_1 _1815_ (.VDD(VPWR),
    .Y(_1142_),
    .A(_1141_),
    .VSS(VGND));
 sg13g2_nand2_1 _1816_ (.Y(_1143_),
    .A(_1140_),
    .B(_1142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1817_ (.A(_1108_),
    .B(_1114_),
    .Y(_1144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1818_ (.B(_1144_),
    .A(_1143_),
    .X(_0071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _1819_ (.A2(_1132_),
    .A1(_1127_),
    .B1(_1134_),
    .X(_1145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1820_ (.Y(_1146_),
    .B1(net499),
    .B2(net406),
    .A2(net460),
    .A1(net405),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _1821_ (.Y(_1147_),
    .A(net405),
    .B(net498),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1822_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1148_),
    .B(_1147_),
    .A(_1094_));
 sg13g2_nand2b_1 _1823_ (.Y(_1149_),
    .B(_1148_),
    .A_N(_1146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1824_ (.B1(_1130_),
    .VDD(VPWR),
    .Y(_1150_),
    .VSS(VGND),
    .A1(_1128_),
    .A2(_1131_));
 sg13g2_o21ai_1 _1825_ (.B1(_1120_),
    .VDD(VPWR),
    .Y(_1151_),
    .VSS(VGND),
    .A1(_1118_),
    .A2(_1121_));
 sg13g2_nand2_1 _1826_ (.Y(_1152_),
    .A(net467),
    .B(net494),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1827_ (.Y(_1153_),
    .A(net462),
    .B(net401),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _1828_ (.A(net465),
    .B(net462),
    .C(net403),
    .D(net401),
    .X(_1154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1829_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1155_),
    .B(_1153_),
    .A(_1129_));
 sg13g2_a22oi_1 _1830_ (.Y(_1156_),
    .B1(net401),
    .B2(net465),
    .A2(net403),
    .A1(net462),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1831_ (.A(_1154_),
    .B(_1156_),
    .Y(_1157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1832_ (.Y(_1158_),
    .A(_1152_),
    .B(_1157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1833_ (.Y(_1159_),
    .A(_1151_),
    .B(_1158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1834_ (.A(_1159_),
    .B_N(_1150_),
    .Y(_1160_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1835_ (.B(_1159_),
    .A(_1150_),
    .X(_1161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1836_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1162_),
    .B(_1161_),
    .A(_1149_));
 sg13g2_xor2_1 _1837_ (.B(_1161_),
    .A(_1149_),
    .X(_1163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1838_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1124_),
    .A2(_1135_),
    .Y(_1164_),
    .B1(_1123_));
 sg13g2_nor2b_1 _1839_ (.A(_1164_),
    .B_N(_1163_),
    .Y(_1165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1840_ (.B(_1164_),
    .A(_1163_),
    .X(_1166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1841_ (.A(_1166_),
    .B_N(_1145_),
    .Y(_1167_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1842_ (.B(_1166_),
    .A(_1145_),
    .X(_1168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1843_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1116_),
    .A2(_1136_),
    .Y(_1169_),
    .B1(_1138_));
 sg13g2_nor2_1 _1844_ (.A(_1168_),
    .B(_1169_),
    .Y(_1170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1845_ (.B(_1169_),
    .A(_1168_),
    .X(_1171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1846_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1108_),
    .A2(_1140_),
    .Y(_1172_),
    .B1(_1141_));
 sg13g2_nor2b_1 _1847_ (.A(_1112_),
    .B_N(_1172_),
    .Y(_1173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1848_ (.Y(_1174_),
    .A(_1109_),
    .B(_1140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _1849_ (.Y(_1175_),
    .B1(_1174_),
    .B2(_1142_),
    .A2(_1173_),
    .A1(_1111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1850_ (.B(_1175_),
    .A(_1171_),
    .X(_0072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _1851_ (.A2(_1158_),
    .A1(_1151_),
    .B1(_1160_),
    .X(_1176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1852_ (.B1(_1155_),
    .VDD(VPWR),
    .Y(_1177_),
    .VSS(VGND),
    .A1(_1152_),
    .A2(_1156_));
 sg13g2_nand2_1 _1853_ (.Y(_1178_),
    .A(net465),
    .B(net494),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1854_ (.Y(_1179_),
    .A(net459),
    .B(net402),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1855_ (.Y(_1180_),
    .A(net403),
    .B(net460),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1856_ (.B(_1180_),
    .A(_1153_),
    .X(_1181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1857_ (.Y(_1182_),
    .B(_1181_),
    .A_N(_1178_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1858_ (.Y(_1183_),
    .A(_1178_),
    .B(_1181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1859_ (.A(_1148_),
    .B_N(_1183_),
    .Y(_1184_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1860_ (.Y(_1185_),
    .A(_1148_),
    .B(_1183_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1861_ (.Y(_1186_),
    .A(_1177_),
    .B(_1185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1862_ (.A(_1147_),
    .B(_1186_),
    .Y(_1187_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1863_ (.Y(_1188_),
    .A(_1147_),
    .B(_1186_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1864_ (.A(_1162_),
    .B(_1188_),
    .Y(_1189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1865_ (.B(_1188_),
    .A(_1162_),
    .X(_1190_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1866_ (.B(_1190_),
    .A(_1176_),
    .X(_1191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1867_ (.B1(_1191_),
    .VDD(VPWR),
    .Y(_1192_),
    .VSS(VGND),
    .A1(_1165_),
    .A2(_1167_));
 sg13g2_or3_1 _1868_ (.A(_1165_),
    .B(_1167_),
    .C(_1191_),
    .X(_1193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1869_ (.A(_1192_),
    .B(_1193_),
    .X(_1194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1870_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1171_),
    .A2(_1175_),
    .Y(_1195_),
    .B1(_1170_));
 sg13g2_xnor2_1 _1871_ (.Y(_0073_),
    .A(_1194_),
    .B(_1195_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1872_ (.Y(_1196_),
    .A(_1171_),
    .B(_1194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1873_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1142_),
    .C1(_1196_),
    .B1(_1174_),
    .A1(_1111_),
    .Y(_1197_),
    .A2(_1173_));
 sg13g2_nand2_1 _1874_ (.Y(_1198_),
    .A(_1170_),
    .B(_1193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1875_ (.Y(_1199_),
    .A(_1192_),
    .B(_1198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1876_ (.A(_1197_),
    .B(_1199_),
    .Y(_1200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1877_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1176_),
    .A2(_1190_),
    .Y(_1201_),
    .B1(_1189_));
 sg13g2_a21o_1 _1878_ (.A2(_1185_),
    .A1(_1177_),
    .B1(_1184_),
    .X(_1202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1879_ (.B1(_1182_),
    .VDD(VPWR),
    .Y(_1203_),
    .VSS(VGND),
    .A1(_1153_),
    .A2(_1180_));
 sg13g2_nand2_1 _1880_ (.Y(_1204_),
    .A(net462),
    .B(net494),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1881_ (.Y(_1205_),
    .A(net402),
    .B(net499),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1882_ (.Y(_1206_),
    .A(net404),
    .B(net498),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1883_ (.B(_1206_),
    .A(_1179_),
    .X(_1207_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1884_ (.Y(_1208_),
    .B(_1207_),
    .A_N(_1204_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1885_ (.Y(_1209_),
    .A(_1204_),
    .B(_1207_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1886_ (.Y(_1210_),
    .A(_1203_),
    .B(_1209_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1887_ (.B(_1209_),
    .A(_1203_),
    .X(_1211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1888_ (.Y(_1212_),
    .A(_1187_),
    .B(_1211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _1889_ (.A(_1212_),
    .B_N(_1202_),
    .Y(_1213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1890_ (.B(_1212_),
    .A(_1202_),
    .X(_1214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1891_ (.B(_1214_),
    .A(_1201_),
    .X(_1215_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1892_ (.B1(_1215_),
    .VDD(VPWR),
    .Y(_1216_),
    .VSS(VGND),
    .A1(_1197_),
    .A2(_1199_));
 sg13g2_xnor2_1 _1893_ (.Y(_0074_),
    .A(_1200_),
    .B(_1215_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1894_ (.B1(_1216_),
    .VDD(VPWR),
    .Y(_1217_),
    .VSS(VGND),
    .A1(_1201_),
    .A2(_1214_));
 sg13g2_a21oi_1 _1895_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1187_),
    .A2(_1211_),
    .Y(_1218_),
    .B1(_1213_));
 sg13g2_o21ai_1 _1896_ (.B1(_1208_),
    .VDD(VPWR),
    .Y(_1219_),
    .VSS(VGND),
    .A1(_1179_),
    .A2(_1206_));
 sg13g2_nand2_1 _1897_ (.Y(_1220_),
    .A(net460),
    .B(net494),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1898_ (.B(_1220_),
    .A(_1205_),
    .X(_1221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1899_ (.Y(_1222_),
    .A(_1219_),
    .B(_1221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1900_ (.Y(_1223_),
    .A(_1210_),
    .B(_1222_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1901_ (.Y(_1224_),
    .A(_1218_),
    .B(_1223_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1902_ (.Y(_0075_),
    .A(_1217_),
    .B(_1224_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1903_ (.A(net457),
    .B(net397),
    .X(_0032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1904_ (.A(net492),
    .B(net437),
    .X(_0037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1905_ (.Y(_1225_),
    .A(net235),
    .B(net161),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1906_ (.Y(_1226_),
    .A(\mac1.sum_lvl2_ff[20] ),
    .B(\mac1.sum_lvl2_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1907_ (.A(\mac1.sum_lvl2_ff[20] ),
    .B(\mac1.sum_lvl2_ff[1] ),
    .Y(_1227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1908_ (.B(\mac1.sum_lvl2_ff[1] ),
    .A(\mac1.sum_lvl2_ff[20] ),
    .X(_1228_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1909_ (.Y(_0007_),
    .A(_1225_),
    .B(_1228_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1910_ (.B1(_1226_),
    .VDD(VPWR),
    .Y(_1229_),
    .VSS(VGND),
    .A1(_1225_),
    .A2(_1227_));
 sg13g2_and2_1 _1911_ (.A(\mac1.sum_lvl2_ff[21] ),
    .B(\mac1.sum_lvl2_ff[2] ),
    .X(_1230_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1912_ (.B(net254),
    .A(\mac1.sum_lvl2_ff[21] ),
    .X(_1231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1913_ (.B(net255),
    .A(_1229_),
    .X(_0008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1914_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1229_),
    .A2(_1231_),
    .Y(_1232_),
    .B1(_1230_));
 sg13g2_nand2_1 _1915_ (.Y(_1233_),
    .A(\mac1.sum_lvl2_ff[22] ),
    .B(net243),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1916_ (.Y(_1234_),
    .A(\mac1.sum_lvl2_ff[22] ),
    .B(net243),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1917_ (.B(net244),
    .A(_1232_),
    .X(_0009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1918_ (.B1(_1233_),
    .VDD(VPWR),
    .Y(_1235_),
    .VSS(VGND),
    .A1(_1232_),
    .A2(_1234_));
 sg13g2_and2_1 _1919_ (.A(\mac1.sum_lvl2_ff[23] ),
    .B(\mac1.sum_lvl2_ff[4] ),
    .X(_1236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1920_ (.B(net265),
    .A(\mac1.sum_lvl2_ff[23] ),
    .X(_1237_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1921_ (.B(net266),
    .A(_1235_),
    .X(_0010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1922_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1235_),
    .A2(_1237_),
    .Y(_1238_),
    .B1(_1236_));
 sg13g2_nor2_1 _1923_ (.A(\mac1.sum_lvl2_ff[24] ),
    .B(net257),
    .Y(_1239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1924_ (.B(net257),
    .A(\mac1.sum_lvl2_ff[24] ),
    .X(_1240_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1925_ (.Y(_0011_),
    .A(_1238_),
    .B(net258),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1926_ (.A(\mac1.sum_lvl2_ff[25] ),
    .B(\mac1.sum_lvl2_ff[6] ),
    .X(_1241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1927_ (.Y(_1242_),
    .A(\mac1.sum_lvl2_ff[25] ),
    .B(net296),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _1928_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1237_),
    .C1(_1236_),
    .B1(_1235_),
    .A1(\mac1.sum_lvl2_ff[24] ),
    .Y(_1243_),
    .A2(net257));
 sg13g2_nor3_2 _1929_ (.A(_1239_),
    .B(net297),
    .C(_1243_),
    .Y(_1244_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1930_ (.B1(net297),
    .VDD(VPWR),
    .Y(_1245_),
    .VSS(VGND),
    .A1(_1239_),
    .A2(_1243_));
 sg13g2_nor2b_2 _1931_ (.A(_1244_),
    .B_N(net298),
    .Y(_0012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1932_ (.Y(_1246_),
    .A(net283),
    .B(\mac1.sum_lvl2_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1933_ (.B(net304),
    .A(\mac1.sum_lvl2_ff[26] ),
    .X(_1247_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1934_ (.B1(_1247_),
    .VDD(VPWR),
    .Y(_1248_),
    .VSS(VGND),
    .A1(_1241_),
    .A2(_1244_));
 sg13g2_or3_1 _1935_ (.A(_1241_),
    .B(_1244_),
    .C(net305),
    .X(_1249_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1936_ (.A(_1248_),
    .B(_1249_),
    .X(_0013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1937_ (.A(\mac1.sum_lvl2_ff[27] ),
    .B(\mac1.sum_lvl2_ff[8] ),
    .X(_1250_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1938_ (.Y(_1251_),
    .A(\mac1.sum_lvl2_ff[27] ),
    .B(\mac1.sum_lvl2_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _1939_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_1251_),
    .Y(_1252_),
    .A2(_1248_),
    .A1(net284));
 sg13g2_nand3_1 _1940_ (.B(_1248_),
    .C(_1251_),
    .A(net284),
    .Y(_1253_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _1941_ (.A(_1252_),
    .B_N(_1253_),
    .Y(_0014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1942_ (.A(_1250_),
    .B(_1252_),
    .Y(_1254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1943_ (.Y(_1255_),
    .A(\mac1.sum_lvl2_ff[28] ),
    .B(\mac1.sum_lvl2_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1944_ (.B(net294),
    .A(\mac1.sum_lvl2_ff[28] ),
    .X(_1256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1945_ (.B1(_1256_),
    .VDD(VPWR),
    .Y(_1257_),
    .VSS(VGND),
    .A1(_1250_),
    .A2(_1252_));
 sg13g2_xnor2_1 _1946_ (.Y(_0015_),
    .A(_1254_),
    .B(net295),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1947_ (.Y(_1258_),
    .A(_1255_),
    .B(_1257_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1948_ (.Y(_1259_),
    .A(net301),
    .B(\mac1.sum_lvl2_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1949_ (.B(\mac1.sum_lvl2_ff[10] ),
    .A(net301),
    .X(_1260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1950_ (.Y(_1261_),
    .A(_1258_),
    .B(_1260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1951_ (.B(net302),
    .A(_1258_),
    .X(_0001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1952_ (.A(\mac1.sum_lvl2_ff[30] ),
    .B(\mac1.sum_lvl2_ff[11] ),
    .Y(_1262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1953_ (.Y(_1263_),
    .A(\mac1.sum_lvl2_ff[30] ),
    .B(\mac1.sum_lvl2_ff[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _1954_ (.Y(_1264_),
    .B(_1263_),
    .A_N(_1262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1955_ (.Y(_1265_),
    .A(_1259_),
    .B(_1261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1956_ (.Y(_0002_),
    .A(_1264_),
    .B(_1265_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1957_ (.Y(_1266_),
    .A(net278),
    .B(\mac1.sum_lvl2_ff[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1958_ (.B(\mac1.sum_lvl2_ff[12] ),
    .A(\mac1.sum_lvl2_ff[31] ),
    .X(_1267_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1959_ (.B1(_1263_),
    .VDD(VPWR),
    .Y(_1268_),
    .VSS(VGND),
    .A1(_1259_),
    .A2(_1262_));
 sg13g2_nand3b_1 _1960_ (.B(_1263_),
    .C(_1260_),
    .Y(_1269_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1262_));
 sg13g2_a21oi_1 _1961_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1255_),
    .A2(_1257_),
    .Y(_1270_),
    .B1(_1269_));
 sg13g2_o21ai_1 _1962_ (.B1(_1267_),
    .VDD(VPWR),
    .Y(_1271_),
    .VSS(VGND),
    .A1(_1268_),
    .A2(_1270_));
 sg13g2_or3_1 _1963_ (.A(_1267_),
    .B(_1268_),
    .C(_1270_),
    .X(_1272_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1964_ (.A(_1271_),
    .B(_1272_),
    .X(_0003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1965_ (.Y(_1273_),
    .A(\mac1.sum_lvl2_ff[32] ),
    .B(\mac1.sum_lvl2_ff[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1966_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net279),
    .A2(_1271_),
    .Y(_1274_),
    .B1(_1273_));
 sg13g2_nand3_1 _1967_ (.B(_1271_),
    .C(_1273_),
    .A(net279),
    .Y(_1275_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _1968_ (.A(_1274_),
    .B_N(net280),
    .Y(_0004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1969_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mac1.sum_lvl2_ff[32] ),
    .A2(\mac1.sum_lvl2_ff[13] ),
    .Y(_1276_),
    .B1(_1274_));
 sg13g2_nand2_1 _1970_ (.Y(_1277_),
    .A(\mac1.sum_lvl2_ff[33] ),
    .B(\mac1.sum_lvl2_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1971_ (.A(\mac1.sum_lvl2_ff[33] ),
    .B(\mac1.sum_lvl2_ff[14] ),
    .Y(_1278_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1972_ (.B(net171),
    .A(\mac1.sum_lvl2_ff[33] ),
    .X(_1279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1973_ (.Y(_0005_),
    .A(_1276_),
    .B(net172),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1974_ (.B1(_1277_),
    .VDD(VPWR),
    .Y(_1280_),
    .VSS(VGND),
    .A1(_1276_),
    .A2(_1278_));
 sg13g2_xnor2_1 _1975_ (.Y(_1281_),
    .A(net168),
    .B(\mac1.sum_lvl2_ff[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1976_ (.Y(_0006_),
    .A(_1280_),
    .B(net169),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1977_ (.B(net161),
    .A(\mac1.sum_lvl2_ff[19] ),
    .X(_0000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1978_ (.Y(_1282_),
    .A(net166),
    .B(net153),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1979_ (.Y(_1283_),
    .A(\mac1.sum_lvl3_ff[1] ),
    .B(\mac1.sum_lvl3_ff[21] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1980_ (.A(\mac1.sum_lvl3_ff[1] ),
    .B(\mac1.sum_lvl3_ff[21] ),
    .Y(_1284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1981_ (.B(\mac1.sum_lvl3_ff[21] ),
    .A(\mac1.sum_lvl3_ff[1] ),
    .X(_1285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1982_ (.Y(_0023_),
    .A(_1282_),
    .B(_1285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1983_ (.B1(_1283_),
    .VDD(VPWR),
    .Y(_1286_),
    .VSS(VGND),
    .A1(_1282_),
    .A2(_1284_));
 sg13g2_and2_1 _1984_ (.A(\mac1.sum_lvl3_ff[2] ),
    .B(net174),
    .X(_1287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1985_ (.B(net174),
    .A(\mac1.sum_lvl3_ff[2] ),
    .X(_1288_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1986_ (.B(net175),
    .A(_1286_),
    .X(_0024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1987_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1286_),
    .A2(net175),
    .Y(_1289_),
    .B1(_1287_));
 sg13g2_nand2_1 _1988_ (.Y(_1290_),
    .A(\mac1.sum_lvl3_ff[3] ),
    .B(net200),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1989_ (.Y(_1291_),
    .A(\mac1.sum_lvl3_ff[3] ),
    .B(net200),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1990_ (.B(net201),
    .A(_1289_),
    .X(_0025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _1991_ (.B1(_1290_),
    .VDD(VPWR),
    .Y(_1292_),
    .VSS(VGND),
    .A1(_1289_),
    .A2(net201));
 sg13g2_and2_1 _1992_ (.A(\mac1.sum_lvl3_ff[4] ),
    .B(net217),
    .X(_1293_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1993_ (.B(net217),
    .A(\mac1.sum_lvl3_ff[4] ),
    .X(_1294_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1994_ (.B(net218),
    .A(_1292_),
    .X(_0026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1995_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1292_),
    .A2(_1294_),
    .Y(_1295_),
    .B1(_1293_));
 sg13g2_nor2_1 _1996_ (.A(net178),
    .B(\mac1.sum_lvl3_ff[25] ),
    .Y(_1296_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _1997_ (.B(\mac1.sum_lvl3_ff[25] ),
    .A(net178),
    .X(_1297_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _1998_ (.Y(_0027_),
    .A(_1295_),
    .B(net179),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _1999_ (.A(\mac1.sum_lvl3_ff[6] ),
    .B(net261),
    .X(_1298_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2000_ (.Y(_1299_),
    .A(\mac1.sum_lvl3_ff[6] ),
    .B(net261),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2001_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1294_),
    .C1(_1293_),
    .B1(_1292_),
    .A1(net178),
    .Y(_1300_),
    .A2(\mac1.sum_lvl3_ff[25] ));
 sg13g2_nor3_1 _2002_ (.A(_1296_),
    .B(net262),
    .C(_1300_),
    .Y(_1301_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2003_ (.B1(net262),
    .VDD(VPWR),
    .Y(_1302_),
    .VSS(VGND),
    .A1(_1296_),
    .A2(_1300_));
 sg13g2_nor2b_1 _2004_ (.A(_1301_),
    .B_N(net263),
    .Y(_0028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2005_ (.Y(_1303_),
    .A(\mac1.sum_lvl3_ff[7] ),
    .B(net239),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2006_ (.B(net239),
    .A(net287),
    .X(_1304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2007_ (.B1(_1304_),
    .VDD(VPWR),
    .Y(_1305_),
    .VSS(VGND),
    .A1(_1298_),
    .A2(_1301_));
 sg13g2_or3_1 _2008_ (.A(_1298_),
    .B(_1301_),
    .C(_1304_),
    .X(_1306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2009_ (.A(net288),
    .B(_1306_),
    .X(_0029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2010_ (.A(\mac1.sum_lvl3_ff[8] ),
    .B(\mac1.sum_lvl3_ff[28] ),
    .X(_1307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2011_ (.Y(_1308_),
    .A(\mac1.sum_lvl3_ff[8] ),
    .B(\mac1.sum_lvl3_ff[28] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2012_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net240),
    .A2(_1305_),
    .Y(_1309_),
    .B1(_1308_));
 sg13g2_nand3_1 _2013_ (.B(_1305_),
    .C(_1308_),
    .A(net240),
    .Y(_1310_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2014_ (.A(_1309_),
    .B_N(net241),
    .Y(_0030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2015_ (.A(_1307_),
    .B(_1309_),
    .Y(_1311_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2016_ (.Y(_1312_),
    .A(\mac1.sum_lvl3_ff[9] ),
    .B(net181),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2017_ (.B(net181),
    .A(\mac1.sum_lvl3_ff[9] ),
    .X(_1313_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2018_ (.B1(net182),
    .VDD(VPWR),
    .Y(_1314_),
    .VSS(VGND),
    .A1(_1307_),
    .A2(_1309_));
 sg13g2_xnor2_1 _2019_ (.Y(_0031_),
    .A(_1311_),
    .B(net182),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2020_ (.Y(_1315_),
    .A(_1312_),
    .B(_1314_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2021_ (.Y(_1316_),
    .A(net206),
    .B(\mac1.sum_lvl3_ff[30] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2022_ (.B(net213),
    .A(net206),
    .X(_1317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2023_ (.Y(_1318_),
    .A(_1315_),
    .B(_1317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2024_ (.B(_1317_),
    .A(_1315_),
    .X(_0017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2025_ (.A(\mac1.sum_lvl3_ff[11] ),
    .B(\mac1.sum_lvl3_ff[31] ),
    .Y(_1319_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2026_ (.Y(_1320_),
    .A(\mac1.sum_lvl3_ff[11] ),
    .B(\mac1.sum_lvl3_ff[31] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2027_ (.Y(_1321_),
    .B(_1320_),
    .A_N(_1319_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2028_ (.Y(_1322_),
    .A(net207),
    .B(_1318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2029_ (.Y(_0018_),
    .A(_1321_),
    .B(net208),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2030_ (.Y(_1323_),
    .A(\mac1.sum_lvl3_ff[12] ),
    .B(\mac1.sum_lvl3_ff[32] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2031_ (.B(net291),
    .A(\mac1.sum_lvl3_ff[12] ),
    .X(_1324_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2032_ (.B1(_1320_),
    .VDD(VPWR),
    .Y(_1325_),
    .VSS(VGND),
    .A1(_1316_),
    .A2(_1319_));
 sg13g2_nand3b_1 _2033_ (.B(_1320_),
    .C(_1317_),
    .Y(_1326_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1319_));
 sg13g2_a21oi_1 _2034_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1312_),
    .A2(_1314_),
    .Y(_1327_),
    .B1(_1326_));
 sg13g2_o21ai_1 _2035_ (.B1(net292),
    .VDD(VPWR),
    .Y(_1328_),
    .VSS(VGND),
    .A1(_1325_),
    .A2(_1327_));
 sg13g2_or3_1 _2036_ (.A(net292),
    .B(_1325_),
    .C(_1327_),
    .X(_1329_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2037_ (.A(_1328_),
    .B(_1329_),
    .X(_0019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2038_ (.Y(_1330_),
    .A(\mac1.sum_lvl3_ff[13] ),
    .B(net231),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2039_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1323_),
    .A2(_1328_),
    .Y(_1331_),
    .B1(net232));
 sg13g2_nand3_1 _2040_ (.B(_1328_),
    .C(net232),
    .A(_1323_),
    .Y(_1332_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2041_ (.A(net233),
    .B_N(_1332_),
    .Y(_0020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2042_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\mac1.sum_lvl3_ff[13] ),
    .A2(\mac1.sum_lvl3_ff[33] ),
    .Y(_1333_),
    .B1(_1331_));
 sg13g2_nand2_1 _2043_ (.Y(_1334_),
    .A(\mac1.sum_lvl3_ff[14] ),
    .B(\mac1.sum_lvl3_ff[34] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2044_ (.A(\mac1.sum_lvl3_ff[14] ),
    .B(\mac1.sum_lvl3_ff[34] ),
    .Y(_1335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2045_ (.B(net186),
    .A(\mac1.sum_lvl3_ff[14] ),
    .X(_1336_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2046_ (.Y(_0021_),
    .A(_1333_),
    .B(net187),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2047_ (.B1(_1334_),
    .VDD(VPWR),
    .Y(_1337_),
    .VSS(VGND),
    .A1(_1333_),
    .A2(_1335_));
 sg13g2_xnor2_1 _2048_ (.Y(_1338_),
    .A(\mac1.sum_lvl3_ff[15] ),
    .B(net163),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2049_ (.Y(_0022_),
    .A(_1337_),
    .B(net164),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2050_ (.B(net153),
    .A(\mac1.sum_lvl3_ff[0] ),
    .X(_0016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _2051_ (.X(_1339_),
    .A(net454),
    .B(net392),
    .C(_0032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2052_ (.Y(_1340_),
    .B1(net392),
    .B2(net457),
    .A2(net454),
    .A1(net397),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2053_ (.A(_1339_),
    .B(_1340_),
    .Y(_0033_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2054_ (.Y(_1341_),
    .A(net457),
    .B(net390),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2055_ (.A(net397),
    .B(net454),
    .C(net452),
    .D(net392),
    .X(_1342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2056_ (.Y(_1343_),
    .B1(net392),
    .B2(net454),
    .A2(net452),
    .A1(net397),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2057_ (.A(_1341_),
    .B(_1342_),
    .C(_1343_),
    .Y(_1344_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2058_ (.B1(_1341_),
    .VDD(VPWR),
    .Y(_1345_),
    .VSS(VGND),
    .A1(_1342_),
    .A2(_1343_));
 sg13g2_nor2b_1 _2059_ (.A(_1344_),
    .B_N(_1345_),
    .Y(_1346_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2060_ (.Y(_1347_),
    .A(_1339_),
    .B(_1346_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2061_ (.B(_1346_),
    .A(_1339_),
    .X(_0034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2062_ (.Y(_1348_),
    .A(net457),
    .B(net388),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2063_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1349_),
    .B(_1344_),
    .A(_1342_));
 sg13g2_nand2_1 _2064_ (.Y(_1350_),
    .A(net454),
    .B(net390),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2065_ (.A(net397),
    .B(net452),
    .C(net450),
    .D(net392),
    .X(_1351_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2066_ (.B(net452),
    .C(net450),
    .A(net398),
    .Y(_1352_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net392));
 sg13g2_a22oi_1 _2067_ (.Y(_1353_),
    .B1(net392),
    .B2(net452),
    .A2(net450),
    .A1(net397),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2068_ (.A(_1350_),
    .B(_1351_),
    .C(_1353_),
    .Y(_1354_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2069_ (.B1(_1350_),
    .VDD(VPWR),
    .Y(_1355_),
    .VSS(VGND),
    .A1(_1351_),
    .A2(_1353_));
 sg13g2_nor2b_1 _2070_ (.A(_1354_),
    .B_N(_1355_),
    .Y(_1356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2071_ (.Y(_1357_),
    .A(_1349_),
    .B(_1356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2072_ (.Y(_1358_),
    .A(_1349_),
    .B(_1356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2073_ (.B(_1358_),
    .A(_1348_),
    .X(_1359_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2074_ (.Y(_1360_),
    .B(_1359_),
    .A_N(_1347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2075_ (.Y(_0035_),
    .A(_1347_),
    .B(_1359_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2076_ (.Y(_1361_),
    .B1(net386),
    .B2(net457),
    .A2(net388),
    .A1(net454),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2077_ (.Y(_1362_),
    .A(net455),
    .B(net386),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2078_ (.A(net457),
    .B(net454),
    .C(net388),
    .D(net386),
    .X(_1363_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2079_ (.A(_1361_),
    .B(_1363_),
    .Y(_1364_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2080_ (.VDD(VPWR),
    .Y(_1365_),
    .A(_1364_),
    .VSS(VGND));
 sg13g2_o21ai_1 _2081_ (.B1(_1352_),
    .VDD(VPWR),
    .Y(_1366_),
    .VSS(VGND),
    .A1(_1350_),
    .A2(_1353_));
 sg13g2_nand2_1 _2082_ (.Y(_1367_),
    .A(net452),
    .B(net390),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2083_ (.A(net397),
    .B(net450),
    .C(net447),
    .D(net393),
    .X(_1368_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2084_ (.B(net450),
    .C(net447),
    .A(net397),
    .Y(_1369_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net392));
 sg13g2_a22oi_1 _2085_ (.Y(_1370_),
    .B1(net393),
    .B2(net450),
    .A2(net447),
    .A1(net398),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2086_ (.A(_1367_),
    .B(_1368_),
    .C(_1370_),
    .X(_1371_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2087_ (.B1(_1367_),
    .VDD(VPWR),
    .Y(_1372_),
    .VSS(VGND),
    .A1(_1368_),
    .A2(_1370_));
 sg13g2_nand3_1 _2088_ (.B(_1371_),
    .C(_1372_),
    .A(_1366_),
    .Y(_1373_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2089_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1371_),
    .A2(_1372_),
    .Y(_1374_),
    .B1(_1366_));
 sg13g2_a21o_1 _2090_ (.A2(_1372_),
    .A1(_1371_),
    .B1(_1366_),
    .X(_1375_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2091_ (.Y(_1376_),
    .A(_1373_),
    .B(_1375_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2092_ (.Y(_1377_),
    .A(_1365_),
    .B(_1376_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2093_ (.B1(_1357_),
    .VDD(VPWR),
    .Y(_1378_),
    .VSS(VGND),
    .A1(_1348_),
    .A2(_1358_));
 sg13g2_nor2b_2 _2094_ (.A(_1377_),
    .B_N(_1378_),
    .Y(_1379_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2095_ (.B(_1378_),
    .A(_1377_),
    .X(_1380_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2096_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1381_),
    .B(_1380_),
    .A(_1360_));
 sg13g2_xor2_1 _2097_ (.B(_1380_),
    .A(_1360_),
    .X(_0036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2098_ (.B1(_1373_),
    .VDD(VPWR),
    .Y(_1382_),
    .VSS(VGND),
    .A1(_1365_),
    .A2(_1374_));
 sg13g2_nand2_1 _2099_ (.Y(_1383_),
    .A(net458),
    .B(net384),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2100_ (.Y(_1384_),
    .A(net452),
    .B(net386),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2101_ (.Y(_1385_),
    .A(net452),
    .B(net388),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2102_ (.B(_1385_),
    .A(_1362_),
    .X(_1386_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2103_ (.Y(_1387_),
    .B(_1386_),
    .A_N(_1383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2104_ (.B(_1386_),
    .A(_1383_),
    .X(_1388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2105_ (.B1(_1369_),
    .VDD(VPWR),
    .Y(_1389_),
    .VSS(VGND),
    .A1(_1367_),
    .A2(_1370_));
 sg13g2_nand2_1 _2106_ (.Y(_1390_),
    .A(net450),
    .B(net390),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2107_ (.A(net398),
    .B(net447),
    .C(net444),
    .D(net393),
    .X(_1391_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2108_ (.B(net447),
    .C(net444),
    .A(net398),
    .Y(_1392_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net393));
 sg13g2_a22oi_1 _2109_ (.Y(_1393_),
    .B1(net393),
    .B2(net447),
    .A2(net444),
    .A1(net398),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2110_ (.A(_1390_),
    .B(_1391_),
    .C(_1393_),
    .X(_1394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2111_ (.B1(_1390_),
    .VDD(VPWR),
    .Y(_1395_),
    .VSS(VGND),
    .A1(_1391_),
    .A2(_1393_));
 sg13g2_and3_1 _2112_ (.X(_1396_),
    .A(_1389_),
    .B(_1394_),
    .C(_1395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2113_ (.B(_1394_),
    .C(_1395_),
    .A(_1389_),
    .Y(_1397_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2114_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1394_),
    .A2(_1395_),
    .Y(_1398_),
    .B1(_1389_));
 sg13g2_or3_1 _2115_ (.A(_1388_),
    .B(_1396_),
    .C(_1398_),
    .X(_1399_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2116_ (.B1(_1388_),
    .VDD(VPWR),
    .Y(_1400_),
    .VSS(VGND),
    .A1(_1396_),
    .A2(_1398_));
 sg13g2_nand3_1 _2117_ (.B(_1399_),
    .C(_1400_),
    .A(_1382_),
    .Y(_1401_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2118_ (.A2(_1400_),
    .A1(_1399_),
    .B1(_1382_),
    .X(_1402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2119_ (.B(_1401_),
    .C(_1402_),
    .A(_1363_),
    .Y(_1403_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2120_ (.A2(_1402_),
    .A1(_1401_),
    .B1(_1363_),
    .X(_1404_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2121_ (.A(_1403_),
    .B(_1404_),
    .X(_1405_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2122_ (.B(_1403_),
    .C(_1404_),
    .A(_1379_),
    .Y(_1406_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2123_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1403_),
    .A2(_1404_),
    .Y(_1407_),
    .B1(_1379_));
 sg13g2_xor2_1 _2124_ (.B(_1405_),
    .A(_1379_),
    .X(_1408_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2125_ (.Y(_0047_),
    .A(_1381_),
    .B(_1408_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2126_ (.Y(_1409_),
    .A(_1401_),
    .B(_1403_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2127_ (.B1(_1387_),
    .VDD(VPWR),
    .Y(_1410_),
    .VSS(VGND),
    .A1(_1362_),
    .A2(_1385_));
 sg13g2_nand2_1 _2128_ (.Y(_1411_),
    .A(net457),
    .B(net382),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2129_ (.Y(_1412_),
    .B(_1410_),
    .A_N(_1411_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2130_ (.B(_1411_),
    .A(_1410_),
    .X(_1413_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2131_ (.B1(_1397_),
    .VDD(VPWR),
    .Y(_1414_),
    .VSS(VGND),
    .A1(_1388_),
    .A2(_1398_));
 sg13g2_nand2_1 _2132_ (.Y(_1415_),
    .A(net455),
    .B(net384),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2133_ (.Y(_1416_),
    .A(net450),
    .B(net386),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2134_ (.Y(_1417_),
    .A(net451),
    .B(net388),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2135_ (.B(_1417_),
    .A(_1384_),
    .X(_1418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2136_ (.Y(_1419_),
    .B(_1418_),
    .A_N(_1415_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2137_ (.Y(_1420_),
    .A(_1415_),
    .B(_1418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2138_ (.B1(_1392_),
    .VDD(VPWR),
    .Y(_1421_),
    .VSS(VGND),
    .A1(_1390_),
    .A2(_1393_));
 sg13g2_nand2_1 _2139_ (.Y(_1422_),
    .A(net447),
    .B(net390),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2140_ (.A(net399),
    .B(net444),
    .C(net442),
    .D(net394),
    .X(_1423_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2141_ (.B(net444),
    .C(net442),
    .A(net399),
    .Y(_1424_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net394));
 sg13g2_a22oi_1 _2142_ (.Y(_1425_),
    .B1(net394),
    .B2(net444),
    .A2(net442),
    .A1(net399),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2143_ (.A(_1422_),
    .B(_1423_),
    .C(_1425_),
    .X(_1426_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2144_ (.B1(_1422_),
    .VDD(VPWR),
    .Y(_1427_),
    .VSS(VGND),
    .A1(_1423_),
    .A2(_1425_));
 sg13g2_and3_1 _2145_ (.X(_1428_),
    .A(_1421_),
    .B(_1426_),
    .C(_1427_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2146_ (.B(_1426_),
    .C(_1427_),
    .A(_1421_),
    .Y(_1429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2147_ (.A2(_1427_),
    .A1(_1426_),
    .B1(_1421_),
    .X(_1430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2148_ (.B(_1429_),
    .C(_1430_),
    .A(_1420_),
    .Y(_1431_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2149_ (.A2(_1430_),
    .A1(_1429_),
    .B1(_1420_),
    .X(_1432_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2150_ (.B(_1431_),
    .C(_1432_),
    .A(_1414_),
    .Y(_1433_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2151_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1431_),
    .A2(_1432_),
    .Y(_1434_),
    .B1(_1414_));
 sg13g2_a21o_1 _2152_ (.A2(_1432_),
    .A1(_1431_),
    .B1(_1414_),
    .X(_1435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2153_ (.Y(_1436_),
    .A(_1433_),
    .B(_1435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2154_ (.Y(_1437_),
    .A(_1413_),
    .B(_1436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2155_ (.A(_1437_),
    .B_N(_1409_),
    .Y(_1438_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2156_ (.Y(_1439_),
    .A(_1409_),
    .B(_1437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2157_ (.B1(_1406_),
    .VDD(VPWR),
    .Y(_1440_),
    .VSS(VGND),
    .A1(_1381_),
    .A2(_1407_));
 sg13g2_xor2_1 _2158_ (.B(_1440_),
    .A(_1439_),
    .X(_0054_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2159_ (.B1(_1433_),
    .VDD(VPWR),
    .Y(_1441_),
    .VSS(VGND),
    .A1(_1413_),
    .A2(_1434_));
 sg13g2_o21ai_1 _2160_ (.B1(_1419_),
    .VDD(VPWR),
    .Y(_1442_),
    .VSS(VGND),
    .A1(_1384_),
    .A2(_1417_));
 sg13g2_a22oi_1 _2161_ (.Y(_1443_),
    .B1(net380),
    .B2(net458),
    .A2(net382),
    .A1(net455),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2162_ (.B(net455),
    .C(net382),
    .A(net458),
    .Y(_1444_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net380));
 sg13g2_nor2b_1 _2163_ (.A(_1443_),
    .B_N(_1444_),
    .Y(_1445_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2164_ (.Y(_1446_),
    .A(_1442_),
    .B(_1445_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2165_ (.Y(_1447_),
    .A(_1442_),
    .B(_1445_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2166_ (.A2(_1430_),
    .A1(_1420_),
    .B1(_1428_),
    .X(_1448_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2167_ (.Y(_1449_),
    .A(net453),
    .B(net384),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2168_ (.Y(_1450_),
    .A(net447),
    .B(net386),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2169_ (.Y(_1451_),
    .A(net448),
    .B(net388),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2170_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1452_),
    .B(_1450_),
    .A(_1417_));
 sg13g2_and2_1 _2171_ (.A(_1416_),
    .B(_1451_),
    .X(_1453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2172_ (.Y(_1454_),
    .A(_1416_),
    .B(_1451_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2173_ (.Y(_1455_),
    .A(_1449_),
    .B(_1454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2174_ (.B1(_1424_),
    .VDD(VPWR),
    .Y(_1456_),
    .VSS(VGND),
    .A1(_1422_),
    .A2(_1425_));
 sg13g2_nand2_1 _2175_ (.Y(_1457_),
    .A(net444),
    .B(net391),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2176_ (.A(net399),
    .B(net442),
    .C(net440),
    .D(net394),
    .X(_1458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2177_ (.B(net442),
    .C(net440),
    .A(net399),
    .Y(_1459_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net395));
 sg13g2_a22oi_1 _2178_ (.Y(_1460_),
    .B1(net395),
    .B2(net442),
    .A2(net440),
    .A1(net399),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2179_ (.A(_1457_),
    .B(_1458_),
    .C(_1460_),
    .X(_1461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2180_ (.B1(_1457_),
    .VDD(VPWR),
    .Y(_1462_),
    .VSS(VGND),
    .A1(_1458_),
    .A2(_1460_));
 sg13g2_and3_1 _2181_ (.X(_1463_),
    .A(_1456_),
    .B(_1461_),
    .C(_1462_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2182_ (.B(_1461_),
    .C(_1462_),
    .A(_1456_),
    .Y(_1464_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2183_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1461_),
    .A2(_1462_),
    .Y(_1465_),
    .B1(_1456_));
 sg13g2_or3_1 _2184_ (.A(_1455_),
    .B(_1463_),
    .C(_1465_),
    .X(_1466_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2185_ (.B1(_1455_),
    .VDD(VPWR),
    .Y(_1467_),
    .VSS(VGND),
    .A1(_1463_),
    .A2(_1465_));
 sg13g2_and3_1 _2186_ (.X(_1468_),
    .A(_1448_),
    .B(_1466_),
    .C(_1467_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2187_ (.B(_1466_),
    .C(_1467_),
    .A(_1448_),
    .Y(_1469_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2188_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1466_),
    .A2(_1467_),
    .Y(_1470_),
    .B1(_1448_));
 sg13g2_or3_1 _2189_ (.A(_1447_),
    .B(_1468_),
    .C(_1470_),
    .X(_1471_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2190_ (.B1(_1447_),
    .VDD(VPWR),
    .Y(_1472_),
    .VSS(VGND),
    .A1(_1468_),
    .A2(_1470_));
 sg13g2_nand3_1 _2191_ (.B(_1471_),
    .C(_1472_),
    .A(_1441_),
    .Y(_1473_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2192_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1471_),
    .A2(_1472_),
    .Y(_1474_),
    .B1(_1441_));
 sg13g2_a21o_1 _2193_ (.A2(_1472_),
    .A1(_1471_),
    .B1(_1441_),
    .X(_1475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2194_ (.Y(_1476_),
    .A(_1473_),
    .B(_1475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2195_ (.B(_1476_),
    .A(_1412_),
    .X(_1477_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _2196_ (.A2(_1440_),
    .A1(_1439_),
    .B1(_1438_),
    .X(_1478_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2197_ (.Y(_1479_),
    .A(_1477_),
    .B(_1478_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2198_ (.B(_1478_),
    .A(_1477_),
    .X(_0055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2199_ (.B1(_1469_),
    .VDD(VPWR),
    .Y(_1480_),
    .VSS(VGND),
    .A1(_1447_),
    .A2(_1470_));
 sg13g2_o21ai_1 _2200_ (.B1(_1452_),
    .VDD(VPWR),
    .Y(_1481_),
    .VSS(VGND),
    .A1(_1449_),
    .A2(_1453_));
 sg13g2_nand2_1 _2201_ (.Y(_1482_),
    .A(net458),
    .B(net502),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2202_ (.Y(_1483_),
    .A(net453),
    .B(net380),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2203_ (.A(net456),
    .B(net453),
    .C(net382),
    .D(net380),
    .X(_1484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2204_ (.Y(_1485_),
    .B1(net380),
    .B2(net456),
    .A2(net382),
    .A1(net453),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2205_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1486_),
    .B(_1485_),
    .A(_1484_));
 sg13g2_nor2_1 _2206_ (.A(_1482_),
    .B(_1486_),
    .Y(_1487_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2207_ (.B(_1486_),
    .A(_1482_),
    .X(_1488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2208_ (.Y(_1489_),
    .A(_1481_),
    .B(_1488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2209_ (.Y(_1490_),
    .A(_1481_),
    .B(_1488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2210_ (.Y(_1491_),
    .A(_1444_),
    .B(_1490_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2211_ (.B1(_1464_),
    .VDD(VPWR),
    .Y(_1492_),
    .VSS(VGND),
    .A1(_1455_),
    .A2(_1465_));
 sg13g2_nand2_1 _2212_ (.Y(_1493_),
    .A(net451),
    .B(net384),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2213_ (.Y(_1494_),
    .A(net445),
    .B(net386),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2214_ (.Y(_1495_),
    .A(net444),
    .B(net388),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2215_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1496_),
    .B(_1494_),
    .A(_1451_));
 sg13g2_xnor2_1 _2216_ (.Y(_1497_),
    .A(_1450_),
    .B(_1495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2217_ (.Y(_1498_),
    .A(_1493_),
    .B(_1497_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2218_ (.B1(_1459_),
    .VDD(VPWR),
    .Y(_1499_),
    .VSS(VGND),
    .A1(_1457_),
    .A2(_1460_));
 sg13g2_nand2_1 _2219_ (.Y(_1500_),
    .A(net442),
    .B(net390),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2220_ (.A(net400),
    .B(net440),
    .C(net496),
    .D(net394),
    .X(_0134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2221_ (.B(net440),
    .C(net496),
    .A(net399),
    .Y(_0135_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net394));
 sg13g2_a22oi_1 _2222_ (.Y(_0136_),
    .B1(net394),
    .B2(net440),
    .A2(net496),
    .A1(net400),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2223_ (.A(_1500_),
    .B(_0134_),
    .C(_0136_),
    .X(_0137_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2224_ (.B1(_1500_),
    .VDD(VPWR),
    .Y(_0138_),
    .VSS(VGND),
    .A1(_0134_),
    .A2(_0136_));
 sg13g2_and3_1 _2225_ (.X(_0139_),
    .A(_1499_),
    .B(_0137_),
    .C(_0138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2226_ (.B(_0137_),
    .C(_0138_),
    .A(_1499_),
    .Y(_0140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2227_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0137_),
    .A2(_0138_),
    .Y(_0141_),
    .B1(_1499_));
 sg13g2_or3_1 _2228_ (.A(_1498_),
    .B(_0139_),
    .C(_0141_),
    .X(_0142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2229_ (.B1(_1498_),
    .VDD(VPWR),
    .Y(_0143_),
    .VSS(VGND),
    .A1(_0139_),
    .A2(_0141_));
 sg13g2_and3_1 _2230_ (.X(_0144_),
    .A(_1492_),
    .B(_0142_),
    .C(_0143_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2231_ (.B(_0142_),
    .C(_0143_),
    .A(_1492_),
    .Y(_0145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2232_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0142_),
    .A2(_0143_),
    .Y(_0146_),
    .B1(_1492_));
 sg13g2_or3_1 _2233_ (.A(_1491_),
    .B(_0144_),
    .C(_0146_),
    .X(_0147_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2234_ (.B1(_1491_),
    .VDD(VPWR),
    .Y(_0148_),
    .VSS(VGND),
    .A1(_0144_),
    .A2(_0146_));
 sg13g2_and3_1 _2235_ (.X(_0149_),
    .A(_1480_),
    .B(_0147_),
    .C(_0148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2236_ (.B(_0147_),
    .C(_0148_),
    .A(_1480_),
    .Y(_0150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2237_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0147_),
    .A2(_0148_),
    .Y(_0151_),
    .B1(_1480_));
 sg13g2_or3_1 _2238_ (.A(_1446_),
    .B(_0149_),
    .C(_0151_),
    .X(_0152_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2239_ (.B1(_1446_),
    .VDD(VPWR),
    .Y(_0153_),
    .VSS(VGND),
    .A1(_0149_),
    .A2(_0151_));
 sg13g2_o21ai_1 _2240_ (.B1(_1473_),
    .VDD(VPWR),
    .Y(_0154_),
    .VSS(VGND),
    .A1(_1412_),
    .A2(_1474_));
 sg13g2_nand3_1 _2241_ (.B(_0153_),
    .C(_0154_),
    .A(_0152_),
    .Y(_0155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2242_ (.A2(_0153_),
    .A1(_0152_),
    .B1(_0154_),
    .X(_0156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2243_ (.Y(_0157_),
    .A(_0155_),
    .B(_0156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2244_ (.A(_1477_),
    .B(_1478_),
    .C(_0155_),
    .D(_0156_),
    .X(_0158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2245_ (.B(_0157_),
    .A(_1479_),
    .X(_0056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2246_ (.B1(_0155_),
    .VDD(VPWR),
    .Y(_0159_),
    .VSS(VGND),
    .A1(_1479_),
    .A2(_0157_));
 sg13g2_o21ai_1 _2247_ (.B1(_0150_),
    .VDD(VPWR),
    .Y(_0160_),
    .VSS(VGND),
    .A1(_1446_),
    .A2(_0151_));
 sg13g2_o21ai_1 _2248_ (.B1(_1489_),
    .VDD(VPWR),
    .Y(_0161_),
    .VSS(VGND),
    .A1(_1444_),
    .A2(_1490_));
 sg13g2_o21ai_1 _2249_ (.B1(_0145_),
    .VDD(VPWR),
    .Y(_0162_),
    .VSS(VGND),
    .A1(_1491_),
    .A2(_0146_));
 sg13g2_nor2_1 _2250_ (.A(_1484_),
    .B(_1487_),
    .Y(_0163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2251_ (.B1(_1496_),
    .VDD(VPWR),
    .Y(_0164_),
    .VSS(VGND),
    .A1(_1493_),
    .A2(_1497_));
 sg13g2_nand2_1 _2252_ (.Y(_0165_),
    .A(net456),
    .B(net502),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2253_ (.Y(_0166_),
    .A(net451),
    .B(net380),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2254_ (.Y(_0167_),
    .A(net451),
    .B(net382),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2255_ (.B(_0167_),
    .A(_1483_),
    .X(_0168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2256_ (.Y(_0169_),
    .B(_0168_),
    .A_N(_0165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2257_ (.Y(_0170_),
    .A(_0165_),
    .B(_0168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2258_ (.Y(_0171_),
    .A(_0164_),
    .B(_0170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2259_ (.A(_0163_),
    .B(_0171_),
    .Y(_0172_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2260_ (.Y(_0173_),
    .A(_0163_),
    .B(_0171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2261_ (.B1(_0140_),
    .VDD(VPWR),
    .Y(_0174_),
    .VSS(VGND),
    .A1(_1498_),
    .A2(_0141_));
 sg13g2_nand2_1 _2262_ (.Y(_0175_),
    .A(net448),
    .B(net384),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2263_ (.Y(_0176_),
    .A(net442),
    .B(net389),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2264_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0177_),
    .B(_0176_),
    .A(_1494_));
 sg13g2_and2_1 _2265_ (.A(_1494_),
    .B(_0176_),
    .X(_0178_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2266_ (.Y(_0179_),
    .A(_1494_),
    .B(_0176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2267_ (.Y(_0180_),
    .A(_0175_),
    .B(_0179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2268_ (.B1(_0135_),
    .VDD(VPWR),
    .Y(_0181_),
    .VSS(VGND),
    .A1(_1500_),
    .A2(_0136_));
 sg13g2_nand2_1 _2269_ (.Y(_0182_),
    .A(net496),
    .B(net390),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2270_ (.A(net440),
    .B(net496),
    .C(net396),
    .D(net390),
    .X(_0183_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2271_ (.Y(_0184_),
    .B1(net391),
    .B2(net440),
    .A2(net396),
    .A1(net496),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2272_ (.A(_0183_),
    .B(_0184_),
    .Y(_0185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2273_ (.Y(_0186_),
    .A(_0181_),
    .B(_0185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2274_ (.Y(_0187_),
    .A(_0181_),
    .B(_0185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2275_ (.B(_0187_),
    .A(_0180_),
    .X(_0188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2276_ (.Y(_0189_),
    .A(_0174_),
    .B(_0188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2277_ (.Y(_0190_),
    .A(_0174_),
    .B(_0188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2278_ (.B(_0190_),
    .A(_0173_),
    .X(_0191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2279_ (.Y(_0192_),
    .A(_0162_),
    .B(_0191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2280_ (.Y(_0193_),
    .A(_0162_),
    .B(_0191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2281_ (.Y(_0194_),
    .B(_0161_),
    .A_N(_0193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2282_ (.Y(_0195_),
    .A(_0161_),
    .B(_0193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2283_ (.A(_0160_),
    .B(_0195_),
    .Y(_0196_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2284_ (.Y(_0197_),
    .A(_0160_),
    .B(_0195_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2285_ (.A(_0196_),
    .B_N(_0197_),
    .Y(_0198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2286_ (.B(_0198_),
    .A(_0159_),
    .X(_0057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2287_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0164_),
    .A2(_0170_),
    .Y(_0199_),
    .B1(_0172_));
 sg13g2_o21ai_1 _2288_ (.B1(_0189_),
    .VDD(VPWR),
    .Y(_0200_),
    .VSS(VGND),
    .A1(_0173_),
    .A2(_0190_));
 sg13g2_o21ai_1 _2289_ (.B1(_0169_),
    .VDD(VPWR),
    .Y(_0201_),
    .VSS(VGND),
    .A1(_1483_),
    .A2(_0167_));
 sg13g2_o21ai_1 _2290_ (.B1(_0177_),
    .VDD(VPWR),
    .Y(_0202_),
    .VSS(VGND),
    .A1(_0175_),
    .A2(_0178_));
 sg13g2_nand2_1 _2291_ (.Y(_0203_),
    .A(\DP_1.matrix[74] ),
    .B(net502),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2292_ (.Y(_0204_),
    .A(net449),
    .B(net380),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2293_ (.Y(_0205_),
    .A(net448),
    .B(net382),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2294_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0206_),
    .B(_0204_),
    .A(_0167_));
 sg13g2_xnor2_1 _2295_ (.Y(_0207_),
    .A(_0166_),
    .B(_0205_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2296_ (.B(_0207_),
    .A(_0203_),
    .X(_0208_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2297_ (.Y(_0209_),
    .A(_0202_),
    .B(_0208_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2298_ (.A(_0209_),
    .B_N(_0201_),
    .Y(_0210_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2299_ (.B(_0209_),
    .A(_0201_),
    .X(_0211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2300_ (.B1(_0186_),
    .VDD(VPWR),
    .Y(_0212_),
    .VSS(VGND),
    .A1(_0180_),
    .A2(_0187_));
 sg13g2_a21oi_1 _2301_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net441),
    .A2(net396),
    .Y(_0213_),
    .B1(_0182_));
 sg13g2_nand2_1 _2302_ (.Y(_0214_),
    .A(net445),
    .B(net384),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2303_ (.Y(_0215_),
    .A(net441),
    .B(net387),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2304_ (.A(net443),
    .B(net441),
    .C(net389),
    .D(net387),
    .X(_0216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2305_ (.Y(_0217_),
    .B1(net387),
    .B2(net443),
    .A2(net389),
    .A1(net441),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2306_ (.A(_0214_),
    .B(_0216_),
    .C(_0217_),
    .Y(_0218_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2307_ (.B1(_0214_),
    .VDD(VPWR),
    .Y(_0219_),
    .VSS(VGND),
    .A1(_0216_),
    .A2(_0217_));
 sg13g2_nor2b_1 _2308_ (.A(_0218_),
    .B_N(_0219_),
    .Y(_0220_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2309_ (.Y(_0221_),
    .A(_0213_),
    .B(_0220_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2310_ (.Y(_0222_),
    .B(_0212_),
    .A_N(_0221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2311_ (.B(_0221_),
    .A(_0212_),
    .X(_0223_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2312_ (.B(_0223_),
    .A(_0211_),
    .X(_0224_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2313_ (.Y(_0225_),
    .A(_0200_),
    .B(_0224_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2314_ (.B(_0224_),
    .A(_0200_),
    .X(_0226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2315_ (.Y(_0227_),
    .B(_0226_),
    .A_N(_0199_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2316_ (.B(_0226_),
    .A(_0199_),
    .X(_0228_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2317_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0192_),
    .A2(_0194_),
    .Y(_0229_),
    .B1(_0228_));
 sg13g2_nand3_1 _2318_ (.B(_0194_),
    .C(_0228_),
    .A(_0192_),
    .Y(_0230_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2319_ (.Y(_0231_),
    .B(_0230_),
    .A_N(_0229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2320_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0155_),
    .A2(_0197_),
    .Y(_0232_),
    .B1(_0196_));
 sg13g2_a21oi_2 _2321_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0232_),
    .Y(_0233_),
    .A2(_0198_),
    .A1(_0158_));
 sg13g2_nor2_1 _2322_ (.A(_0231_),
    .B(_0233_),
    .Y(_0234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2323_ (.B(_0233_),
    .A(_0231_),
    .X(_0048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2324_ (.A2(_0208_),
    .A1(_0202_),
    .B1(_0210_),
    .X(_0235_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2325_ (.B1(_0222_),
    .VDD(VPWR),
    .Y(_0236_),
    .VSS(VGND),
    .A1(_0211_),
    .A2(_0223_));
 sg13g2_a21o_1 _2326_ (.A2(_0220_),
    .A1(_0213_),
    .B1(_0183_),
    .X(_0237_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2327_ (.Y(_0238_),
    .A(net443),
    .B(net384),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2328_ (.Y(_0239_),
    .A(net497),
    .B(net389),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2329_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0240_),
    .B(_0239_),
    .A(_0215_));
 sg13g2_xnor2_1 _2330_ (.Y(_0241_),
    .A(_0215_),
    .B(_0239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2331_ (.B(_0241_),
    .A(_0238_),
    .X(_0242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2332_ (.Y(_0243_),
    .A(_0237_),
    .B(_0242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2333_ (.B1(_0206_),
    .VDD(VPWR),
    .Y(_0244_),
    .VSS(VGND),
    .A1(_0203_),
    .A2(_0207_));
 sg13g2_or2_1 _2334_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0245_),
    .B(_0218_),
    .A(_0216_));
 sg13g2_nand2_1 _2335_ (.Y(_0246_),
    .A(\DP_1.matrix[75] ),
    .B(net502),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2336_ (.Y(_0247_),
    .A(net446),
    .B(net382),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2337_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0248_),
    .B(_0247_),
    .A(_0204_));
 sg13g2_xnor2_1 _2338_ (.Y(_0249_),
    .A(_0204_),
    .B(_0247_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2339_ (.B(_0249_),
    .A(_0246_),
    .X(_0250_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2340_ (.Y(_0251_),
    .A(_0245_),
    .B(_0250_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2341_ (.A(_0251_),
    .B_N(_0244_),
    .Y(_0252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2342_ (.B(_0251_),
    .A(_0244_),
    .X(_0253_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2343_ (.A(_0243_),
    .B(_0253_),
    .Y(_0254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2344_ (.B(_0253_),
    .A(_0243_),
    .X(_0255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2345_ (.Y(_0256_),
    .A(_0236_),
    .B(_0255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2346_ (.A(_0256_),
    .B_N(_0235_),
    .Y(_0257_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2347_ (.B(_0256_),
    .A(_0235_),
    .X(_0258_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2348_ (.B(_0227_),
    .C(_0258_),
    .A(_0225_),
    .Y(_0259_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2349_ (.VDD(VPWR),
    .Y(_0260_),
    .A(_0259_),
    .VSS(VGND));
 sg13g2_a21oi_1 _2350_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0225_),
    .A2(_0227_),
    .Y(_0261_),
    .B1(_0258_));
 sg13g2_nor2_1 _2351_ (.A(_0260_),
    .B(_0261_),
    .Y(_0262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2352_ (.A(_0229_),
    .B(_0234_),
    .Y(_0263_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2353_ (.Y(_0049_),
    .A(_0262_),
    .B(_0263_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2354_ (.A2(_0250_),
    .A1(_0245_),
    .B1(_0252_),
    .X(_0264_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2355_ (.Y(_0265_),
    .B1(net384),
    .B2(net441),
    .A2(net387),
    .A1(net497),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2356_ (.Y(_0266_),
    .A(net496),
    .B(net385),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2357_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0267_),
    .B(_0266_),
    .A(_0215_));
 sg13g2_nand2b_1 _2358_ (.Y(_0268_),
    .B(_0267_),
    .A_N(_0265_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2359_ (.B1(_0248_),
    .VDD(VPWR),
    .Y(_0269_),
    .VSS(VGND),
    .A1(_0246_),
    .A2(_0249_));
 sg13g2_o21ai_1 _2360_ (.B1(_0240_),
    .VDD(VPWR),
    .Y(_0270_),
    .VSS(VGND),
    .A1(_0238_),
    .A2(_0241_));
 sg13g2_nand2_1 _2361_ (.Y(_0271_),
    .A(net449),
    .B(net502),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2362_ (.Y(_0272_),
    .A(net443),
    .B(net380),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2363_ (.A(_0247_),
    .B(_0272_),
    .Y(_0273_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2364_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0274_),
    .B(_0272_),
    .A(_0247_));
 sg13g2_a22oi_1 _2365_ (.Y(_0275_),
    .B1(net381),
    .B2(net446),
    .A2(net383),
    .A1(net443),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2366_ (.A(_0273_),
    .B(_0275_),
    .Y(_0276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2367_ (.Y(_0277_),
    .A(_0271_),
    .B(_0276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2368_ (.Y(_0278_),
    .A(_0270_),
    .B(_0277_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2369_ (.A(_0278_),
    .B_N(_0269_),
    .Y(_0279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2370_ (.B(_0278_),
    .A(_0269_),
    .X(_0280_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2371_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0281_),
    .B(_0280_),
    .A(_0268_));
 sg13g2_xor2_1 _2372_ (.B(_0280_),
    .A(_0268_),
    .X(_0282_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2373_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0237_),
    .A2(_0242_),
    .Y(_0283_),
    .B1(_0254_));
 sg13g2_nor2b_1 _2374_ (.A(_0283_),
    .B_N(_0282_),
    .Y(_0284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2375_ (.B(_0283_),
    .A(_0282_),
    .X(_0285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2376_ (.A(_0285_),
    .B_N(_0264_),
    .Y(_0286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2377_ (.B(_0285_),
    .A(_0264_),
    .X(_0287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2378_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0236_),
    .A2(_0255_),
    .Y(_0288_),
    .B1(_0257_));
 sg13g2_nor2_1 _2379_ (.A(_0287_),
    .B(_0288_),
    .Y(_0289_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2380_ (.B(_0288_),
    .A(_0287_),
    .X(_0290_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2381_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0229_),
    .A2(_0259_),
    .Y(_0291_),
    .B1(_0261_));
 sg13g2_a21oi_1 _2382_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0230_),
    .A2(_0259_),
    .Y(_0292_),
    .B1(_0261_));
 sg13g2_a21oi_2 _2383_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0292_),
    .Y(_0293_),
    .A2(_0291_),
    .A1(_0233_));
 sg13g2_xor2_1 _2384_ (.B(_0293_),
    .A(_0290_),
    .X(_0050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2385_ (.A2(_0277_),
    .A1(_0270_),
    .B1(_0279_),
    .X(_0294_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2386_ (.B1(_0274_),
    .VDD(VPWR),
    .Y(_0295_),
    .VSS(VGND),
    .A1(_0271_),
    .A2(_0275_));
 sg13g2_nand2_1 _2387_ (.Y(_0296_),
    .A(net446),
    .B(net502),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2388_ (.Y(_0297_),
    .A(\DP_1.matrix[79] ),
    .B(net381),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2389_ (.Y(_0298_),
    .A(\DP_1.matrix[79] ),
    .B(net383),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2390_ (.B(_0298_),
    .A(_0272_),
    .X(_0299_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2391_ (.Y(_0300_),
    .B(_0299_),
    .A_N(_0296_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2392_ (.Y(_0301_),
    .A(_0296_),
    .B(_0299_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2393_ (.A(_0267_),
    .B_N(_0301_),
    .Y(_0302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2394_ (.Y(_0303_),
    .A(_0267_),
    .B(_0301_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2395_ (.Y(_0304_),
    .A(_0295_),
    .B(_0303_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2396_ (.A(_0266_),
    .B(_0304_),
    .Y(_0305_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2397_ (.B(_0304_),
    .A(_0266_),
    .X(_0306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2398_ (.Y(_0307_),
    .B(_0306_),
    .A_N(_0281_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2399_ (.Y(_0308_),
    .A(_0281_),
    .B(_0306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2400_ (.Y(_0309_),
    .A(_0294_),
    .B(_0308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2401_ (.B(_0308_),
    .A(_0294_),
    .X(_0310_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2402_ (.B1(_0310_),
    .VDD(VPWR),
    .Y(_0311_),
    .VSS(VGND),
    .A1(_0284_),
    .A2(_0286_));
 sg13g2_or3_1 _2403_ (.A(_0284_),
    .B(_0286_),
    .C(_0310_),
    .X(_0312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2404_ (.A(_0311_),
    .B(_0312_),
    .X(_0313_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2405_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0290_),
    .A2(_0293_),
    .Y(_0314_),
    .B1(_0289_));
 sg13g2_xnor2_1 _2406_ (.Y(_0051_),
    .A(_0313_),
    .B(_0314_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2407_ (.A(_0290_),
    .B(_0313_),
    .X(_0315_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2408_ (.Y(_0316_),
    .A(_0289_),
    .B(_0312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2409_ (.Y(_0317_),
    .A(_0311_),
    .B(_0316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2410_ (.A2(_0315_),
    .A1(_0293_),
    .B1(_0317_),
    .X(_0318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2411_ (.A(_0307_),
    .B(_0309_),
    .X(_0319_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2412_ (.A2(_0303_),
    .A1(_0295_),
    .B1(_0302_),
    .X(_0320_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2413_ (.B1(_0300_),
    .VDD(VPWR),
    .Y(_0321_),
    .VSS(VGND),
    .A1(_0272_),
    .A2(_0298_));
 sg13g2_nand2_1 _2414_ (.Y(_0322_),
    .A(net443),
    .B(\DP_2.matrix[80] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2415_ (.Y(_0323_),
    .A(net497),
    .B(net381),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2416_ (.Y(_0324_),
    .A(net497),
    .B(net383),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2417_ (.B(_0324_),
    .A(_0297_),
    .X(_0325_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2418_ (.Y(_0326_),
    .B(_0325_),
    .A_N(_0322_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2419_ (.Y(_0327_),
    .A(_0322_),
    .B(_0325_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2420_ (.Y(_0328_),
    .A(_0321_),
    .B(_0327_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2421_ (.B(_0327_),
    .A(_0321_),
    .X(_0329_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2422_ (.Y(_0330_),
    .A(_0305_),
    .B(_0329_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2423_ (.A(_0330_),
    .B_N(_0320_),
    .Y(_0331_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2424_ (.B(_0330_),
    .A(_0320_),
    .X(_0332_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2425_ (.A(_0319_),
    .B(_0332_),
    .Y(_0333_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2426_ (.B(_0332_),
    .A(_0319_),
    .X(_0334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2427_ (.B(_0334_),
    .A(_0318_),
    .X(_0052_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2428_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0318_),
    .A2(_0334_),
    .Y(_0335_),
    .B1(_0333_));
 sg13g2_a21oi_1 _2429_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0305_),
    .A2(_0329_),
    .Y(_0336_),
    .B1(_0331_));
 sg13g2_o21ai_1 _2430_ (.B1(_0326_),
    .VDD(VPWR),
    .Y(_0337_),
    .VSS(VGND),
    .A1(_0297_),
    .A2(_0324_));
 sg13g2_nand2_1 _2431_ (.Y(_0338_),
    .A(net441),
    .B(net502),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2432_ (.Y(_0339_),
    .A(_0323_),
    .B(_0338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2433_ (.Y(_0340_),
    .A(_0337_),
    .B(_0339_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2434_ (.Y(_0341_),
    .A(_0328_),
    .B(_0340_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2435_ (.Y(_0342_),
    .A(_0336_),
    .B(_0341_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2436_ (.Y(_0053_),
    .A(_0335_),
    .B(_0342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _2437_ (.X(_0343_),
    .A(net490),
    .B(net433),
    .C(_0037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2438_ (.Y(_0344_),
    .B1(net433),
    .B2(net492),
    .A2(net490),
    .A1(net437),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2439_ (.A(_0343_),
    .B(_0344_),
    .Y(_0038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2440_ (.Y(_0345_),
    .A(net492),
    .B(net431),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2441_ (.A(net437),
    .B(net490),
    .C(net488),
    .D(net433),
    .X(_0346_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2442_ (.Y(_0347_),
    .B1(net433),
    .B2(net490),
    .A2(net488),
    .A1(net437),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2443_ (.A(_0345_),
    .B(_0346_),
    .C(_0347_),
    .Y(_0348_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2444_ (.B1(_0345_),
    .VDD(VPWR),
    .Y(_0349_),
    .VSS(VGND),
    .A1(_0346_),
    .A2(_0347_));
 sg13g2_nor2b_1 _2445_ (.A(_0348_),
    .B_N(_0349_),
    .Y(_0350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2446_ (.Y(_0351_),
    .A(_0343_),
    .B(_0350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2447_ (.B(_0350_),
    .A(_0343_),
    .X(_0039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2448_ (.Y(_0352_),
    .A(net492),
    .B(net429),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2449_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0353_),
    .B(_0348_),
    .A(_0346_));
 sg13g2_nand2_1 _2450_ (.Y(_0354_),
    .A(net490),
    .B(net431),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2451_ (.A(net437),
    .B(net488),
    .C(net486),
    .D(net433),
    .X(_0355_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2452_ (.B(net488),
    .C(net486),
    .A(net437),
    .Y(_0356_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net433));
 sg13g2_a22oi_1 _2453_ (.Y(_0357_),
    .B1(\DP_2.matrix[1] ),
    .B2(net488),
    .A2(net486),
    .A1(\DP_2.matrix[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2454_ (.A(_0354_),
    .B(_0355_),
    .C(_0357_),
    .Y(_0358_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2455_ (.B1(_0354_),
    .VDD(VPWR),
    .Y(_0359_),
    .VSS(VGND),
    .A1(_0355_),
    .A2(_0357_));
 sg13g2_nor2b_1 _2456_ (.A(_0358_),
    .B_N(_0359_),
    .Y(_0360_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2457_ (.Y(_0361_),
    .A(_0353_),
    .B(_0360_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2458_ (.Y(_0362_),
    .A(_0353_),
    .B(_0360_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2459_ (.Y(_0363_),
    .A(_0352_),
    .B(_0362_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2460_ (.A(_0351_),
    .B(_0363_),
    .Y(_0364_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2461_ (.B(_0363_),
    .A(_0351_),
    .X(_0040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2462_ (.Y(_0365_),
    .B1(net427),
    .B2(net492),
    .A2(net429),
    .A1(net490),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2463_ (.Y(_0366_),
    .A(net491),
    .B(net427),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2464_ (.A(_0352_),
    .B(_0366_),
    .Y(_0367_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2465_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0368_),
    .B(_0366_),
    .A(_0352_));
 sg13g2_nand2b_1 _2466_ (.Y(_0369_),
    .B(_0368_),
    .A_N(_0365_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2467_ (.B1(_0356_),
    .VDD(VPWR),
    .Y(_0370_),
    .VSS(VGND),
    .A1(_0354_),
    .A2(_0357_));
 sg13g2_nand2_1 _2468_ (.Y(_0371_),
    .A(net488),
    .B(net431),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2469_ (.A(net439),
    .B(net486),
    .C(net485),
    .D(net436),
    .X(_0372_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2470_ (.B(net486),
    .C(net485),
    .A(net439),
    .Y(_0373_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net436));
 sg13g2_a22oi_1 _2471_ (.Y(_0374_),
    .B1(net436),
    .B2(net486),
    .A2(net485),
    .A1(net439),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2472_ (.A(_0371_),
    .B(_0372_),
    .C(_0374_),
    .X(_0375_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2473_ (.B1(_0371_),
    .VDD(VPWR),
    .Y(_0376_),
    .VSS(VGND),
    .A1(_0372_),
    .A2(_0374_));
 sg13g2_nand3_1 _2474_ (.B(_0375_),
    .C(_0376_),
    .A(_0370_),
    .Y(_0377_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2475_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0375_),
    .A2(_0376_),
    .Y(_0378_),
    .B1(_0370_));
 sg13g2_a21o_1 _2476_ (.A2(_0376_),
    .A1(_0375_),
    .B1(_0370_),
    .X(_0379_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2477_ (.Y(_0380_),
    .A(_0377_),
    .B(_0379_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2478_ (.Y(_0381_),
    .A(_0369_),
    .B(_0380_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2479_ (.B1(_0361_),
    .VDD(VPWR),
    .Y(_0382_),
    .VSS(VGND),
    .A1(_0352_),
    .A2(_0362_));
 sg13g2_nand2b_1 _2480_ (.Y(_0383_),
    .B(_0382_),
    .A_N(_0381_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2481_ (.Y(_0384_),
    .A(_0381_),
    .B(_0382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2482_ (.Y(_0385_),
    .A(_0364_),
    .B(_0384_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2483_ (.B(_0384_),
    .A(_0364_),
    .X(_0041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2484_ (.B1(_0377_),
    .VDD(VPWR),
    .Y(_0386_),
    .VSS(VGND),
    .A1(_0369_),
    .A2(_0378_));
 sg13g2_nand2_1 _2485_ (.Y(_0387_),
    .A(net492),
    .B(net426),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2486_ (.Y(_0388_),
    .A(net489),
    .B(net427),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2487_ (.Y(_0389_),
    .A(net489),
    .B(net429),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2488_ (.B(_0389_),
    .A(_0366_),
    .X(_0390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2489_ (.Y(_0391_),
    .B(_0390_),
    .A_N(_0387_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2490_ (.Y(_0392_),
    .A(_0387_),
    .B(_0390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2491_ (.B1(_0373_),
    .VDD(VPWR),
    .Y(_0393_),
    .VSS(VGND),
    .A1(_0371_),
    .A2(_0374_));
 sg13g2_nand2_1 _2492_ (.Y(_0394_),
    .A(net487),
    .B(net431),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2493_ (.A(net439),
    .B(net485),
    .C(net481),
    .D(net436),
    .X(_0395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2494_ (.B(net484),
    .C(net481),
    .A(net439),
    .Y(_0396_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net436));
 sg13g2_a22oi_1 _2495_ (.Y(_0397_),
    .B1(net436),
    .B2(net484),
    .A2(net481),
    .A1(net439),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2496_ (.A(_0394_),
    .B(_0395_),
    .C(_0397_),
    .X(_0398_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2497_ (.B1(_0394_),
    .VDD(VPWR),
    .Y(_0399_),
    .VSS(VGND),
    .A1(_0395_),
    .A2(_0397_));
 sg13g2_and3_1 _2498_ (.X(_0400_),
    .A(_0393_),
    .B(_0398_),
    .C(_0399_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2499_ (.B(_0398_),
    .C(_0399_),
    .A(_0393_),
    .Y(_0401_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2500_ (.A2(_0399_),
    .A1(_0398_),
    .B1(_0393_),
    .X(_0402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2501_ (.B(_0401_),
    .C(_0402_),
    .A(_0392_),
    .Y(_0403_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2502_ (.A2(_0402_),
    .A1(_0401_),
    .B1(_0392_),
    .X(_0404_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2503_ (.B(_0403_),
    .C(_0404_),
    .A(_0386_),
    .Y(_0405_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2504_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0403_),
    .A2(_0404_),
    .Y(_0406_),
    .B1(_0386_));
 sg13g2_a21o_1 _2505_ (.A2(_0404_),
    .A1(_0403_),
    .B1(_0386_),
    .X(_0407_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2506_ (.B(_0405_),
    .C(_0407_),
    .A(_0367_),
    .Y(_0408_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2507_ (.A2(_0407_),
    .A1(_0405_),
    .B1(_0367_),
    .X(_0409_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2508_ (.A(_0408_),
    .B(_0409_),
    .X(_0410_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2509_ (.Y(_0411_),
    .A(_0383_),
    .B(_0385_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2510_ (.B(_0411_),
    .A(_0410_),
    .X(_0058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2511_ (.A(_0385_),
    .B_N(_0410_),
    .Y(_0412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _2512_ (.B(_0408_),
    .C(_0409_),
    .Y(_0413_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0383_));
 sg13g2_o21ai_1 _2513_ (.B1(_0405_),
    .VDD(VPWR),
    .Y(_0414_),
    .VSS(VGND),
    .A1(_0368_),
    .A2(_0406_));
 sg13g2_o21ai_1 _2514_ (.B1(_0391_),
    .VDD(VPWR),
    .Y(_0415_),
    .VSS(VGND),
    .A1(_0366_),
    .A2(_0389_));
 sg13g2_nand2_2 _2515_ (.Y(_0416_),
    .A(net493),
    .B(net425),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2516_ (.Y(_0417_),
    .B(_0415_),
    .A_N(_0416_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2517_ (.Y(_0418_),
    .A(_0415_),
    .B(_0416_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2518_ (.B(_0416_),
    .A(_0415_),
    .X(_0419_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2519_ (.A2(_0402_),
    .A1(_0392_),
    .B1(_0400_),
    .X(_0420_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2520_ (.Y(_0421_),
    .A(net491),
    .B(\DP_2.matrix[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2521_ (.Y(_0422_),
    .A(net487),
    .B(net427),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2522_ (.Y(_0423_),
    .A(net487),
    .B(net429),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2523_ (.B(_0423_),
    .A(_0388_),
    .X(_0424_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2524_ (.Y(_0425_),
    .B(_0424_),
    .A_N(_0421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2525_ (.Y(_0426_),
    .A(_0421_),
    .B(_0424_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2526_ (.B1(_0396_),
    .VDD(VPWR),
    .Y(_0427_),
    .VSS(VGND),
    .A1(_0394_),
    .A2(_0397_));
 sg13g2_nand2_1 _2527_ (.Y(_0428_),
    .A(net484),
    .B(net431),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2528_ (.A(net438),
    .B(net481),
    .C(net480),
    .D(net435),
    .X(_0429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2529_ (.B(net481),
    .C(net480),
    .A(net439),
    .Y(_0430_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net435));
 sg13g2_a22oi_1 _2530_ (.Y(_0431_),
    .B1(net435),
    .B2(net481),
    .A2(net480),
    .A1(net438),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2531_ (.A(_0428_),
    .B(_0429_),
    .C(_0431_),
    .X(_0432_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2532_ (.B1(_0428_),
    .VDD(VPWR),
    .Y(_0433_),
    .VSS(VGND),
    .A1(_0429_),
    .A2(_0431_));
 sg13g2_and3_1 _2533_ (.X(_0434_),
    .A(_0427_),
    .B(_0432_),
    .C(_0433_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2534_ (.B(_0432_),
    .C(_0433_),
    .A(_0427_),
    .Y(_0435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2535_ (.A2(_0433_),
    .A1(_0432_),
    .B1(_0427_),
    .X(_0436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2536_ (.B(_0435_),
    .C(_0436_),
    .A(_0426_),
    .Y(_0437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2537_ (.A2(_0436_),
    .A1(_0435_),
    .B1(_0426_),
    .X(_0438_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2538_ (.B(_0437_),
    .C(_0438_),
    .A(_0420_),
    .Y(_0439_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2539_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0437_),
    .A2(_0438_),
    .Y(_0440_),
    .B1(_0420_));
 sg13g2_a21o_1 _2540_ (.A2(_0438_),
    .A1(_0437_),
    .B1(_0420_),
    .X(_0441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2541_ (.B(_0439_),
    .C(_0441_),
    .A(_0418_),
    .Y(_0442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2542_ (.A2(_0441_),
    .A1(_0439_),
    .B1(_0418_),
    .X(_0443_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _2543_ (.X(_0444_),
    .A(_0414_),
    .B(_0442_),
    .C(_0443_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2544_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0442_),
    .A2(_0443_),
    .Y(_0445_),
    .B1(_0414_));
 sg13g2_nor3_1 _2545_ (.A(_0413_),
    .B(_0444_),
    .C(_0445_),
    .Y(_0446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2546_ (.B1(_0413_),
    .VDD(VPWR),
    .Y(_0447_),
    .VSS(VGND),
    .A1(_0444_),
    .A2(_0445_));
 sg13g2_nor2b_1 _2547_ (.A(_0446_),
    .B_N(_0447_),
    .Y(_0448_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2548_ (.B(_0448_),
    .A(_0412_),
    .X(_0065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2549_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0412_),
    .A2(_0447_),
    .Y(_0449_),
    .B1(_0446_));
 sg13g2_o21ai_1 _2550_ (.B1(_0439_),
    .VDD(VPWR),
    .Y(_0450_),
    .VSS(VGND),
    .A1(_0419_),
    .A2(_0440_));
 sg13g2_o21ai_1 _2551_ (.B1(_0425_),
    .VDD(VPWR),
    .Y(_0451_),
    .VSS(VGND),
    .A1(_0388_),
    .A2(_0423_));
 sg13g2_a22oi_1 _2552_ (.Y(_0452_),
    .B1(net421),
    .B2(net493),
    .A2(net425),
    .A1(net491),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2553_ (.B(net491),
    .C(net425),
    .A(net493),
    .Y(_0453_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net421));
 sg13g2_nor2b_1 _2554_ (.A(_0452_),
    .B_N(_0453_),
    .Y(_0454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2555_ (.Y(_0455_),
    .A(_0451_),
    .B(_0454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2556_ (.Y(_0456_),
    .A(_0451_),
    .B(_0454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2557_ (.A2(_0436_),
    .A1(_0426_),
    .B1(_0434_),
    .X(_0457_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2558_ (.Y(_0458_),
    .A(net489),
    .B(net426),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2559_ (.Y(_0459_),
    .A(net484),
    .B(net427),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2560_ (.Y(_0460_),
    .A(net485),
    .B(net429),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2561_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0461_),
    .B(_0459_),
    .A(_0423_));
 sg13g2_and2_1 _2562_ (.A(_0422_),
    .B(_0460_),
    .X(_0462_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2563_ (.Y(_0463_),
    .A(_0422_),
    .B(_0460_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2564_ (.Y(_0464_),
    .A(_0458_),
    .B(_0463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2565_ (.B1(_0430_),
    .VDD(VPWR),
    .Y(_0465_),
    .VSS(VGND),
    .A1(_0428_),
    .A2(_0431_));
 sg13g2_nand2_1 _2566_ (.Y(_0466_),
    .A(net482),
    .B(net431),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2567_ (.A(net438),
    .B(net480),
    .C(net477),
    .D(net434),
    .X(_0467_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2568_ (.B(net479),
    .C(net477),
    .A(net438),
    .Y(_0468_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net434));
 sg13g2_a22oi_1 _2569_ (.Y(_0469_),
    .B1(net434),
    .B2(net479),
    .A2(net477),
    .A1(net438),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2570_ (.A(_0466_),
    .B(_0467_),
    .C(_0469_),
    .X(_0470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2571_ (.B1(_0466_),
    .VDD(VPWR),
    .Y(_0471_),
    .VSS(VGND),
    .A1(_0467_),
    .A2(_0469_));
 sg13g2_and3_1 _2572_ (.X(_0472_),
    .A(_0465_),
    .B(_0470_),
    .C(_0471_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2573_ (.B(_0470_),
    .C(_0471_),
    .A(_0465_),
    .Y(_0473_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2574_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0470_),
    .A2(_0471_),
    .Y(_0474_),
    .B1(_0465_));
 sg13g2_or3_1 _2575_ (.A(_0464_),
    .B(_0472_),
    .C(_0474_),
    .X(_0475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2576_ (.B1(_0464_),
    .VDD(VPWR),
    .Y(_0476_),
    .VSS(VGND),
    .A1(_0472_),
    .A2(_0474_));
 sg13g2_and3_1 _2577_ (.X(_0477_),
    .A(_0457_),
    .B(_0475_),
    .C(_0476_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2578_ (.B(_0475_),
    .C(_0476_),
    .A(_0457_),
    .Y(_0478_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2579_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0475_),
    .A2(_0476_),
    .Y(_0479_),
    .B1(_0457_));
 sg13g2_or3_1 _2580_ (.A(_0456_),
    .B(_0477_),
    .C(_0479_),
    .X(_0480_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2581_ (.B1(_0456_),
    .VDD(VPWR),
    .Y(_0481_),
    .VSS(VGND),
    .A1(_0477_),
    .A2(_0479_));
 sg13g2_and3_1 _2582_ (.X(_0482_),
    .A(_0450_),
    .B(_0480_),
    .C(_0481_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2583_ (.B(_0480_),
    .C(_0481_),
    .A(_0450_),
    .Y(_0483_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2584_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0480_),
    .A2(_0481_),
    .Y(_0484_),
    .B1(_0450_));
 sg13g2_or3_1 _2585_ (.A(_0417_),
    .B(_0482_),
    .C(_0484_),
    .X(_0485_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2586_ (.B1(_0417_),
    .VDD(VPWR),
    .Y(_0486_),
    .VSS(VGND),
    .A1(_0482_),
    .A2(_0484_));
 sg13g2_and3_1 _2587_ (.X(_0487_),
    .A(_0444_),
    .B(_0485_),
    .C(_0486_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2588_ (.B(_0485_),
    .C(_0486_),
    .A(_0444_),
    .Y(_0488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2589_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0485_),
    .A2(_0486_),
    .Y(_0489_),
    .B1(_0444_));
 sg13g2_nor2_1 _2590_ (.A(_0487_),
    .B(_0489_),
    .Y(_0490_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2591_ (.Y(_0066_),
    .A(_0449_),
    .B(_0490_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2592_ (.B1(_0478_),
    .VDD(VPWR),
    .Y(_0491_),
    .VSS(VGND),
    .A1(_0456_),
    .A2(_0479_));
 sg13g2_o21ai_1 _2593_ (.B1(_0461_),
    .VDD(VPWR),
    .Y(_0492_),
    .VSS(VGND),
    .A1(_0458_),
    .A2(_0462_));
 sg13g2_nand2_1 _2594_ (.Y(_0493_),
    .A(net493),
    .B(net495),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2595_ (.Y(_0494_),
    .A(net489),
    .B(net421),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2596_ (.A(net491),
    .B(net489),
    .C(net425),
    .D(net421),
    .X(_0495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2597_ (.Y(_0496_),
    .B1(net421),
    .B2(net491),
    .A2(net425),
    .A1(net489),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2598_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0497_),
    .B(_0496_),
    .A(_0495_));
 sg13g2_nor2_1 _2599_ (.A(_0493_),
    .B(_0497_),
    .Y(_0498_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2600_ (.B(_0497_),
    .A(_0493_),
    .X(_0499_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2601_ (.Y(_0500_),
    .A(_0492_),
    .B(_0499_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2602_ (.Y(_0501_),
    .A(_0492_),
    .B(_0499_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2603_ (.Y(_0502_),
    .A(_0453_),
    .B(_0501_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2604_ (.B1(_0473_),
    .VDD(VPWR),
    .Y(_0503_),
    .VSS(VGND),
    .A1(_0464_),
    .A2(_0474_));
 sg13g2_nand2_1 _2605_ (.Y(_0504_),
    .A(net487),
    .B(net426),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2606_ (.Y(_0505_),
    .A(net482),
    .B(net427),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2607_ (.Y(_0506_),
    .A(net482),
    .B(net429),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2608_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0507_),
    .B(_0505_),
    .A(_0460_));
 sg13g2_xnor2_1 _2609_ (.Y(_0508_),
    .A(_0459_),
    .B(_0506_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2610_ (.Y(_0509_),
    .A(_0504_),
    .B(_0508_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2611_ (.B1(_0468_),
    .VDD(VPWR),
    .Y(_0510_),
    .VSS(VGND),
    .A1(_0466_),
    .A2(_0469_));
 sg13g2_nand2_1 _2612_ (.Y(_0511_),
    .A(net479),
    .B(net432),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2613_ (.A(net438),
    .B(net477),
    .C(net500),
    .D(net434),
    .X(_0512_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2614_ (.B(net477),
    .C(net500),
    .A(net438),
    .Y(_0513_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net434));
 sg13g2_a22oi_1 _2615_ (.Y(_0514_),
    .B1(net434),
    .B2(net477),
    .A2(net500),
    .A1(net438),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2616_ (.A(_0511_),
    .B(_0512_),
    .C(_0514_),
    .X(_0515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2617_ (.B1(_0511_),
    .VDD(VPWR),
    .Y(_0516_),
    .VSS(VGND),
    .A1(_0512_),
    .A2(_0514_));
 sg13g2_and3_1 _2618_ (.X(_0517_),
    .A(_0510_),
    .B(_0515_),
    .C(_0516_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2619_ (.B(_0515_),
    .C(_0516_),
    .A(_0510_),
    .Y(_0518_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2620_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0515_),
    .A2(_0516_),
    .Y(_0519_),
    .B1(_0510_));
 sg13g2_or3_1 _2621_ (.A(_0509_),
    .B(_0517_),
    .C(_0519_),
    .X(_0520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2622_ (.B1(_0509_),
    .VDD(VPWR),
    .Y(_0521_),
    .VSS(VGND),
    .A1(_0517_),
    .A2(_0519_));
 sg13g2_and3_1 _2623_ (.X(_0522_),
    .A(_0503_),
    .B(_0520_),
    .C(_0521_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2624_ (.B(_0520_),
    .C(_0521_),
    .A(_0503_),
    .Y(_0523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2625_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0520_),
    .A2(_0521_),
    .Y(_0524_),
    .B1(_0503_));
 sg13g2_or3_1 _2626_ (.A(_0502_),
    .B(_0522_),
    .C(_0524_),
    .X(_0525_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2627_ (.B1(_0502_),
    .VDD(VPWR),
    .Y(_0526_),
    .VSS(VGND),
    .A1(_0522_),
    .A2(_0524_));
 sg13g2_and3_1 _2628_ (.X(_0527_),
    .A(_0491_),
    .B(_0525_),
    .C(_0526_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2629_ (.B(_0525_),
    .C(_0526_),
    .A(_0491_),
    .Y(_0528_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2630_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0525_),
    .A2(_0526_),
    .Y(_0529_),
    .B1(_0491_));
 sg13g2_or3_1 _2631_ (.A(_0455_),
    .B(_0527_),
    .C(_0529_),
    .X(_0530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2632_ (.B1(_0455_),
    .VDD(VPWR),
    .Y(_0531_),
    .VSS(VGND),
    .A1(_0527_),
    .A2(_0529_));
 sg13g2_o21ai_1 _2633_ (.B1(_0483_),
    .VDD(VPWR),
    .Y(_0532_),
    .VSS(VGND),
    .A1(_0417_),
    .A2(_0484_));
 sg13g2_nand3_1 _2634_ (.B(_0531_),
    .C(_0532_),
    .A(_0530_),
    .Y(_0533_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2635_ (.A2(_0531_),
    .A1(_0530_),
    .B1(_0532_),
    .X(_0534_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2636_ (.A(_0533_),
    .B(_0534_),
    .X(_0535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2637_ (.B1(_0488_),
    .VDD(VPWR),
    .Y(_0536_),
    .VSS(VGND),
    .A1(_0449_),
    .A2(_0489_));
 sg13g2_nand2_1 _2638_ (.Y(_0537_),
    .A(_0535_),
    .B(_0536_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2639_ (.B(_0536_),
    .A(_0535_),
    .X(_0067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2640_ (.Y(_0538_),
    .A(_0533_),
    .B(_0537_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2641_ (.B1(_0528_),
    .VDD(VPWR),
    .Y(_0539_),
    .VSS(VGND),
    .A1(_0455_),
    .A2(_0529_));
 sg13g2_o21ai_1 _2642_ (.B1(_0500_),
    .VDD(VPWR),
    .Y(_0540_),
    .VSS(VGND),
    .A1(_0453_),
    .A2(_0501_));
 sg13g2_o21ai_1 _2643_ (.B1(_0523_),
    .VDD(VPWR),
    .Y(_0541_),
    .VSS(VGND),
    .A1(_0502_),
    .A2(_0524_));
 sg13g2_nor2_1 _2644_ (.A(_0495_),
    .B(_0498_),
    .Y(_0542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2645_ (.B1(_0507_),
    .VDD(VPWR),
    .Y(_0543_),
    .VSS(VGND),
    .A1(_0504_),
    .A2(_0508_));
 sg13g2_nand2_1 _2646_ (.Y(_0544_),
    .A(net491),
    .B(net495),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2647_ (.Y(_0545_),
    .A(net487),
    .B(net421),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2648_ (.Y(_0546_),
    .A(net487),
    .B(net424),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2649_ (.B(_0546_),
    .A(_0494_),
    .X(_0547_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2650_ (.Y(_0548_),
    .B(_0547_),
    .A_N(_0544_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2651_ (.Y(_0549_),
    .A(_0544_),
    .B(_0547_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2652_ (.Y(_0550_),
    .A(_0543_),
    .B(_0549_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2653_ (.A(_0542_),
    .B(_0550_),
    .Y(_0551_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2654_ (.Y(_0552_),
    .A(_0542_),
    .B(_0550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2655_ (.B1(_0518_),
    .VDD(VPWR),
    .Y(_0553_),
    .VSS(VGND),
    .A1(_0509_),
    .A2(_0519_));
 sg13g2_nand2_1 _2656_ (.Y(_0554_),
    .A(net484),
    .B(net426),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2657_ (.Y(_0555_),
    .A(net479),
    .B(net430),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2658_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0556_),
    .B(_0555_),
    .A(_0505_));
 sg13g2_and2_1 _2659_ (.A(_0505_),
    .B(_0555_),
    .X(_0557_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2660_ (.Y(_0558_),
    .A(_0505_),
    .B(_0555_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2661_ (.Y(_0559_),
    .A(_0554_),
    .B(_0558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2662_ (.B1(_0513_),
    .VDD(VPWR),
    .Y(_0560_),
    .VSS(VGND),
    .A1(_0511_),
    .A2(_0514_));
 sg13g2_nand2_1 _2663_ (.Y(_0561_),
    .A(net501),
    .B(net432),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2664_ (.A(net476),
    .B(net501),
    .C(net435),
    .D(net432),
    .X(_0562_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2665_ (.Y(_0563_),
    .B1(net432),
    .B2(net476),
    .A2(net434),
    .A1(net501),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2666_ (.A(_0562_),
    .B(_0563_),
    .Y(_0564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2667_ (.Y(_0565_),
    .A(_0560_),
    .B(_0564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2668_ (.Y(_0566_),
    .A(_0560_),
    .B(_0564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2669_ (.B(_0566_),
    .A(_0559_),
    .X(_0567_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2670_ (.Y(_0568_),
    .A(_0553_),
    .B(_0567_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2671_ (.Y(_0569_),
    .A(_0553_),
    .B(_0567_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2672_ (.B(_0569_),
    .A(_0552_),
    .X(_0570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2673_ (.Y(_0571_),
    .A(_0541_),
    .B(_0570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2674_ (.Y(_0572_),
    .A(_0541_),
    .B(_0570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2675_ (.Y(_0573_),
    .B(_0540_),
    .A_N(_0572_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2676_ (.Y(_0574_),
    .A(_0540_),
    .B(_0572_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2677_ (.A(_0539_),
    .B(_0574_),
    .Y(_0575_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2678_ (.Y(_0576_),
    .A(_0539_),
    .B(_0574_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2679_ (.Y(_0577_),
    .A(_0539_),
    .B(_0574_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2680_ (.VDD(VPWR),
    .Y(_0578_),
    .A(_0577_),
    .VSS(VGND));
 sg13g2_xnor2_1 _2681_ (.Y(_0068_),
    .A(_0538_),
    .B(_0577_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2682_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0543_),
    .A2(_0549_),
    .Y(_0579_),
    .B1(_0551_));
 sg13g2_o21ai_1 _2683_ (.B1(_0568_),
    .VDD(VPWR),
    .Y(_0580_),
    .VSS(VGND),
    .A1(_0552_),
    .A2(_0569_));
 sg13g2_o21ai_1 _2684_ (.B1(_0548_),
    .VDD(VPWR),
    .Y(_0581_),
    .VSS(VGND),
    .A1(_0494_),
    .A2(_0546_));
 sg13g2_o21ai_1 _2685_ (.B1(_0556_),
    .VDD(VPWR),
    .Y(_0582_),
    .VSS(VGND),
    .A1(_0554_),
    .A2(_0557_));
 sg13g2_nand2_1 _2686_ (.Y(_0583_),
    .A(net489),
    .B(net495),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2687_ (.Y(_0584_),
    .A(net484),
    .B(net421),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2688_ (.Y(_0585_),
    .A(net484),
    .B(net424),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2689_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0586_),
    .B(_0584_),
    .A(_0546_));
 sg13g2_xnor2_1 _2690_ (.Y(_0587_),
    .A(_0545_),
    .B(_0585_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2691_ (.B(_0587_),
    .A(_0583_),
    .X(_0588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2692_ (.Y(_0589_),
    .A(_0582_),
    .B(_0588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2693_ (.A(_0589_),
    .B_N(_0581_),
    .Y(_0590_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2694_ (.B(_0589_),
    .A(_0581_),
    .X(_0591_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2695_ (.B1(_0565_),
    .VDD(VPWR),
    .Y(_0592_),
    .VSS(VGND),
    .A1(_0559_),
    .A2(_0566_));
 sg13g2_a21oi_1 _2696_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net476),
    .A2(net434),
    .Y(_0593_),
    .B1(_0561_));
 sg13g2_nand2_1 _2697_ (.Y(_0594_),
    .A(net481),
    .B(net426),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2698_ (.Y(_0595_),
    .A(net476),
    .B(net428),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2699_ (.A(net479),
    .B(net476),
    .C(net430),
    .D(net428),
    .X(_0596_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2700_ (.Y(_0597_),
    .B1(net428),
    .B2(net479),
    .A2(net430),
    .A1(net476),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2701_ (.A(_0594_),
    .B(_0596_),
    .C(_0597_),
    .Y(_0598_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2702_ (.B1(_0594_),
    .VDD(VPWR),
    .Y(_0599_),
    .VSS(VGND),
    .A1(_0596_),
    .A2(_0597_));
 sg13g2_nor2b_1 _2703_ (.A(_0598_),
    .B_N(_0599_),
    .Y(_0600_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2704_ (.Y(_0601_),
    .A(_0593_),
    .B(_0600_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2705_ (.Y(_0602_),
    .B(_0592_),
    .A_N(_0601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2706_ (.B(_0601_),
    .A(_0592_),
    .X(_0603_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2707_ (.B(_0603_),
    .A(_0591_),
    .X(_0604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2708_ (.Y(_0605_),
    .A(_0580_),
    .B(_0604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2709_ (.B(_0604_),
    .A(_0580_),
    .X(_0606_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2710_ (.Y(_0607_),
    .B(_0606_),
    .A_N(_0579_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2711_ (.B(_0606_),
    .A(_0579_),
    .X(_0608_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2712_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0571_),
    .A2(_0573_),
    .Y(_0609_),
    .B1(_0608_));
 sg13g2_nand3_1 _2713_ (.B(_0573_),
    .C(_0608_),
    .A(_0571_),
    .Y(_0610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2714_ (.Y(_0611_),
    .B(_0610_),
    .A_N(_0609_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2715_ (.B(_0536_),
    .C(_0578_),
    .A(_0535_),
    .Y(_0612_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2716_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0533_),
    .A2(_0576_),
    .Y(_0613_),
    .B1(_0575_));
 sg13g2_inv_1 _2717_ (.VDD(VPWR),
    .Y(_0614_),
    .A(_0613_),
    .VSS(VGND));
 sg13g2_a21oi_1 _2718_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0612_),
    .A2(_0614_),
    .Y(_0615_),
    .B1(_0611_));
 sg13g2_nand3_1 _2719_ (.B(_0612_),
    .C(_0614_),
    .A(_0611_),
    .Y(_0616_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2720_ (.A(_0615_),
    .B_N(_0616_),
    .Y(_0059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2721_ (.A2(_0588_),
    .A1(_0582_),
    .B1(_0590_),
    .X(_0617_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2722_ (.B1(_0602_),
    .VDD(VPWR),
    .Y(_0618_),
    .VSS(VGND),
    .A1(_0591_),
    .A2(_0603_));
 sg13g2_a21o_2 _2723_ (.A2(_0600_),
    .A1(_0593_),
    .B1(_0562_),
    .X(_0619_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2724_ (.Y(_0620_),
    .A(net479),
    .B(net426),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2725_ (.Y(_0621_),
    .A(net500),
    .B(net430),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2726_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0622_),
    .B(_0621_),
    .A(_0595_));
 sg13g2_xnor2_1 _2727_ (.Y(_0623_),
    .A(_0595_),
    .B(_0621_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2728_ (.B(_0623_),
    .A(_0620_),
    .X(_0624_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2729_ (.A(_0619_),
    .B(_0624_),
    .X(_0625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2730_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0626_),
    .B(_0624_),
    .A(_0619_));
 sg13g2_xnor2_1 _2731_ (.Y(_0627_),
    .A(_0619_),
    .B(_0624_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2732_ (.B1(_0586_),
    .VDD(VPWR),
    .Y(_0628_),
    .VSS(VGND),
    .A1(_0583_),
    .A2(_0587_));
 sg13g2_or2_1 _2733_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0629_),
    .B(_0598_),
    .A(_0596_));
 sg13g2_nand2_1 _2734_ (.Y(_0630_),
    .A(net487),
    .B(net495),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2735_ (.Y(_0631_),
    .A(net481),
    .B(net424),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2736_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0632_),
    .B(_0631_),
    .A(_0584_));
 sg13g2_xnor2_1 _2737_ (.Y(_0633_),
    .A(_0584_),
    .B(_0631_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2738_ (.B(_0633_),
    .A(_0630_),
    .X(_0634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2739_ (.Y(_0635_),
    .A(_0629_),
    .B(_0634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2740_ (.A(_0635_),
    .B_N(_0628_),
    .Y(_0636_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2741_ (.Y(_0637_),
    .A(_0628_),
    .B(_0635_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2742_ (.Y(_0638_),
    .A(_0627_),
    .B(_0637_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2743_ (.Y(_0639_),
    .A(_0618_),
    .B(_0638_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2744_ (.A(_0639_),
    .B_N(_0617_),
    .Y(_0640_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2745_ (.B(_0639_),
    .A(_0617_),
    .X(_0641_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2746_ (.B(_0607_),
    .C(_0641_),
    .A(_0605_),
    .Y(_0642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2747_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0605_),
    .A2(_0607_),
    .Y(_0643_),
    .B1(_0641_));
 sg13g2_inv_1 _2748_ (.VDD(VPWR),
    .Y(_0644_),
    .A(_0643_),
    .VSS(VGND));
 sg13g2_nand2_1 _2749_ (.Y(_0645_),
    .A(_0642_),
    .B(_0644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2750_ (.A(_0609_),
    .B(_0615_),
    .Y(_0646_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2751_ (.B(_0646_),
    .A(_0645_),
    .X(_0060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2752_ (.A2(_0634_),
    .A1(_0629_),
    .B1(_0636_),
    .X(_0647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2753_ (.Y(_0648_),
    .B1(\DP_2.matrix[5] ),
    .B2(net476),
    .A2(net428),
    .A1(net500),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2754_ (.Y(_0649_),
    .A(net500),
    .B(\DP_2.matrix[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2755_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0650_),
    .B(_0649_),
    .A(_0595_));
 sg13g2_nand2b_1 _2756_ (.Y(_0651_),
    .B(_0650_),
    .A_N(_0648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2757_ (.B1(_0632_),
    .VDD(VPWR),
    .Y(_0652_),
    .VSS(VGND),
    .A1(_0630_),
    .A2(_0633_));
 sg13g2_o21ai_1 _2758_ (.B1(_0622_),
    .VDD(VPWR),
    .Y(_0653_),
    .VSS(VGND),
    .A1(_0620_),
    .A2(_0623_));
 sg13g2_nand2_1 _2759_ (.Y(_0654_),
    .A(net484),
    .B(net495),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2760_ (.Y(_0655_),
    .A(net480),
    .B(net422),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2761_ (.A(net482),
    .B(net480),
    .C(net424),
    .D(net422),
    .X(_0656_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2762_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0657_),
    .B(_0655_),
    .A(_0631_));
 sg13g2_a22oi_1 _2763_ (.Y(_0658_),
    .B1(net422),
    .B2(net482),
    .A2(net424),
    .A1(net479),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2764_ (.A(_0656_),
    .B(_0658_),
    .Y(_0659_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2765_ (.Y(_0660_),
    .A(_0654_),
    .B(_0659_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2766_ (.Y(_0661_),
    .A(_0653_),
    .B(_0660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2767_ (.A(_0661_),
    .B_N(_0652_),
    .Y(_0662_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2768_ (.B(_0661_),
    .A(_0652_),
    .X(_0663_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2769_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0664_),
    .B(_0663_),
    .A(_0651_));
 sg13g2_xor2_1 _2770_ (.B(_0663_),
    .A(_0651_),
    .X(_0665_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2771_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0626_),
    .A2(_0637_),
    .Y(_0666_),
    .B1(_0625_));
 sg13g2_nor2b_1 _2772_ (.A(_0666_),
    .B_N(_0665_),
    .Y(_0667_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2773_ (.B(_0666_),
    .A(_0665_),
    .X(_0668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2774_ (.A(_0668_),
    .B_N(_0647_),
    .Y(_0669_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2775_ (.B(_0668_),
    .A(_0647_),
    .X(_0670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2776_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0618_),
    .A2(_0638_),
    .Y(_0671_),
    .B1(_0640_));
 sg13g2_nor2_1 _2777_ (.A(_0670_),
    .B(_0671_),
    .Y(_0672_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2778_ (.B(_0671_),
    .A(_0670_),
    .X(_0673_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2779_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0609_),
    .A2(_0642_),
    .Y(_0674_),
    .B1(_0643_));
 sg13g2_nor2b_1 _2780_ (.A(_0613_),
    .B_N(_0674_),
    .Y(_0675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2781_ (.Y(_0676_),
    .A(_0610_),
    .B(_0642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2782_ (.Y(_0677_),
    .B1(_0676_),
    .B2(_0644_),
    .A2(_0675_),
    .A1(_0612_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2783_ (.B(_0677_),
    .A(_0673_),
    .X(_0061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2784_ (.A2(_0660_),
    .A1(_0653_),
    .B1(_0662_),
    .X(_0678_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2785_ (.B1(_0657_),
    .VDD(VPWR),
    .Y(_0679_),
    .VSS(VGND),
    .A1(_0654_),
    .A2(_0658_));
 sg13g2_nand2_1 _2786_ (.Y(_0680_),
    .A(net482),
    .B(net495),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2787_ (.Y(_0681_),
    .A(net477),
    .B(net422),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2788_ (.Y(_0682_),
    .A(net476),
    .B(net424),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2789_ (.B(_0682_),
    .A(_0655_),
    .X(_0683_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2790_ (.Y(_0684_),
    .B(_0683_),
    .A_N(_0680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2791_ (.Y(_0685_),
    .A(_0680_),
    .B(_0683_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2792_ (.A(_0650_),
    .B_N(_0685_),
    .Y(_0686_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2793_ (.Y(_0687_),
    .A(_0650_),
    .B(_0685_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2794_ (.Y(_0688_),
    .A(_0679_),
    .B(_0687_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2795_ (.A(_0649_),
    .B(_0688_),
    .Y(_0689_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2796_ (.Y(_0690_),
    .A(_0649_),
    .B(_0688_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2797_ (.A(_0664_),
    .B(_0690_),
    .Y(_0691_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2798_ (.B(_0690_),
    .A(_0664_),
    .X(_0692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2799_ (.B(_0692_),
    .A(_0678_),
    .X(_0693_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2800_ (.B1(_0693_),
    .VDD(VPWR),
    .Y(_0694_),
    .VSS(VGND),
    .A1(_0667_),
    .A2(_0669_));
 sg13g2_or3_1 _2801_ (.A(_0667_),
    .B(_0669_),
    .C(_0693_),
    .X(_0695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2802_ (.A(_0694_),
    .B(_0695_),
    .X(_0696_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2803_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0673_),
    .A2(_0677_),
    .Y(_0697_),
    .B1(_0672_));
 sg13g2_xnor2_1 _2804_ (.Y(_0062_),
    .A(_0696_),
    .B(_0697_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2805_ (.Y(_0698_),
    .A(_0673_),
    .B(_0696_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2806_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0644_),
    .C1(_0698_),
    .B1(_0676_),
    .A1(_0612_),
    .Y(_0699_),
    .A2(_0675_));
 sg13g2_nand2_1 _2807_ (.Y(_0700_),
    .A(_0672_),
    .B(_0695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2808_ (.Y(_0701_),
    .A(_0694_),
    .B(_0700_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2809_ (.A(_0699_),
    .B(_0701_),
    .Y(_0702_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2810_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0678_),
    .A2(_0692_),
    .Y(_0703_),
    .B1(_0691_));
 sg13g2_a21o_1 _2811_ (.A2(_0687_),
    .A1(_0679_),
    .B1(_0686_),
    .X(_0704_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2812_ (.B1(_0684_),
    .VDD(VPWR),
    .Y(_0705_),
    .VSS(VGND),
    .A1(_0655_),
    .A2(_0682_));
 sg13g2_nand2_1 _2813_ (.Y(_0706_),
    .A(net480),
    .B(\DP_2.matrix[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2814_ (.Y(_0707_),
    .A(net500),
    .B(net421),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2815_ (.Y(_0708_),
    .A(net500),
    .B(net425),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2816_ (.B(_0708_),
    .A(_0681_),
    .X(_0709_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2817_ (.Y(_0710_),
    .B(_0709_),
    .A_N(_0706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2818_ (.Y(_0711_),
    .A(_0706_),
    .B(_0709_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2819_ (.Y(_0712_),
    .A(_0705_),
    .B(_0711_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2820_ (.B(_0711_),
    .A(_0705_),
    .X(_0713_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2821_ (.Y(_0714_),
    .A(_0689_),
    .B(_0713_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2822_ (.A(_0714_),
    .B_N(_0704_),
    .Y(_0715_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2823_ (.B(_0714_),
    .A(_0704_),
    .X(_0716_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2824_ (.B(_0716_),
    .A(_0703_),
    .X(_0717_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2825_ (.B1(_0717_),
    .VDD(VPWR),
    .Y(_0718_),
    .VSS(VGND),
    .A1(_0699_),
    .A2(_0701_));
 sg13g2_xnor2_1 _2826_ (.Y(_0063_),
    .A(_0702_),
    .B(_0717_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2827_ (.B1(_0718_),
    .VDD(VPWR),
    .Y(_0719_),
    .VSS(VGND),
    .A1(_0703_),
    .A2(_0716_));
 sg13g2_a21oi_1 _2828_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0689_),
    .A2(_0713_),
    .Y(_0720_),
    .B1(_0715_));
 sg13g2_o21ai_1 _2829_ (.B1(_0710_),
    .VDD(VPWR),
    .Y(_0721_),
    .VSS(VGND),
    .A1(_0681_),
    .A2(_0708_));
 sg13g2_nand2_1 _2830_ (.Y(_0722_),
    .A(net477),
    .B(\DP_2.matrix[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2831_ (.B(_0722_),
    .A(_0707_),
    .X(_0723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2832_ (.Y(_0724_),
    .A(_0721_),
    .B(_0723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2833_ (.Y(_0725_),
    .A(_0712_),
    .B(_0724_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2834_ (.Y(_0726_),
    .A(_0720_),
    .B(_0725_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2835_ (.Y(_0064_),
    .A(_0719_),
    .B(_0726_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2836_ (.Y(_0727_),
    .A(net474),
    .B(net412),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2837_ (.Y(_0043_),
    .B1(_0727_),
    .B2(_0844_),
    .A2(_0042_),
    .A1(_0845_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2838_ (.Y(_0728_),
    .A(\DP_1.I_range.out_data[3] ),
    .B(\DP_1.Q_range.out_data[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2839_ (.Y(_0729_),
    .B(\DP_1.I_range.out_data[2] ),
    .A_N(\DP_1.Q_range.out_data[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2840_ (.Y(_0730_),
    .A(\DP_1.I_range.out_data[2] ),
    .B(\DP_1.Q_range.out_data[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2841_ (.B(\DP_1.Q_range.out_data[2] ),
    .A(\DP_1.I_range.out_data[2] ),
    .X(_0731_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2842_ (.A(_0728_),
    .B(net379),
    .X(_0732_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2843_ (.Y(_0733_),
    .A(net446),
    .B(_0732_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2844_ (.Y(_0734_),
    .A(_0728_),
    .B(_0729_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2845_ (.VDD(VPWR),
    .Y(_0735_),
    .A(_0734_),
    .VSS(VGND));
 sg13g2_nor2_1 _2846_ (.A(net464),
    .B(net379),
    .Y(_0736_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2847_ (.B1(net376),
    .VDD(VPWR),
    .Y(_0737_),
    .VSS(VGND),
    .A1(net483),
    .A2(_0731_));
 sg13g2_o21ai_1 _2848_ (.B1(_0733_),
    .VDD(VPWR),
    .Y(_0738_),
    .VSS(VGND),
    .A1(_0736_),
    .A2(_0737_));
 sg13g2_mux2_1 _2849_ (.A0(net468),
    .A1(net486),
    .S(net379),
    .X(_0739_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2850_ (.Y(_0740_),
    .B1(net376),
    .B2(_0739_),
    .A2(_0732_),
    .A1(net220),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2851_ (.A0(net474),
    .A1(net492),
    .S(net379),
    .X(_0741_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2852_ (.Y(_0742_),
    .B1(net376),
    .B2(_0741_),
    .A2(_0732_),
    .A1(net458),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2853_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net472),
    .A2(net376),
    .Y(_0743_),
    .B1(net379));
 sg13g2_nor2_1 _2854_ (.A(net456),
    .B(net376),
    .Y(_0744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2855_ (.A(net490),
    .B(_0728_),
    .C(_0731_),
    .Y(_0745_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2856_ (.A(_0743_),
    .B(_0744_),
    .C(_0745_),
    .Y(_0746_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2857_ (.A(_0742_),
    .B_N(_0746_),
    .Y(_0747_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2858_ (.A0(net470),
    .A1(net488),
    .S(net379),
    .X(_0748_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2859_ (.Y(_0749_),
    .B1(net376),
    .B2(_0748_),
    .A2(_0732_),
    .A1(net215),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2860_ (.A(_0749_),
    .B_N(_0747_),
    .Y(_0750_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2861_ (.Y(_0751_),
    .B(_0750_),
    .A_N(_0740_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2862_ (.Y(_0752_),
    .A(net449),
    .B(_0732_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2863_ (.A(net466),
    .B(net379),
    .Y(_0753_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2864_ (.B1(net376),
    .VDD(VPWR),
    .Y(_0754_),
    .VSS(VGND),
    .A1(net485),
    .A2(_0731_));
 sg13g2_o21ai_1 _2865_ (.B1(_0752_),
    .VDD(VPWR),
    .Y(_0755_),
    .VSS(VGND),
    .A1(_0753_),
    .A2(_0754_));
 sg13g2_nand2b_1 _2866_ (.Y(_0756_),
    .B(_0755_),
    .A_N(_0751_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2867_ (.Y(_0757_),
    .B(_0738_),
    .A_N(_0756_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2868_ (.Y(_0758_),
    .A(net443),
    .B(_0732_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2869_ (.A(net463),
    .B(_0730_),
    .Y(_0759_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2870_ (.B1(net376),
    .VDD(VPWR),
    .Y(_0760_),
    .VSS(VGND),
    .A1(\DP_1.matrix[6] ),
    .A2(_0731_));
 sg13g2_o21ai_1 _2871_ (.B1(_0758_),
    .VDD(VPWR),
    .Y(_0761_),
    .VSS(VGND),
    .A1(_0759_),
    .A2(_0760_));
 sg13g2_nor2b_1 _2872_ (.A(_0757_),
    .B_N(_0761_),
    .Y(_0762_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2873_ (.A0(net461),
    .A1(net478),
    .S(_0730_),
    .X(_0763_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2874_ (.Y(_0764_),
    .B1(_0735_),
    .B2(_0763_),
    .A2(_0732_),
    .A1(net441),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2875_ (.Y(_0765_),
    .B(_0762_),
    .A_N(_0764_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2876_ (.A(\DP_1.Q_range.out_data[4] ),
    .B(\DP_1.Q_range.out_data[6] ),
    .Y(_0766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2877_ (.A(\DP_1.I_range.out_data[6] ),
    .B(\DP_1.I_range.out_data[3] ),
    .Y(_0767_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2878_ (.Y(_0768_),
    .A(\DP_1.I_range.out_data[5] ),
    .B(_0767_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2879_ (.A(\DP_1.I_range.out_data[2] ),
    .B(\DP_1.I_range.out_data[4] ),
    .C(\DP_1.Q_range.out_data[2] ),
    .D(_0768_),
    .Y(_0769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _2880_ (.A(\DP_1.Q_range.out_data[3] ),
    .B(\DP_1.Q_range.out_data[5] ),
    .C(_0766_),
    .D(_0769_),
    .X(_0770_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2881_ (.A(net499),
    .B(net379),
    .Y(_0771_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2882_ (.A(net253),
    .B(_0731_),
    .Y(_0772_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2883_ (.A(_0734_),
    .B(_0771_),
    .C(_0772_),
    .Y(_0773_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2884_ (.A(_0773_),
    .B_N(net372),
    .Y(_0774_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2885_ (.Y(_0775_),
    .A(_0765_),
    .B(net372),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2886_ (.A(net371),
    .B_N(net253),
    .Y(_0776_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2887_ (.A(_0774_),
    .B(_0776_),
    .Y(_0777_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2888_ (.Y(_0081_),
    .B1(_0775_),
    .B2(_0777_),
    .A2(_0774_),
    .A1(_0765_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2889_ (.A(\DP_2.Q_range.out_data[2] ),
    .B(_0842_),
    .C(\DP_2.Q_range.out_data[4] ),
    .D(\DP_2.Q_range.out_data[6] ),
    .Y(_0778_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2890_ (.A(\DP_2.I_range.out_data[3] ),
    .B_N(\DP_2.Q_range.out_data[3] ),
    .Y(_0779_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2891_ (.A(\DP_2.Q_range.out_data[2] ),
    .B_N(\DP_2.I_range.out_data[2] ),
    .Y(_0780_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2892_ (.Y(_0781_),
    .A(\DP_2.I_range.out_data[2] ),
    .B(\DP_2.Q_range.out_data[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2893_ (.Y(_0782_),
    .A(\DP_2.I_range.out_data[3] ),
    .B(\DP_2.Q_range.out_data[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2894_ (.A(net378),
    .B(_0782_),
    .X(_0783_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2895_ (.Y(_0784_),
    .A(_0780_),
    .B(_0782_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2896_ (.A0(net402),
    .A1(net423),
    .S(net378),
    .X(_0785_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2897_ (.Y(_0786_),
    .B1(net377),
    .B2(_0785_),
    .A2(_0783_),
    .A1(net381),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2898_ (.A0(net405),
    .A1(net426),
    .S(net378),
    .X(_0787_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2899_ (.Y(_0788_),
    .B1(net377),
    .B2(_0787_),
    .A2(_0783_),
    .A1(net385),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2900_ (.A0(net408),
    .A1(net429),
    .S(net378),
    .X(_0789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2901_ (.Y(_0790_),
    .B1(net377),
    .B2(_0789_),
    .A2(_0783_),
    .A1(net389),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2902_ (.A0(net418),
    .A1(net437),
    .S(net378),
    .X(_0791_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2903_ (.Y(_0792_),
    .B1(net377),
    .B2(_0791_),
    .A2(_0783_),
    .A1(\DP_2.matrix[72] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2904_ (.A(net396),
    .B(net377),
    .Y(_0793_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2905_ (.B1(net378),
    .VDD(VPWR),
    .Y(_0794_),
    .VSS(VGND),
    .A1(net433),
    .A2(_0782_));
 sg13g2_nand3b_1 _2906_ (.B(net377),
    .C(net416),
    .Y(_0795_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net378));
 sg13g2_o21ai_1 _2907_ (.B1(_0795_),
    .VDD(VPWR),
    .Y(_0796_),
    .VSS(VGND),
    .A1(_0793_),
    .A2(_0794_));
 sg13g2_nor2b_1 _2908_ (.A(_0792_),
    .B_N(_0796_),
    .Y(_0797_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2909_ (.A0(net410),
    .A1(net431),
    .S(net378),
    .X(_0798_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2910_ (.Y(_0799_),
    .B1(net377),
    .B2(_0798_),
    .A2(_0783_),
    .A1(net391),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2911_ (.A(_0799_),
    .B_N(_0797_),
    .Y(_0800_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2912_ (.Y(_0801_),
    .B(_0800_),
    .A_N(_0790_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2913_ (.A0(net406),
    .A1(net427),
    .S(_0781_),
    .X(_0802_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2914_ (.Y(_0803_),
    .B1(net377),
    .B2(_0802_),
    .A2(_0783_),
    .A1(net387),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2915_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0804_),
    .B(_0803_),
    .A(_0801_));
 sg13g2_or2_1 _2916_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0805_),
    .B(_0804_),
    .A(_0788_));
 sg13g2_mux2_1 _2917_ (.A0(net404),
    .A1(net424),
    .S(_0781_),
    .X(_0806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2918_ (.Y(_0807_),
    .B1(_0784_),
    .B2(_0806_),
    .A2(_0783_),
    .A1(net383),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2919_ (.A(_0805_),
    .B(_0807_),
    .Y(_0808_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2920_ (.A(_0786_),
    .B(_0805_),
    .C(_0807_),
    .Y(_0809_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2921_ (.A0(\DP_2.matrix[44] ),
    .A1(net495),
    .S(_0781_),
    .X(_0810_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2922_ (.Y(_0811_),
    .B1(_0784_),
    .B2(_0810_),
    .A2(_0783_),
    .A1(net502),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2923_ (.B(_0811_),
    .A(_0809_),
    .X(_0812_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2924_ (.A(\DP_2.I_range.out_data[2] ),
    .B(\DP_2.I_range.out_data[4] ),
    .Y(_0813_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2925_ (.A(\DP_2.I_range.out_data[6] ),
    .B_N(\DP_2.I_range.out_data[5] ),
    .Y(_0814_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2926_ (.B(_0779_),
    .C(_0813_),
    .A(_0778_),
    .Y(_0815_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0814_));
 sg13g2_nand2_1 _2927_ (.Y(_0816_),
    .A(net495),
    .B(net374),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2928_ (.B1(_0816_),
    .VDD(VPWR),
    .Y(_0084_),
    .VSS(VGND),
    .A1(_0812_),
    .A2(net374));
 sg13g2_xor2_1 _2929_ (.B(net373),
    .A(net492),
    .X(_0086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2930_ (.A(net490),
    .B(net373),
    .Y(_0817_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2931_ (.B(_0746_),
    .A(_0742_),
    .X(_0818_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2932_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net373),
    .A2(_0818_),
    .Y(_0087_),
    .B1(net247));
 sg13g2_nor2_1 _2933_ (.A(net488),
    .B(net373),
    .Y(_0819_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2934_ (.B(_0749_),
    .A(_0747_),
    .X(_0820_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2935_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net373),
    .A2(_0820_),
    .Y(_0088_),
    .B1(net250));
 sg13g2_nor2_1 _2936_ (.A(net486),
    .B(net372),
    .Y(_0821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2937_ (.B(_0750_),
    .A(_0740_),
    .X(_0822_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2938_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net372),
    .A2(_0822_),
    .Y(_0089_),
    .B1(_0821_));
 sg13g2_nor2_1 _2939_ (.A(net485),
    .B(net371),
    .Y(_0823_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2940_ (.B(_0755_),
    .A(_0751_),
    .X(_0824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2941_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net371),
    .A2(_0824_),
    .Y(_0090_),
    .B1(_0823_));
 sg13g2_xor2_1 _2942_ (.B(_0756_),
    .A(_0738_),
    .X(_0825_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2943_ (.A(net483),
    .B(net371),
    .Y(_0826_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2944_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net371),
    .A2(_0825_),
    .Y(_0091_),
    .B1(_0826_));
 sg13g2_xor2_1 _2945_ (.B(_0761_),
    .A(_0757_),
    .X(_0827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2946_ (.A(net160),
    .B(net371),
    .Y(_0828_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2947_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net371),
    .A2(_0827_),
    .Y(_0092_),
    .B1(_0828_));
 sg13g2_nand2b_1 _2948_ (.Y(_0829_),
    .B(net478),
    .A_N(net371),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2949_ (.A(_0762_),
    .B_N(_0764_),
    .Y(_0830_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2950_ (.B1(_0829_),
    .VDD(VPWR),
    .Y(_0093_),
    .VSS(VGND),
    .A1(_0775_),
    .A2(_0830_));
 sg13g2_xnor2_1 _2951_ (.Y(_0110_),
    .A(net437),
    .B(net374),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2952_ (.B(_0796_),
    .A(_0792_),
    .X(_0831_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2953_ (.Y(_0832_),
    .A(net433),
    .B(net374),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2954_ (.B1(_0832_),
    .VDD(VPWR),
    .Y(_0111_),
    .VSS(VGND),
    .A1(net374),
    .A2(_0831_));
 sg13g2_xor2_1 _2955_ (.B(_0799_),
    .A(_0797_),
    .X(_0833_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2956_ (.Y(_0834_),
    .A(net431),
    .B(net374),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2957_ (.B1(_0834_),
    .VDD(VPWR),
    .Y(_0112_),
    .VSS(VGND),
    .A1(net374),
    .A2(_0833_));
 sg13g2_xor2_1 _2958_ (.B(_0800_),
    .A(_0790_),
    .X(_0835_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2959_ (.Y(_0836_),
    .A(net429),
    .B(net375),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2960_ (.B1(_0836_),
    .VDD(VPWR),
    .Y(_0113_),
    .VSS(VGND),
    .A1(net374),
    .A2(_0835_));
 sg13g2_xnor2_1 _2961_ (.Y(_0837_),
    .A(_0801_),
    .B(_0803_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2962_ (.Y(_0838_),
    .A(net427),
    .B(net375),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2963_ (.B1(_0838_),
    .VDD(VPWR),
    .Y(_0114_),
    .VSS(VGND),
    .A1(net375),
    .A2(_0837_));
 sg13g2_xor2_1 _2964_ (.B(_0804_),
    .A(_0788_),
    .X(_0839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2965_ (.A0(_0839_),
    .A1(net426),
    .S(net375),
    .X(_0115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2966_ (.B(_0807_),
    .A(_0805_),
    .X(_0840_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2967_ (.A0(_0840_),
    .A1(net424),
    .S(net375),
    .X(_0116_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2968_ (.Y(_0841_),
    .A(_0786_),
    .B(_0808_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2969_ (.A0(_0841_),
    .A1(net423),
    .S(net375),
    .X(_0117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2970_ (.A(net156),
    .X(_0080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2971_ (.A(net499),
    .X(_0082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2972_ (.A(net496),
    .X(_0083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2973_ (.A(net159),
    .X(_0085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2974_ (.A(net474),
    .X(_0094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2975_ (.A(net472),
    .X(_0095_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2976_ (.A(net470),
    .X(_0096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2977_ (.A(net468),
    .X(_0097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2978_ (.A(net467),
    .X(_0098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2979_ (.A(net464),
    .X(_0099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2980_ (.A(net463),
    .X(_0100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2981_ (.A(net459),
    .X(_0101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2982_ (.A(net457),
    .X(_0102_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2983_ (.A(net454),
    .X(_0103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2984_ (.A(net453),
    .X(_0104_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2985_ (.A(net451),
    .X(_0105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2986_ (.A(net448),
    .X(_0106_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2987_ (.A(net445),
    .X(_0107_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2988_ (.A(net155),
    .X(_0108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2989_ (.A(net157),
    .X(_0109_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2990_ (.A(net417),
    .X(_0118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2991_ (.A(net412),
    .X(_0119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2992_ (.A(net410),
    .X(_0120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2993_ (.A(net408),
    .X(_0121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2994_ (.A(net407),
    .X(_0122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2995_ (.A(net158),
    .X(_0123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2996_ (.A(net404),
    .X(_0124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2997_ (.A(net402),
    .X(_0125_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2998_ (.A(net399),
    .X(_0126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2999_ (.A(net394),
    .X(_0127_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3000_ (.A(net391),
    .X(_0128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3001_ (.A(net388),
    .X(_0129_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3002_ (.A(net386),
    .X(_0130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3003_ (.A(net385),
    .X(_0131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3004_ (.A(net383),
    .X(_0132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _3005_ (.A(net381),
    .X(_0133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbpq_1 _3006_ (.RESET_B(net521),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0037_),
    .Q(\mac1.products_ff[0] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _3007_ (.RESET_B(net524),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0038_),
    .Q(\mac1.products_ff[1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _3008_ (.RESET_B(net523),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0039_),
    .Q(\mac1.products_ff[2] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _3009_ (.RESET_B(net525),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0040_),
    .Q(\mac1.products_ff[3] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _3010_ (.RESET_B(net526),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0041_),
    .Q(\mac1.products_ff[4] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _3011_ (.RESET_B(net534),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0058_),
    .Q(\mac1.products_ff[5] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _3012_ (.RESET_B(net535),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0065_),
    .Q(\mac1.products_ff[6] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _3013_ (.RESET_B(net536),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0066_),
    .Q(\mac1.products_ff[7] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _3014_ (.RESET_B(net543),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0067_),
    .Q(\mac1.products_ff[8] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _3015_ (.RESET_B(net546),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0068_),
    .Q(\mac1.products_ff[9] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _3016_ (.RESET_B(net546),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0059_),
    .Q(\mac1.products_ff[10] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _3017_ (.RESET_B(net546),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0060_),
    .Q(\mac1.products_ff[11] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _3018_ (.RESET_B(net546),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0061_),
    .Q(\mac1.products_ff[12] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _3019_ (.RESET_B(net547),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0062_),
    .Q(\mac1.products_ff[13] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _3020_ (.RESET_B(net547),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0063_),
    .Q(\mac1.products_ff[14] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _3021_ (.RESET_B(net547),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0064_),
    .Q(\mac1.products_ff[15] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _3022_ (.RESET_B(net514),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1),
    .Q(\DP_1.I_range.out_data[2] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3023_ (.RESET_B(net514),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2),
    .Q(\DP_1.I_range.out_data[3] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _3024_ (.RESET_B(net514),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3),
    .Q(\DP_1.I_range.out_data[4] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _3025_ (.RESET_B(net514),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\DP_1.I_range.data_plus_4[6] ),
    .Q(\DP_1.I_range.out_data[5] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _3026_ (.RESET_B(net514),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net4),
    .Q(\DP_1.I_range.out_data[6] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _3027_ (.RESET_B(net538),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0080_),
    .Q(\DP_2.matrix[80] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _3028_ (.RESET_B(net531),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0081_),
    .Q(\DP_1.matrix[8] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _3029_ (.RESET_B(net527),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0082_),
    .Q(\DP_1.matrix[44] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _3030_ (.RESET_B(net532),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0083_),
    .Q(\DP_1.matrix[80] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _3031_ (.RESET_B(net538),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net228),
    .Q(\DP_2.matrix[8] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _3032_ (.RESET_B(net548),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0085_),
    .Q(\DP_2.matrix[44] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _3033_ (.RESET_B(net531),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net195),
    .Q(\DP_1.matrix[0] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _3034_ (.RESET_B(net531),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net248),
    .Q(\DP_1.matrix[1] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _3035_ (.RESET_B(net531),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net251),
    .Q(\DP_1.matrix[2] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _3036_ (.RESET_B(net531),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0089_),
    .Q(\DP_1.matrix[3] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3037_ (.RESET_B(net539),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0090_),
    .Q(\DP_1.matrix[4] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3038_ (.RESET_B(net539),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0091_),
    .Q(\DP_1.matrix[5] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _3039_ (.RESET_B(net539),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0092_),
    .Q(\DP_1.matrix[6] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3040_ (.RESET_B(net539),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0093_),
    .Q(\DP_1.matrix[7] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3041_ (.RESET_B(net528),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0094_),
    .Q(\DP_1.matrix[36] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _3042_ (.RESET_B(net527),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0095_),
    .Q(\DP_1.matrix[37] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _3043_ (.RESET_B(net527),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0096_),
    .Q(\DP_1.matrix[38] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _3044_ (.RESET_B(net535),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0097_),
    .Q(\DP_1.matrix[39] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _3045_ (.RESET_B(net543),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0098_),
    .Q(\DP_1.matrix[40] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _3046_ (.RESET_B(net527),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0099_),
    .Q(\DP_1.matrix[41] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _3047_ (.RESET_B(net535),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0100_),
    .Q(\DP_1.matrix[42] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _3048_ (.RESET_B(net537),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0101_),
    .Q(\DP_1.matrix[43] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _3049_ (.RESET_B(net515),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0102_),
    .Q(\DP_1.matrix[72] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _3050_ (.RESET_B(net517),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0103_),
    .Q(\DP_1.matrix[73] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _3051_ (.RESET_B(net517),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0104_),
    .Q(\DP_1.matrix[74] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _3052_ (.RESET_B(net517),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0105_),
    .Q(\DP_1.matrix[75] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _3053_ (.RESET_B(net517),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0106_),
    .Q(\DP_1.matrix[76] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _3054_ (.RESET_B(net519),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0107_),
    .Q(\DP_1.matrix[77] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _3055_ (.RESET_B(net532),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0108_),
    .Q(\DP_1.matrix[78] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _3056_ (.RESET_B(net532),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0109_),
    .Q(\DP_1.matrix[79] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _3057_ (.RESET_B(net531),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net199),
    .Q(\DP_2.matrix[0] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _3058_ (.RESET_B(net531),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net222),
    .Q(\DP_2.matrix[1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3059_ (.RESET_B(net531),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net224),
    .Q(\DP_2.matrix[2] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3060_ (.RESET_B(net538),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net230),
    .Q(\DP_2.matrix[3] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3061_ (.RESET_B(net538),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0114_),
    .Q(\DP_2.matrix[4] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_2 _3062_ (.RESET_B(net539),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0115_),
    .Q(\DP_2.matrix[5] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3063_ (.RESET_B(net538),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0116_),
    .Q(\DP_2.matrix[6] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3064_ (.RESET_B(net539),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0117_),
    .Q(\DP_2.matrix[7] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _3065_ (.RESET_B(net527),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0118_),
    .Q(\DP_2.matrix[36] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _3066_ (.RESET_B(net528),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0119_),
    .Q(\DP_2.matrix[37] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _3067_ (.RESET_B(net527),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0120_),
    .Q(\DP_2.matrix[38] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _3068_ (.RESET_B(net535),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0121_),
    .Q(\DP_2.matrix[39] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _3069_ (.RESET_B(net548),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0122_),
    .Q(\DP_2.matrix[40] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _3070_ (.RESET_B(net548),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0123_),
    .Q(\DP_2.matrix[41] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _3071_ (.RESET_B(net548),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0124_),
    .Q(\DP_2.matrix[42] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _3072_ (.RESET_B(net548),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0125_),
    .Q(\DP_2.matrix[43] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _3073_ (.RESET_B(net518),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0126_),
    .Q(\DP_2.matrix[72] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _3074_ (.RESET_B(net518),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0127_),
    .Q(\DP_2.matrix[73] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _3075_ (.RESET_B(net517),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0128_),
    .Q(\DP_2.matrix[74] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3076_ (.RESET_B(net519),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0129_),
    .Q(\DP_2.matrix[75] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _3077_ (.RESET_B(net519),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0130_),
    .Q(\DP_2.matrix[76] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _3078_ (.RESET_B(net538),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0131_),
    .Q(\DP_2.matrix[77] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _3079_ (.RESET_B(net538),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0132_),
    .Q(\DP_2.matrix[78] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3080_ (.RESET_B(net538),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0133_),
    .Q(\DP_2.matrix[79] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _3081_ (.RESET_B(net521),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0042_),
    .Q(\mac1.products_ff[68] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _3082_ (.RESET_B(net520),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net269),
    .Q(\mac1.products_ff[69] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _3083_ (.RESET_B(net520),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0044_),
    .Q(\mac1.products_ff[70] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _3084_ (.RESET_B(net525),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0045_),
    .Q(\mac1.products_ff[71] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _3085_ (.RESET_B(net525),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0046_),
    .Q(\mac1.products_ff[72] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _3086_ (.RESET_B(net526),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0069_),
    .Q(\mac1.products_ff[73] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _3087_ (.RESET_B(net534),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0076_),
    .Q(\mac1.products_ff[74] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _3088_ (.RESET_B(net536),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0077_),
    .Q(\mac1.products_ff[75] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _3089_ (.RESET_B(net543),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0078_),
    .Q(\mac1.products_ff[76] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _3090_ (.RESET_B(net543),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0079_),
    .Q(\mac1.products_ff[77] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _3091_ (.RESET_B(net542),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0070_),
    .Q(\mac1.products_ff[78] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _3092_ (.RESET_B(net541),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0071_),
    .Q(\mac1.products_ff[79] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _3093_ (.RESET_B(net541),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0072_),
    .Q(\mac1.products_ff[80] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _3094_ (.RESET_B(net541),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0073_),
    .Q(\mac1.products_ff[81] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _3095_ (.RESET_B(net546),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0074_),
    .Q(\mac1.products_ff[82] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _3096_ (.RESET_B(net546),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0075_),
    .Q(\mac1.products_ff[83] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _3097_ (.RESET_B(net507),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0032_),
    .Q(\mac1.products_ff[136] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3098_ (.RESET_B(net503),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0033_),
    .Q(\mac1.products_ff[137] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3099_ (.RESET_B(net508),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0034_),
    .Q(\mac1.products_ff[138] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3100_ (.RESET_B(net508),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0035_),
    .Q(\mac1.products_ff[139] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _3101_ (.RESET_B(net508),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0036_),
    .Q(\mac1.products_ff[140] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _3102_ (.RESET_B(net507),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0047_),
    .Q(\mac1.products_ff[141] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _3103_ (.RESET_B(net512),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0054_),
    .Q(\mac1.products_ff[142] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _3104_ (.RESET_B(net512),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0055_),
    .Q(\mac1.products_ff[143] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3105_ (.RESET_B(net512),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0056_),
    .Q(\mac1.products_ff[144] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3106_ (.RESET_B(net511),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0057_),
    .Q(\mac1.products_ff[145] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3107_ (.RESET_B(net511),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0048_),
    .Q(\mac1.products_ff[146] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3108_ (.RESET_B(net519),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0049_),
    .Q(\mac1.products_ff[147] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _3109_ (.RESET_B(net529),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0050_),
    .Q(\mac1.products_ff[148] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3110_ (.RESET_B(net529),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0051_),
    .Q(\mac1.products_ff[149] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3111_ (.RESET_B(net529),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0052_),
    .Q(\mac1.products_ff[150] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3112_ (.RESET_B(net529),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0053_),
    .Q(\mac1.products_ff[151] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _3113_ (.RESET_B(net521),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net140),
    .Q(\mac1.sum_lvl1_ff[0] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _3114_ (.RESET_B(net520),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net123),
    .Q(\mac1.sum_lvl1_ff[1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _3115_ (.RESET_B(net525),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net150),
    .Q(\mac1.sum_lvl1_ff[2] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _3116_ (.RESET_B(net525),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net133),
    .Q(\mac1.sum_lvl1_ff[3] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _3117_ (.RESET_B(net534),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net95),
    .Q(\mac1.sum_lvl1_ff[4] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _3118_ (.RESET_B(net535),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net61),
    .Q(\mac1.sum_lvl1_ff[5] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _3119_ (.RESET_B(net536),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net87),
    .Q(\mac1.sum_lvl1_ff[6] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _3120_ (.RESET_B(net536),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net106),
    .Q(\mac1.sum_lvl1_ff[7] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _3121_ (.RESET_B(net542),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net96),
    .Q(\mac1.sum_lvl1_ff[8] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _3122_ (.RESET_B(net541),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net152),
    .Q(\mac1.sum_lvl1_ff[9] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _3123_ (.RESET_B(net544),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net151),
    .Q(\mac1.sum_lvl1_ff[10] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _3124_ (.RESET_B(net544),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net45),
    .Q(\mac1.sum_lvl1_ff[11] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _3125_ (.RESET_B(net545),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net130),
    .Q(\mac1.sum_lvl1_ff[12] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _3126_ (.RESET_B(net545),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net117),
    .Q(\mac1.sum_lvl1_ff[13] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _3127_ (.RESET_B(net547),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net121),
    .Q(\mac1.sum_lvl1_ff[14] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _3128_ (.RESET_B(net547),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net127),
    .Q(\mac1.sum_lvl1_ff[15] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _3129_ (.RESET_B(net521),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net137),
    .Q(\mac1.sum_lvl1_ff[36] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _3130_ (.RESET_B(net520),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net143),
    .Q(\mac1.sum_lvl1_ff[37] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _3131_ (.RESET_B(net520),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net74),
    .Q(\mac1.sum_lvl1_ff[38] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _3132_ (.RESET_B(net525),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net69),
    .Q(\mac1.sum_lvl1_ff[39] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _3133_ (.RESET_B(net526),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net135),
    .Q(\mac1.sum_lvl1_ff[40] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _3134_ (.RESET_B(net534),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net73),
    .Q(\mac1.sum_lvl1_ff[41] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _3135_ (.RESET_B(net534),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net62),
    .Q(\mac1.sum_lvl1_ff[42] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _3136_ (.RESET_B(net536),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net43),
    .Q(\mac1.sum_lvl1_ff[43] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _3137_ (.RESET_B(net543),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net81),
    .Q(\mac1.sum_lvl1_ff[44] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _3138_ (.RESET_B(net542),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net84),
    .Q(\mac1.sum_lvl1_ff[45] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _3139_ (.RESET_B(net542),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net82),
    .Q(\mac1.sum_lvl1_ff[46] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _3140_ (.RESET_B(net540),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net67),
    .Q(\mac1.sum_lvl1_ff[47] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _3141_ (.RESET_B(net540),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net53),
    .Q(\mac1.sum_lvl1_ff[48] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _3142_ (.RESET_B(net540),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net47),
    .Q(\mac1.sum_lvl1_ff[49] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _3143_ (.RESET_B(net544),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net63),
    .Q(\mac1.sum_lvl1_ff[50] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _3144_ (.RESET_B(net544),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net85),
    .Q(\mac1.sum_lvl1_ff[51] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _3145_ (.RESET_B(net520),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net118),
    .Q(\mac1.sum_lvl2_ff[0] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _3146_ (.RESET_B(net520),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net145),
    .Q(\mac1.sum_lvl2_ff[1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _3147_ (.RESET_B(net525),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net49),
    .Q(\mac1.sum_lvl2_ff[2] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _3148_ (.RESET_B(net526),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net116),
    .Q(\mac1.sum_lvl2_ff[3] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _3149_ (.RESET_B(net534),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net60),
    .Q(\mac1.sum_lvl2_ff[4] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _3150_ (.RESET_B(net535),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net101),
    .Q(\mac1.sum_lvl2_ff[5] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _3151_ (.RESET_B(net536),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net44),
    .Q(\mac1.sum_lvl2_ff[6] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _3152_ (.RESET_B(net536),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net100),
    .Q(\mac1.sum_lvl2_ff[7] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _3153_ (.RESET_B(net542),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net86),
    .Q(\mac1.sum_lvl2_ff[8] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _3154_ (.RESET_B(net540),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net68),
    .Q(\mac1.sum_lvl2_ff[9] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _3155_ (.RESET_B(net540),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net103),
    .Q(\mac1.sum_lvl2_ff[10] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _3156_ (.RESET_B(net544),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net72),
    .Q(\mac1.sum_lvl2_ff[11] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _3157_ (.RESET_B(net545),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net97),
    .Q(\mac1.sum_lvl2_ff[12] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _3158_ (.RESET_B(net545),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net99),
    .Q(\mac1.sum_lvl2_ff[13] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _3159_ (.RESET_B(net545),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net120),
    .Q(\mac1.sum_lvl2_ff[14] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _3160_ (.RESET_B(net547),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net79),
    .Q(\mac1.sum_lvl2_ff[15] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _3161_ (.RESET_B(net521),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net94),
    .Q(\mac1.sum_lvl2_ff[19] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _3162_ (.RESET_B(net520),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net64),
    .Q(\mac1.sum_lvl2_ff[20] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _3163_ (.RESET_B(net525),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net105),
    .Q(\mac1.sum_lvl2_ff[21] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _3164_ (.RESET_B(net526),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net104),
    .Q(\mac1.sum_lvl2_ff[22] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _3165_ (.RESET_B(net534),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net55),
    .Q(\mac1.sum_lvl2_ff[23] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _3166_ (.RESET_B(net534),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net98),
    .Q(\mac1.sum_lvl2_ff[24] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _3167_ (.RESET_B(net536),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net122),
    .Q(\mac1.sum_lvl2_ff[25] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _3168_ (.RESET_B(net537),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net129),
    .Q(\mac1.sum_lvl2_ff[26] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _3169_ (.RESET_B(net542),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net93),
    .Q(\mac1.sum_lvl2_ff[27] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _3170_ (.RESET_B(net542),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net77),
    .Q(\mac1.sum_lvl2_ff[28] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _3171_ (.RESET_B(net540),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net102),
    .Q(\mac1.sum_lvl2_ff[29] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _3172_ (.RESET_B(net540),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net58),
    .Q(\mac1.sum_lvl2_ff[30] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _3173_ (.RESET_B(net541),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net52),
    .Q(\mac1.sum_lvl2_ff[31] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _3174_ (.RESET_B(net540),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net59),
    .Q(\mac1.sum_lvl2_ff[32] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _3175_ (.RESET_B(net544),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net42),
    .Q(\mac1.sum_lvl2_ff[33] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _3176_ (.RESET_B(net545),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net149),
    .Q(\mac1.sum_lvl2_ff[34] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _3177_ (.RESET_B(net505),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net56),
    .Q(\mac1.sum_lvl2_ff[38] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3178_ (.RESET_B(net505),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net70),
    .Q(\mac1.sum_lvl2_ff[39] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3179_ (.RESET_B(net506),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net147),
    .Q(\mac1.sum_lvl2_ff[40] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3180_ (.RESET_B(net506),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net126),
    .Q(\mac1.sum_lvl2_ff[41] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3181_ (.RESET_B(net509),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net139),
    .Q(\mac1.sum_lvl2_ff[42] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3182_ (.RESET_B(net509),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net134),
    .Q(\mac1.sum_lvl2_ff[43] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3183_ (.RESET_B(net512),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net54),
    .Q(\mac1.sum_lvl2_ff[44] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3184_ (.RESET_B(net511),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net109),
    .Q(\mac1.sum_lvl2_ff[45] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _3185_ (.RESET_B(net511),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net112),
    .Q(\mac1.sum_lvl2_ff[46] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3186_ (.RESET_B(net511),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net78),
    .Q(\mac1.sum_lvl2_ff[47] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3187_ (.RESET_B(net522),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net57),
    .Q(\mac1.sum_lvl2_ff[48] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3188_ (.RESET_B(net522),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net71),
    .Q(\mac1.sum_lvl2_ff[49] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3189_ (.RESET_B(net523),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net132),
    .Q(\mac1.sum_lvl2_ff[50] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _3190_ (.RESET_B(net530),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net83),
    .Q(\mac1.sum_lvl2_ff[51] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3191_ (.RESET_B(net530),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net80),
    .Q(\mac1.sum_lvl2_ff[52] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3192_ (.RESET_B(net529),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net41),
    .Q(\mac1.sum_lvl2_ff[53] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3193_ (.RESET_B(net503),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net131),
    .Q(\mac1.sum_lvl1_ff[72] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3194_ (.RESET_B(net505),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net48),
    .Q(\mac1.sum_lvl1_ff[73] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3195_ (.RESET_B(net505),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net91),
    .Q(\mac1.sum_lvl1_ff[74] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3196_ (.RESET_B(net505),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net128),
    .Q(\mac1.sum_lvl1_ff[75] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3197_ (.RESET_B(net506),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net119),
    .Q(\mac1.sum_lvl1_ff[76] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3198_ (.RESET_B(net512),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net108),
    .Q(\mac1.sum_lvl1_ff[77] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _3199_ (.RESET_B(net512),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net125),
    .Q(\mac1.sum_lvl1_ff[78] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _3200_ (.RESET_B(net512),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net113),
    .Q(\mac1.sum_lvl1_ff[79] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _3201_ (.RESET_B(net512),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net46),
    .Q(\mac1.sum_lvl1_ff[80] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3202_ (.RESET_B(net513),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net88),
    .Q(\mac1.sum_lvl1_ff[81] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3203_ (.RESET_B(net511),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net66),
    .Q(\mac1.sum_lvl1_ff[82] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3204_ (.RESET_B(net522),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net146),
    .Q(\mac1.sum_lvl1_ff[83] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3205_ (.RESET_B(net522),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net107),
    .Q(\mac1.sum_lvl1_ff[84] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3206_ (.RESET_B(net529),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net148),
    .Q(\mac1.sum_lvl1_ff[85] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3207_ (.RESET_B(net530),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net110),
    .Q(\mac1.sum_lvl1_ff[86] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3208_ (.RESET_B(net529),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net51),
    .Q(\mac1.sum_lvl1_ff[87] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _3209_ (.RESET_B(net505),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net50),
    .Q(\mac1.sum_lvl3_ff[20] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3210_ (.RESET_B(net505),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net89),
    .Q(\mac1.sum_lvl3_ff[21] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3211_ (.RESET_B(net509),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net115),
    .Q(\mac1.sum_lvl3_ff[22] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3212_ (.RESET_B(net509),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net141),
    .Q(\mac1.sum_lvl3_ff[23] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3213_ (.RESET_B(net509),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net114),
    .Q(\mac1.sum_lvl3_ff[24] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3214_ (.RESET_B(net509),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net111),
    .Q(\mac1.sum_lvl3_ff[25] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3215_ (.RESET_B(net510),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net138),
    .Q(\mac1.sum_lvl3_ff[26] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3216_ (.RESET_B(net511),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net124),
    .Q(\mac1.sum_lvl3_ff[27] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _3217_ (.RESET_B(net511),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net136),
    .Q(\mac1.sum_lvl3_ff[28] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _3218_ (.RESET_B(net522),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net144),
    .Q(\mac1.sum_lvl3_ff[29] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _3219_ (.RESET_B(net522),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net92),
    .Q(\mac1.sum_lvl3_ff[30] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3220_ (.RESET_B(net522),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net65),
    .Q(\mac1.sum_lvl3_ff[31] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3221_ (.RESET_B(net523),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net90),
    .Q(\mac1.sum_lvl3_ff[32] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _3222_ (.RESET_B(net523),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net142),
    .Q(\mac1.sum_lvl3_ff[33] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _3223_ (.RESET_B(net530),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net75),
    .Q(\mac1.sum_lvl3_ff[34] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3224_ (.RESET_B(net529),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net76),
    .Q(\mac1.sum_lvl3_ff[35] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3225_ (.RESET_B(net505),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net162),
    .Q(\mac1.sum_lvl3_ff[0] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _3226_ (.RESET_B(net509),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net236),
    .Q(\mac1.sum_lvl3_ff[1] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3227_ (.RESET_B(net509),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net256),
    .Q(\mac1.sum_lvl3_ff[2] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3228_ (.RESET_B(net510),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net245),
    .Q(\mac1.sum_lvl3_ff[3] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _3229_ (.RESET_B(net510),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net267),
    .Q(\mac1.sum_lvl3_ff[4] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _3230_ (.RESET_B(net510),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net259),
    .Q(\mac1.sum_lvl3_ff[5] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3231_ (.RESET_B(net510),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net299),
    .Q(\mac1.sum_lvl3_ff[6] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _3232_ (.RESET_B(net521),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0013_),
    .Q(\mac1.sum_lvl3_ff[7] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _3233_ (.RESET_B(net521),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net285),
    .Q(\mac1.sum_lvl3_ff[8] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _3234_ (.RESET_B(net521),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0015_),
    .Q(\mac1.sum_lvl3_ff[9] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _3235_ (.RESET_B(net523),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net303),
    .Q(\mac1.sum_lvl3_ff[10] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _3236_ (.RESET_B(net522),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0002_),
    .Q(\mac1.sum_lvl3_ff[11] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _3237_ (.RESET_B(net527),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0003_),
    .Q(\mac1.sum_lvl3_ff[12] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _3238_ (.RESET_B(net527),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net281),
    .Q(\mac1.sum_lvl3_ff[13] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _3239_ (.RESET_B(net544),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net173),
    .Q(\mac1.sum_lvl3_ff[14] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _3240_ (.RESET_B(net544),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net170),
    .Q(\mac1.sum_lvl3_ff[15] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _3241_ (.RESET_B(net503),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net154),
    .Q(net25),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3242_ (.RESET_B(net503),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net167),
    .Q(net26),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _3243_ (.RESET_B(net503),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net176),
    .Q(net27),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _3244_ (.RESET_B(net503),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net202),
    .Q(net28),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _3245_ (.RESET_B(net503),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net219),
    .Q(net29),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _3246_ (.RESET_B(net503),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net180),
    .Q(net30),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _3247_ (.RESET_B(net504),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net264),
    .Q(net31),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _3248_ (.RESET_B(net504),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net289),
    .Q(net32),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _3249_ (.RESET_B(net504),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net242),
    .Q(net17),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _3250_ (.RESET_B(net504),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net183),
    .Q(net18),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _3251_ (.RESET_B(net507),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net214),
    .Q(net19),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _3252_ (.RESET_B(net507),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net209),
    .Q(net20),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _3253_ (.RESET_B(net507),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net293),
    .Q(net21),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _3254_ (.RESET_B(net507),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net234),
    .Q(net22),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _3255_ (.RESET_B(net507),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net188),
    .Q(net23),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _3256_ (.RESET_B(net507),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net165),
    .Q(net24),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _3257_ (.RESET_B(net514),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net5),
    .Q(\DP_1.Q_range.out_data[2] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _3258_ (.RESET_B(net514),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net6),
    .Q(\DP_1.Q_range.out_data[3] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3259_ (.RESET_B(net514),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net7),
    .Q(\DP_1.Q_range.out_data[4] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3260_ (.RESET_B(net515),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\DP_1.Q_range.data_plus_4[6] ),
    .Q(\DP_1.Q_range.out_data[5] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3261_ (.RESET_B(net515),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net8),
    .Q(\DP_1.Q_range.out_data[6] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _3262_ (.RESET_B(net516),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net13),
    .Q(\DP_2.I_range.out_data[2] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3263_ (.RESET_B(net516),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net14),
    .Q(\DP_2.I_range.out_data[3] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3264_ (.RESET_B(net516),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net15),
    .Q(\DP_2.I_range.out_data[4] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3265_ (.RESET_B(net516),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\DP_2.I_range.data_plus_4[6] ),
    .Q(\DP_2.I_range.out_data[5] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3266_ (.RESET_B(net516),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net16),
    .Q(\DP_2.I_range.out_data[6] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3267_ (.RESET_B(net516),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net9),
    .Q(\DP_2.Q_range.out_data[2] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3268_ (.RESET_B(net516),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net10),
    .Q(\DP_2.Q_range.out_data[3] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3269_ (.RESET_B(net516),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net11),
    .Q(\DP_2.Q_range.out_data[4] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3270_ (.RESET_B(net517),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\DP_2.Q_range.data_plus_4[6] ),
    .Q(\DP_2.Q_range.out_data[5] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3271_ (.RESET_B(net517),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net12),
    .Q(\DP_2.Q_range.out_data[6] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_tiehi heichips25_template_34 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net34));
 sg13g2_tiehi heichips25_template_35 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net35));
 sg13g2_tiehi heichips25_template_36 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net36));
 sg13g2_tiehi heichips25_template_37 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net37));
 sg13g2_tiehi heichips25_template_38 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net38));
 sg13g2_tiehi heichips25_template_39 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net39));
 sg13g2_tiehi heichips25_template_40 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net40));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout371 (.A(net372),
    .X(net371),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout372 (.A(net373),
    .X(net372),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout373 (.A(_0770_),
    .X(net373),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout374 (.A(_0815_),
    .X(net374),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout375 (.A(_0815_),
    .X(net375),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout376 (.A(_0735_),
    .X(net376),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout377 (.A(_0784_),
    .X(net377),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout378 (.A(_0781_),
    .X(net378),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout379 (.A(_0730_),
    .X(net379),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout380 (.A(net381),
    .X(net380),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout381 (.A(net185),
    .X(net381),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout382 (.A(net383),
    .X(net382),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout383 (.A(net184),
    .X(net383),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout384 (.A(net385),
    .X(net384),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout385 (.A(net177),
    .X(net385),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout386 (.A(net387),
    .X(net386),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout387 (.A(net275),
    .X(net387),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout388 (.A(net389),
    .X(net388),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout389 (.A(net273),
    .X(net389),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout390 (.A(net391),
    .X(net390),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout391 (.A(net190),
    .X(net391),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout392 (.A(net393),
    .X(net392),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout393 (.A(net395),
    .X(net393),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout394 (.A(net395),
    .X(net394),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout395 (.A(net396),
    .X(net395),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout396 (.A(\DP_2.matrix[73] ),
    .X(net396),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout397 (.A(net398),
    .X(net397),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout398 (.A(net400),
    .X(net398),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout399 (.A(net400),
    .X(net399),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout400 (.A(net290),
    .X(net400),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout401 (.A(net402),
    .X(net401),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout402 (.A(net192),
    .X(net402),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout403 (.A(net404),
    .X(net403),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout404 (.A(net191),
    .X(net404),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout405 (.A(\DP_2.matrix[41] ),
    .X(net405),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout406 (.A(\DP_2.matrix[40] ),
    .X(net406),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout407 (.A(net238),
    .X(net407),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout408 (.A(net203),
    .X(net408),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout409 (.A(\DP_2.matrix[39] ),
    .X(net409),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout410 (.A(net197),
    .X(net410),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout411 (.A(\DP_2.matrix[38] ),
    .X(net411),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout412 (.A(net416),
    .X(net412),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout413 (.A(net416),
    .X(net413),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout414 (.A(net416),
    .X(net414),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout415 (.A(net416),
    .X(net415),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout416 (.A(net268),
    .X(net416),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout417 (.A(net418),
    .X(net417),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout418 (.A(net270),
    .X(net418),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout419 (.A(\DP_2.matrix[36] ),
    .X(net419),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout420 (.A(\DP_2.matrix[36] ),
    .X(net420),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout421 (.A(net423),
    .X(net421),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout422 (.A(net423),
    .X(net422),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout423 (.A(net252),
    .X(net423),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout424 (.A(net425),
    .X(net424),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout425 (.A(net300),
    .X(net425),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout426 (.A(net282),
    .X(net426),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout427 (.A(net237),
    .X(net427),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout428 (.A(\DP_2.matrix[4] ),
    .X(net428),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout429 (.A(net229),
    .X(net429),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout430 (.A(\DP_2.matrix[3] ),
    .X(net430),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout431 (.A(net223),
    .X(net431),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout432 (.A(\DP_2.matrix[2] ),
    .X(net432),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout433 (.A(net221),
    .X(net433),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout434 (.A(net435),
    .X(net434),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout435 (.A(net436),
    .X(net435),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout436 (.A(\DP_2.matrix[1] ),
    .X(net436),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout437 (.A(net198),
    .X(net437),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout438 (.A(net439),
    .X(net438),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout439 (.A(\DP_2.matrix[0] ),
    .X(net439),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout440 (.A(net441),
    .X(net440),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout441 (.A(\DP_1.matrix[79] ),
    .X(net441),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout442 (.A(net443),
    .X(net442),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout443 (.A(\DP_1.matrix[78] ),
    .X(net443),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout444 (.A(net445),
    .X(net444),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout445 (.A(net446),
    .X(net445),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout446 (.A(net286),
    .X(net446),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout447 (.A(net448),
    .X(net447),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout448 (.A(net449),
    .X(net448),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout449 (.A(net272),
    .X(net449),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout450 (.A(net451),
    .X(net450),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout451 (.A(net220),
    .X(net451),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout452 (.A(net453),
    .X(net452),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout453 (.A(net215),
    .X(net453),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout454 (.A(net456),
    .X(net454),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout455 (.A(net456),
    .X(net455),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout456 (.A(net271),
    .X(net456),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout457 (.A(net458),
    .X(net457),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout458 (.A(net277),
    .X(net458),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout459 (.A(net461),
    .X(net459),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout460 (.A(net461),
    .X(net460),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout461 (.A(net274),
    .X(net461),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout462 (.A(net463),
    .X(net462),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout463 (.A(net211),
    .X(net463),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout464 (.A(net204),
    .X(net464),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout465 (.A(\DP_1.matrix[41] ),
    .X(net465),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout466 (.A(\DP_1.matrix[40] ),
    .X(net466),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout467 (.A(net210),
    .X(net467),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout468 (.A(net212),
    .X(net468),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout469 (.A(\DP_1.matrix[39] ),
    .X(net469),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout470 (.A(net205),
    .X(net470),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout471 (.A(\DP_1.matrix[38] ),
    .X(net471),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout472 (.A(net473),
    .X(net472),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout473 (.A(net276),
    .X(net473),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout474 (.A(net196),
    .X(net474),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout475 (.A(\DP_1.matrix[36] ),
    .X(net475),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout476 (.A(net478),
    .X(net476),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout477 (.A(net478),
    .X(net477),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout478 (.A(net216),
    .X(net478),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout479 (.A(net480),
    .X(net479),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout480 (.A(\DP_1.matrix[6] ),
    .X(net480),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout481 (.A(net483),
    .X(net481),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout482 (.A(net483),
    .X(net482),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout483 (.A(net225),
    .X(net483),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout484 (.A(net485),
    .X(net484),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout485 (.A(net226),
    .X(net485),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout486 (.A(net260),
    .X(net486),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout487 (.A(\DP_1.matrix[3] ),
    .X(net487),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout488 (.A(net249),
    .X(net488),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout489 (.A(\DP_1.matrix[2] ),
    .X(net489),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout490 (.A(net246),
    .X(net490),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout491 (.A(\DP_1.matrix[1] ),
    .X(net491),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout492 (.A(net194),
    .X(net492),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout493 (.A(\DP_1.matrix[0] ),
    .X(net493),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout494 (.A(\DP_2.matrix[44] ),
    .X(net494),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout495 (.A(net227),
    .X(net495),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout496 (.A(net193),
    .X(net496),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout497 (.A(\DP_1.matrix[80] ),
    .X(net497),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout498 (.A(net499),
    .X(net498),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout499 (.A(net189),
    .X(net499),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout500 (.A(net501),
    .X(net500),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout501 (.A(\DP_1.matrix[8] ),
    .X(net501),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout502 (.A(\DP_2.matrix[80] ),
    .X(net502),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout503 (.A(net506),
    .X(net503),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout504 (.A(net506),
    .X(net504),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout505 (.A(net506),
    .X(net505),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout506 (.A(net508),
    .X(net506),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout507 (.A(net508),
    .X(net507),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout508 (.A(net533),
    .X(net508),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout509 (.A(net513),
    .X(net509),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout510 (.A(net513),
    .X(net510),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout511 (.A(net513),
    .X(net511),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout512 (.A(net513),
    .X(net512),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout513 (.A(net533),
    .X(net513),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout514 (.A(net515),
    .X(net514),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout515 (.A(net518),
    .X(net515),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout516 (.A(net517),
    .X(net516),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout517 (.A(net518),
    .X(net517),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout518 (.A(net519),
    .X(net518),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout519 (.A(net533),
    .X(net519),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout520 (.A(net524),
    .X(net520),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout521 (.A(net524),
    .X(net521),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout522 (.A(net524),
    .X(net522),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout523 (.A(net524),
    .X(net523),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout524 (.A(net533),
    .X(net524),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout525 (.A(net528),
    .X(net525),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout526 (.A(net528),
    .X(net526),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout527 (.A(net528),
    .X(net527),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout528 (.A(net533),
    .X(net528),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout529 (.A(net532),
    .X(net529),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout530 (.A(net532),
    .X(net530),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout531 (.A(net532),
    .X(net531),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout532 (.A(net533),
    .X(net532),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout533 (.A(rst_n),
    .X(net533),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout534 (.A(net535),
    .X(net534),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout535 (.A(net537),
    .X(net535),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout536 (.A(net537),
    .X(net536),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout537 (.A(net549),
    .X(net537),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout538 (.A(net539),
    .X(net538),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout539 (.A(net549),
    .X(net539),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout540 (.A(net541),
    .X(net540),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout541 (.A(net542),
    .X(net541),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout542 (.A(net543),
    .X(net542),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout543 (.A(net549),
    .X(net543),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout544 (.A(net546),
    .X(net544),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout545 (.A(net546),
    .X(net545),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout546 (.A(net547),
    .X(net546),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout547 (.A(net548),
    .X(net547),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout548 (.A(net549),
    .X(net548),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout549 (.A(rst_n),
    .X(net549),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input14 (.A(uio_in[5]),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input16 (.A(uio_in[7]),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uio_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uio_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uio_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uio_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uo_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uo_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uo_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output30 (.A(net30),
    .X(uo_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output31 (.A(net31),
    .X(uo_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output32 (.A(net32),
    .X(uo_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tiehi heichips25_template_33 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net33));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_2_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_3_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_4_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_6_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_7_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_8_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_9_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_10_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_11_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_12_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_13_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_14_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_16_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_22_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_23_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_24_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_25_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_26_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_27_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_28_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_29_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_30_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_31_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_32_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_33_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_34_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_35_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_36_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_37_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_38_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload0 (.A(clknet_3_6__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload1 (.A(clknet_3_7__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_8 clkload2 (.A(clknet_leaf_1_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload3 (.A(clknet_leaf_38_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_8 clkload4 (.A(clknet_leaf_2_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload5 (.VDD(VPWR),
    .A(clknet_leaf_8_clk),
    .VSS(VGND));
 sg13g2_inv_4 clkload6 (.A(clknet_leaf_7_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_12_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload8 (.VDD(VPWR),
    .A(clknet_leaf_22_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload9 (.VDD(VPWR),
    .A(clknet_leaf_25_clk),
    .VSS(VGND));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_29_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload11 (.VDD(VPWR),
    .A(clknet_leaf_18_clk),
    .VSS(VGND));
 sg13g2_inv_4 clkload12 (.A(clknet_leaf_21_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_20_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd3_1 hold1 (.A(\mac1.sum_lvl1_ff[87] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold2 (.A(\mac1.sum_lvl1_ff[50] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold3 (.A(\mac1.products_ff[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold4 (.A(\mac1.sum_lvl1_ff[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold5 (.A(\mac1.products_ff[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold6 (.A(\mac1.products_ff[144] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold7 (.A(\mac1.products_ff[81] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold8 (.A(\mac1.products_ff[137] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold9 (.A(\mac1.sum_lvl1_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold10 (.A(\mac1.sum_lvl2_ff[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold11 (.A(\mac1.products_ff[151] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold12 (.A(\mac1.sum_lvl1_ff[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold13 (.A(\mac1.products_ff[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold14 (.A(\mac1.sum_lvl1_ff[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold15 (.A(\mac1.sum_lvl1_ff[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold16 (.A(\mac1.sum_lvl1_ff[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold17 (.A(\mac1.sum_lvl1_ff[82] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold18 (.A(\mac1.sum_lvl1_ff[47] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold19 (.A(\mac1.sum_lvl1_ff[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold20 (.A(\mac1.sum_lvl1_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold21 (.A(\mac1.products_ff[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold22 (.A(\mac1.products_ff[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold23 (.A(\mac1.products_ff[82] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold24 (.A(\mac1.sum_lvl1_ff[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold25 (.A(\mac1.sum_lvl2_ff[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold26 (.A(\mac1.products_ff[146] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold27 (.A(\mac1.products_ff[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold28 (.A(\mac1.sum_lvl1_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold29 (.A(\mac1.products_ff[71] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold30 (.A(\mac1.sum_lvl1_ff[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold31 (.A(\mac1.sum_lvl1_ff[83] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold32 (.A(\mac1.sum_lvl1_ff[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold33 (.A(\mac1.products_ff[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold34 (.A(\mac1.products_ff[70] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold35 (.A(\mac1.sum_lvl2_ff[52] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold36 (.A(\mac1.sum_lvl2_ff[53] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold37 (.A(\mac1.sum_lvl1_ff[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold38 (.A(\mac1.sum_lvl1_ff[81] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold39 (.A(\mac1.sum_lvl1_ff[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold40 (.A(\mac1.sum_lvl1_ff[86] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold41 (.A(\mac1.products_ff[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold42 (.A(\mac1.products_ff[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold43 (.A(\mac1.sum_lvl1_ff[85] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold44 (.A(\mac1.products_ff[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold45 (.A(\mac1.products_ff[83] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold46 (.A(\mac1.sum_lvl1_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold47 (.A(\mac1.products_ff[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold48 (.A(\mac1.products_ff[145] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold49 (.A(\mac1.sum_lvl2_ff[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold50 (.A(\mac1.sum_lvl2_ff[50] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold51 (.A(\mac1.products_ff[138] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold52 (.A(\mac1.sum_lvl2_ff[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold53 (.A(\mac1.sum_lvl1_ff[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold54 (.A(\mac1.sum_lvl1_ff[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold55 (.A(\mac1.products_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold56 (.A(\mac1.products_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold57 (.A(\mac1.sum_lvl1_ff[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold58 (.A(\mac1.sum_lvl1_ff[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold59 (.A(\mac1.sum_lvl1_ff[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold60 (.A(\mac1.sum_lvl1_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold61 (.A(\mac1.sum_lvl1_ff[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold62 (.A(\mac1.sum_lvl1_ff[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold63 (.A(\mac1.sum_lvl1_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold64 (.A(\mac1.sum_lvl1_ff[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold65 (.A(\mac1.sum_lvl1_ff[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold66 (.A(\mac1.products_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold67 (.A(\mac1.products_ff[148] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold68 (.A(\mac1.products_ff[141] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold69 (.A(\mac1.sum_lvl1_ff[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold70 (.A(\mac1.products_ff[150] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold71 (.A(\mac1.sum_lvl2_ff[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold72 (.A(\mac1.sum_lvl1_ff[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold73 (.A(\mac1.products_ff[143] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold74 (.A(\mac1.sum_lvl2_ff[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold75 (.A(\mac1.sum_lvl2_ff[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold76 (.A(\mac1.sum_lvl1_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold77 (.A(\mac1.products_ff[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold78 (.A(\mac1.sum_lvl1_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold79 (.A(\mac1.products_ff[140] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold80 (.A(\mac1.sum_lvl1_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold81 (.A(\mac1.products_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold82 (.A(\mac1.sum_lvl1_ff[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold83 (.A(\mac1.products_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold84 (.A(\mac1.sum_lvl2_ff[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold85 (.A(\mac1.products_ff[142] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold86 (.A(\mac1.sum_lvl1_ff[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold87 (.A(\mac1.products_ff[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold88 (.A(\mac1.products_ff[139] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold89 (.A(\mac1.sum_lvl1_ff[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold90 (.A(\mac1.products_ff[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold91 (.A(\mac1.products_ff[136] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold92 (.A(\mac1.sum_lvl1_ff[84] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold93 (.A(\mac1.products_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold94 (.A(\mac1.sum_lvl1_ff[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold95 (.A(\mac1.products_ff[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold96 (.A(\mac1.sum_lvl2_ff[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold97 (.A(\mac1.products_ff[68] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold98 (.A(\mac1.sum_lvl2_ff[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold99 (.A(\mac1.sum_lvl1_ff[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold100 (.A(\mac1.products_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold101 (.A(\mac1.sum_lvl2_ff[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold102 (.A(\mac1.sum_lvl2_ff[51] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold103 (.A(\mac1.products_ff[69] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold104 (.A(\mac1.sum_lvl2_ff[47] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold105 (.A(\mac1.sum_lvl1_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold106 (.A(\mac1.products_ff[147] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold107 (.A(\mac1.sum_lvl1_ff[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold108 (.A(\mac1.products_ff[149] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold109 (.A(\mac1.sum_lvl1_ff[51] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold110 (.A(\mac1.products_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold111 (.A(\mac1.products_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold112 (.A(\mac1.products_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold113 (.A(\mac1.sum_lvl3_ff[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0016_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold115 (.A(\DP_1.matrix[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold116 (.A(\DP_2.matrix[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold117 (.A(\DP_1.matrix[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold118 (.A(\DP_2.matrix[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold119 (.A(\DP_2.matrix[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold120 (.A(\DP_1.matrix[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold121 (.A(\mac1.sum_lvl2_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0000_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold123 (.A(\mac1.sum_lvl3_ff[35] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold124 (.A(_1338_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0022_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold126 (.A(\mac1.sum_lvl3_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0023_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold128 (.A(\mac1.sum_lvl2_ff[34] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold129 (.A(_1281_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0006_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold131 (.A(\mac1.sum_lvl2_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold132 (.A(_1279_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0005_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold134 (.A(\mac1.sum_lvl3_ff[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold135 (.A(_1288_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0024_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold137 (.A(\DP_2.matrix[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold138 (.A(\mac1.sum_lvl3_ff[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold139 (.A(_1297_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0027_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold141 (.A(\mac1.sum_lvl3_ff[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold142 (.A(_1313_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0031_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold144 (.A(\DP_2.matrix[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold145 (.A(\DP_2.matrix[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold146 (.A(\mac1.sum_lvl3_ff[34] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold147 (.A(_1336_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0021_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold149 (.A(\DP_1.matrix[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold150 (.A(\DP_2.matrix[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold151 (.A(\DP_2.matrix[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold152 (.A(\DP_2.matrix[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold153 (.A(\DP_1.matrix[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold154 (.A(\DP_1.matrix[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0086_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold156 (.A(\DP_1.matrix[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold157 (.A(\DP_2.matrix[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold158 (.A(\DP_2.matrix[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0110_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold160 (.A(\mac1.sum_lvl3_ff[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold161 (.A(_1291_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0025_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold163 (.A(\DP_2.matrix[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold164 (.A(\DP_1.matrix[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold165 (.A(\DP_1.matrix[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold166 (.A(\mac1.sum_lvl3_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold167 (.A(_1316_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold168 (.A(_1322_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0018_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold170 (.A(\DP_1.matrix[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold171 (.A(\DP_1.matrix[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold172 (.A(\DP_1.matrix[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold173 (.A(\mac1.sum_lvl3_ff[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0017_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold175 (.A(\DP_1.matrix[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold176 (.A(\DP_1.matrix[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold177 (.A(\mac1.sum_lvl3_ff[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold178 (.A(_1294_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0026_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold180 (.A(\DP_1.matrix[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold181 (.A(\DP_2.matrix[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0111_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold183 (.A(\DP_2.matrix[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0112_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold185 (.A(\DP_1.matrix[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold186 (.A(\DP_1.matrix[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold187 (.A(\DP_2.matrix[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0084_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold189 (.A(\DP_2.matrix[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0113_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold191 (.A(\mac1.sum_lvl3_ff[33] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold192 (.A(_1330_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold193 (.A(_1331_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0020_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold195 (.A(\mac1.sum_lvl2_ff[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0007_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold197 (.A(\DP_2.matrix[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold198 (.A(\DP_2.matrix[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold199 (.A(\mac1.sum_lvl3_ff[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold200 (.A(_1303_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold201 (.A(_1310_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0030_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold203 (.A(\mac1.sum_lvl2_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold204 (.A(_1234_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0009_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold206 (.A(\DP_1.matrix[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0817_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0087_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold209 (.A(\DP_1.matrix[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0819_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0088_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold212 (.A(\DP_2.matrix[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold213 (.A(\DP_1.matrix[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold214 (.A(\mac1.sum_lvl2_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold215 (.A(_1231_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0008_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold217 (.A(\mac1.sum_lvl2_ff[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold218 (.A(_1240_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0011_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold220 (.A(\DP_1.matrix[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold221 (.A(\mac1.sum_lvl3_ff[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold222 (.A(_1299_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold223 (.A(_1302_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0028_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold225 (.A(\mac1.sum_lvl2_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold226 (.A(_1237_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0010_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold228 (.A(\DP_2.matrix[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0043_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold230 (.A(\DP_2.matrix[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold231 (.A(\DP_1.matrix[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold232 (.A(\DP_1.matrix[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold233 (.A(\DP_2.matrix[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold234 (.A(\DP_1.matrix[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold235 (.A(\DP_2.matrix[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold236 (.A(\DP_1.matrix[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold237 (.A(\DP_1.matrix[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold238 (.A(\mac1.sum_lvl2_ff[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold239 (.A(_1266_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold240 (.A(_1275_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0004_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold242 (.A(\DP_2.matrix[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold243 (.A(\mac1.sum_lvl2_ff[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold244 (.A(_1246_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0014_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold246 (.A(\DP_1.matrix[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold247 (.A(\mac1.sum_lvl3_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold248 (.A(_1305_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0029_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold250 (.A(\DP_2.matrix[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold251 (.A(\mac1.sum_lvl3_ff[32] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold252 (.A(_1324_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0019_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold254 (.A(\mac1.sum_lvl2_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold255 (.A(_1256_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold256 (.A(\mac1.sum_lvl2_ff[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold257 (.A(_1242_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold258 (.A(_1245_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold259 (.A(_0012_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold260 (.A(\DP_2.matrix[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold261 (.A(\mac1.sum_lvl2_ff[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold262 (.A(_1260_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0001_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold264 (.A(\mac1.sum_lvl2_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold265 (.A(_1247_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net305));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_6 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_1028 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net33;
 assign uio_oe[1] = net34;
 assign uio_oe[2] = net35;
 assign uio_oe[3] = net36;
 assign uio_oe[4] = net37;
 assign uio_oe[5] = net38;
 assign uio_oe[6] = net39;
 assign uio_oe[7] = net40;
endmodule
