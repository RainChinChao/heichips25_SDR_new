module heichips25_template (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \DP_1.I_range.data_plus_4[6] ;
 wire \DP_1.I_range.out_data[2] ;
 wire \DP_1.I_range.out_data[3] ;
 wire \DP_1.I_range.out_data[4] ;
 wire \DP_1.I_range.out_data[5] ;
 wire \DP_1.I_range.out_data[6] ;
 wire \DP_1.Q_range.data_plus_4[6] ;
 wire \DP_1.Q_range.out_data[2] ;
 wire \DP_1.Q_range.out_data[3] ;
 wire \DP_1.Q_range.out_data[4] ;
 wire \DP_1.Q_range.out_data[5] ;
 wire \DP_1.Q_range.out_data[6] ;
 wire \DP_1.matrix[0] ;
 wire \DP_1.matrix[1] ;
 wire \DP_1.matrix[2] ;
 wire \DP_1.matrix[36] ;
 wire \DP_1.matrix[37] ;
 wire \DP_1.matrix[38] ;
 wire \DP_1.matrix[39] ;
 wire \DP_1.matrix[3] ;
 wire \DP_1.matrix[40] ;
 wire \DP_1.matrix[41] ;
 wire \DP_1.matrix[42] ;
 wire \DP_1.matrix[43] ;
 wire \DP_1.matrix[44] ;
 wire \DP_1.matrix[4] ;
 wire \DP_1.matrix[5] ;
 wire \DP_1.matrix[6] ;
 wire \DP_1.matrix[72] ;
 wire \DP_1.matrix[73] ;
 wire \DP_1.matrix[74] ;
 wire \DP_1.matrix[75] ;
 wire \DP_1.matrix[76] ;
 wire \DP_1.matrix[77] ;
 wire \DP_1.matrix[78] ;
 wire \DP_1.matrix[79] ;
 wire \DP_1.matrix[7] ;
 wire \DP_1.matrix[80] ;
 wire \DP_1.matrix[8] ;
 wire \DP_2.matrix[0] ;
 wire \DP_2.matrix[1] ;
 wire \DP_2.matrix[2] ;
 wire \DP_2.matrix[36] ;
 wire \DP_2.matrix[37] ;
 wire \DP_2.matrix[38] ;
 wire \DP_2.matrix[39] ;
 wire \DP_2.matrix[3] ;
 wire \DP_2.matrix[40] ;
 wire \DP_2.matrix[41] ;
 wire \DP_2.matrix[42] ;
 wire \DP_2.matrix[43] ;
 wire \DP_2.matrix[44] ;
 wire \DP_2.matrix[4] ;
 wire \DP_2.matrix[5] ;
 wire \DP_2.matrix[6] ;
 wire \DP_2.matrix[72] ;
 wire \DP_2.matrix[73] ;
 wire \DP_2.matrix[74] ;
 wire \DP_2.matrix[75] ;
 wire \DP_2.matrix[76] ;
 wire \DP_2.matrix[77] ;
 wire \DP_2.matrix[78] ;
 wire \DP_2.matrix[79] ;
 wire \DP_2.matrix[7] ;
 wire \DP_2.matrix[80] ;
 wire \DP_2.matrix[8] ;
 wire \DP_3.I_range.data_plus_4[6] ;
 wire \DP_3.I_range.out_data[2] ;
 wire \DP_3.I_range.out_data[3] ;
 wire \DP_3.I_range.out_data[4] ;
 wire \DP_3.I_range.out_data[5] ;
 wire \DP_3.I_range.out_data[6] ;
 wire \DP_3.Q_range.data_plus_4[6] ;
 wire \DP_3.Q_range.out_data[2] ;
 wire \DP_3.Q_range.out_data[3] ;
 wire \DP_3.Q_range.out_data[4] ;
 wire \DP_3.Q_range.out_data[5] ;
 wire \DP_3.Q_range.out_data[6] ;
 wire \DP_3.matrix[0] ;
 wire \DP_3.matrix[1] ;
 wire \DP_3.matrix[2] ;
 wire \DP_3.matrix[36] ;
 wire \DP_3.matrix[37] ;
 wire \DP_3.matrix[38] ;
 wire \DP_3.matrix[39] ;
 wire \DP_3.matrix[3] ;
 wire \DP_3.matrix[40] ;
 wire \DP_3.matrix[41] ;
 wire \DP_3.matrix[42] ;
 wire \DP_3.matrix[43] ;
 wire \DP_3.matrix[44] ;
 wire \DP_3.matrix[4] ;
 wire \DP_3.matrix[5] ;
 wire \DP_3.matrix[6] ;
 wire \DP_3.matrix[72] ;
 wire \DP_3.matrix[73] ;
 wire \DP_3.matrix[74] ;
 wire \DP_3.matrix[75] ;
 wire \DP_3.matrix[76] ;
 wire \DP_3.matrix[77] ;
 wire \DP_3.matrix[78] ;
 wire \DP_3.matrix[79] ;
 wire \DP_3.matrix[7] ;
 wire \DP_3.matrix[80] ;
 wire \DP_3.matrix[8] ;
 wire \DP_4.matrix[0] ;
 wire \DP_4.matrix[1] ;
 wire \DP_4.matrix[2] ;
 wire \DP_4.matrix[36] ;
 wire \DP_4.matrix[37] ;
 wire \DP_4.matrix[38] ;
 wire \DP_4.matrix[39] ;
 wire \DP_4.matrix[3] ;
 wire \DP_4.matrix[40] ;
 wire \DP_4.matrix[41] ;
 wire \DP_4.matrix[42] ;
 wire \DP_4.matrix[43] ;
 wire \DP_4.matrix[44] ;
 wire \DP_4.matrix[4] ;
 wire \DP_4.matrix[5] ;
 wire \DP_4.matrix[6] ;
 wire \DP_4.matrix[72] ;
 wire \DP_4.matrix[73] ;
 wire \DP_4.matrix[74] ;
 wire \DP_4.matrix[75] ;
 wire \DP_4.matrix[76] ;
 wire \DP_4.matrix[77] ;
 wire \DP_4.matrix[78] ;
 wire \DP_4.matrix[79] ;
 wire \DP_4.matrix[7] ;
 wire \DP_4.matrix[80] ;
 wire \DP_4.matrix[8] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire \mac1.products_ff[0] ;
 wire \mac1.products_ff[10] ;
 wire \mac1.products_ff[11] ;
 wire \mac1.products_ff[12] ;
 wire \mac1.products_ff[136] ;
 wire \mac1.products_ff[137] ;
 wire \mac1.products_ff[138] ;
 wire \mac1.products_ff[139] ;
 wire \mac1.products_ff[13] ;
 wire \mac1.products_ff[140] ;
 wire \mac1.products_ff[141] ;
 wire \mac1.products_ff[142] ;
 wire \mac1.products_ff[143] ;
 wire \mac1.products_ff[144] ;
 wire \mac1.products_ff[145] ;
 wire \mac1.products_ff[146] ;
 wire \mac1.products_ff[147] ;
 wire \mac1.products_ff[148] ;
 wire \mac1.products_ff[149] ;
 wire \mac1.products_ff[14] ;
 wire \mac1.products_ff[150] ;
 wire \mac1.products_ff[151] ;
 wire \mac1.products_ff[15] ;
 wire \mac1.products_ff[1] ;
 wire \mac1.products_ff[2] ;
 wire \mac1.products_ff[3] ;
 wire \mac1.products_ff[4] ;
 wire \mac1.products_ff[5] ;
 wire \mac1.products_ff[68] ;
 wire \mac1.products_ff[69] ;
 wire \mac1.products_ff[6] ;
 wire \mac1.products_ff[70] ;
 wire \mac1.products_ff[71] ;
 wire \mac1.products_ff[72] ;
 wire \mac1.products_ff[73] ;
 wire \mac1.products_ff[74] ;
 wire \mac1.products_ff[75] ;
 wire \mac1.products_ff[76] ;
 wire \mac1.products_ff[77] ;
 wire \mac1.products_ff[78] ;
 wire \mac1.products_ff[79] ;
 wire \mac1.products_ff[7] ;
 wire \mac1.products_ff[80] ;
 wire \mac1.products_ff[81] ;
 wire \mac1.products_ff[82] ;
 wire \mac1.products_ff[83] ;
 wire \mac1.products_ff[8] ;
 wire \mac1.products_ff[9] ;
 wire \mac1.sum_lvl1_ff[0] ;
 wire \mac1.sum_lvl1_ff[10] ;
 wire \mac1.sum_lvl1_ff[11] ;
 wire \mac1.sum_lvl1_ff[12] ;
 wire \mac1.sum_lvl1_ff[13] ;
 wire \mac1.sum_lvl1_ff[14] ;
 wire \mac1.sum_lvl1_ff[15] ;
 wire \mac1.sum_lvl1_ff[1] ;
 wire \mac1.sum_lvl1_ff[2] ;
 wire \mac1.sum_lvl1_ff[36] ;
 wire \mac1.sum_lvl1_ff[37] ;
 wire \mac1.sum_lvl1_ff[38] ;
 wire \mac1.sum_lvl1_ff[39] ;
 wire \mac1.sum_lvl1_ff[3] ;
 wire \mac1.sum_lvl1_ff[40] ;
 wire \mac1.sum_lvl1_ff[41] ;
 wire \mac1.sum_lvl1_ff[42] ;
 wire \mac1.sum_lvl1_ff[43] ;
 wire \mac1.sum_lvl1_ff[44] ;
 wire \mac1.sum_lvl1_ff[45] ;
 wire \mac1.sum_lvl1_ff[46] ;
 wire \mac1.sum_lvl1_ff[47] ;
 wire \mac1.sum_lvl1_ff[48] ;
 wire \mac1.sum_lvl1_ff[49] ;
 wire \mac1.sum_lvl1_ff[4] ;
 wire \mac1.sum_lvl1_ff[50] ;
 wire \mac1.sum_lvl1_ff[51] ;
 wire \mac1.sum_lvl1_ff[5] ;
 wire \mac1.sum_lvl1_ff[6] ;
 wire \mac1.sum_lvl1_ff[72] ;
 wire \mac1.sum_lvl1_ff[73] ;
 wire \mac1.sum_lvl1_ff[74] ;
 wire \mac1.sum_lvl1_ff[75] ;
 wire \mac1.sum_lvl1_ff[76] ;
 wire \mac1.sum_lvl1_ff[77] ;
 wire \mac1.sum_lvl1_ff[78] ;
 wire \mac1.sum_lvl1_ff[79] ;
 wire \mac1.sum_lvl1_ff[7] ;
 wire \mac1.sum_lvl1_ff[80] ;
 wire \mac1.sum_lvl1_ff[81] ;
 wire \mac1.sum_lvl1_ff[82] ;
 wire \mac1.sum_lvl1_ff[83] ;
 wire \mac1.sum_lvl1_ff[84] ;
 wire \mac1.sum_lvl1_ff[85] ;
 wire \mac1.sum_lvl1_ff[86] ;
 wire \mac1.sum_lvl1_ff[87] ;
 wire \mac1.sum_lvl1_ff[8] ;
 wire \mac1.sum_lvl1_ff[9] ;
 wire \mac1.sum_lvl2_ff[0] ;
 wire \mac1.sum_lvl2_ff[10] ;
 wire \mac1.sum_lvl2_ff[11] ;
 wire \mac1.sum_lvl2_ff[12] ;
 wire \mac1.sum_lvl2_ff[13] ;
 wire \mac1.sum_lvl2_ff[14] ;
 wire \mac1.sum_lvl2_ff[15] ;
 wire \mac1.sum_lvl2_ff[19] ;
 wire \mac1.sum_lvl2_ff[1] ;
 wire \mac1.sum_lvl2_ff[20] ;
 wire \mac1.sum_lvl2_ff[21] ;
 wire \mac1.sum_lvl2_ff[22] ;
 wire \mac1.sum_lvl2_ff[23] ;
 wire \mac1.sum_lvl2_ff[24] ;
 wire \mac1.sum_lvl2_ff[25] ;
 wire \mac1.sum_lvl2_ff[26] ;
 wire \mac1.sum_lvl2_ff[27] ;
 wire \mac1.sum_lvl2_ff[28] ;
 wire \mac1.sum_lvl2_ff[29] ;
 wire \mac1.sum_lvl2_ff[2] ;
 wire \mac1.sum_lvl2_ff[30] ;
 wire \mac1.sum_lvl2_ff[31] ;
 wire \mac1.sum_lvl2_ff[32] ;
 wire \mac1.sum_lvl2_ff[33] ;
 wire \mac1.sum_lvl2_ff[34] ;
 wire \mac1.sum_lvl2_ff[38] ;
 wire \mac1.sum_lvl2_ff[39] ;
 wire \mac1.sum_lvl2_ff[3] ;
 wire \mac1.sum_lvl2_ff[40] ;
 wire \mac1.sum_lvl2_ff[41] ;
 wire \mac1.sum_lvl2_ff[42] ;
 wire \mac1.sum_lvl2_ff[43] ;
 wire \mac1.sum_lvl2_ff[44] ;
 wire \mac1.sum_lvl2_ff[45] ;
 wire \mac1.sum_lvl2_ff[46] ;
 wire \mac1.sum_lvl2_ff[47] ;
 wire \mac1.sum_lvl2_ff[48] ;
 wire \mac1.sum_lvl2_ff[49] ;
 wire \mac1.sum_lvl2_ff[4] ;
 wire \mac1.sum_lvl2_ff[50] ;
 wire \mac1.sum_lvl2_ff[51] ;
 wire \mac1.sum_lvl2_ff[52] ;
 wire \mac1.sum_lvl2_ff[53] ;
 wire \mac1.sum_lvl2_ff[5] ;
 wire \mac1.sum_lvl2_ff[6] ;
 wire \mac1.sum_lvl2_ff[7] ;
 wire \mac1.sum_lvl2_ff[8] ;
 wire \mac1.sum_lvl2_ff[9] ;
 wire \mac1.sum_lvl3_ff[0] ;
 wire \mac1.sum_lvl3_ff[10] ;
 wire \mac1.sum_lvl3_ff[11] ;
 wire \mac1.sum_lvl3_ff[12] ;
 wire \mac1.sum_lvl3_ff[13] ;
 wire \mac1.sum_lvl3_ff[14] ;
 wire \mac1.sum_lvl3_ff[15] ;
 wire \mac1.sum_lvl3_ff[1] ;
 wire \mac1.sum_lvl3_ff[20] ;
 wire \mac1.sum_lvl3_ff[21] ;
 wire \mac1.sum_lvl3_ff[22] ;
 wire \mac1.sum_lvl3_ff[23] ;
 wire \mac1.sum_lvl3_ff[24] ;
 wire \mac1.sum_lvl3_ff[25] ;
 wire \mac1.sum_lvl3_ff[26] ;
 wire \mac1.sum_lvl3_ff[27] ;
 wire \mac1.sum_lvl3_ff[28] ;
 wire \mac1.sum_lvl3_ff[29] ;
 wire \mac1.sum_lvl3_ff[2] ;
 wire \mac1.sum_lvl3_ff[30] ;
 wire \mac1.sum_lvl3_ff[31] ;
 wire \mac1.sum_lvl3_ff[32] ;
 wire \mac1.sum_lvl3_ff[33] ;
 wire \mac1.sum_lvl3_ff[34] ;
 wire \mac1.sum_lvl3_ff[35] ;
 wire \mac1.sum_lvl3_ff[3] ;
 wire \mac1.sum_lvl3_ff[4] ;
 wire \mac1.sum_lvl3_ff[5] ;
 wire \mac1.sum_lvl3_ff[6] ;
 wire \mac1.sum_lvl3_ff[7] ;
 wire \mac1.sum_lvl3_ff[8] ;
 wire \mac1.sum_lvl3_ff[9] ;
 wire \mac1.total_sum[0] ;
 wire \mac1.total_sum[10] ;
 wire \mac1.total_sum[11] ;
 wire \mac1.total_sum[12] ;
 wire \mac1.total_sum[13] ;
 wire \mac1.total_sum[14] ;
 wire \mac1.total_sum[15] ;
 wire \mac1.total_sum[1] ;
 wire \mac1.total_sum[2] ;
 wire \mac1.total_sum[3] ;
 wire \mac1.total_sum[4] ;
 wire \mac1.total_sum[5] ;
 wire \mac1.total_sum[6] ;
 wire \mac1.total_sum[7] ;
 wire \mac1.total_sum[8] ;
 wire \mac1.total_sum[9] ;
 wire \mac2.products_ff[0] ;
 wire \mac2.products_ff[10] ;
 wire \mac2.products_ff[11] ;
 wire \mac2.products_ff[12] ;
 wire \mac2.products_ff[136] ;
 wire \mac2.products_ff[137] ;
 wire \mac2.products_ff[138] ;
 wire \mac2.products_ff[139] ;
 wire \mac2.products_ff[13] ;
 wire \mac2.products_ff[140] ;
 wire \mac2.products_ff[141] ;
 wire \mac2.products_ff[142] ;
 wire \mac2.products_ff[143] ;
 wire \mac2.products_ff[144] ;
 wire \mac2.products_ff[145] ;
 wire \mac2.products_ff[146] ;
 wire \mac2.products_ff[147] ;
 wire \mac2.products_ff[148] ;
 wire \mac2.products_ff[149] ;
 wire \mac2.products_ff[14] ;
 wire \mac2.products_ff[150] ;
 wire \mac2.products_ff[151] ;
 wire \mac2.products_ff[15] ;
 wire \mac2.products_ff[1] ;
 wire \mac2.products_ff[2] ;
 wire \mac2.products_ff[3] ;
 wire \mac2.products_ff[4] ;
 wire \mac2.products_ff[5] ;
 wire \mac2.products_ff[68] ;
 wire \mac2.products_ff[69] ;
 wire \mac2.products_ff[6] ;
 wire \mac2.products_ff[70] ;
 wire \mac2.products_ff[71] ;
 wire \mac2.products_ff[72] ;
 wire \mac2.products_ff[73] ;
 wire \mac2.products_ff[74] ;
 wire \mac2.products_ff[75] ;
 wire \mac2.products_ff[76] ;
 wire \mac2.products_ff[77] ;
 wire \mac2.products_ff[78] ;
 wire \mac2.products_ff[79] ;
 wire \mac2.products_ff[7] ;
 wire \mac2.products_ff[80] ;
 wire \mac2.products_ff[81] ;
 wire \mac2.products_ff[82] ;
 wire \mac2.products_ff[83] ;
 wire \mac2.products_ff[8] ;
 wire \mac2.products_ff[9] ;
 wire \mac2.sum_lvl1_ff[0] ;
 wire \mac2.sum_lvl1_ff[10] ;
 wire \mac2.sum_lvl1_ff[11] ;
 wire \mac2.sum_lvl1_ff[12] ;
 wire \mac2.sum_lvl1_ff[13] ;
 wire \mac2.sum_lvl1_ff[14] ;
 wire \mac2.sum_lvl1_ff[15] ;
 wire \mac2.sum_lvl1_ff[1] ;
 wire \mac2.sum_lvl1_ff[2] ;
 wire \mac2.sum_lvl1_ff[36] ;
 wire \mac2.sum_lvl1_ff[37] ;
 wire \mac2.sum_lvl1_ff[38] ;
 wire \mac2.sum_lvl1_ff[39] ;
 wire \mac2.sum_lvl1_ff[3] ;
 wire \mac2.sum_lvl1_ff[40] ;
 wire \mac2.sum_lvl1_ff[41] ;
 wire \mac2.sum_lvl1_ff[42] ;
 wire \mac2.sum_lvl1_ff[43] ;
 wire \mac2.sum_lvl1_ff[44] ;
 wire \mac2.sum_lvl1_ff[45] ;
 wire \mac2.sum_lvl1_ff[46] ;
 wire \mac2.sum_lvl1_ff[47] ;
 wire \mac2.sum_lvl1_ff[48] ;
 wire \mac2.sum_lvl1_ff[49] ;
 wire \mac2.sum_lvl1_ff[4] ;
 wire \mac2.sum_lvl1_ff[50] ;
 wire \mac2.sum_lvl1_ff[51] ;
 wire \mac2.sum_lvl1_ff[5] ;
 wire \mac2.sum_lvl1_ff[6] ;
 wire \mac2.sum_lvl1_ff[72] ;
 wire \mac2.sum_lvl1_ff[73] ;
 wire \mac2.sum_lvl1_ff[74] ;
 wire \mac2.sum_lvl1_ff[75] ;
 wire \mac2.sum_lvl1_ff[76] ;
 wire \mac2.sum_lvl1_ff[77] ;
 wire \mac2.sum_lvl1_ff[78] ;
 wire \mac2.sum_lvl1_ff[79] ;
 wire \mac2.sum_lvl1_ff[7] ;
 wire \mac2.sum_lvl1_ff[80] ;
 wire \mac2.sum_lvl1_ff[81] ;
 wire \mac2.sum_lvl1_ff[82] ;
 wire \mac2.sum_lvl1_ff[83] ;
 wire \mac2.sum_lvl1_ff[84] ;
 wire \mac2.sum_lvl1_ff[85] ;
 wire \mac2.sum_lvl1_ff[86] ;
 wire \mac2.sum_lvl1_ff[87] ;
 wire \mac2.sum_lvl1_ff[8] ;
 wire \mac2.sum_lvl1_ff[9] ;
 wire \mac2.sum_lvl2_ff[0] ;
 wire \mac2.sum_lvl2_ff[10] ;
 wire \mac2.sum_lvl2_ff[11] ;
 wire \mac2.sum_lvl2_ff[12] ;
 wire \mac2.sum_lvl2_ff[13] ;
 wire \mac2.sum_lvl2_ff[14] ;
 wire \mac2.sum_lvl2_ff[15] ;
 wire \mac2.sum_lvl2_ff[19] ;
 wire \mac2.sum_lvl2_ff[1] ;
 wire \mac2.sum_lvl2_ff[20] ;
 wire \mac2.sum_lvl2_ff[21] ;
 wire \mac2.sum_lvl2_ff[22] ;
 wire \mac2.sum_lvl2_ff[23] ;
 wire \mac2.sum_lvl2_ff[24] ;
 wire \mac2.sum_lvl2_ff[25] ;
 wire \mac2.sum_lvl2_ff[26] ;
 wire \mac2.sum_lvl2_ff[27] ;
 wire \mac2.sum_lvl2_ff[28] ;
 wire \mac2.sum_lvl2_ff[29] ;
 wire \mac2.sum_lvl2_ff[2] ;
 wire \mac2.sum_lvl2_ff[30] ;
 wire \mac2.sum_lvl2_ff[31] ;
 wire \mac2.sum_lvl2_ff[32] ;
 wire \mac2.sum_lvl2_ff[33] ;
 wire \mac2.sum_lvl2_ff[34] ;
 wire \mac2.sum_lvl2_ff[38] ;
 wire \mac2.sum_lvl2_ff[39] ;
 wire \mac2.sum_lvl2_ff[3] ;
 wire \mac2.sum_lvl2_ff[40] ;
 wire \mac2.sum_lvl2_ff[41] ;
 wire \mac2.sum_lvl2_ff[42] ;
 wire \mac2.sum_lvl2_ff[43] ;
 wire \mac2.sum_lvl2_ff[44] ;
 wire \mac2.sum_lvl2_ff[45] ;
 wire \mac2.sum_lvl2_ff[46] ;
 wire \mac2.sum_lvl2_ff[47] ;
 wire \mac2.sum_lvl2_ff[48] ;
 wire \mac2.sum_lvl2_ff[49] ;
 wire \mac2.sum_lvl2_ff[4] ;
 wire \mac2.sum_lvl2_ff[50] ;
 wire \mac2.sum_lvl2_ff[51] ;
 wire \mac2.sum_lvl2_ff[52] ;
 wire \mac2.sum_lvl2_ff[53] ;
 wire \mac2.sum_lvl2_ff[5] ;
 wire \mac2.sum_lvl2_ff[6] ;
 wire \mac2.sum_lvl2_ff[7] ;
 wire \mac2.sum_lvl2_ff[8] ;
 wire \mac2.sum_lvl2_ff[9] ;
 wire \mac2.sum_lvl3_ff[0] ;
 wire \mac2.sum_lvl3_ff[10] ;
 wire \mac2.sum_lvl3_ff[11] ;
 wire \mac2.sum_lvl3_ff[12] ;
 wire \mac2.sum_lvl3_ff[13] ;
 wire \mac2.sum_lvl3_ff[14] ;
 wire \mac2.sum_lvl3_ff[15] ;
 wire \mac2.sum_lvl3_ff[1] ;
 wire \mac2.sum_lvl3_ff[20] ;
 wire \mac2.sum_lvl3_ff[21] ;
 wire \mac2.sum_lvl3_ff[22] ;
 wire \mac2.sum_lvl3_ff[23] ;
 wire \mac2.sum_lvl3_ff[24] ;
 wire \mac2.sum_lvl3_ff[25] ;
 wire \mac2.sum_lvl3_ff[26] ;
 wire \mac2.sum_lvl3_ff[27] ;
 wire \mac2.sum_lvl3_ff[28] ;
 wire \mac2.sum_lvl3_ff[29] ;
 wire \mac2.sum_lvl3_ff[2] ;
 wire \mac2.sum_lvl3_ff[30] ;
 wire \mac2.sum_lvl3_ff[31] ;
 wire \mac2.sum_lvl3_ff[32] ;
 wire \mac2.sum_lvl3_ff[33] ;
 wire \mac2.sum_lvl3_ff[34] ;
 wire \mac2.sum_lvl3_ff[35] ;
 wire \mac2.sum_lvl3_ff[3] ;
 wire \mac2.sum_lvl3_ff[4] ;
 wire \mac2.sum_lvl3_ff[5] ;
 wire \mac2.sum_lvl3_ff[6] ;
 wire \mac2.sum_lvl3_ff[7] ;
 wire \mac2.sum_lvl3_ff[8] ;
 wire \mac2.sum_lvl3_ff[9] ;
 wire \mac2.total_sum[0] ;
 wire \mac2.total_sum[10] ;
 wire \mac2.total_sum[11] ;
 wire \mac2.total_sum[12] ;
 wire \mac2.total_sum[13] ;
 wire \mac2.total_sum[14] ;
 wire \mac2.total_sum[15] ;
 wire \mac2.total_sum[1] ;
 wire \mac2.total_sum[2] ;
 wire \mac2.total_sum[3] ;
 wire \mac2.total_sum[4] ;
 wire \mac2.total_sum[5] ;
 wire \mac2.total_sum[6] ;
 wire \mac2.total_sum[7] ;
 wire \mac2.total_sum[8] ;
 wire \mac2.total_sum[9] ;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire clknet_leaf_0_clk;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net33;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;

 sg13g2_inv_1 _2996_ (.VDD(VPWR),
    .Y(_2600_),
    .A(\DP_1.Q_range.out_data[3] ),
    .VSS(VGND));
 sg13g2_inv_1 _2997_ (.VDD(VPWR),
    .Y(_2601_),
    .A(\DP_1.I_range.out_data[5] ),
    .VSS(VGND));
 sg13g2_inv_1 _2998_ (.VDD(VPWR),
    .Y(_2602_),
    .A(\DP_1.Q_range.out_data[5] ),
    .VSS(VGND));
 sg13g2_inv_1 _2999_ (.VDD(VPWR),
    .Y(_2603_),
    .A(\DP_3.I_range.out_data[5] ),
    .VSS(VGND));
 sg13g2_inv_1 _3000_ (.VDD(VPWR),
    .Y(_2604_),
    .A(\DP_3.Q_range.out_data[5] ),
    .VSS(VGND));
 sg13g2_inv_1 _3001_ (.VDD(VPWR),
    .Y(\DP_1.I_range.data_plus_4[6] ),
    .A(net4),
    .VSS(VGND));
 sg13g2_inv_1 _3002_ (.VDD(VPWR),
    .Y(\DP_3.I_range.data_plus_4[6] ),
    .A(net16),
    .VSS(VGND));
 sg13g2_inv_1 _3003_ (.VDD(VPWR),
    .Y(\DP_3.Q_range.data_plus_4[6] ),
    .A(net12),
    .VSS(VGND));
 sg13g2_inv_1 _3004_ (.VDD(VPWR),
    .Y(\DP_1.Q_range.data_plus_4[6] ),
    .A(net8),
    .VSS(VGND));
 sg13g2_inv_1 _3005_ (.VDD(VPWR),
    .Y(_2605_),
    .A(net1006),
    .VSS(VGND));
 sg13g2_inv_1 _3006_ (.VDD(VPWR),
    .Y(_2606_),
    .A(net292),
    .VSS(VGND));
 sg13g2_inv_1 _3007_ (.VDD(VPWR),
    .Y(_2607_),
    .A(net1026),
    .VSS(VGND));
 sg13g2_and2_1 _3008_ (.A(net984),
    .B(net923),
    .X(_0064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _3009_ (.X(_2608_),
    .A(net981),
    .B(net917),
    .C(_0064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3010_ (.Y(_2609_),
    .B1(net917),
    .B2(net984),
    .A2(net981),
    .A1(net923),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3011_ (.A(_2608_),
    .B(_2609_),
    .Y(_0065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3012_ (.Y(_2610_),
    .A(net984),
    .B(net915),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3013_ (.A(net923),
    .B(net981),
    .C(net917),
    .D(net978),
    .X(_2611_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3014_ (.Y(_2612_),
    .B1(net978),
    .B2(net923),
    .A2(net917),
    .A1(net981),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3015_ (.A(_2610_),
    .B(_2611_),
    .C(_2612_),
    .Y(_2613_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3016_ (.B1(_2610_),
    .VDD(VPWR),
    .Y(_2614_),
    .VSS(VGND),
    .A1(_2611_),
    .A2(_2612_));
 sg13g2_nor2b_1 _3017_ (.A(_2613_),
    .B_N(_2614_),
    .Y(_2615_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3018_ (.Y(_2616_),
    .A(_2608_),
    .B(_2615_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3019_ (.B(_2615_),
    .A(_2608_),
    .X(_0066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3020_ (.Y(_2617_),
    .A(net984),
    .B(net913),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3021_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2618_),
    .B(_2613_),
    .A(_2611_));
 sg13g2_nand2_1 _3022_ (.Y(_2619_),
    .A(net983),
    .B(net916),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3023_ (.A(net923),
    .B(net920),
    .C(net978),
    .D(net976),
    .X(_2620_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3024_ (.B(net920),
    .C(net978),
    .A(net924),
    .Y(_2621_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net976));
 sg13g2_a22oi_1 _3025_ (.Y(_2622_),
    .B1(net976),
    .B2(net924),
    .A2(net980),
    .A1(net920),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3026_ (.A(_2619_),
    .B(_2620_),
    .C(_2622_),
    .Y(_2623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3027_ (.B1(_2619_),
    .VDD(VPWR),
    .Y(_2624_),
    .VSS(VGND),
    .A1(_2620_),
    .A2(_2622_));
 sg13g2_nor2b_2 _3028_ (.A(_2623_),
    .B_N(_2624_),
    .Y(_2625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3029_ (.Y(_2626_),
    .A(_2618_),
    .B(_2625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3030_ (.Y(_2627_),
    .A(_2618_),
    .B(_2625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3031_ (.B(_2627_),
    .A(_2617_),
    .X(_2628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3032_ (.Y(_2629_),
    .B(_2628_),
    .A_N(_2616_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3033_ (.Y(_0067_),
    .A(_2616_),
    .B(_2628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3034_ (.Y(_2630_),
    .B1(net911),
    .B2(net984),
    .A2(net913),
    .A1(net981),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3035_ (.Y(_2631_),
    .A(net982),
    .B(net911),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3036_ (.A(net984),
    .B(net981),
    .C(net913),
    .D(net911),
    .X(_2632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3037_ (.A(_2630_),
    .B(_2632_),
    .Y(_2633_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3038_ (.VDD(VPWR),
    .Y(_2634_),
    .A(_2633_),
    .VSS(VGND));
 sg13g2_o21ai_1 _3039_ (.B1(_2621_),
    .VDD(VPWR),
    .Y(_2635_),
    .VSS(VGND),
    .A1(_2619_),
    .A2(_2622_));
 sg13g2_nand2_1 _3040_ (.Y(_2636_),
    .A(net978),
    .B(net915),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3041_ (.A(net922),
    .B(net917),
    .C(net975),
    .D(net972),
    .X(_2637_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3042_ (.B(net919),
    .C(net975),
    .A(net922),
    .Y(_2638_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net972));
 sg13g2_a22oi_1 _3043_ (.Y(_2639_),
    .B1(net972),
    .B2(net922),
    .A2(net976),
    .A1(net919),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3044_ (.A(_2636_),
    .B(_2637_),
    .C(_2639_),
    .X(_2640_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3045_ (.B1(_2636_),
    .VDD(VPWR),
    .Y(_2641_),
    .VSS(VGND),
    .A1(_2637_),
    .A2(_2639_));
 sg13g2_nand3_1 _3046_ (.B(_2640_),
    .C(_2641_),
    .A(_2635_),
    .Y(_2642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3047_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2640_),
    .A2(_2641_),
    .Y(_2643_),
    .B1(_2635_));
 sg13g2_a21o_1 _3048_ (.A2(_2641_),
    .A1(_2640_),
    .B1(_2635_),
    .X(_2644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3049_ (.Y(_2645_),
    .A(_2642_),
    .B(_2644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3050_ (.Y(_2646_),
    .A(_2634_),
    .B(_2645_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3051_ (.B1(_2626_),
    .VDD(VPWR),
    .Y(_2647_),
    .VSS(VGND),
    .A1(_2617_),
    .A2(_2627_));
 sg13g2_nor2b_2 _3052_ (.A(_2646_),
    .B_N(_2647_),
    .Y(_2648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3053_ (.B(_2647_),
    .A(_2646_),
    .X(_2649_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3054_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2650_),
    .B(_2649_),
    .A(_2629_));
 sg13g2_xor2_1 _3055_ (.B(_2649_),
    .A(_2629_),
    .X(_0068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3056_ (.B1(_2642_),
    .VDD(VPWR),
    .Y(_2651_),
    .VSS(VGND),
    .A1(_2634_),
    .A2(_2643_));
 sg13g2_nand2_1 _3057_ (.Y(_2652_),
    .A(net984),
    .B(net909),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3058_ (.Y(_2653_),
    .A(net979),
    .B(net911),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3059_ (.Y(_2654_),
    .A(net978),
    .B(net913),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3060_ (.B(_2654_),
    .A(_2631_),
    .X(_2655_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3061_ (.Y(_2656_),
    .B(_2655_),
    .A_N(_2652_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3062_ (.B(_2655_),
    .A(_2652_),
    .X(_2657_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3063_ (.B1(_2638_),
    .VDD(VPWR),
    .Y(_2658_),
    .VSS(VGND),
    .A1(_2636_),
    .A2(_2639_));
 sg13g2_nand2_1 _3064_ (.Y(_2659_),
    .A(net915),
    .B(net975),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3065_ (.A(net921),
    .B(net917),
    .C(net972),
    .D(net969),
    .X(_2660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3066_ (.B(net917),
    .C(net972),
    .A(net921),
    .Y(_2661_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net969));
 sg13g2_a22oi_1 _3067_ (.Y(_2662_),
    .B1(net969),
    .B2(net921),
    .A2(net972),
    .A1(net917),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3068_ (.A(_2659_),
    .B(_2660_),
    .C(_2662_),
    .X(_2663_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3069_ (.B1(_2659_),
    .VDD(VPWR),
    .Y(_2664_),
    .VSS(VGND),
    .A1(_2660_),
    .A2(_2662_));
 sg13g2_and3_1 _3070_ (.X(_2665_),
    .A(_2658_),
    .B(_2663_),
    .C(_2664_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3071_ (.B(_2663_),
    .C(_2664_),
    .A(_2658_),
    .Y(_2666_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3072_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2663_),
    .A2(_2664_),
    .Y(_2667_),
    .B1(_2658_));
 sg13g2_or3_1 _3073_ (.A(_2657_),
    .B(_2665_),
    .C(_2667_),
    .X(_2668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3074_ (.B1(_2657_),
    .VDD(VPWR),
    .Y(_2669_),
    .VSS(VGND),
    .A1(_2665_),
    .A2(_2667_));
 sg13g2_nand3_1 _3075_ (.B(_2668_),
    .C(_2669_),
    .A(_2651_),
    .Y(_2670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3076_ (.A2(_2669_),
    .A1(_2668_),
    .B1(_2651_),
    .X(_2671_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3077_ (.B(_2670_),
    .C(_2671_),
    .A(_2632_),
    .Y(_2672_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3078_ (.A2(_2671_),
    .A1(_2670_),
    .B1(_2632_),
    .X(_2673_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3079_ (.A(_2672_),
    .B(_2673_),
    .X(_2674_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3080_ (.B(_2672_),
    .C(_2673_),
    .A(_2648_),
    .Y(_2675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3081_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2672_),
    .A2(_2673_),
    .Y(_2676_),
    .B1(_2648_));
 sg13g2_xor2_1 _3082_ (.B(_2674_),
    .A(_2648_),
    .X(_2677_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3083_ (.Y(_0094_),
    .A(_2650_),
    .B(_2677_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3084_ (.Y(_2678_),
    .A(_2670_),
    .B(_2672_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3085_ (.B1(_2656_),
    .VDD(VPWR),
    .Y(_2679_),
    .VSS(VGND),
    .A1(_2631_),
    .A2(_2654_));
 sg13g2_nand2_1 _3086_ (.Y(_2680_),
    .A(net985),
    .B(net907),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3087_ (.Y(_2681_),
    .B(_2679_),
    .A_N(_2680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3088_ (.B(_2680_),
    .A(_2679_),
    .X(_2682_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3089_ (.B1(_2666_),
    .VDD(VPWR),
    .Y(_2683_),
    .VSS(VGND),
    .A1(_2657_),
    .A2(_2667_));
 sg13g2_nand2_1 _3090_ (.Y(_2684_),
    .A(net982),
    .B(net909),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3091_ (.Y(_2685_),
    .A(net975),
    .B(net911),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3092_ (.Y(_2686_),
    .A(net975),
    .B(net913),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3093_ (.B(_2686_),
    .A(_2653_),
    .X(_2687_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3094_ (.Y(_2688_),
    .B(_2687_),
    .A_N(_2684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3095_ (.Y(_2689_),
    .A(_2684_),
    .B(_2687_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3096_ (.B1(_2661_),
    .VDD(VPWR),
    .Y(_2690_),
    .VSS(VGND),
    .A1(_2659_),
    .A2(_2662_));
 sg13g2_nand2_1 _3097_ (.Y(_2691_),
    .A(net915),
    .B(net972),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3098_ (.A(net921),
    .B(net918),
    .C(net969),
    .D(net967),
    .X(_2692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3099_ (.B(net918),
    .C(net969),
    .A(net921),
    .Y(_2693_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net967));
 sg13g2_a22oi_1 _3100_ (.Y(_2694_),
    .B1(net967),
    .B2(net921),
    .A2(net969),
    .A1(net918),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3101_ (.A(_2691_),
    .B(_2692_),
    .C(_2694_),
    .X(_2695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3102_ (.B1(_2691_),
    .VDD(VPWR),
    .Y(_2696_),
    .VSS(VGND),
    .A1(_2692_),
    .A2(_2694_));
 sg13g2_and3_1 _3103_ (.X(_2697_),
    .A(_2690_),
    .B(_2695_),
    .C(_2696_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3104_ (.B(_2695_),
    .C(_2696_),
    .A(_2690_),
    .Y(_2698_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3105_ (.A2(_2696_),
    .A1(_2695_),
    .B1(_2690_),
    .X(_2699_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3106_ (.B(_2698_),
    .C(_2699_),
    .A(_2689_),
    .Y(_2700_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3107_ (.A2(_2699_),
    .A1(_2698_),
    .B1(_2689_),
    .X(_2701_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3108_ (.B(_2700_),
    .C(_2701_),
    .A(_2683_),
    .Y(_2702_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3109_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2700_),
    .A2(_2701_),
    .Y(_2703_),
    .B1(_2683_));
 sg13g2_a21o_1 _3110_ (.A2(_2701_),
    .A1(_2700_),
    .B1(_2683_),
    .X(_2704_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3111_ (.Y(_2705_),
    .A(_2702_),
    .B(_2704_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3112_ (.Y(_2706_),
    .A(_2682_),
    .B(_2705_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3113_ (.A(_2706_),
    .B_N(_2678_),
    .Y(_2707_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3114_ (.Y(_2708_),
    .A(_2678_),
    .B(_2706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3115_ (.B1(_2675_),
    .VDD(VPWR),
    .Y(_2709_),
    .VSS(VGND),
    .A1(_2650_),
    .A2(_2676_));
 sg13g2_xor2_1 _3116_ (.B(_2709_),
    .A(_2708_),
    .X(_0101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3117_ (.B1(_2702_),
    .VDD(VPWR),
    .Y(_2710_),
    .VSS(VGND),
    .A1(_2682_),
    .A2(_2703_));
 sg13g2_o21ai_1 _3118_ (.B1(_2688_),
    .VDD(VPWR),
    .Y(_2711_),
    .VSS(VGND),
    .A1(_2653_),
    .A2(_2686_));
 sg13g2_a22oi_1 _3119_ (.Y(_2712_),
    .B1(net905),
    .B2(net984),
    .A2(net907),
    .A1(net982),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3120_ (.B(net982),
    .C(net907),
    .A(net985),
    .Y(_2713_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net905));
 sg13g2_nor2b_1 _3121_ (.A(_2712_),
    .B_N(_2713_),
    .Y(_2714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3122_ (.Y(_2715_),
    .A(_2711_),
    .B(_2714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3123_ (.Y(_2716_),
    .A(_2711_),
    .B(_2714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3124_ (.A2(_2699_),
    .A1(_2689_),
    .B1(_2697_),
    .X(_2717_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3125_ (.Y(_2718_),
    .A(net979),
    .B(net909),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3126_ (.Y(_2719_),
    .A(net973),
    .B(net911),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3127_ (.Y(_2720_),
    .A(net913),
    .B(net973),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3128_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2721_),
    .B(_2719_),
    .A(_2686_));
 sg13g2_and2_1 _3129_ (.A(_2685_),
    .B(_2720_),
    .X(_2722_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3130_ (.Y(_2723_),
    .A(_2685_),
    .B(_2720_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3131_ (.Y(_2724_),
    .A(_2718_),
    .B(_2723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3132_ (.B1(_2693_),
    .VDD(VPWR),
    .Y(_2725_),
    .VSS(VGND),
    .A1(_2691_),
    .A2(_2694_));
 sg13g2_nand2_1 _3133_ (.Y(_2726_),
    .A(net915),
    .B(net969),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3134_ (.A(net921),
    .B(net918),
    .C(net967),
    .D(net964),
    .X(_2727_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3135_ (.B(net918),
    .C(net967),
    .A(net922),
    .Y(_2728_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net964));
 sg13g2_a22oi_1 _3136_ (.Y(_2729_),
    .B1(net964),
    .B2(net921),
    .A2(net967),
    .A1(net918),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3137_ (.A(_2726_),
    .B(_2727_),
    .C(_2729_),
    .X(_2730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3138_ (.B1(_2726_),
    .VDD(VPWR),
    .Y(_2731_),
    .VSS(VGND),
    .A1(_2727_),
    .A2(_2729_));
 sg13g2_and3_1 _3139_ (.X(_2732_),
    .A(_2725_),
    .B(_2730_),
    .C(_2731_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3140_ (.B(_2730_),
    .C(_2731_),
    .A(_2725_),
    .Y(_2733_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3141_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2730_),
    .A2(_2731_),
    .Y(_2734_),
    .B1(_2725_));
 sg13g2_or3_1 _3142_ (.A(_2724_),
    .B(_2732_),
    .C(_2734_),
    .X(_2735_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3143_ (.B1(_2724_),
    .VDD(VPWR),
    .Y(_2736_),
    .VSS(VGND),
    .A1(_2732_),
    .A2(_2734_));
 sg13g2_and3_1 _3144_ (.X(_2737_),
    .A(_2717_),
    .B(_2735_),
    .C(_2736_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3145_ (.B(_2735_),
    .C(_2736_),
    .A(_2717_),
    .Y(_2738_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3146_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2735_),
    .A2(_2736_),
    .Y(_2739_),
    .B1(_2717_));
 sg13g2_or3_1 _3147_ (.A(_2716_),
    .B(_2737_),
    .C(_2739_),
    .X(_2740_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3148_ (.B1(_2716_),
    .VDD(VPWR),
    .Y(_2741_),
    .VSS(VGND),
    .A1(_2737_),
    .A2(_2739_));
 sg13g2_nand3_1 _3149_ (.B(_2740_),
    .C(_2741_),
    .A(_2710_),
    .Y(_2742_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3150_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2740_),
    .A2(_2741_),
    .Y(_2743_),
    .B1(_2710_));
 sg13g2_a21o_1 _3151_ (.A2(_2741_),
    .A1(_2740_),
    .B1(_2710_),
    .X(_2744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3152_ (.Y(_2745_),
    .A(_2742_),
    .B(_2744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3153_ (.B(_2745_),
    .A(_2681_),
    .X(_2746_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _3154_ (.A2(_2709_),
    .A1(_2708_),
    .B1(_2707_),
    .X(_2747_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3155_ (.Y(_2748_),
    .A(_2746_),
    .B(_2747_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3156_ (.B(_2747_),
    .A(_2746_),
    .X(_0102_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3157_ (.B1(_2738_),
    .VDD(VPWR),
    .Y(_2749_),
    .VSS(VGND),
    .A1(_2716_),
    .A2(_2739_));
 sg13g2_o21ai_1 _3158_ (.B1(_2721_),
    .VDD(VPWR),
    .Y(_2750_),
    .VSS(VGND),
    .A1(_2718_),
    .A2(_2722_));
 sg13g2_nand2_1 _3159_ (.Y(_2751_),
    .A(net985),
    .B(net1030),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3160_ (.Y(_2752_),
    .A(net978),
    .B(net905),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3161_ (.A(net981),
    .B(net979),
    .C(net907),
    .D(net905),
    .X(_2753_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3162_ (.Y(_2754_),
    .B1(net905),
    .B2(net982),
    .A2(net907),
    .A1(net979),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3163_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2755_),
    .B(_2754_),
    .A(_2753_));
 sg13g2_nor2_1 _3164_ (.A(_2751_),
    .B(_2755_),
    .Y(_2756_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3165_ (.B(_2755_),
    .A(_2751_),
    .X(_2757_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3166_ (.Y(_2758_),
    .A(_2750_),
    .B(_2757_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3167_ (.Y(_2759_),
    .A(_2750_),
    .B(_2757_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3168_ (.Y(_2760_),
    .A(_2713_),
    .B(_2759_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3169_ (.B1(_2733_),
    .VDD(VPWR),
    .Y(_2761_),
    .VSS(VGND),
    .A1(_2724_),
    .A2(_2734_));
 sg13g2_nand2_1 _3170_ (.Y(_2762_),
    .A(net975),
    .B(net909),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3171_ (.Y(_2763_),
    .A(net911),
    .B(net969),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3172_ (.Y(_2764_),
    .A(net913),
    .B(net970),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3173_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2765_),
    .B(_2763_),
    .A(_2720_));
 sg13g2_xnor2_1 _3174_ (.Y(_2766_),
    .A(_2719_),
    .B(_2764_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3175_ (.Y(_2767_),
    .A(_2762_),
    .B(_2766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3176_ (.B1(_2728_),
    .VDD(VPWR),
    .Y(_2768_),
    .VSS(VGND),
    .A1(_2726_),
    .A2(_2729_));
 sg13g2_nand2_1 _3177_ (.Y(_2769_),
    .A(net915),
    .B(net967),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3178_ (.A(net922),
    .B(net919),
    .C(net964),
    .D(net1033),
    .X(_2770_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3179_ (.B(net919),
    .C(net964),
    .A(net922),
    .Y(_2771_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net1033));
 sg13g2_a22oi_1 _3180_ (.Y(_2772_),
    .B1(net1033),
    .B2(net922),
    .A2(net964),
    .A1(net919),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3181_ (.A(_2769_),
    .B(_2770_),
    .C(_2772_),
    .X(_2773_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3182_ (.B1(_2769_),
    .VDD(VPWR),
    .Y(_2774_),
    .VSS(VGND),
    .A1(_2770_),
    .A2(_2772_));
 sg13g2_and3_1 _3183_ (.X(_2775_),
    .A(_2768_),
    .B(_2773_),
    .C(_2774_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3184_ (.B(_2773_),
    .C(_2774_),
    .A(_2768_),
    .Y(_2776_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3185_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2773_),
    .A2(_2774_),
    .Y(_2777_),
    .B1(_2768_));
 sg13g2_or3_1 _3186_ (.A(_2767_),
    .B(_2775_),
    .C(_2777_),
    .X(_2778_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3187_ (.B1(_2767_),
    .VDD(VPWR),
    .Y(_2779_),
    .VSS(VGND),
    .A1(_2775_),
    .A2(_2777_));
 sg13g2_and3_1 _3188_ (.X(_2780_),
    .A(_2761_),
    .B(_2778_),
    .C(_2779_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3189_ (.B(_2778_),
    .C(_2779_),
    .A(_2761_),
    .Y(_2781_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3190_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2778_),
    .A2(_2779_),
    .Y(_2782_),
    .B1(_2761_));
 sg13g2_or3_1 _3191_ (.A(_2760_),
    .B(_2780_),
    .C(_2782_),
    .X(_2783_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3192_ (.B1(_2760_),
    .VDD(VPWR),
    .Y(_2784_),
    .VSS(VGND),
    .A1(_2780_),
    .A2(_2782_));
 sg13g2_and3_1 _3193_ (.X(_2785_),
    .A(_2749_),
    .B(_2783_),
    .C(_2784_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3194_ (.B(_2783_),
    .C(_2784_),
    .A(_2749_),
    .Y(_2786_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3195_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2783_),
    .A2(_2784_),
    .Y(_2787_),
    .B1(_2749_));
 sg13g2_or3_1 _3196_ (.A(_2715_),
    .B(_2785_),
    .C(_2787_),
    .X(_2788_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3197_ (.B1(_2715_),
    .VDD(VPWR),
    .Y(_2789_),
    .VSS(VGND),
    .A1(_2785_),
    .A2(_2787_));
 sg13g2_o21ai_1 _3198_ (.B1(_2742_),
    .VDD(VPWR),
    .Y(_2790_),
    .VSS(VGND),
    .A1(_2681_),
    .A2(_2743_));
 sg13g2_nand3_1 _3199_ (.B(_2789_),
    .C(_2790_),
    .A(_2788_),
    .Y(_2791_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3200_ (.A2(_2789_),
    .A1(_2788_),
    .B1(_2790_),
    .X(_2792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3201_ (.Y(_2793_),
    .A(_2791_),
    .B(_2792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3202_ (.A(_2746_),
    .B(_2747_),
    .C(_2791_),
    .D(_2792_),
    .X(_2794_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3203_ (.B(_2793_),
    .A(_2748_),
    .X(_0103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3204_ (.B1(_2791_),
    .VDD(VPWR),
    .Y(_2795_),
    .VSS(VGND),
    .A1(_2748_),
    .A2(_2793_));
 sg13g2_o21ai_1 _3205_ (.B1(_2786_),
    .VDD(VPWR),
    .Y(_2796_),
    .VSS(VGND),
    .A1(_2715_),
    .A2(_2787_));
 sg13g2_o21ai_1 _3206_ (.B1(_2758_),
    .VDD(VPWR),
    .Y(_2797_),
    .VSS(VGND),
    .A1(_2713_),
    .A2(_2759_));
 sg13g2_o21ai_1 _3207_ (.B1(_2781_),
    .VDD(VPWR),
    .Y(_2798_),
    .VSS(VGND),
    .A1(_2760_),
    .A2(_2782_));
 sg13g2_nor2_1 _3208_ (.A(_2753_),
    .B(_2756_),
    .Y(_2799_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3209_ (.B1(_2765_),
    .VDD(VPWR),
    .Y(_2800_),
    .VSS(VGND),
    .A1(_2762_),
    .A2(_2766_));
 sg13g2_nand2_1 _3210_ (.Y(_2801_),
    .A(net981),
    .B(net1030),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3211_ (.Y(_2802_),
    .A(net976),
    .B(net905),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3212_ (.Y(_2803_),
    .A(net975),
    .B(net907),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3213_ (.B(_2803_),
    .A(_2752_),
    .X(_2804_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3214_ (.Y(_2805_),
    .B(_2804_),
    .A_N(_2801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3215_ (.Y(_2806_),
    .A(_2801_),
    .B(_2804_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3216_ (.Y(_2807_),
    .A(_2800_),
    .B(_2806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3217_ (.A(_2799_),
    .B(_2807_),
    .Y(_2808_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3218_ (.Y(_2809_),
    .A(_2799_),
    .B(_2807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3219_ (.B1(_2776_),
    .VDD(VPWR),
    .Y(_2810_),
    .VSS(VGND),
    .A1(_2767_),
    .A2(_2777_));
 sg13g2_nand2_1 _3220_ (.Y(_2811_),
    .A(net972),
    .B(net909),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3221_ (.Y(_2812_),
    .A(net913),
    .B(net967),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3222_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2813_),
    .B(_2812_),
    .A(_2763_));
 sg13g2_and2_1 _3223_ (.A(_2763_),
    .B(_2812_),
    .X(_2814_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3224_ (.Y(_2815_),
    .A(_2763_),
    .B(_2812_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3225_ (.Y(_2816_),
    .A(_2811_),
    .B(_2815_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3226_ (.B1(_2771_),
    .VDD(VPWR),
    .Y(_2817_),
    .VSS(VGND),
    .A1(_2769_),
    .A2(_2772_));
 sg13g2_nand2_1 _3227_ (.Y(_2818_),
    .A(net916),
    .B(net1033),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3228_ (.A(net918),
    .B(net915),
    .C(net964),
    .D(net1033),
    .X(_2819_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3229_ (.Y(_2820_),
    .B1(net1033),
    .B2(net918),
    .A2(net964),
    .A1(net915),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3230_ (.A(_2819_),
    .B(_2820_),
    .Y(_2821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3231_ (.Y(_2822_),
    .A(_2817_),
    .B(_2821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3232_ (.Y(_2823_),
    .A(_2817_),
    .B(_2821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3233_ (.B(_2823_),
    .A(_2816_),
    .X(_2824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3234_ (.Y(_2825_),
    .A(_2810_),
    .B(_2824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3235_ (.Y(_2826_),
    .A(_2810_),
    .B(_2824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3236_ (.B(_2826_),
    .A(_2809_),
    .X(_2827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3237_ (.Y(_2828_),
    .A(_2798_),
    .B(_2827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3238_ (.Y(_2829_),
    .A(_2798_),
    .B(_2827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3239_ (.Y(_2830_),
    .B(_2797_),
    .A_N(_2829_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3240_ (.Y(_2831_),
    .A(_2797_),
    .B(_2829_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3241_ (.A(_2796_),
    .B(_2831_),
    .Y(_2832_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3242_ (.Y(_2833_),
    .A(_2796_),
    .B(_2831_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3243_ (.A(_2832_),
    .B_N(_2833_),
    .Y(_2834_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3244_ (.B(_2834_),
    .A(_2795_),
    .X(_0104_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3245_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2800_),
    .A2(_2806_),
    .Y(_2835_),
    .B1(_2808_));
 sg13g2_o21ai_1 _3246_ (.B1(_2825_),
    .VDD(VPWR),
    .Y(_2836_),
    .VSS(VGND),
    .A1(_2809_),
    .A2(_2826_));
 sg13g2_o21ai_1 _3247_ (.B1(_2805_),
    .VDD(VPWR),
    .Y(_2837_),
    .VSS(VGND),
    .A1(_2752_),
    .A2(_2803_));
 sg13g2_o21ai_1 _3248_ (.B1(_2813_),
    .VDD(VPWR),
    .Y(_2838_),
    .VSS(VGND),
    .A1(_2811_),
    .A2(_2814_));
 sg13g2_nand2_1 _3249_ (.Y(_2839_),
    .A(net978),
    .B(net1030),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3250_ (.Y(_2840_),
    .A(net973),
    .B(net905),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3251_ (.Y(_2841_),
    .A(net973),
    .B(net907),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3252_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2842_),
    .B(_2840_),
    .A(_2803_));
 sg13g2_xnor2_1 _3253_ (.Y(_2843_),
    .A(_2802_),
    .B(_2841_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3254_ (.B(_2843_),
    .A(_2839_),
    .X(_2844_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3255_ (.Y(_2845_),
    .A(_2838_),
    .B(_2844_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3256_ (.A(_2845_),
    .B_N(_2837_),
    .Y(_2846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3257_ (.B(_2845_),
    .A(_2837_),
    .X(_2847_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3258_ (.B1(_2822_),
    .VDD(VPWR),
    .Y(_2848_),
    .VSS(VGND),
    .A1(_2816_),
    .A2(_2823_));
 sg13g2_a21oi_1 _3259_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net920),
    .A2(net965),
    .Y(_2849_),
    .B1(_2818_));
 sg13g2_nand2_1 _3260_ (.Y(_2850_),
    .A(net970),
    .B(net909),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3261_ (.Y(_2851_),
    .A(net912),
    .B(net965),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3262_ (.A(net914),
    .B(net911),
    .C(net968),
    .D(net965),
    .X(_2852_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3263_ (.Y(_2853_),
    .B1(net965),
    .B2(net914),
    .A2(net968),
    .A1(net912),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3264_ (.A(_2850_),
    .B(_2852_),
    .C(_2853_),
    .Y(_2854_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3265_ (.B1(_2850_),
    .VDD(VPWR),
    .Y(_2855_),
    .VSS(VGND),
    .A1(_2852_),
    .A2(_2853_));
 sg13g2_nor2b_1 _3266_ (.A(_2854_),
    .B_N(_2855_),
    .Y(_2856_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3267_ (.Y(_2857_),
    .A(_2849_),
    .B(_2856_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3268_ (.Y(_2858_),
    .B(_2848_),
    .A_N(_2857_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3269_ (.B(_2857_),
    .A(_2848_),
    .X(_2859_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3270_ (.B(_2859_),
    .A(_2847_),
    .X(_2860_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3271_ (.Y(_2861_),
    .A(_2836_),
    .B(_2860_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3272_ (.B(_2860_),
    .A(_2836_),
    .X(_2862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3273_ (.Y(_2863_),
    .B(_2862_),
    .A_N(_2835_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3274_ (.B(_2862_),
    .A(_2835_),
    .X(_2864_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3275_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2828_),
    .A2(_2830_),
    .Y(_2865_),
    .B1(_2864_));
 sg13g2_nand3_1 _3276_ (.B(_2830_),
    .C(_2864_),
    .A(_2828_),
    .Y(_2866_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3277_ (.Y(_2867_),
    .B(_2866_),
    .A_N(_2865_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3278_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2791_),
    .A2(_2833_),
    .Y(_2868_),
    .B1(_2832_));
 sg13g2_a21oi_2 _3279_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_2868_),
    .Y(_2869_),
    .A2(_2834_),
    .A1(_2794_));
 sg13g2_nor2_1 _3280_ (.A(_2867_),
    .B(_2869_),
    .Y(_2870_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3281_ (.B(_2869_),
    .A(_2867_),
    .X(_0095_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3282_ (.A2(_2844_),
    .A1(_2838_),
    .B1(_2846_),
    .X(_2871_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3283_ (.B1(_2858_),
    .VDD(VPWR),
    .Y(_2872_),
    .VSS(VGND),
    .A1(_2847_),
    .A2(_2859_));
 sg13g2_a21o_2 _3284_ (.A2(_2856_),
    .A1(_2849_),
    .B1(_2819_),
    .X(_2873_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3285_ (.Y(_2874_),
    .A(net909),
    .B(net968),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3286_ (.Y(_2875_),
    .A(net914),
    .B(net1034),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3287_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2876_),
    .B(_2875_),
    .A(_2851_));
 sg13g2_xnor2_1 _3288_ (.Y(_2877_),
    .A(_2851_),
    .B(_2875_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3289_ (.B(_2877_),
    .A(_2874_),
    .X(_2878_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3290_ (.A(_2873_),
    .B(_2878_),
    .X(_2879_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3291_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2880_),
    .B(_2878_),
    .A(_2873_));
 sg13g2_xnor2_1 _3292_ (.Y(_2881_),
    .A(_2873_),
    .B(_2878_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3293_ (.B1(_2842_),
    .VDD(VPWR),
    .Y(_2882_),
    .VSS(VGND),
    .A1(_2839_),
    .A2(_2843_));
 sg13g2_or2_1 _3294_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2883_),
    .B(_2854_),
    .A(_2852_));
 sg13g2_nand2_1 _3295_ (.Y(_2884_),
    .A(net975),
    .B(net1030),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3296_ (.Y(_2885_),
    .A(net971),
    .B(net905),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3297_ (.Y(_2886_),
    .A(net970),
    .B(net907),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3298_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2887_),
    .B(_2885_),
    .A(_2841_));
 sg13g2_xnor2_1 _3299_ (.Y(_2888_),
    .A(_2840_),
    .B(_2886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3300_ (.B(_2888_),
    .A(_2884_),
    .X(_2889_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3301_ (.Y(_2890_),
    .A(_2883_),
    .B(_2889_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3302_ (.A(_2890_),
    .B_N(_2882_),
    .Y(_2891_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3303_ (.Y(_2892_),
    .A(_2882_),
    .B(_2890_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3304_ (.Y(_2893_),
    .A(_2881_),
    .B(_2892_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3305_ (.Y(_2894_),
    .A(_2872_),
    .B(_2893_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3306_ (.A(_2894_),
    .B_N(_2871_),
    .Y(_2895_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3307_ (.B(_2894_),
    .A(_2871_),
    .X(_2896_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3308_ (.B(_2863_),
    .C(_2896_),
    .A(_2861_),
    .Y(_2897_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3309_ (.VDD(VPWR),
    .Y(_2898_),
    .A(_2897_),
    .VSS(VGND));
 sg13g2_a21oi_1 _3310_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2861_),
    .A2(_2863_),
    .Y(_2899_),
    .B1(_2896_));
 sg13g2_nor2_1 _3311_ (.A(_2898_),
    .B(_2899_),
    .Y(_2900_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3312_ (.A(_2865_),
    .B(_2870_),
    .Y(_2901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3313_ (.Y(_0096_),
    .A(_2900_),
    .B(_2901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3314_ (.A2(_2889_),
    .A1(_2883_),
    .B1(_2891_),
    .X(_2902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3315_ (.Y(_2903_),
    .B1(net1033),
    .B2(net912),
    .A2(net966),
    .A1(net910),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3316_ (.Y(_2904_),
    .A(net909),
    .B(net1034),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3317_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2905_),
    .B(_2904_),
    .A(_2851_));
 sg13g2_nand2b_1 _3318_ (.Y(_2906_),
    .B(_2905_),
    .A_N(_2903_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3319_ (.B1(_2887_),
    .VDD(VPWR),
    .Y(_2907_),
    .VSS(VGND),
    .A1(_2884_),
    .A2(_2888_));
 sg13g2_o21ai_1 _3320_ (.B1(_2876_),
    .VDD(VPWR),
    .Y(_2908_),
    .VSS(VGND),
    .A1(_2874_),
    .A2(_2877_));
 sg13g2_nand2_1 _3321_ (.Y(_2909_),
    .A(net974),
    .B(net1030),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3322_ (.Y(_2910_),
    .A(net968),
    .B(net906),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3323_ (.Y(_2911_),
    .A(net968),
    .B(net908),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3324_ (.B(_2911_),
    .A(_2885_),
    .X(_2912_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3325_ (.Y(_2913_),
    .B(_2912_),
    .A_N(_2909_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3326_ (.Y(_2914_),
    .A(_2909_),
    .B(_2912_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3327_ (.Y(_2915_),
    .A(_2908_),
    .B(_2914_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3328_ (.A(_2915_),
    .B_N(_2907_),
    .Y(_2916_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3329_ (.B(_2915_),
    .A(_2907_),
    .X(_2917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3330_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2918_),
    .B(_2917_),
    .A(_2906_));
 sg13g2_xor2_1 _3331_ (.B(_2917_),
    .A(_2906_),
    .X(_2919_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3332_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2880_),
    .A2(_2892_),
    .Y(_2920_),
    .B1(_2879_));
 sg13g2_nor2b_1 _3333_ (.A(_2920_),
    .B_N(_2919_),
    .Y(_2921_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3334_ (.B(_2920_),
    .A(_2919_),
    .X(_2922_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3335_ (.A(_2922_),
    .B_N(_2902_),
    .Y(_2923_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3336_ (.B(_2922_),
    .A(_2902_),
    .X(_2924_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3337_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2872_),
    .A2(_2893_),
    .Y(_2925_),
    .B1(_2895_));
 sg13g2_nor2_1 _3338_ (.A(_2924_),
    .B(_2925_),
    .Y(_2926_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3339_ (.B(_2925_),
    .A(_2924_),
    .X(_2927_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3340_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2865_),
    .A2(_2897_),
    .Y(_2928_),
    .B1(_2899_));
 sg13g2_a21oi_1 _3341_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2866_),
    .A2(_2897_),
    .Y(_2929_),
    .B1(_2899_));
 sg13g2_a21oi_1 _3342_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2869_),
    .A2(_2928_),
    .Y(_2930_),
    .B1(_2929_));
 sg13g2_xor2_1 _3343_ (.B(_2930_),
    .A(_2927_),
    .X(_0097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3344_ (.A2(_2914_),
    .A1(_2908_),
    .B1(_2916_),
    .X(_2931_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3345_ (.B1(_2913_),
    .VDD(VPWR),
    .Y(_2932_),
    .VSS(VGND),
    .A1(_2885_),
    .A2(_2911_));
 sg13g2_nand2_1 _3346_ (.Y(_2933_),
    .A(net971),
    .B(net1030),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3347_ (.Y(_2934_),
    .A(net965),
    .B(net906),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3348_ (.Y(_2935_),
    .A(net908),
    .B(net965),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3349_ (.B(_2935_),
    .A(_2910_),
    .X(_2936_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3350_ (.Y(_2937_),
    .B(_2936_),
    .A_N(_2933_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3351_ (.Y(_2938_),
    .A(_2933_),
    .B(_2936_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3352_ (.A(_2905_),
    .B_N(_2938_),
    .Y(_2939_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3353_ (.Y(_2940_),
    .A(_2905_),
    .B(_2938_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3354_ (.Y(_2941_),
    .A(_2932_),
    .B(_2940_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3355_ (.A(_2904_),
    .B(_2941_),
    .Y(_2942_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3356_ (.Y(_2943_),
    .A(_2904_),
    .B(_2941_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3357_ (.A(_2918_),
    .B(_2943_),
    .Y(_2944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3358_ (.B(_2943_),
    .A(_2918_),
    .X(_2945_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3359_ (.B(_2945_),
    .A(_2931_),
    .X(_2946_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3360_ (.B1(_2946_),
    .VDD(VPWR),
    .Y(_2947_),
    .VSS(VGND),
    .A1(_2921_),
    .A2(_2923_));
 sg13g2_or3_1 _3361_ (.A(_2921_),
    .B(_2923_),
    .C(_2946_),
    .X(_2948_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3362_ (.A(_2947_),
    .B(_2948_),
    .X(_2949_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3363_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2927_),
    .A2(_2930_),
    .Y(_2950_),
    .B1(_2926_));
 sg13g2_xnor2_1 _3364_ (.Y(_0098_),
    .A(_2949_),
    .B(_2950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3365_ (.Y(_2951_),
    .A(_2927_),
    .B(_2949_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3366_ (.VDD(VPWR),
    .Y(_2952_),
    .A(_2951_),
    .VSS(VGND));
 sg13g2_o21ai_1 _3367_ (.B1(_2947_),
    .VDD(VPWR),
    .Y(_2953_),
    .VSS(VGND),
    .A1(_2924_),
    .A2(_2925_));
 sg13g2_a22oi_1 _3368_ (.Y(_2954_),
    .B1(_2953_),
    .B2(_2948_),
    .A2(_2952_),
    .A1(_2930_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3369_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2931_),
    .A2(_2945_),
    .Y(_2955_),
    .B1(_2944_));
 sg13g2_a21o_1 _3370_ (.A2(_2940_),
    .A1(_2932_),
    .B1(_2939_),
    .X(_2956_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3371_ (.Y(_2957_),
    .A(net968),
    .B(net1030),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3372_ (.Y(_2958_),
    .A(net906),
    .B(net1034),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3373_ (.Y(_2959_),
    .A(net908),
    .B(net1034),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3374_ (.B(_2959_),
    .A(_2934_),
    .X(_2960_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3375_ (.Y(_2961_),
    .B(_2960_),
    .A_N(_2957_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3376_ (.Y(_2962_),
    .A(_2957_),
    .B(_2960_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3377_ (.B1(_2937_),
    .VDD(VPWR),
    .Y(_2963_),
    .VSS(VGND),
    .A1(_2910_),
    .A2(_2935_));
 sg13g2_nand2_1 _3378_ (.Y(_2964_),
    .A(_2962_),
    .B(_2963_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3379_ (.B(_2963_),
    .A(_2962_),
    .X(_2965_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3380_ (.Y(_2966_),
    .A(_2942_),
    .B(_2965_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3381_ (.A(_2966_),
    .B_N(_2956_),
    .Y(_2967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3382_ (.B(_2966_),
    .A(_2956_),
    .X(_2968_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3383_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2969_),
    .B(_2968_),
    .A(_2955_));
 sg13g2_xor2_1 _3384_ (.B(_2968_),
    .A(_2955_),
    .X(_2970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3385_ (.VDD(VPWR),
    .Y(_2971_),
    .A(_2970_),
    .VSS(VGND));
 sg13g2_xnor2_1 _3386_ (.Y(_0099_),
    .A(_2954_),
    .B(_2970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3387_ (.B1(_2969_),
    .VDD(VPWR),
    .Y(_2972_),
    .VSS(VGND),
    .A1(_2954_),
    .A2(_2971_));
 sg13g2_a21oi_1 _3388_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2942_),
    .A2(_2965_),
    .Y(_2973_),
    .B1(_2967_));
 sg13g2_o21ai_1 _3389_ (.B1(_2961_),
    .VDD(VPWR),
    .Y(_2974_),
    .VSS(VGND),
    .A1(_2934_),
    .A2(_2959_));
 sg13g2_nand2_1 _3390_ (.Y(_2975_),
    .A(net965),
    .B(net1030),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3391_ (.B(_2975_),
    .A(_2958_),
    .X(_2976_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3392_ (.Y(_2977_),
    .A(_2974_),
    .B(_2976_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3393_ (.Y(_2978_),
    .A(_2964_),
    .B(_2977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3394_ (.Y(_2979_),
    .A(_2973_),
    .B(_2978_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3395_ (.Y(_0100_),
    .A(_2972_),
    .B(_2979_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3396_ (.A(net1019),
    .B(net960),
    .X(_0069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _3397_ (.X(_2980_),
    .A(net1018),
    .B(net956),
    .C(_0069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3398_ (.Y(_2981_),
    .B1(net956),
    .B2(net1019),
    .A2(net1018),
    .A1(net960),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3399_ (.A(_2980_),
    .B(net442),
    .Y(_0070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3400_ (.Y(_2982_),
    .A(net1019),
    .B(net954),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3401_ (.A(net960),
    .B(net1018),
    .C(net956),
    .D(net1015),
    .X(_2983_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3402_ (.Y(_2984_),
    .B1(net1015),
    .B2(net960),
    .A2(net956),
    .A1(net1018),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3403_ (.A(_2982_),
    .B(_2983_),
    .C(_2984_),
    .Y(_2985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3404_ (.B1(_2982_),
    .VDD(VPWR),
    .Y(_2986_),
    .VSS(VGND),
    .A1(_2983_),
    .A2(_2984_));
 sg13g2_nor2b_1 _3405_ (.A(_2985_),
    .B_N(_2986_),
    .Y(_2987_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3406_ (.Y(_2988_),
    .A(_2980_),
    .B(_2987_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3407_ (.B(_2987_),
    .A(_2980_),
    .X(_0071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3408_ (.Y(_2989_),
    .A(net1019),
    .B(net952),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3409_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2990_),
    .B(_2985_),
    .A(_2983_));
 sg13g2_nand2_1 _3410_ (.Y(_2991_),
    .A(net1018),
    .B(net954),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3411_ (.A(\DP_2.matrix[0] ),
    .B(net956),
    .C(net1015),
    .D(net1013),
    .X(_2992_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3412_ (.B(net956),
    .C(net1015),
    .A(net960),
    .Y(_2993_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net1013));
 sg13g2_a22oi_1 _3413_ (.Y(_2994_),
    .B1(net1013),
    .B2(net960),
    .A2(net1015),
    .A1(net959),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3414_ (.A(_2991_),
    .B(_2992_),
    .C(_2994_),
    .Y(_2995_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3415_ (.B1(_2991_),
    .VDD(VPWR),
    .Y(_0268_),
    .VSS(VGND),
    .A1(_2992_),
    .A2(_2994_));
 sg13g2_nor2b_1 _3416_ (.A(_2995_),
    .B_N(_0268_),
    .Y(_0269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3417_ (.Y(_0270_),
    .A(_2990_),
    .B(_0269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3418_ (.Y(_0271_),
    .A(_2990_),
    .B(_0269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3419_ (.B(_0271_),
    .A(_2989_),
    .X(_0272_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3420_ (.Y(_0273_),
    .B(_0272_),
    .A_N(_2988_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3421_ (.Y(_0072_),
    .A(_2988_),
    .B(_0272_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3422_ (.Y(_0274_),
    .B1(net951),
    .B2(net1019),
    .A2(net952),
    .A1(net1017),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3423_ (.Y(_0275_),
    .A(net1017),
    .B(net950),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3424_ (.A(net1019),
    .B(net1017),
    .C(net952),
    .D(net951),
    .X(_0276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3425_ (.A(_0274_),
    .B(_0276_),
    .Y(_0277_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3426_ (.VDD(VPWR),
    .Y(_0278_),
    .A(_0277_),
    .VSS(VGND));
 sg13g2_o21ai_1 _3427_ (.B1(_2993_),
    .VDD(VPWR),
    .Y(_0279_),
    .VSS(VGND),
    .A1(_2991_),
    .A2(_2994_));
 sg13g2_nand2_1 _3428_ (.Y(_0280_),
    .A(net1015),
    .B(net954),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3429_ (.A(net963),
    .B(net959),
    .C(net1013),
    .D(net1011),
    .X(_0281_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3430_ (.B(net958),
    .C(net1013),
    .A(net963),
    .Y(_0282_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net1011));
 sg13g2_a22oi_1 _3431_ (.Y(_0283_),
    .B1(net1011),
    .B2(net963),
    .A2(net1013),
    .A1(net959),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3432_ (.A(_0280_),
    .B(_0281_),
    .C(_0283_),
    .X(_0284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3433_ (.B1(_0280_),
    .VDD(VPWR),
    .Y(_0285_),
    .VSS(VGND),
    .A1(_0281_),
    .A2(_0283_));
 sg13g2_nand3_1 _3434_ (.B(_0284_),
    .C(_0285_),
    .A(_0279_),
    .Y(_0286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3435_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0284_),
    .A2(_0285_),
    .Y(_0287_),
    .B1(_0279_));
 sg13g2_a21o_1 _3436_ (.A2(_0285_),
    .A1(_0284_),
    .B1(_0279_),
    .X(_0288_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3437_ (.Y(_0289_),
    .A(_0286_),
    .B(_0288_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3438_ (.Y(_0290_),
    .A(_0278_),
    .B(_0289_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3439_ (.B1(_0270_),
    .VDD(VPWR),
    .Y(_0291_),
    .VSS(VGND),
    .A1(_2989_),
    .A2(_0271_));
 sg13g2_nor2b_2 _3440_ (.A(_0290_),
    .B_N(_0291_),
    .Y(_0292_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3441_ (.B(_0291_),
    .A(_0290_),
    .X(_0293_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3442_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0294_),
    .B(_0293_),
    .A(_0273_));
 sg13g2_xor2_1 _3443_ (.B(_0293_),
    .A(_0273_),
    .X(_0073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3444_ (.B1(_0286_),
    .VDD(VPWR),
    .Y(_0295_),
    .VSS(VGND),
    .A1(_0278_),
    .A2(_0287_));
 sg13g2_nand2_1 _3445_ (.Y(_0296_),
    .A(net1020),
    .B(net949),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3446_ (.Y(_0297_),
    .A(net1016),
    .B(net950),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3447_ (.Y(_0298_),
    .A(net1016),
    .B(net952),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3448_ (.B(_0298_),
    .A(_0275_),
    .X(_0299_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3449_ (.Y(_0300_),
    .B(_0299_),
    .A_N(_0296_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3450_ (.B(_0299_),
    .A(_0296_),
    .X(_0301_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3451_ (.B1(_0282_),
    .VDD(VPWR),
    .Y(_0302_),
    .VSS(VGND),
    .A1(_0280_),
    .A2(_0283_));
 sg13g2_nand2_1 _3452_ (.Y(_0303_),
    .A(net954),
    .B(net1014),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3453_ (.A(net963),
    .B(net958),
    .C(net1011),
    .D(net1009),
    .X(_0304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3454_ (.B(net958),
    .C(net1011),
    .A(net962),
    .Y(_0305_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net1009));
 sg13g2_a22oi_1 _3455_ (.Y(_0306_),
    .B1(net1009),
    .B2(net962),
    .A2(net1011),
    .A1(net958),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3456_ (.A(_0303_),
    .B(_0304_),
    .C(_0306_),
    .X(_0307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3457_ (.B1(_0303_),
    .VDD(VPWR),
    .Y(_0308_),
    .VSS(VGND),
    .A1(_0304_),
    .A2(_0306_));
 sg13g2_and3_1 _3458_ (.X(_0309_),
    .A(_0302_),
    .B(_0307_),
    .C(_0308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3459_ (.B(_0307_),
    .C(_0308_),
    .A(_0302_),
    .Y(_0310_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3460_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0307_),
    .A2(_0308_),
    .Y(_0311_),
    .B1(_0302_));
 sg13g2_or3_1 _3461_ (.A(_0301_),
    .B(_0309_),
    .C(_0311_),
    .X(_0312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3462_ (.B1(_0301_),
    .VDD(VPWR),
    .Y(_0313_),
    .VSS(VGND),
    .A1(_0309_),
    .A2(_0311_));
 sg13g2_nand3_1 _3463_ (.B(_0312_),
    .C(_0313_),
    .A(_0295_),
    .Y(_0314_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3464_ (.A2(_0313_),
    .A1(_0312_),
    .B1(_0295_),
    .X(_0315_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3465_ (.B(_0314_),
    .C(_0315_),
    .A(_0276_),
    .Y(_0316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3466_ (.A2(_0315_),
    .A1(_0314_),
    .B1(_0276_),
    .X(_0317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3467_ (.A(_0316_),
    .B(_0317_),
    .X(_0318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3468_ (.B(_0316_),
    .C(_0317_),
    .A(_0292_),
    .Y(_0319_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3469_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0316_),
    .A2(_0317_),
    .Y(_0320_),
    .B1(_0292_));
 sg13g2_xor2_1 _3470_ (.B(_0318_),
    .A(_0292_),
    .X(_0321_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3471_ (.Y(_0105_),
    .A(_0294_),
    .B(_0321_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3472_ (.Y(_0322_),
    .A(_0314_),
    .B(_0316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3473_ (.B1(_0300_),
    .VDD(VPWR),
    .Y(_0323_),
    .VSS(VGND),
    .A1(_0275_),
    .A2(_0298_));
 sg13g2_nand2_1 _3474_ (.Y(_0324_),
    .A(net1020),
    .B(net946),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3475_ (.Y(_0325_),
    .B(_0323_),
    .A_N(_0324_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3476_ (.B(_0324_),
    .A(_0323_),
    .X(_0326_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3477_ (.B1(_0310_),
    .VDD(VPWR),
    .Y(_0327_),
    .VSS(VGND),
    .A1(_0301_),
    .A2(_0311_));
 sg13g2_nand2_1 _3478_ (.Y(_0328_),
    .A(net1017),
    .B(net949),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3479_ (.Y(_0329_),
    .A(net1014),
    .B(net950),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3480_ (.Y(_0330_),
    .A(net1014),
    .B(net953),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3481_ (.B(_0330_),
    .A(_0297_),
    .X(_0331_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3482_ (.Y(_0332_),
    .B(_0331_),
    .A_N(_0328_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3483_ (.Y(_0333_),
    .A(_0328_),
    .B(_0331_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3484_ (.B1(_0305_),
    .VDD(VPWR),
    .Y(_0334_),
    .VSS(VGND),
    .A1(_0303_),
    .A2(_0306_));
 sg13g2_nand2_1 _3485_ (.Y(_0335_),
    .A(net954),
    .B(net1012),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3486_ (.A(net961),
    .B(net958),
    .C(net1009),
    .D(net1007),
    .X(_0336_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3487_ (.B(net957),
    .C(net1009),
    .A(net961),
    .Y(_0337_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net1007));
 sg13g2_a22oi_1 _3488_ (.Y(_0338_),
    .B1(net1007),
    .B2(net961),
    .A2(net1009),
    .A1(net958),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3489_ (.A(_0335_),
    .B(_0336_),
    .C(_0338_),
    .X(_0339_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3490_ (.B1(_0335_),
    .VDD(VPWR),
    .Y(_0340_),
    .VSS(VGND),
    .A1(_0336_),
    .A2(_0338_));
 sg13g2_and3_1 _3491_ (.X(_0341_),
    .A(_0334_),
    .B(_0339_),
    .C(_0340_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3492_ (.B(_0339_),
    .C(_0340_),
    .A(_0334_),
    .Y(_0342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3493_ (.A2(_0340_),
    .A1(_0339_),
    .B1(_0334_),
    .X(_0343_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3494_ (.B(_0342_),
    .C(_0343_),
    .A(_0333_),
    .Y(_0344_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3495_ (.A2(_0343_),
    .A1(_0342_),
    .B1(_0333_),
    .X(_0345_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3496_ (.B(_0344_),
    .C(_0345_),
    .A(_0327_),
    .Y(_0346_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3497_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0344_),
    .A2(_0345_),
    .Y(_0347_),
    .B1(_0327_));
 sg13g2_a21o_1 _3498_ (.A2(_0345_),
    .A1(_0344_),
    .B1(_0327_),
    .X(_0348_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3499_ (.Y(_0349_),
    .A(_0346_),
    .B(_0348_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3500_ (.Y(_0350_),
    .A(_0326_),
    .B(_0349_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3501_ (.A(_0350_),
    .B_N(_0322_),
    .Y(_0351_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3502_ (.Y(_0352_),
    .A(_0322_),
    .B(_0350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3503_ (.B1(_0319_),
    .VDD(VPWR),
    .Y(_0353_),
    .VSS(VGND),
    .A1(_0294_),
    .A2(_0320_));
 sg13g2_xor2_1 _3504_ (.B(_0353_),
    .A(_0352_),
    .X(_0112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3505_ (.B1(_0346_),
    .VDD(VPWR),
    .Y(_0354_),
    .VSS(VGND),
    .A1(_0326_),
    .A2(_0347_));
 sg13g2_o21ai_1 _3506_ (.B1(_0332_),
    .VDD(VPWR),
    .Y(_0355_),
    .VSS(VGND),
    .A1(_0297_),
    .A2(_0330_));
 sg13g2_a22oi_1 _3507_ (.Y(_0356_),
    .B1(net944),
    .B2(net1020),
    .A2(net946),
    .A1(net1017),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3508_ (.B(net1017),
    .C(net946),
    .A(net1020),
    .Y(_0357_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net944));
 sg13g2_nor2b_1 _3509_ (.A(_0356_),
    .B_N(_0357_),
    .Y(_0358_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3510_ (.Y(_0359_),
    .A(_0355_),
    .B(_0358_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3511_ (.Y(_0360_),
    .A(_0355_),
    .B(_0358_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3512_ (.A2(_0343_),
    .A1(_0333_),
    .B1(_0341_),
    .X(_0361_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3513_ (.Y(_0362_),
    .A(net1016),
    .B(net949),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3514_ (.Y(_0363_),
    .A(net1012),
    .B(net950),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3515_ (.Y(_0364_),
    .A(net953),
    .B(net1012),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3516_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0365_),
    .B(_0363_),
    .A(_0330_));
 sg13g2_and2_1 _3517_ (.A(_0329_),
    .B(_0364_),
    .X(_0366_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3518_ (.Y(_0367_),
    .A(_0329_),
    .B(_0364_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3519_ (.Y(_0368_),
    .A(_0362_),
    .B(_0367_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3520_ (.B1(_0337_),
    .VDD(VPWR),
    .Y(_0369_),
    .VSS(VGND),
    .A1(_0335_),
    .A2(_0338_));
 sg13g2_nand2_1 _3521_ (.Y(_0370_),
    .A(net954),
    .B(net1009),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3522_ (.A(net961),
    .B(net957),
    .C(net1007),
    .D(net1006),
    .X(_0371_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3523_ (.B(net957),
    .C(net1007),
    .A(net961),
    .Y(_0372_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net1006));
 sg13g2_a22oi_1 _3524_ (.Y(_0373_),
    .B1(net1006),
    .B2(net962),
    .A2(net1007),
    .A1(net957),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3525_ (.A(_0370_),
    .B(_0371_),
    .C(_0373_),
    .X(_0374_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3526_ (.B1(_0370_),
    .VDD(VPWR),
    .Y(_0375_),
    .VSS(VGND),
    .A1(_0371_),
    .A2(_0373_));
 sg13g2_and3_1 _3527_ (.X(_0376_),
    .A(_0369_),
    .B(_0374_),
    .C(_0375_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3528_ (.B(_0374_),
    .C(_0375_),
    .A(_0369_),
    .Y(_0377_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3529_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0374_),
    .A2(_0375_),
    .Y(_0378_),
    .B1(_0369_));
 sg13g2_or3_1 _3530_ (.A(_0368_),
    .B(_0376_),
    .C(_0378_),
    .X(_0379_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3531_ (.B1(_0368_),
    .VDD(VPWR),
    .Y(_0380_),
    .VSS(VGND),
    .A1(_0376_),
    .A2(_0378_));
 sg13g2_and3_1 _3532_ (.X(_0381_),
    .A(_0361_),
    .B(_0379_),
    .C(_0380_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3533_ (.B(_0379_),
    .C(_0380_),
    .A(_0361_),
    .Y(_0382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3534_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0379_),
    .A2(_0380_),
    .Y(_0383_),
    .B1(_0361_));
 sg13g2_or3_1 _3535_ (.A(_0360_),
    .B(_0381_),
    .C(_0383_),
    .X(_0384_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3536_ (.B1(_0360_),
    .VDD(VPWR),
    .Y(_0385_),
    .VSS(VGND),
    .A1(_0381_),
    .A2(_0383_));
 sg13g2_nand3_1 _3537_ (.B(_0384_),
    .C(_0385_),
    .A(_0354_),
    .Y(_0386_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3538_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0384_),
    .A2(_0385_),
    .Y(_0387_),
    .B1(_0354_));
 sg13g2_a21o_1 _3539_ (.A2(_0385_),
    .A1(_0384_),
    .B1(_0354_),
    .X(_0388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3540_ (.Y(_0389_),
    .A(_0386_),
    .B(_0388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3541_ (.B(_0389_),
    .A(_0325_),
    .X(_0390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _3542_ (.A2(_0353_),
    .A1(_0352_),
    .B1(_0351_),
    .X(_0391_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3543_ (.Y(_0392_),
    .A(_0390_),
    .B(_0391_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3544_ (.B(_0391_),
    .A(_0390_),
    .X(_0113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3545_ (.B1(_0382_),
    .VDD(VPWR),
    .Y(_0393_),
    .VSS(VGND),
    .A1(_0360_),
    .A2(_0383_));
 sg13g2_o21ai_1 _3546_ (.B1(_0365_),
    .VDD(VPWR),
    .Y(_0394_),
    .VSS(VGND),
    .A1(_0362_),
    .A2(_0366_));
 sg13g2_nand2_1 _3547_ (.Y(_0395_),
    .A(net1020),
    .B(net1032),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3548_ (.Y(_0396_),
    .A(net1016),
    .B(net944),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3549_ (.A(net1017),
    .B(net1016),
    .C(net946),
    .D(net944),
    .X(_0397_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3550_ (.Y(_0398_),
    .B1(net944),
    .B2(net1017),
    .A2(net946),
    .A1(net1016),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3551_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0399_),
    .B(_0398_),
    .A(_0397_));
 sg13g2_nor2_1 _3552_ (.A(_0395_),
    .B(_0399_),
    .Y(_0400_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3553_ (.B(_0399_),
    .A(_0395_),
    .X(_0401_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3554_ (.Y(_0402_),
    .A(_0394_),
    .B(_0401_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3555_ (.Y(_0403_),
    .A(_0394_),
    .B(_0401_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3556_ (.Y(_0404_),
    .A(_0357_),
    .B(_0403_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3557_ (.B1(_0377_),
    .VDD(VPWR),
    .Y(_0405_),
    .VSS(VGND),
    .A1(_0368_),
    .A2(_0378_));
 sg13g2_nand2_1 _3558_ (.Y(_0406_),
    .A(net1014),
    .B(net949),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3559_ (.Y(_0407_),
    .A(net950),
    .B(net1010),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3560_ (.Y(_0408_),
    .A(net952),
    .B(net1010),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3561_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0409_),
    .B(_0407_),
    .A(_0364_));
 sg13g2_xnor2_1 _3562_ (.Y(_0410_),
    .A(_0363_),
    .B(_0408_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3563_ (.Y(_0411_),
    .A(_0406_),
    .B(_0410_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3564_ (.B1(_0372_),
    .VDD(VPWR),
    .Y(_0412_),
    .VSS(VGND),
    .A1(_0370_),
    .A2(_0373_));
 sg13g2_nand2_1 _3565_ (.Y(_0413_),
    .A(net955),
    .B(net1007),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3566_ (.A(net961),
    .B(net957),
    .C(net1006),
    .D(net1037),
    .X(_0414_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3567_ (.B(net957),
    .C(net1006),
    .A(net961),
    .Y(_0415_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net1037));
 sg13g2_a22oi_1 _3568_ (.Y(_0416_),
    .B1(net1037),
    .B2(net961),
    .A2(net1006),
    .A1(net957),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3569_ (.A(_0413_),
    .B(_0414_),
    .C(_0416_),
    .X(_0417_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3570_ (.B1(_0413_),
    .VDD(VPWR),
    .Y(_0418_),
    .VSS(VGND),
    .A1(_0414_),
    .A2(_0416_));
 sg13g2_and3_1 _3571_ (.X(_0419_),
    .A(_0412_),
    .B(_0417_),
    .C(_0418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3572_ (.B(_0417_),
    .C(_0418_),
    .A(_0412_),
    .Y(_0420_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3573_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0417_),
    .A2(_0418_),
    .Y(_0421_),
    .B1(_0412_));
 sg13g2_or3_1 _3574_ (.A(_0411_),
    .B(_0419_),
    .C(_0421_),
    .X(_0422_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3575_ (.B1(_0411_),
    .VDD(VPWR),
    .Y(_0423_),
    .VSS(VGND),
    .A1(_0419_),
    .A2(_0421_));
 sg13g2_and3_1 _3576_ (.X(_0424_),
    .A(_0405_),
    .B(_0422_),
    .C(_0423_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3577_ (.B(_0422_),
    .C(_0423_),
    .A(_0405_),
    .Y(_0425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3578_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0422_),
    .A2(_0423_),
    .Y(_0426_),
    .B1(_0405_));
 sg13g2_or3_1 _3579_ (.A(_0404_),
    .B(_0424_),
    .C(_0426_),
    .X(_0427_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3580_ (.B1(_0404_),
    .VDD(VPWR),
    .Y(_0428_),
    .VSS(VGND),
    .A1(_0424_),
    .A2(_0426_));
 sg13g2_and3_1 _3581_ (.X(_0429_),
    .A(_0393_),
    .B(_0427_),
    .C(_0428_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3582_ (.B(_0427_),
    .C(_0428_),
    .A(_0393_),
    .Y(_0430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3583_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0427_),
    .A2(_0428_),
    .Y(_0431_),
    .B1(_0393_));
 sg13g2_or3_1 _3584_ (.A(_0359_),
    .B(_0429_),
    .C(_0431_),
    .X(_0432_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3585_ (.B1(_0359_),
    .VDD(VPWR),
    .Y(_0433_),
    .VSS(VGND),
    .A1(_0429_),
    .A2(_0431_));
 sg13g2_o21ai_1 _3586_ (.B1(_0386_),
    .VDD(VPWR),
    .Y(_0434_),
    .VSS(VGND),
    .A1(_0325_),
    .A2(_0387_));
 sg13g2_nand3_1 _3587_ (.B(_0433_),
    .C(_0434_),
    .A(_0432_),
    .Y(_0435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3588_ (.A2(_0433_),
    .A1(_0432_),
    .B1(_0434_),
    .X(_0436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3589_ (.Y(_0437_),
    .A(_0435_),
    .B(_0436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3590_ (.A(_0390_),
    .B(_0391_),
    .C(_0435_),
    .D(_0436_),
    .X(_0438_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3591_ (.B(_0437_),
    .A(_0392_),
    .X(_0114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3592_ (.B1(_0435_),
    .VDD(VPWR),
    .Y(_0439_),
    .VSS(VGND),
    .A1(_0392_),
    .A2(_0437_));
 sg13g2_o21ai_1 _3593_ (.B1(_0430_),
    .VDD(VPWR),
    .Y(_0440_),
    .VSS(VGND),
    .A1(_0359_),
    .A2(_0431_));
 sg13g2_o21ai_1 _3594_ (.B1(_0402_),
    .VDD(VPWR),
    .Y(_0441_),
    .VSS(VGND),
    .A1(_0357_),
    .A2(_0403_));
 sg13g2_o21ai_1 _3595_ (.B1(_0425_),
    .VDD(VPWR),
    .Y(_0442_),
    .VSS(VGND),
    .A1(_0404_),
    .A2(_0426_));
 sg13g2_nor2_1 _3596_ (.A(_0397_),
    .B(_0400_),
    .Y(_0443_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3597_ (.B1(_0409_),
    .VDD(VPWR),
    .Y(_0444_),
    .VSS(VGND),
    .A1(_0406_),
    .A2(_0410_));
 sg13g2_nand2_1 _3598_ (.Y(_0445_),
    .A(\DP_1.matrix[1] ),
    .B(net1032),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3599_ (.Y(_0446_),
    .A(net1014),
    .B(net944),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3600_ (.Y(_0447_),
    .A(net1014),
    .B(net946),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3601_ (.B(_0447_),
    .A(_0396_),
    .X(_0448_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3602_ (.Y(_0449_),
    .B(_0448_),
    .A_N(_0445_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3603_ (.Y(_0450_),
    .A(_0445_),
    .B(_0448_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3604_ (.Y(_0451_),
    .A(_0444_),
    .B(_0450_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3605_ (.A(_0443_),
    .B(_0451_),
    .Y(_0452_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3606_ (.Y(_0453_),
    .A(_0443_),
    .B(_0451_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3607_ (.B1(_0420_),
    .VDD(VPWR),
    .Y(_0454_),
    .VSS(VGND),
    .A1(_0411_),
    .A2(_0421_));
 sg13g2_nand2_1 _3608_ (.Y(_0455_),
    .A(net1012),
    .B(net949),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3609_ (.Y(_0456_),
    .A(net952),
    .B(net1008),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3610_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0457_),
    .B(_0456_),
    .A(_0407_));
 sg13g2_and2_1 _3611_ (.A(_0407_),
    .B(_0456_),
    .X(_0458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3612_ (.Y(_0459_),
    .A(_0407_),
    .B(_0456_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3613_ (.Y(_0460_),
    .A(_0455_),
    .B(_0459_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3614_ (.B1(_0415_),
    .VDD(VPWR),
    .Y(_0461_),
    .VSS(VGND),
    .A1(_0413_),
    .A2(_0416_));
 sg13g2_nand2_1 _3615_ (.Y(_0462_),
    .A(net955),
    .B(net1038),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3616_ (.A(net957),
    .B(net955),
    .C(net1005),
    .D(net1038),
    .X(_0463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3617_ (.Y(_0464_),
    .B1(net1038),
    .B2(net958),
    .A2(net1005),
    .A1(net955),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3618_ (.A(_0463_),
    .B(_0464_),
    .Y(_0465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3619_ (.Y(_0466_),
    .A(_0461_),
    .B(_0465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3620_ (.Y(_0467_),
    .A(_0461_),
    .B(_0465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3621_ (.B(_0467_),
    .A(_0460_),
    .X(_0468_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3622_ (.Y(_0469_),
    .A(_0454_),
    .B(_0468_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3623_ (.Y(_0470_),
    .A(_0454_),
    .B(_0468_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3624_ (.B(_0470_),
    .A(_0453_),
    .X(_0471_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3625_ (.Y(_0472_),
    .A(_0442_),
    .B(_0471_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3626_ (.Y(_0473_),
    .A(_0442_),
    .B(_0471_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3627_ (.Y(_0474_),
    .B(_0441_),
    .A_N(_0473_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3628_ (.Y(_0475_),
    .A(_0441_),
    .B(_0473_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3629_ (.A(_0440_),
    .B(_0475_),
    .Y(_0476_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3630_ (.Y(_0477_),
    .A(_0440_),
    .B(_0475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3631_ (.A(_0476_),
    .B_N(_0477_),
    .Y(_0478_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3632_ (.B(_0478_),
    .A(_0439_),
    .X(_0115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3633_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0444_),
    .A2(_0450_),
    .Y(_0479_),
    .B1(_0452_));
 sg13g2_o21ai_1 _3634_ (.B1(_0469_),
    .VDD(VPWR),
    .Y(_0480_),
    .VSS(VGND),
    .A1(_0453_),
    .A2(_0470_));
 sg13g2_o21ai_1 _3635_ (.B1(_0449_),
    .VDD(VPWR),
    .Y(_0481_),
    .VSS(VGND),
    .A1(_0396_),
    .A2(_0447_));
 sg13g2_o21ai_1 _3636_ (.B1(_0457_),
    .VDD(VPWR),
    .Y(_0482_),
    .VSS(VGND),
    .A1(_0455_),
    .A2(_0458_));
 sg13g2_nand2_1 _3637_ (.Y(_0483_),
    .A(net1016),
    .B(net1032),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3638_ (.Y(_0484_),
    .A(net1012),
    .B(net945),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3639_ (.Y(_0485_),
    .A(net1012),
    .B(net946),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3640_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0486_),
    .B(_0484_),
    .A(_0447_));
 sg13g2_xnor2_1 _3641_ (.Y(_0487_),
    .A(_0446_),
    .B(_0485_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3642_ (.B(_0487_),
    .A(_0483_),
    .X(_0488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3643_ (.Y(_0489_),
    .A(_0482_),
    .B(_0488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3644_ (.A(_0489_),
    .B_N(_0481_),
    .Y(_0490_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3645_ (.B(_0489_),
    .A(_0481_),
    .X(_0491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3646_ (.B1(_0466_),
    .VDD(VPWR),
    .Y(_0492_),
    .VSS(VGND),
    .A1(_0460_),
    .A2(_0467_));
 sg13g2_a21oi_1 _3647_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net958),
    .A2(net1005),
    .Y(_0493_),
    .B1(_0462_));
 sg13g2_nand2_1 _3648_ (.Y(_0494_),
    .A(net1010),
    .B(\DP_2.matrix[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3649_ (.Y(_0495_),
    .A(net950),
    .B(\DP_1.matrix[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3650_ (.A(net953),
    .B(net950),
    .C(net1008),
    .D(net1005),
    .X(_0496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3651_ (.Y(_0497_),
    .B1(net1005),
    .B2(net953),
    .A2(net1008),
    .A1(net950),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3652_ (.A(_0494_),
    .B(_0496_),
    .C(_0497_),
    .Y(_0498_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3653_ (.B1(_0494_),
    .VDD(VPWR),
    .Y(_0499_),
    .VSS(VGND),
    .A1(_0496_),
    .A2(_0497_));
 sg13g2_nor2b_1 _3654_ (.A(_0498_),
    .B_N(_0499_),
    .Y(_0500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3655_ (.Y(_0501_),
    .A(_0493_),
    .B(_0500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3656_ (.Y(_0502_),
    .B(_0492_),
    .A_N(_0501_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3657_ (.B(_0501_),
    .A(_0492_),
    .X(_0503_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3658_ (.B(_0503_),
    .A(_0491_),
    .X(_0504_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3659_ (.Y(_0505_),
    .A(_0480_),
    .B(_0504_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3660_ (.B(_0504_),
    .A(_0480_),
    .X(_0506_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3661_ (.Y(_0507_),
    .B(_0506_),
    .A_N(_0479_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3662_ (.B(_0506_),
    .A(_0479_),
    .X(_0508_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3663_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0472_),
    .A2(_0474_),
    .Y(_0509_),
    .B1(_0508_));
 sg13g2_nand3_1 _3664_ (.B(_0474_),
    .C(_0508_),
    .A(_0472_),
    .Y(_0510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3665_ (.Y(_0511_),
    .B(_0510_),
    .A_N(_0509_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3666_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0435_),
    .A2(_0477_),
    .Y(_0512_),
    .B1(_0476_));
 sg13g2_a21oi_2 _3667_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0512_),
    .Y(_0513_),
    .A2(_0478_),
    .A1(_0438_));
 sg13g2_nor2_1 _3668_ (.A(_0511_),
    .B(_0513_),
    .Y(_0514_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3669_ (.B(_0513_),
    .A(_0511_),
    .X(_0106_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3670_ (.A2(_0488_),
    .A1(_0482_),
    .B1(_0490_),
    .X(_0515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3671_ (.B1(_0502_),
    .VDD(VPWR),
    .Y(_0516_),
    .VSS(VGND),
    .A1(_0491_),
    .A2(_0503_));
 sg13g2_a21o_2 _3672_ (.A2(_0500_),
    .A1(_0493_),
    .B1(_0463_),
    .X(_0517_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3673_ (.Y(_0518_),
    .A(\DP_2.matrix[5] ),
    .B(net1008),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3674_ (.Y(_0519_),
    .A(net953),
    .B(net1037),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3675_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0520_),
    .B(_0519_),
    .A(_0495_));
 sg13g2_xnor2_1 _3676_ (.Y(_0521_),
    .A(_0495_),
    .B(_0519_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3677_ (.B(_0521_),
    .A(_0518_),
    .X(_0522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3678_ (.A(_0517_),
    .B(_0522_),
    .X(_0523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3679_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0524_),
    .B(_0522_),
    .A(_0517_));
 sg13g2_xnor2_1 _3680_ (.Y(_0525_),
    .A(_0517_),
    .B(_0522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3681_ (.B1(_0486_),
    .VDD(VPWR),
    .Y(_0526_),
    .VSS(VGND),
    .A1(_0483_),
    .A2(_0487_));
 sg13g2_or2_1 _3682_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0527_),
    .B(_0498_),
    .A(_0496_));
 sg13g2_nand2_1 _3683_ (.Y(_0528_),
    .A(net1014),
    .B(net1032),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3684_ (.Y(_0529_),
    .A(net1010),
    .B(net946),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3685_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0530_),
    .B(_0529_),
    .A(_0484_));
 sg13g2_xnor2_1 _3686_ (.Y(_0531_),
    .A(_0484_),
    .B(_0529_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3687_ (.B(_0531_),
    .A(_0528_),
    .X(_0532_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3688_ (.Y(_0533_),
    .A(_0527_),
    .B(_0532_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3689_ (.A(_0533_),
    .B_N(_0526_),
    .Y(_0534_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3690_ (.Y(_0535_),
    .A(_0526_),
    .B(_0533_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3691_ (.Y(_0536_),
    .A(_0525_),
    .B(_0535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3692_ (.Y(_0537_),
    .A(_0516_),
    .B(_0536_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3693_ (.A(_0537_),
    .B_N(_0515_),
    .Y(_0538_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3694_ (.B(_0537_),
    .A(_0515_),
    .X(_0539_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3695_ (.B(_0507_),
    .C(_0539_),
    .A(_0505_),
    .Y(_0540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3696_ (.VDD(VPWR),
    .Y(_0541_),
    .A(_0540_),
    .VSS(VGND));
 sg13g2_a21oi_1 _3697_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0505_),
    .A2(_0507_),
    .Y(_0542_),
    .B1(_0539_));
 sg13g2_nor2_1 _3698_ (.A(_0541_),
    .B(_0542_),
    .Y(_0543_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3699_ (.A(_0509_),
    .B(_0514_),
    .Y(_0544_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3700_ (.Y(_0107_),
    .A(_0543_),
    .B(_0544_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3701_ (.A2(_0532_),
    .A1(_0527_),
    .B1(_0534_),
    .X(_0545_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3702_ (.Y(_0546_),
    .B1(net1037),
    .B2(net951),
    .A2(\DP_1.matrix[7] ),
    .A1(\DP_2.matrix[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3703_ (.Y(_0547_),
    .A(net949),
    .B(net1038),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3704_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0548_),
    .B(_0547_),
    .A(_0495_));
 sg13g2_nand2b_1 _3705_ (.Y(_0549_),
    .B(_0548_),
    .A_N(_0546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3706_ (.B1(_0530_),
    .VDD(VPWR),
    .Y(_0550_),
    .VSS(VGND),
    .A1(_0528_),
    .A2(_0531_));
 sg13g2_o21ai_1 _3707_ (.B1(_0520_),
    .VDD(VPWR),
    .Y(_0551_),
    .VSS(VGND),
    .A1(_0518_),
    .A2(_0521_));
 sg13g2_nand2_1 _3708_ (.Y(_0552_),
    .A(net1012),
    .B(net1032),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3709_ (.Y(_0553_),
    .A(net1008),
    .B(net945),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3710_ (.A(net1010),
    .B(\DP_1.matrix[6] ),
    .C(net947),
    .D(net945),
    .X(_0554_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3711_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0555_),
    .B(_0553_),
    .A(_0529_));
 sg13g2_a22oi_1 _3712_ (.Y(_0556_),
    .B1(net945),
    .B2(\DP_1.matrix[5] ),
    .A2(net947),
    .A1(net1008),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3713_ (.A(_0554_),
    .B(_0556_),
    .Y(_0557_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3714_ (.Y(_0558_),
    .A(_0552_),
    .B(_0557_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3715_ (.Y(_0559_),
    .A(_0551_),
    .B(_0558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3716_ (.A(_0559_),
    .B_N(_0550_),
    .Y(_0560_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3717_ (.B(_0559_),
    .A(_0550_),
    .X(_0561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3718_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0562_),
    .B(_0561_),
    .A(_0549_));
 sg13g2_xor2_1 _3719_ (.B(_0561_),
    .A(_0549_),
    .X(_0563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3720_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0524_),
    .A2(_0535_),
    .Y(_0564_),
    .B1(_0523_));
 sg13g2_nor2b_1 _3721_ (.A(_0564_),
    .B_N(_0563_),
    .Y(_0565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3722_ (.B(_0564_),
    .A(_0563_),
    .X(_0566_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3723_ (.A(_0566_),
    .B_N(_0545_),
    .Y(_0567_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3724_ (.B(_0566_),
    .A(_0545_),
    .X(_0568_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3725_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0516_),
    .A2(_0536_),
    .Y(_0569_),
    .B1(_0538_));
 sg13g2_nor2_1 _3726_ (.A(_0568_),
    .B(_0569_),
    .Y(_0570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3727_ (.B(_0569_),
    .A(_0568_),
    .X(_0571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3728_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0509_),
    .A2(_0540_),
    .Y(_0572_),
    .B1(_0542_));
 sg13g2_a21oi_1 _3729_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0510_),
    .A2(_0540_),
    .Y(_0573_),
    .B1(_0542_));
 sg13g2_a21oi_1 _3730_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0513_),
    .A2(_0572_),
    .Y(_0574_),
    .B1(_0573_));
 sg13g2_xor2_1 _3731_ (.B(_0574_),
    .A(_0571_),
    .X(_0108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3732_ (.A2(_0558_),
    .A1(_0551_),
    .B1(_0560_),
    .X(_0575_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3733_ (.B1(_0555_),
    .VDD(VPWR),
    .Y(_0576_),
    .VSS(VGND),
    .A1(_0552_),
    .A2(_0556_));
 sg13g2_nand2_1 _3734_ (.Y(_0577_),
    .A(net1010),
    .B(net1032),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3735_ (.Y(_0578_),
    .A(net1005),
    .B(net944),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3736_ (.Y(_0579_),
    .A(net947),
    .B(net1005),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3737_ (.B(_0579_),
    .A(_0553_),
    .X(_0580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3738_ (.Y(_0581_),
    .B(_0580_),
    .A_N(_0577_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3739_ (.Y(_0582_),
    .A(_0577_),
    .B(_0580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3740_ (.A(_0548_),
    .B_N(_0582_),
    .Y(_0583_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3741_ (.Y(_0584_),
    .A(_0548_),
    .B(_0582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3742_ (.Y(_0585_),
    .A(_0576_),
    .B(_0584_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3743_ (.A(_0547_),
    .B(_0585_),
    .Y(_0586_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3744_ (.Y(_0587_),
    .A(_0547_),
    .B(_0585_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3745_ (.A(_0562_),
    .B(_0587_),
    .Y(_0588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3746_ (.B(_0587_),
    .A(_0562_),
    .X(_0589_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3747_ (.B(_0589_),
    .A(_0575_),
    .X(_0590_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3748_ (.B1(_0590_),
    .VDD(VPWR),
    .Y(_0591_),
    .VSS(VGND),
    .A1(_0565_),
    .A2(_0567_));
 sg13g2_or3_1 _3749_ (.A(_0565_),
    .B(_0567_),
    .C(_0590_),
    .X(_0592_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3750_ (.A(_0591_),
    .B(_0592_),
    .X(_0593_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3751_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0571_),
    .A2(_0574_),
    .Y(_0594_),
    .B1(_0570_));
 sg13g2_xnor2_1 _3752_ (.Y(_0109_),
    .A(_0593_),
    .B(_0594_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3753_ (.Y(_0595_),
    .A(_0571_),
    .B(_0593_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3754_ (.VDD(VPWR),
    .Y(_0596_),
    .A(_0595_),
    .VSS(VGND));
 sg13g2_o21ai_1 _3755_ (.B1(_0591_),
    .VDD(VPWR),
    .Y(_0597_),
    .VSS(VGND),
    .A1(_0568_),
    .A2(_0569_));
 sg13g2_a22oi_1 _3756_ (.Y(_0598_),
    .B1(_0597_),
    .B2(_0592_),
    .A2(_0596_),
    .A1(_0574_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3757_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0575_),
    .A2(_0589_),
    .Y(_0599_),
    .B1(_0588_));
 sg13g2_a21o_1 _3758_ (.A2(_0584_),
    .A1(_0576_),
    .B1(_0583_),
    .X(_0600_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3759_ (.B1(_0581_),
    .VDD(VPWR),
    .Y(_0601_),
    .VSS(VGND),
    .A1(_0553_),
    .A2(_0579_));
 sg13g2_nand2_1 _3760_ (.Y(_0602_),
    .A(\DP_1.matrix[6] ),
    .B(\DP_2.matrix[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3761_ (.Y(_0603_),
    .A(net944),
    .B(net1038),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3762_ (.Y(_0604_),
    .A(net947),
    .B(net1037),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3763_ (.B(_0604_),
    .A(_0578_),
    .X(_0605_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3764_ (.Y(_0606_),
    .B(_0605_),
    .A_N(_0602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3765_ (.Y(_0607_),
    .A(_0602_),
    .B(_0605_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3766_ (.Y(_0608_),
    .A(_0601_),
    .B(_0607_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3767_ (.B(_0607_),
    .A(_0601_),
    .X(_0609_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3768_ (.Y(_0610_),
    .A(_0586_),
    .B(_0609_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3769_ (.A(_0610_),
    .B_N(_0600_),
    .Y(_0611_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3770_ (.B(_0610_),
    .A(_0600_),
    .X(_0612_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3771_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0613_),
    .B(_0612_),
    .A(_0599_));
 sg13g2_xor2_1 _3772_ (.B(_0612_),
    .A(_0599_),
    .X(_0614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3773_ (.VDD(VPWR),
    .Y(_0615_),
    .A(_0614_),
    .VSS(VGND));
 sg13g2_xnor2_1 _3774_ (.Y(_0110_),
    .A(_0598_),
    .B(_0614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3775_ (.B1(_0613_),
    .VDD(VPWR),
    .Y(_0616_),
    .VSS(VGND),
    .A1(_0598_),
    .A2(_0615_));
 sg13g2_a21oi_1 _3776_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0586_),
    .A2(_0609_),
    .Y(_0617_),
    .B1(_0611_));
 sg13g2_o21ai_1 _3777_ (.B1(_0606_),
    .VDD(VPWR),
    .Y(_0618_),
    .VSS(VGND),
    .A1(_0578_),
    .A2(_0604_));
 sg13g2_nand2_1 _3778_ (.Y(_0619_),
    .A(net1005),
    .B(\DP_2.matrix[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3779_ (.B(_0619_),
    .A(_0603_),
    .X(_0620_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3780_ (.Y(_0621_),
    .A(_0618_),
    .B(_0620_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3781_ (.Y(_0622_),
    .A(_0608_),
    .B(_0621_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3782_ (.Y(_0623_),
    .A(_0617_),
    .B(_0622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3783_ (.Y(_0111_),
    .A(_0616_),
    .B(_0623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3784_ (.A(net1003),
    .B(net943),
    .X(_0074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _3785_ (.X(_0624_),
    .A(net1002),
    .B(net940),
    .C(_0074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3786_ (.Y(_0625_),
    .B1(net940),
    .B2(net1003),
    .A2(net1002),
    .A1(net943),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3787_ (.A(_0624_),
    .B(net432),
    .Y(_0075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3788_ (.Y(_0626_),
    .A(net1003),
    .B(net936),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3789_ (.A(net943),
    .B(net1002),
    .C(net940),
    .D(net1000),
    .X(_0627_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3790_ (.Y(_0628_),
    .B1(net1000),
    .B2(net943),
    .A2(net940),
    .A1(net1002),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3791_ (.A(_0626_),
    .B(_0627_),
    .C(_0628_),
    .Y(_0629_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3792_ (.B1(_0626_),
    .VDD(VPWR),
    .Y(_0630_),
    .VSS(VGND),
    .A1(_0627_),
    .A2(_0628_));
 sg13g2_nor2b_2 _3793_ (.A(_0629_),
    .B_N(_0630_),
    .Y(_0631_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3794_ (.Y(_0632_),
    .A(_0624_),
    .B(_0631_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3795_ (.B(_0631_),
    .A(_0624_),
    .X(_0076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3796_ (.Y(_0633_),
    .A(net1003),
    .B(net934),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3797_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0634_),
    .B(_0629_),
    .A(_0627_));
 sg13g2_nand2_1 _3798_ (.Y(_0635_),
    .A(net1002),
    .B(net936),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3799_ (.A(net943),
    .B(net940),
    .C(net1000),
    .D(net998),
    .X(_0636_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3800_ (.B(net940),
    .C(net1000),
    .A(net943),
    .Y(_0637_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net998));
 sg13g2_a22oi_1 _3801_ (.Y(_0638_),
    .B1(net998),
    .B2(net943),
    .A2(net1000),
    .A1(net940),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3802_ (.A(_0635_),
    .B(_0636_),
    .C(_0638_),
    .Y(_0639_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3803_ (.B1(_0635_),
    .VDD(VPWR),
    .Y(_0640_),
    .VSS(VGND),
    .A1(_0636_),
    .A2(_0638_));
 sg13g2_nor2b_1 _3804_ (.A(_0639_),
    .B_N(_0640_),
    .Y(_0641_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3805_ (.Y(_0642_),
    .A(_0634_),
    .B(_0641_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3806_ (.Y(_0643_),
    .A(_0634_),
    .B(_0641_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3807_ (.B(_0643_),
    .A(_0633_),
    .X(_0644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3808_ (.Y(_0645_),
    .B(_0644_),
    .A_N(_0632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3809_ (.Y(_0077_),
    .A(_0632_),
    .B(_0644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3810_ (.Y(_0646_),
    .B1(net932),
    .B2(net1003),
    .A2(net933),
    .A1(net1001),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3811_ (.Y(_0647_),
    .A(net1001),
    .B(net932),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3812_ (.A(net1003),
    .B(net1001),
    .C(net933),
    .D(net932),
    .X(_0648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3813_ (.A(_0646_),
    .B(_0648_),
    .Y(_0649_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3814_ (.VDD(VPWR),
    .Y(_0650_),
    .A(_0649_),
    .VSS(VGND));
 sg13g2_o21ai_1 _3815_ (.B1(_0637_),
    .VDD(VPWR),
    .Y(_0651_),
    .VSS(VGND),
    .A1(_0635_),
    .A2(_0638_));
 sg13g2_nand2_1 _3816_ (.Y(_0652_),
    .A(net999),
    .B(net935),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3817_ (.A(net942),
    .B(net939),
    .C(net998),
    .D(net996),
    .X(_0653_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3818_ (.B(net939),
    .C(net997),
    .A(net942),
    .Y(_0654_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net994));
 sg13g2_a22oi_1 _3819_ (.Y(_0655_),
    .B1(net996),
    .B2(net942),
    .A2(net997),
    .A1(net939),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3820_ (.A(_0652_),
    .B(_0653_),
    .C(_0655_),
    .X(_0656_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3821_ (.B1(_0652_),
    .VDD(VPWR),
    .Y(_0657_),
    .VSS(VGND),
    .A1(_0653_),
    .A2(_0655_));
 sg13g2_nand3_1 _3822_ (.B(_0656_),
    .C(_0657_),
    .A(_0651_),
    .Y(_0658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3823_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0656_),
    .A2(_0657_),
    .Y(_0659_),
    .B1(_0651_));
 sg13g2_a21o_1 _3824_ (.A2(_0657_),
    .A1(_0656_),
    .B1(_0651_),
    .X(_0660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3825_ (.Y(_0661_),
    .A(_0658_),
    .B(_0660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3826_ (.Y(_0662_),
    .A(_0650_),
    .B(_0661_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3827_ (.B1(_0642_),
    .VDD(VPWR),
    .Y(_0663_),
    .VSS(VGND),
    .A1(_0633_),
    .A2(_0643_));
 sg13g2_nor2b_2 _3828_ (.A(_0662_),
    .B_N(_0663_),
    .Y(_0664_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3829_ (.B(_0663_),
    .A(_0662_),
    .X(_0665_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3830_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0666_),
    .B(_0665_),
    .A(_0645_));
 sg13g2_xor2_1 _3831_ (.B(_0665_),
    .A(_0645_),
    .X(_0078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3832_ (.B1(_0658_),
    .VDD(VPWR),
    .Y(_0667_),
    .VSS(VGND),
    .A1(_0650_),
    .A2(_0659_));
 sg13g2_nand2_1 _3833_ (.Y(_0668_),
    .A(net1003),
    .B(net929),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3834_ (.Y(_0669_),
    .A(net999),
    .B(net931),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3835_ (.Y(_0670_),
    .A(net1000),
    .B(net933),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3836_ (.B(_0670_),
    .A(_0647_),
    .X(_0671_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3837_ (.Y(_0672_),
    .B(_0671_),
    .A_N(_0668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3838_ (.B(_0671_),
    .A(_0668_),
    .X(_0673_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3839_ (.B1(_0654_),
    .VDD(VPWR),
    .Y(_0674_),
    .VSS(VGND),
    .A1(_0652_),
    .A2(_0655_));
 sg13g2_nand2_1 _3840_ (.Y(_0675_),
    .A(net935),
    .B(net997),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3841_ (.A(net942),
    .B(net939),
    .C(net994),
    .D(net993),
    .X(_0676_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3842_ (.B(net939),
    .C(net994),
    .A(net941),
    .Y(_0677_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net993));
 sg13g2_a22oi_1 _3843_ (.Y(_0678_),
    .B1(net993),
    .B2(net942),
    .A2(net994),
    .A1(net939),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3844_ (.A(_0675_),
    .B(_0676_),
    .C(_0678_),
    .X(_0679_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3845_ (.B1(_0675_),
    .VDD(VPWR),
    .Y(_0680_),
    .VSS(VGND),
    .A1(_0676_),
    .A2(_0678_));
 sg13g2_and3_1 _3846_ (.X(_0681_),
    .A(_0674_),
    .B(_0679_),
    .C(_0680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3847_ (.B(_0679_),
    .C(_0680_),
    .A(_0674_),
    .Y(_0682_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3848_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0679_),
    .A2(_0680_),
    .Y(_0683_),
    .B1(_0674_));
 sg13g2_or3_1 _3849_ (.A(_0673_),
    .B(_0681_),
    .C(_0683_),
    .X(_0684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3850_ (.B1(_0673_),
    .VDD(VPWR),
    .Y(_0685_),
    .VSS(VGND),
    .A1(_0681_),
    .A2(_0683_));
 sg13g2_nand3_1 _3851_ (.B(_0684_),
    .C(_0685_),
    .A(_0667_),
    .Y(_0686_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3852_ (.A2(_0685_),
    .A1(_0684_),
    .B1(_0667_),
    .X(_0687_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3853_ (.B(_0686_),
    .C(_0687_),
    .A(_0648_),
    .Y(_0688_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3854_ (.A2(_0687_),
    .A1(_0686_),
    .B1(_0648_),
    .X(_0689_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3855_ (.A(_0688_),
    .B(_0689_),
    .X(_0690_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3856_ (.B(_0688_),
    .C(_0689_),
    .A(_0664_),
    .Y(_0691_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3857_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0688_),
    .A2(_0689_),
    .Y(_0692_),
    .B1(_0664_));
 sg13g2_xor2_1 _3858_ (.B(_0690_),
    .A(_0664_),
    .X(_0693_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3859_ (.Y(_0116_),
    .A(_0666_),
    .B(_0693_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3860_ (.Y(_0694_),
    .A(_0686_),
    .B(_0688_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3861_ (.B1(_0672_),
    .VDD(VPWR),
    .Y(_0695_),
    .VSS(VGND),
    .A1(_0647_),
    .A2(_0670_));
 sg13g2_nand2_1 _3862_ (.Y(_0696_),
    .A(net1004),
    .B(net927),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3863_ (.Y(_0697_),
    .B(_0695_),
    .A_N(_0696_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3864_ (.B(_0696_),
    .A(_0695_),
    .X(_0698_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3865_ (.B1(_0682_),
    .VDD(VPWR),
    .Y(_0699_),
    .VSS(VGND),
    .A1(_0673_),
    .A2(_0683_));
 sg13g2_nand2_1 _3866_ (.Y(_0700_),
    .A(net1001),
    .B(net930),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3867_ (.Y(_0701_),
    .A(net998),
    .B(net931),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3868_ (.Y(_0702_),
    .A(net998),
    .B(net933),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3869_ (.B(_0702_),
    .A(_0669_),
    .X(_0703_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3870_ (.Y(_0704_),
    .B(_0703_),
    .A_N(_0700_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3871_ (.Y(_0705_),
    .A(_0700_),
    .B(_0703_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3872_ (.B1(_0677_),
    .VDD(VPWR),
    .Y(_0706_),
    .VSS(VGND),
    .A1(_0675_),
    .A2(_0678_));
 sg13g2_nand2_1 _3873_ (.Y(_0707_),
    .A(net936),
    .B(net995),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3874_ (.A(net941),
    .B(\DP_2.matrix[37] ),
    .C(net992),
    .D(net990),
    .X(_0708_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3875_ (.B(net938),
    .C(net991),
    .A(net941),
    .Y(_0709_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net990));
 sg13g2_a22oi_1 _3876_ (.Y(_0710_),
    .B1(net990),
    .B2(net941),
    .A2(net991),
    .A1(net939),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3877_ (.A(_0707_),
    .B(_0708_),
    .C(_0710_),
    .X(_0711_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3878_ (.B1(_0707_),
    .VDD(VPWR),
    .Y(_0712_),
    .VSS(VGND),
    .A1(_0708_),
    .A2(_0710_));
 sg13g2_and3_1 _3879_ (.X(_0713_),
    .A(_0706_),
    .B(_0711_),
    .C(_0712_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3880_ (.B(_0711_),
    .C(_0712_),
    .A(_0706_),
    .Y(_0714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3881_ (.A2(_0712_),
    .A1(_0711_),
    .B1(_0706_),
    .X(_0715_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3882_ (.B(_0714_),
    .C(_0715_),
    .A(_0705_),
    .Y(_0716_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3883_ (.A2(_0715_),
    .A1(_0714_),
    .B1(_0705_),
    .X(_0717_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3884_ (.B(_0716_),
    .C(_0717_),
    .A(_0699_),
    .Y(_0718_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3885_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0716_),
    .A2(_0717_),
    .Y(_0719_),
    .B1(_0699_));
 sg13g2_a21o_1 _3886_ (.A2(_0717_),
    .A1(_0716_),
    .B1(_0699_),
    .X(_0720_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3887_ (.Y(_0721_),
    .A(_0718_),
    .B(_0720_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3888_ (.Y(_0722_),
    .A(_0698_),
    .B(_0721_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3889_ (.A(_0722_),
    .B_N(_0694_),
    .Y(_0723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3890_ (.Y(_0724_),
    .A(_0694_),
    .B(_0722_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3891_ (.B1(_0691_),
    .VDD(VPWR),
    .Y(_0725_),
    .VSS(VGND),
    .A1(_0666_),
    .A2(_0692_));
 sg13g2_xor2_1 _3892_ (.B(_0725_),
    .A(_0724_),
    .X(_0123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3893_ (.B1(_0718_),
    .VDD(VPWR),
    .Y(_0726_),
    .VSS(VGND),
    .A1(_0698_),
    .A2(_0719_));
 sg13g2_o21ai_1 _3894_ (.B1(_0704_),
    .VDD(VPWR),
    .Y(_0727_),
    .VSS(VGND),
    .A1(_0669_),
    .A2(_0702_));
 sg13g2_a22oi_1 _3895_ (.Y(_0728_),
    .B1(net925),
    .B2(net1004),
    .A2(net927),
    .A1(net1001),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3896_ (.B(net1001),
    .C(net927),
    .A(net1004),
    .Y(_0729_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net925));
 sg13g2_nor2b_1 _3897_ (.A(_0728_),
    .B_N(_0729_),
    .Y(_0730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3898_ (.Y(_0731_),
    .A(_0727_),
    .B(_0730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3899_ (.Y(_0732_),
    .A(_0727_),
    .B(_0730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3900_ (.A2(_0715_),
    .A1(_0705_),
    .B1(_0713_),
    .X(_0733_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3901_ (.Y(_0734_),
    .A(net999),
    .B(net930),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3902_ (.Y(_0735_),
    .A(net995),
    .B(net931),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3903_ (.Y(_0736_),
    .A(net933),
    .B(net995),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3904_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0737_),
    .B(_0735_),
    .A(_0702_));
 sg13g2_and2_1 _3905_ (.A(_0701_),
    .B(_0736_),
    .X(_0738_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3906_ (.Y(_0739_),
    .A(_0701_),
    .B(_0736_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3907_ (.Y(_0740_),
    .A(_0734_),
    .B(_0739_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3908_ (.B1(_0709_),
    .VDD(VPWR),
    .Y(_0741_),
    .VSS(VGND),
    .A1(_0707_),
    .A2(_0710_));
 sg13g2_nand2_1 _3909_ (.Y(_0742_),
    .A(net935),
    .B(net991),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3910_ (.A(net941),
    .B(net937),
    .C(net989),
    .D(net987),
    .X(_0743_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3911_ (.B(net937),
    .C(net989),
    .A(net941),
    .Y(_0744_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net986));
 sg13g2_a22oi_1 _3912_ (.Y(_0745_),
    .B1(net987),
    .B2(net941),
    .A2(net989),
    .A1(net938),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3913_ (.A(_0742_),
    .B(_0743_),
    .C(_0745_),
    .X(_0746_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3914_ (.B1(_0742_),
    .VDD(VPWR),
    .Y(_0747_),
    .VSS(VGND),
    .A1(_0743_),
    .A2(_0745_));
 sg13g2_and3_1 _3915_ (.X(_0748_),
    .A(_0741_),
    .B(_0746_),
    .C(_0747_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3916_ (.B(_0746_),
    .C(_0747_),
    .A(_0741_),
    .Y(_0749_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3917_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0746_),
    .A2(_0747_),
    .Y(_0750_),
    .B1(_0741_));
 sg13g2_or3_1 _3918_ (.A(_0740_),
    .B(_0748_),
    .C(_0750_),
    .X(_0751_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3919_ (.B1(_0740_),
    .VDD(VPWR),
    .Y(_0752_),
    .VSS(VGND),
    .A1(_0748_),
    .A2(_0750_));
 sg13g2_and3_1 _3920_ (.X(_0753_),
    .A(_0733_),
    .B(_0751_),
    .C(_0752_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3921_ (.B(_0751_),
    .C(_0752_),
    .A(_0733_),
    .Y(_0754_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3922_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0751_),
    .A2(_0752_),
    .Y(_0755_),
    .B1(_0733_));
 sg13g2_or3_1 _3923_ (.A(_0732_),
    .B(_0753_),
    .C(_0755_),
    .X(_0756_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3924_ (.B1(_0732_),
    .VDD(VPWR),
    .Y(_0757_),
    .VSS(VGND),
    .A1(_0753_),
    .A2(_0755_));
 sg13g2_nand3_1 _3925_ (.B(_0756_),
    .C(_0757_),
    .A(_0726_),
    .Y(_0758_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3926_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0756_),
    .A2(_0757_),
    .Y(_0759_),
    .B1(_0726_));
 sg13g2_a21o_1 _3927_ (.A2(_0757_),
    .A1(_0756_),
    .B1(_0726_),
    .X(_0760_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3928_ (.Y(_0761_),
    .A(_0758_),
    .B(_0760_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3929_ (.B(_0761_),
    .A(_0697_),
    .X(_0762_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _3930_ (.A2(_0725_),
    .A1(_0724_),
    .B1(_0723_),
    .X(_0763_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3931_ (.Y(_0764_),
    .A(_0762_),
    .B(_0763_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3932_ (.B(_0763_),
    .A(_0762_),
    .X(_0124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3933_ (.B1(_0754_),
    .VDD(VPWR),
    .Y(_0765_),
    .VSS(VGND),
    .A1(_0732_),
    .A2(_0755_));
 sg13g2_o21ai_1 _3934_ (.B1(_0737_),
    .VDD(VPWR),
    .Y(_0766_),
    .VSS(VGND),
    .A1(_0734_),
    .A2(_0738_));
 sg13g2_nand2_1 _3935_ (.Y(_0767_),
    .A(net1004),
    .B(net1031),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3936_ (.Y(_0768_),
    .A(net999),
    .B(net925),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3937_ (.A(net1001),
    .B(net999),
    .C(net927),
    .D(net925),
    .X(_0769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3938_ (.Y(_0770_),
    .B1(net925),
    .B2(\DP_1.matrix[37] ),
    .A2(net927),
    .A1(net999),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3939_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0771_),
    .B(_0770_),
    .A(_0769_));
 sg13g2_nor2_1 _3940_ (.A(_0767_),
    .B(_0771_),
    .Y(_0772_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3941_ (.B(_0771_),
    .A(_0767_),
    .X(_0773_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3942_ (.Y(_0774_),
    .A(_0766_),
    .B(_0773_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3943_ (.Y(_0775_),
    .A(_0766_),
    .B(_0773_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3944_ (.Y(_0776_),
    .A(_0729_),
    .B(_0775_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3945_ (.B1(_0749_),
    .VDD(VPWR),
    .Y(_0777_),
    .VSS(VGND),
    .A1(_0740_),
    .A2(_0750_));
 sg13g2_nand2_1 _3946_ (.Y(_0778_),
    .A(net997),
    .B(net929),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3947_ (.Y(_0779_),
    .A(net931),
    .B(net991),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3948_ (.Y(_0780_),
    .A(net933),
    .B(net991),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3949_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0781_),
    .B(_0779_),
    .A(_0736_));
 sg13g2_xnor2_1 _3950_ (.Y(_0782_),
    .A(_0735_),
    .B(_0780_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3951_ (.Y(_0783_),
    .A(_0778_),
    .B(_0782_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3952_ (.B1(_0744_),
    .VDD(VPWR),
    .Y(_0784_),
    .VSS(VGND),
    .A1(_0742_),
    .A2(_0745_));
 sg13g2_nand2_1 _3953_ (.Y(_0785_),
    .A(net935),
    .B(net989),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3954_ (.A(\DP_2.matrix[36] ),
    .B(net937),
    .C(net986),
    .D(net1035),
    .X(_0786_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3955_ (.B(net937),
    .C(net986),
    .A(net941),
    .Y(_0787_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net1035));
 sg13g2_a22oi_1 _3956_ (.Y(_0788_),
    .B1(net1035),
    .B2(net942),
    .A2(net986),
    .A1(net937),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3957_ (.A(_0785_),
    .B(_0786_),
    .C(_0788_),
    .X(_0789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3958_ (.B1(_0785_),
    .VDD(VPWR),
    .Y(_0790_),
    .VSS(VGND),
    .A1(_0786_),
    .A2(_0788_));
 sg13g2_and3_1 _3959_ (.X(_0791_),
    .A(_0784_),
    .B(_0789_),
    .C(_0790_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3960_ (.B(_0789_),
    .C(_0790_),
    .A(_0784_),
    .Y(_0792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3961_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0789_),
    .A2(_0790_),
    .Y(_0793_),
    .B1(_0784_));
 sg13g2_or3_1 _3962_ (.A(_0783_),
    .B(_0791_),
    .C(_0793_),
    .X(_0794_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3963_ (.B1(_0783_),
    .VDD(VPWR),
    .Y(_0795_),
    .VSS(VGND),
    .A1(_0791_),
    .A2(_0793_));
 sg13g2_and3_1 _3964_ (.X(_0796_),
    .A(_0777_),
    .B(_0794_),
    .C(_0795_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3965_ (.B(_0794_),
    .C(_0795_),
    .A(_0777_),
    .Y(_0797_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3966_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0794_),
    .A2(_0795_),
    .Y(_0798_),
    .B1(_0777_));
 sg13g2_or3_1 _3967_ (.A(_0776_),
    .B(_0796_),
    .C(_0798_),
    .X(_0799_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3968_ (.B1(_0776_),
    .VDD(VPWR),
    .Y(_0800_),
    .VSS(VGND),
    .A1(_0796_),
    .A2(_0798_));
 sg13g2_and3_1 _3969_ (.X(_0801_),
    .A(_0765_),
    .B(_0799_),
    .C(_0800_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3970_ (.B(_0799_),
    .C(_0800_),
    .A(_0765_),
    .Y(_0802_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3971_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0799_),
    .A2(_0800_),
    .Y(_0803_),
    .B1(_0765_));
 sg13g2_or3_1 _3972_ (.A(_0731_),
    .B(_0801_),
    .C(_0803_),
    .X(_0804_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3973_ (.B1(_0731_),
    .VDD(VPWR),
    .Y(_0805_),
    .VSS(VGND),
    .A1(_0801_),
    .A2(_0803_));
 sg13g2_o21ai_1 _3974_ (.B1(_0758_),
    .VDD(VPWR),
    .Y(_0806_),
    .VSS(VGND),
    .A1(_0697_),
    .A2(_0759_));
 sg13g2_nand3_1 _3975_ (.B(_0805_),
    .C(_0806_),
    .A(_0804_),
    .Y(_0807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3976_ (.A2(_0805_),
    .A1(_0804_),
    .B1(_0806_),
    .X(_0808_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3977_ (.Y(_0809_),
    .A(_0807_),
    .B(_0808_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3978_ (.A(_0762_),
    .B(_0763_),
    .C(_0807_),
    .D(_0808_),
    .X(_0810_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3979_ (.B(_0809_),
    .A(_0764_),
    .X(_0125_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3980_ (.B1(_0807_),
    .VDD(VPWR),
    .Y(_0811_),
    .VSS(VGND),
    .A1(_0764_),
    .A2(_0809_));
 sg13g2_o21ai_1 _3981_ (.B1(_0802_),
    .VDD(VPWR),
    .Y(_0812_),
    .VSS(VGND),
    .A1(_0731_),
    .A2(_0803_));
 sg13g2_o21ai_1 _3982_ (.B1(_0774_),
    .VDD(VPWR),
    .Y(_0813_),
    .VSS(VGND),
    .A1(_0729_),
    .A2(_0775_));
 sg13g2_o21ai_1 _3983_ (.B1(_0797_),
    .VDD(VPWR),
    .Y(_0814_),
    .VSS(VGND),
    .A1(_0776_),
    .A2(_0798_));
 sg13g2_nor2_1 _3984_ (.A(_0769_),
    .B(_0772_),
    .Y(_0815_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3985_ (.B1(_0781_),
    .VDD(VPWR),
    .Y(_0816_),
    .VSS(VGND),
    .A1(_0778_),
    .A2(_0782_));
 sg13g2_nand2_1 _3986_ (.Y(_0817_),
    .A(net1002),
    .B(net1031),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3987_ (.Y(_0818_),
    .A(net997),
    .B(net925),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3988_ (.Y(_0819_),
    .A(net997),
    .B(net927),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3989_ (.B(_0819_),
    .A(_0768_),
    .X(_0820_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3990_ (.Y(_0821_),
    .B(_0820_),
    .A_N(_0817_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3991_ (.Y(_0822_),
    .A(_0817_),
    .B(_0820_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3992_ (.Y(_0823_),
    .A(_0816_),
    .B(_0822_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3993_ (.A(_0815_),
    .B(_0823_),
    .Y(_0824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3994_ (.Y(_0825_),
    .A(_0815_),
    .B(_0823_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3995_ (.B1(_0792_),
    .VDD(VPWR),
    .Y(_0826_),
    .VSS(VGND),
    .A1(_0783_),
    .A2(_0793_));
 sg13g2_nand2_1 _3996_ (.Y(_0827_),
    .A(net994),
    .B(net929),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3997_ (.Y(_0828_),
    .A(net933),
    .B(net989),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3998_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0829_),
    .B(_0828_),
    .A(_0779_));
 sg13g2_and2_1 _3999_ (.A(_0779_),
    .B(_0828_),
    .X(_0830_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4000_ (.Y(_0831_),
    .A(_0779_),
    .B(_0828_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4001_ (.Y(_0832_),
    .A(_0827_),
    .B(_0831_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4002_ (.B1(_0787_),
    .VDD(VPWR),
    .Y(_0833_),
    .VSS(VGND),
    .A1(_0785_),
    .A2(_0788_));
 sg13g2_nand2_1 _4003_ (.Y(_0834_),
    .A(net935),
    .B(net1035),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4004_ (.A(net937),
    .B(net935),
    .C(net986),
    .D(net1035),
    .X(_0835_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4005_ (.Y(_0836_),
    .B1(net1035),
    .B2(net937),
    .A2(net986),
    .A1(net935),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4006_ (.A(_0835_),
    .B(_0836_),
    .Y(_0837_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4007_ (.Y(_0838_),
    .A(_0833_),
    .B(_0837_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4008_ (.Y(_0839_),
    .A(_0833_),
    .B(_0837_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4009_ (.B(_0839_),
    .A(_0832_),
    .X(_0840_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4010_ (.Y(_0841_),
    .A(_0826_),
    .B(_0840_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4011_ (.Y(_0842_),
    .A(_0826_),
    .B(_0840_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4012_ (.B(_0842_),
    .A(_0825_),
    .X(_0843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4013_ (.Y(_0844_),
    .A(_0814_),
    .B(_0843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4014_ (.Y(_0845_),
    .A(_0814_),
    .B(_0843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4015_ (.Y(_0846_),
    .B(_0813_),
    .A_N(_0845_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4016_ (.Y(_0847_),
    .A(_0813_),
    .B(_0845_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4017_ (.A(_0812_),
    .B(_0847_),
    .Y(_0848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4018_ (.Y(_0849_),
    .A(_0812_),
    .B(_0847_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4019_ (.A(_0848_),
    .B_N(_0849_),
    .Y(_0850_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4020_ (.B(_0850_),
    .A(_0811_),
    .X(_0126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4021_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0816_),
    .A2(_0822_),
    .Y(_0851_),
    .B1(_0824_));
 sg13g2_o21ai_1 _4022_ (.B1(_0841_),
    .VDD(VPWR),
    .Y(_0852_),
    .VSS(VGND),
    .A1(_0825_),
    .A2(_0842_));
 sg13g2_o21ai_1 _4023_ (.B1(_0821_),
    .VDD(VPWR),
    .Y(_0853_),
    .VSS(VGND),
    .A1(_0768_),
    .A2(_0819_));
 sg13g2_o21ai_1 _4024_ (.B1(_0829_),
    .VDD(VPWR),
    .Y(_0854_),
    .VSS(VGND),
    .A1(_0827_),
    .A2(_0830_));
 sg13g2_nand2_1 _4025_ (.Y(_0855_),
    .A(net999),
    .B(net1031),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4026_ (.Y(_0856_),
    .A(net994),
    .B(net925),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4027_ (.Y(_0857_),
    .A(net994),
    .B(net927),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4028_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0858_),
    .B(_0856_),
    .A(_0819_));
 sg13g2_xnor2_1 _4029_ (.Y(_0859_),
    .A(_0818_),
    .B(_0857_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4030_ (.B(_0859_),
    .A(_0855_),
    .X(_0860_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4031_ (.Y(_0861_),
    .A(_0854_),
    .B(_0860_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4032_ (.A(_0861_),
    .B_N(_0853_),
    .Y(_0862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4033_ (.B(_0861_),
    .A(_0853_),
    .X(_0863_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4034_ (.B1(_0838_),
    .VDD(VPWR),
    .Y(_0864_),
    .VSS(VGND),
    .A1(_0832_),
    .A2(_0839_));
 sg13g2_a21oi_1 _4035_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net937),
    .A2(net986),
    .Y(_0865_),
    .B1(_0834_));
 sg13g2_nand2_1 _4036_ (.Y(_0866_),
    .A(net991),
    .B(net929),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4037_ (.Y(_0867_),
    .A(net931),
    .B(net988),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4038_ (.A(net934),
    .B(net931),
    .C(net990),
    .D(net987),
    .X(_0868_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4039_ (.Y(_0869_),
    .B1(net986),
    .B2(net934),
    .A2(net990),
    .A1(net931),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4040_ (.A(_0866_),
    .B(_0868_),
    .C(_0869_),
    .Y(_0870_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4041_ (.B1(_0866_),
    .VDD(VPWR),
    .Y(_0871_),
    .VSS(VGND),
    .A1(_0868_),
    .A2(_0869_));
 sg13g2_nor2b_1 _4042_ (.A(_0870_),
    .B_N(_0871_),
    .Y(_0872_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4043_ (.Y(_0873_),
    .A(_0865_),
    .B(_0872_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4044_ (.Y(_0874_),
    .B(_0864_),
    .A_N(_0873_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4045_ (.B(_0873_),
    .A(_0864_),
    .X(_0875_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4046_ (.B(_0875_),
    .A(_0863_),
    .X(_0876_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4047_ (.Y(_0877_),
    .A(_0852_),
    .B(_0876_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4048_ (.B(_0876_),
    .A(_0852_),
    .X(_0878_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4049_ (.Y(_0879_),
    .B(_0878_),
    .A_N(_0851_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4050_ (.B(_0878_),
    .A(_0851_),
    .X(_0880_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4051_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0844_),
    .A2(_0846_),
    .Y(_0881_),
    .B1(_0880_));
 sg13g2_nand3_1 _4052_ (.B(_0846_),
    .C(_0880_),
    .A(_0844_),
    .Y(_0882_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4053_ (.Y(_0883_),
    .B(_0882_),
    .A_N(_0881_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4054_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0807_),
    .A2(_0849_),
    .Y(_0884_),
    .B1(_0848_));
 sg13g2_a21oi_2 _4055_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0884_),
    .Y(_0885_),
    .A2(_0850_),
    .A1(_0810_));
 sg13g2_nor2_1 _4056_ (.A(_0883_),
    .B(_0885_),
    .Y(_0886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4057_ (.B(_0885_),
    .A(_0883_),
    .X(_0117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4058_ (.A2(_0860_),
    .A1(_0854_),
    .B1(_0862_),
    .X(_0887_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4059_ (.B1(_0874_),
    .VDD(VPWR),
    .Y(_0888_),
    .VSS(VGND),
    .A1(_0863_),
    .A2(_0875_));
 sg13g2_a21o_1 _4060_ (.A2(_0872_),
    .A1(_0865_),
    .B1(_0835_),
    .X(_0889_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4061_ (.Y(_0890_),
    .A(net929),
    .B(net989),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4062_ (.Y(_0891_),
    .A(net934),
    .B(net1035),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4063_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0892_),
    .B(_0891_),
    .A(_0867_));
 sg13g2_xnor2_1 _4064_ (.Y(_0893_),
    .A(_0867_),
    .B(_0891_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4065_ (.B(_0893_),
    .A(_0890_),
    .X(_0894_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4066_ (.Y(_0895_),
    .A(_0889_),
    .B(_0894_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4067_ (.B1(_0858_),
    .VDD(VPWR),
    .Y(_0896_),
    .VSS(VGND),
    .A1(_0855_),
    .A2(_0859_));
 sg13g2_or2_1 _4068_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0897_),
    .B(_0870_),
    .A(_0868_));
 sg13g2_nand2_1 _4069_ (.Y(_0898_),
    .A(net997),
    .B(net1031),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4070_ (.Y(_0899_),
    .A(net991),
    .B(net927),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4071_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0900_),
    .B(_0899_),
    .A(_0856_));
 sg13g2_xnor2_1 _4072_ (.Y(_0901_),
    .A(_0856_),
    .B(_0899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4073_ (.B(_0901_),
    .A(_0898_),
    .X(_0902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4074_ (.Y(_0903_),
    .A(_0897_),
    .B(_0902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4075_ (.A(_0903_),
    .B_N(_0896_),
    .Y(_0904_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4076_ (.B(_0903_),
    .A(_0896_),
    .X(_0905_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4077_ (.A(_0895_),
    .B(_0905_),
    .Y(_0906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4078_ (.B(_0905_),
    .A(_0895_),
    .X(_0907_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4079_ (.Y(_0908_),
    .A(_0888_),
    .B(_0907_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4080_ (.A(_0908_),
    .B_N(_0887_),
    .Y(_0909_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4081_ (.B(_0908_),
    .A(_0887_),
    .X(_0910_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4082_ (.B(_0879_),
    .C(_0910_),
    .A(_0877_),
    .Y(_0911_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4083_ (.VDD(VPWR),
    .Y(_0912_),
    .A(_0911_),
    .VSS(VGND));
 sg13g2_a21oi_1 _4084_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0877_),
    .A2(_0879_),
    .Y(_0913_),
    .B1(_0910_));
 sg13g2_nor2_1 _4085_ (.A(_0912_),
    .B(_0913_),
    .Y(_0914_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4086_ (.A(_0881_),
    .B(_0886_),
    .Y(_0915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4087_ (.Y(_0118_),
    .A(_0914_),
    .B(_0915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4088_ (.A2(_0902_),
    .A1(_0897_),
    .B1(_0904_),
    .X(_0916_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4089_ (.Y(_0917_),
    .B1(net1036),
    .B2(net932),
    .A2(net988),
    .A1(net929),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4090_ (.Y(_0918_),
    .A(net929),
    .B(net1036),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4091_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0919_),
    .B(_0918_),
    .A(_0867_));
 sg13g2_nand2b_1 _4092_ (.Y(_0920_),
    .B(_0919_),
    .A_N(_0917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4093_ (.B1(_0900_),
    .VDD(VPWR),
    .Y(_0921_),
    .VSS(VGND),
    .A1(_0898_),
    .A2(_0901_));
 sg13g2_o21ai_1 _4094_ (.B1(_0892_),
    .VDD(VPWR),
    .Y(_0922_),
    .VSS(VGND),
    .A1(_0890_),
    .A2(_0893_));
 sg13g2_nand2_1 _4095_ (.Y(_0923_),
    .A(net995),
    .B(net1031),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4096_ (.Y(_0924_),
    .A(net989),
    .B(net925),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4097_ (.A(_0899_),
    .B(_0924_),
    .Y(_0925_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4098_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0926_),
    .B(_0924_),
    .A(_0899_));
 sg13g2_a22oi_1 _4099_ (.Y(_0927_),
    .B1(net926),
    .B2(net991),
    .A2(net928),
    .A1(net989),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4100_ (.A(_0925_),
    .B(_0927_),
    .Y(_0928_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4101_ (.Y(_0929_),
    .A(_0923_),
    .B(_0928_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4102_ (.Y(_0930_),
    .A(_0922_),
    .B(_0929_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4103_ (.A(_0930_),
    .B_N(_0921_),
    .Y(_0931_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4104_ (.B(_0930_),
    .A(_0921_),
    .X(_0932_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4105_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0933_),
    .B(_0932_),
    .A(_0920_));
 sg13g2_xor2_1 _4106_ (.B(_0932_),
    .A(_0920_),
    .X(_0934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4107_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0889_),
    .A2(_0894_),
    .Y(_0935_),
    .B1(_0906_));
 sg13g2_nor2b_1 _4108_ (.A(_0935_),
    .B_N(_0934_),
    .Y(_0936_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4109_ (.B(_0935_),
    .A(_0934_),
    .X(_0937_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4110_ (.A(_0937_),
    .B_N(_0916_),
    .Y(_0938_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4111_ (.B(_0937_),
    .A(_0916_),
    .X(_0939_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4112_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0888_),
    .A2(_0907_),
    .Y(_0940_),
    .B1(_0909_));
 sg13g2_nor2_1 _4113_ (.A(_0939_),
    .B(_0940_),
    .Y(_0941_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4114_ (.B(_0940_),
    .A(_0939_),
    .X(_0942_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4115_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0881_),
    .A2(_0911_),
    .Y(_0943_),
    .B1(_0913_));
 sg13g2_a21oi_1 _4116_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0882_),
    .A2(_0911_),
    .Y(_0944_),
    .B1(_0913_));
 sg13g2_a21oi_2 _4117_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0944_),
    .Y(_0945_),
    .A2(_0943_),
    .A1(_0885_));
 sg13g2_xor2_1 _4118_ (.B(_0945_),
    .A(_0942_),
    .X(_0119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4119_ (.A2(_0929_),
    .A1(_0922_),
    .B1(_0931_),
    .X(_0946_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4120_ (.B1(_0926_),
    .VDD(VPWR),
    .Y(_0947_),
    .VSS(VGND),
    .A1(_0923_),
    .A2(_0927_));
 sg13g2_nand2_1 _4121_ (.Y(_0948_),
    .A(net992),
    .B(net1031),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4122_ (.Y(_0949_),
    .A(net988),
    .B(net926),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4123_ (.Y(_0950_),
    .A(net928),
    .B(net988),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4124_ (.B(_0950_),
    .A(_0924_),
    .X(_0951_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4125_ (.Y(_0952_),
    .B(_0951_),
    .A_N(_0948_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4126_ (.Y(_0953_),
    .A(_0948_),
    .B(_0951_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4127_ (.A(_0919_),
    .B_N(_0953_),
    .Y(_0954_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4128_ (.Y(_0955_),
    .A(_0919_),
    .B(_0953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4129_ (.Y(_0956_),
    .A(_0947_),
    .B(_0955_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4130_ (.A(_0918_),
    .B(_0956_),
    .Y(_0957_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4131_ (.B(_0956_),
    .A(_0918_),
    .X(_0958_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4132_ (.Y(_0959_),
    .B(_0958_),
    .A_N(_0933_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4133_ (.Y(_0960_),
    .A(_0933_),
    .B(_0958_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4134_ (.Y(_0961_),
    .A(_0946_),
    .B(_0960_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4135_ (.B(_0960_),
    .A(_0946_),
    .X(_0962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4136_ (.B1(_0962_),
    .VDD(VPWR),
    .Y(_0963_),
    .VSS(VGND),
    .A1(_0936_),
    .A2(_0938_));
 sg13g2_or3_1 _4137_ (.A(_0936_),
    .B(_0938_),
    .C(_0962_),
    .X(_0964_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4138_ (.A(_0963_),
    .B(_0964_),
    .X(_0965_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4139_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0942_),
    .A2(_0945_),
    .Y(_0966_),
    .B1(_0941_));
 sg13g2_xnor2_1 _4140_ (.Y(_0120_),
    .A(_0965_),
    .B(_0966_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4141_ (.A(_0942_),
    .B(_0965_),
    .X(_0967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4142_ (.Y(_0968_),
    .A(_0941_),
    .B(_0964_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4143_ (.Y(_0969_),
    .A(_0963_),
    .B(_0968_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4144_ (.A2(_0967_),
    .A1(_0945_),
    .B1(_0969_),
    .X(_0970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4145_ (.A(_0959_),
    .B(_0961_),
    .X(_0971_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4146_ (.A2(_0955_),
    .A1(_0947_),
    .B1(_0954_),
    .X(_0972_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4147_ (.B1(_0952_),
    .VDD(VPWR),
    .Y(_0973_),
    .VSS(VGND),
    .A1(_0924_),
    .A2(_0950_));
 sg13g2_nand2_1 _4148_ (.Y(_0974_),
    .A(net990),
    .B(\DP_2.matrix[44] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4149_ (.Y(_0975_),
    .A(net926),
    .B(net1035),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4150_ (.Y(_0976_),
    .A(net928),
    .B(net1036),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4151_ (.B(_0976_),
    .A(_0949_),
    .X(_0977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4152_ (.Y(_0978_),
    .B(_0977_),
    .A_N(_0974_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4153_ (.Y(_0979_),
    .A(_0974_),
    .B(_0977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4154_ (.Y(_0980_),
    .A(_0973_),
    .B(_0979_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4155_ (.B(_0979_),
    .A(_0973_),
    .X(_0981_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4156_ (.Y(_0982_),
    .A(_0957_),
    .B(_0981_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4157_ (.A(_0982_),
    .B_N(_0972_),
    .Y(_0983_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4158_ (.B(_0982_),
    .A(_0972_),
    .X(_0984_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4159_ (.A(_0971_),
    .B(_0984_),
    .Y(_0985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4160_ (.B(_0984_),
    .A(_0971_),
    .X(_0986_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4161_ (.B(_0986_),
    .A(_0970_),
    .X(_0121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4162_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0970_),
    .A2(_0986_),
    .Y(_0987_),
    .B1(_0985_));
 sg13g2_a21oi_1 _4163_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0957_),
    .A2(_0981_),
    .Y(_0988_),
    .B1(_0983_));
 sg13g2_o21ai_1 _4164_ (.B1(_0978_),
    .VDD(VPWR),
    .Y(_0989_),
    .VSS(VGND),
    .A1(_0949_),
    .A2(_0976_));
 sg13g2_nand2_1 _4165_ (.Y(_0990_),
    .A(net988),
    .B(net1031),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4166_ (.Y(_0991_),
    .A(_0975_),
    .B(_0990_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4167_ (.Y(_0992_),
    .A(_0989_),
    .B(_0991_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4168_ (.Y(_0993_),
    .A(_0980_),
    .B(_0992_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4169_ (.Y(_0994_),
    .A(_0988_),
    .B(_0993_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4170_ (.Y(_0122_),
    .A(_0987_),
    .B(_0994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4171_ (.A(net886),
    .B(net831),
    .X(_0079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _4172_ (.X(_0995_),
    .A(net885),
    .B(net825),
    .C(_0079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4173_ (.Y(_0996_),
    .B1(net825),
    .B2(net886),
    .A2(net885),
    .A1(net831),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4174_ (.A(_0995_),
    .B(net401),
    .Y(_0080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4175_ (.Y(_0997_),
    .A(net886),
    .B(net823),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4176_ (.A(net831),
    .B(net885),
    .C(net825),
    .D(net882),
    .X(_0998_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4177_ (.Y(_0999_),
    .B1(net882),
    .B2(net831),
    .A2(net825),
    .A1(net885),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4178_ (.A(_0997_),
    .B(_0998_),
    .C(_0999_),
    .Y(_1000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4179_ (.B1(_0997_),
    .VDD(VPWR),
    .Y(_1001_),
    .VSS(VGND),
    .A1(_0998_),
    .A2(_0999_));
 sg13g2_nor2b_1 _4180_ (.A(_1000_),
    .B_N(_1001_),
    .Y(_1002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4181_ (.Y(_1003_),
    .A(_0995_),
    .B(_1002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4182_ (.B(_1002_),
    .A(_0995_),
    .X(_0081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4183_ (.Y(_1004_),
    .A(net886),
    .B(net822),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4184_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1005_),
    .B(_1000_),
    .A(_0998_));
 sg13g2_nand2_1 _4185_ (.Y(_1006_),
    .A(net885),
    .B(net823),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4186_ (.A(net831),
    .B(net825),
    .C(net882),
    .D(net880),
    .X(_1007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4187_ (.B(net825),
    .C(net882),
    .A(net831),
    .Y(_1008_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net880));
 sg13g2_a22oi_1 _4188_ (.Y(_1009_),
    .B1(net880),
    .B2(net831),
    .A2(net882),
    .A1(net825),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4189_ (.A(_1006_),
    .B(_1007_),
    .C(_1009_),
    .Y(_1010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4190_ (.B1(_1006_),
    .VDD(VPWR),
    .Y(_1011_),
    .VSS(VGND),
    .A1(_1007_),
    .A2(_1009_));
 sg13g2_nor2b_1 _4191_ (.A(_1010_),
    .B_N(_1011_),
    .Y(_1012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4192_ (.Y(_1013_),
    .A(_1005_),
    .B(_1012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4193_ (.Y(_1014_),
    .A(_1005_),
    .B(_1012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4194_ (.B(_1014_),
    .A(_1004_),
    .X(_1015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4195_ (.Y(_1016_),
    .B(_1015_),
    .A_N(_1003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4196_ (.Y(_0082_),
    .A(_1003_),
    .B(_1015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4197_ (.Y(_1017_),
    .B1(net820),
    .B2(net887),
    .A2(net822),
    .A1(net884),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4198_ (.Y(_1018_),
    .A(net884),
    .B(net819),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4199_ (.A(net887),
    .B(net884),
    .C(net822),
    .D(net820),
    .X(_1019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4200_ (.A(_1017_),
    .B(_1019_),
    .Y(_1020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4201_ (.VDD(VPWR),
    .Y(_1021_),
    .A(_1020_),
    .VSS(VGND));
 sg13g2_o21ai_1 _4202_ (.B1(_1008_),
    .VDD(VPWR),
    .Y(_1022_),
    .VSS(VGND),
    .A1(_1006_),
    .A2(_1009_));
 sg13g2_nand2_1 _4203_ (.Y(_1023_),
    .A(net882),
    .B(net823),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4204_ (.A(net830),
    .B(net828),
    .C(net880),
    .D(net878),
    .X(_1024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4205_ (.B(net827),
    .C(net880),
    .A(net830),
    .Y(_1025_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net878));
 sg13g2_a22oi_1 _4206_ (.Y(_1026_),
    .B1(net878),
    .B2(net830),
    .A2(net880),
    .A1(net827),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4207_ (.A(_1023_),
    .B(_1024_),
    .C(_1026_),
    .X(_1027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4208_ (.B1(_1023_),
    .VDD(VPWR),
    .Y(_1028_),
    .VSS(VGND),
    .A1(_1024_),
    .A2(_1026_));
 sg13g2_nand3_1 _4209_ (.B(_1027_),
    .C(_1028_),
    .A(_1022_),
    .Y(_1029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4210_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1027_),
    .A2(_1028_),
    .Y(_1030_),
    .B1(_1022_));
 sg13g2_a21o_1 _4211_ (.A2(_1028_),
    .A1(_1027_),
    .B1(_1022_),
    .X(_1031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4212_ (.Y(_1032_),
    .A(_1029_),
    .B(_1031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4213_ (.Y(_1033_),
    .A(_1021_),
    .B(_1032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4214_ (.B1(_1013_),
    .VDD(VPWR),
    .Y(_1034_),
    .VSS(VGND),
    .A1(_1004_),
    .A2(_1014_));
 sg13g2_nor2b_2 _4215_ (.A(_1033_),
    .B_N(_1034_),
    .Y(_1035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4216_ (.B(_1034_),
    .A(_1033_),
    .X(_1036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4217_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1037_),
    .B(_1036_),
    .A(_1016_));
 sg13g2_xor2_1 _4218_ (.B(_1036_),
    .A(_1016_),
    .X(_0083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4219_ (.B1(_1029_),
    .VDD(VPWR),
    .Y(_1038_),
    .VSS(VGND),
    .A1(_1021_),
    .A2(_1030_));
 sg13g2_nand2_1 _4220_ (.Y(_1039_),
    .A(net886),
    .B(net818),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4221_ (.Y(_1040_),
    .A(net883),
    .B(net819),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4222_ (.Y(_1041_),
    .A(net883),
    .B(net821),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4223_ (.B(_1041_),
    .A(_1018_),
    .X(_1042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4224_ (.Y(_1043_),
    .B(_1042_),
    .A_N(_1039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4225_ (.B(_1042_),
    .A(_1039_),
    .X(_1044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4226_ (.B1(_1025_),
    .VDD(VPWR),
    .Y(_1045_),
    .VSS(VGND),
    .A1(_1023_),
    .A2(_1026_));
 sg13g2_nand2_1 _4227_ (.Y(_1046_),
    .A(net824),
    .B(net881),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4228_ (.A(net830),
    .B(net827),
    .C(net878),
    .D(net876),
    .X(_1047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4229_ (.B(net827),
    .C(net878),
    .A(net830),
    .Y(_1048_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net876));
 sg13g2_a22oi_1 _4230_ (.Y(_1049_),
    .B1(net876),
    .B2(net830),
    .A2(net878),
    .A1(net827),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4231_ (.A(_1046_),
    .B(_1047_),
    .C(_1049_),
    .X(_1050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4232_ (.B1(_1046_),
    .VDD(VPWR),
    .Y(_1051_),
    .VSS(VGND),
    .A1(_1047_),
    .A2(_1049_));
 sg13g2_and3_1 _4233_ (.X(_1052_),
    .A(_1045_),
    .B(_1050_),
    .C(_1051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4234_ (.B(_1050_),
    .C(_1051_),
    .A(_1045_),
    .Y(_1053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4235_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1050_),
    .A2(_1051_),
    .Y(_1054_),
    .B1(_1045_));
 sg13g2_or3_1 _4236_ (.A(_1044_),
    .B(_1052_),
    .C(_1054_),
    .X(_1055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4237_ (.B1(_1044_),
    .VDD(VPWR),
    .Y(_1056_),
    .VSS(VGND),
    .A1(_1052_),
    .A2(_1054_));
 sg13g2_nand3_1 _4238_ (.B(_1055_),
    .C(_1056_),
    .A(_1038_),
    .Y(_1057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4239_ (.A2(_1056_),
    .A1(_1055_),
    .B1(_1038_),
    .X(_1058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4240_ (.B(_1057_),
    .C(_1058_),
    .A(_1019_),
    .Y(_1059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4241_ (.A2(_1058_),
    .A1(_1057_),
    .B1(_1019_),
    .X(_1060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4242_ (.A(_1059_),
    .B(_1060_),
    .X(_1061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4243_ (.B(_1059_),
    .C(_1060_),
    .A(_1035_),
    .Y(_1062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4244_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1059_),
    .A2(_1060_),
    .Y(_1063_),
    .B1(_1035_));
 sg13g2_xor2_1 _4245_ (.B(_1061_),
    .A(_1035_),
    .X(_1064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4246_ (.Y(_0127_),
    .A(_1037_),
    .B(_1064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4247_ (.Y(_1065_),
    .A(_1057_),
    .B(_1059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4248_ (.B1(_1043_),
    .VDD(VPWR),
    .Y(_1066_),
    .VSS(VGND),
    .A1(_1018_),
    .A2(_1041_));
 sg13g2_nand2_1 _4249_ (.Y(_1067_),
    .A(net887),
    .B(net817),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4250_ (.Y(_1068_),
    .B(_1066_),
    .A_N(_1067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4251_ (.B(_1067_),
    .A(_1066_),
    .X(_1069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4252_ (.B1(_1053_),
    .VDD(VPWR),
    .Y(_1070_),
    .VSS(VGND),
    .A1(_1044_),
    .A2(_1054_));
 sg13g2_nand2_1 _4253_ (.Y(_1071_),
    .A(net884),
    .B(net818),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4254_ (.Y(_1072_),
    .A(net881),
    .B(net820),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4255_ (.Y(_1073_),
    .A(net881),
    .B(net822),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4256_ (.B(_1073_),
    .A(_1040_),
    .X(_1074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4257_ (.Y(_1075_),
    .B(_1074_),
    .A_N(_1071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4258_ (.Y(_1076_),
    .A(_1071_),
    .B(_1074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4259_ (.B1(_1048_),
    .VDD(VPWR),
    .Y(_1077_),
    .VSS(VGND),
    .A1(_1046_),
    .A2(_1049_));
 sg13g2_nand2_1 _4260_ (.Y(_1078_),
    .A(net824),
    .B(net879),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4261_ (.A(net829),
    .B(net827),
    .C(net876),
    .D(net875),
    .X(_1079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4262_ (.B(net827),
    .C(net876),
    .A(net829),
    .Y(_1080_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net875));
 sg13g2_a22oi_1 _4263_ (.Y(_1081_),
    .B1(net875),
    .B2(net829),
    .A2(net876),
    .A1(net827),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4264_ (.A(_1078_),
    .B(_1079_),
    .C(_1081_),
    .X(_1082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4265_ (.B1(_1078_),
    .VDD(VPWR),
    .Y(_1083_),
    .VSS(VGND),
    .A1(_1079_),
    .A2(_1081_));
 sg13g2_and3_1 _4266_ (.X(_1084_),
    .A(_1077_),
    .B(_1082_),
    .C(_1083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4267_ (.B(_1082_),
    .C(_1083_),
    .A(_1077_),
    .Y(_1085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4268_ (.A2(_1083_),
    .A1(_1082_),
    .B1(_1077_),
    .X(_1086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4269_ (.B(_1085_),
    .C(_1086_),
    .A(_1076_),
    .Y(_1087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4270_ (.A2(_1086_),
    .A1(_1085_),
    .B1(_1076_),
    .X(_1088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4271_ (.B(_1087_),
    .C(_1088_),
    .A(_1070_),
    .Y(_1089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4272_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1087_),
    .A2(_1088_),
    .Y(_1090_),
    .B1(_1070_));
 sg13g2_a21o_1 _4273_ (.A2(_1088_),
    .A1(_1087_),
    .B1(_1070_),
    .X(_1091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4274_ (.Y(_1092_),
    .A(_1089_),
    .B(_1091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4275_ (.Y(_1093_),
    .A(_1069_),
    .B(_1092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4276_ (.A(_1093_),
    .B_N(_1065_),
    .Y(_1094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4277_ (.Y(_1095_),
    .A(_1065_),
    .B(_1093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4278_ (.B1(_1062_),
    .VDD(VPWR),
    .Y(_1096_),
    .VSS(VGND),
    .A1(_1037_),
    .A2(_1063_));
 sg13g2_xor2_1 _4279_ (.B(_1096_),
    .A(_1095_),
    .X(_0134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4280_ (.B1(_1089_),
    .VDD(VPWR),
    .Y(_1097_),
    .VSS(VGND),
    .A1(_1069_),
    .A2(_1090_));
 sg13g2_o21ai_1 _4281_ (.B1(_1075_),
    .VDD(VPWR),
    .Y(_1098_),
    .VSS(VGND),
    .A1(_1040_),
    .A2(_1073_));
 sg13g2_a22oi_1 _4282_ (.Y(_1099_),
    .B1(net814),
    .B2(net886),
    .A2(net816),
    .A1(net884),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4283_ (.B(\DP_3.matrix[37] ),
    .C(net816),
    .A(net887),
    .Y(_1100_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net814));
 sg13g2_nor2b_1 _4284_ (.A(_1099_),
    .B_N(_1100_),
    .Y(_1101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4285_ (.Y(_1102_),
    .A(_1098_),
    .B(_1101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4286_ (.Y(_1103_),
    .A(_1098_),
    .B(_1101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4287_ (.A2(_1086_),
    .A1(_1076_),
    .B1(_1084_),
    .X(_1104_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4288_ (.Y(_1105_),
    .A(net883),
    .B(\DP_4.matrix[41] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4289_ (.Y(_1106_),
    .A(net879),
    .B(net820),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4290_ (.Y(_1107_),
    .A(net821),
    .B(net879),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4291_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1108_),
    .B(_1106_),
    .A(_1073_));
 sg13g2_and2_1 _4292_ (.A(_1072_),
    .B(_1107_),
    .X(_1109_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4293_ (.Y(_1110_),
    .A(_1072_),
    .B(_1107_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4294_ (.Y(_1111_),
    .A(_1105_),
    .B(_1110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4295_ (.B1(_1080_),
    .VDD(VPWR),
    .Y(_1112_),
    .VSS(VGND),
    .A1(_1078_),
    .A2(_1081_));
 sg13g2_nand2_1 _4296_ (.Y(_1113_),
    .A(net824),
    .B(net877),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4297_ (.A(\DP_4.matrix[36] ),
    .B(net826),
    .C(net874),
    .D(net872),
    .X(_1114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4298_ (.B(net826),
    .C(net874),
    .A(net830),
    .Y(_1115_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net871));
 sg13g2_a22oi_1 _4299_ (.Y(_1116_),
    .B1(net871),
    .B2(net829),
    .A2(net874),
    .A1(net826),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4300_ (.A(_1113_),
    .B(_1114_),
    .C(_1116_),
    .X(_1117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4301_ (.B1(_1113_),
    .VDD(VPWR),
    .Y(_1118_),
    .VSS(VGND),
    .A1(_1114_),
    .A2(_1116_));
 sg13g2_and3_1 _4302_ (.X(_1119_),
    .A(_1112_),
    .B(_1117_),
    .C(_1118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4303_ (.B(_1117_),
    .C(_1118_),
    .A(_1112_),
    .Y(_1120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4304_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1117_),
    .A2(_1118_),
    .Y(_1121_),
    .B1(_1112_));
 sg13g2_or3_1 _4305_ (.A(_1111_),
    .B(_1119_),
    .C(_1121_),
    .X(_1122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4306_ (.B1(_1111_),
    .VDD(VPWR),
    .Y(_1123_),
    .VSS(VGND),
    .A1(_1119_),
    .A2(_1121_));
 sg13g2_and3_1 _4307_ (.X(_1124_),
    .A(_1104_),
    .B(_1122_),
    .C(_1123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4308_ (.B(_1122_),
    .C(_1123_),
    .A(_1104_),
    .Y(_1125_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4309_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1122_),
    .A2(_1123_),
    .Y(_1126_),
    .B1(_1104_));
 sg13g2_or3_1 _4310_ (.A(_1103_),
    .B(_1124_),
    .C(_1126_),
    .X(_1127_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4311_ (.B1(_1103_),
    .VDD(VPWR),
    .Y(_1128_),
    .VSS(VGND),
    .A1(_1124_),
    .A2(_1126_));
 sg13g2_nand3_1 _4312_ (.B(_1127_),
    .C(_1128_),
    .A(_1097_),
    .Y(_1129_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4313_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1127_),
    .A2(_1128_),
    .Y(_1130_),
    .B1(_1097_));
 sg13g2_a21o_1 _4314_ (.A2(_1128_),
    .A1(_1127_),
    .B1(_1097_),
    .X(_1131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4315_ (.Y(_1132_),
    .A(_1129_),
    .B(_1131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4316_ (.B(_1132_),
    .A(_1068_),
    .X(_1133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _4317_ (.A2(_1096_),
    .A1(_1095_),
    .B1(_1094_),
    .X(_1134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4318_ (.Y(_1135_),
    .A(_1133_),
    .B(_1134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4319_ (.B(_1134_),
    .A(_1133_),
    .X(_0135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4320_ (.B1(_1125_),
    .VDD(VPWR),
    .Y(_1136_),
    .VSS(VGND),
    .A1(_1103_),
    .A2(_1126_));
 sg13g2_o21ai_1 _4321_ (.B1(_1108_),
    .VDD(VPWR),
    .Y(_1137_),
    .VSS(VGND),
    .A1(_1105_),
    .A2(_1109_));
 sg13g2_nand2_1 _4322_ (.Y(_1138_),
    .A(net887),
    .B(net1022),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4323_ (.Y(_1139_),
    .A(net883),
    .B(net814),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4324_ (.A(net884),
    .B(net883),
    .C(net817),
    .D(net814),
    .X(_1140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4325_ (.Y(_1141_),
    .B1(net814),
    .B2(net884),
    .A2(net817),
    .A1(net883),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4326_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1142_),
    .B(_1141_),
    .A(_1140_));
 sg13g2_nor2_1 _4327_ (.A(_1138_),
    .B(_1142_),
    .Y(_1143_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4328_ (.B(_1142_),
    .A(_1138_),
    .X(_1144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4329_ (.Y(_1145_),
    .A(_1137_),
    .B(_1144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4330_ (.Y(_1146_),
    .A(_1137_),
    .B(_1144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4331_ (.Y(_1147_),
    .A(_1100_),
    .B(_1146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4332_ (.B1(_1120_),
    .VDD(VPWR),
    .Y(_1148_),
    .VSS(VGND),
    .A1(_1111_),
    .A2(_1121_));
 sg13g2_nand2_1 _4333_ (.Y(_1149_),
    .A(net881),
    .B(\DP_4.matrix[41] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4334_ (.Y(_1150_),
    .A(net819),
    .B(net877),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4335_ (.Y(_1151_),
    .A(net821),
    .B(net877),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4336_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1152_),
    .B(_1150_),
    .A(_1107_));
 sg13g2_xnor2_1 _4337_ (.Y(_1153_),
    .A(_1106_),
    .B(_1151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4338_ (.Y(_1154_),
    .A(_1149_),
    .B(_1153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4339_ (.B1(_1115_),
    .VDD(VPWR),
    .Y(_1155_),
    .VSS(VGND),
    .A1(_1113_),
    .A2(_1116_));
 sg13g2_nand2_1 _4340_ (.Y(_1156_),
    .A(net823),
    .B(net873),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4341_ (.A(net829),
    .B(net826),
    .C(net871),
    .D(net1026),
    .X(_1157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4342_ (.B(net826),
    .C(net871),
    .A(net829),
    .Y(_1158_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net1026));
 sg13g2_a22oi_1 _4343_ (.Y(_1159_),
    .B1(net1026),
    .B2(net829),
    .A2(net871),
    .A1(net828),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4344_ (.A(_1156_),
    .B(_1157_),
    .C(_1159_),
    .X(_1160_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4345_ (.B1(_1156_),
    .VDD(VPWR),
    .Y(_1161_),
    .VSS(VGND),
    .A1(_1157_),
    .A2(_1159_));
 sg13g2_and3_1 _4346_ (.X(_1162_),
    .A(_1155_),
    .B(_1160_),
    .C(_1161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4347_ (.B(_1160_),
    .C(_1161_),
    .A(_1155_),
    .Y(_1163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4348_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1160_),
    .A2(_1161_),
    .Y(_1164_),
    .B1(_1155_));
 sg13g2_or3_1 _4349_ (.A(_1154_),
    .B(_1162_),
    .C(_1164_),
    .X(_1165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4350_ (.B1(_1154_),
    .VDD(VPWR),
    .Y(_1166_),
    .VSS(VGND),
    .A1(_1162_),
    .A2(_1164_));
 sg13g2_and3_1 _4351_ (.X(_1167_),
    .A(_1148_),
    .B(_1165_),
    .C(_1166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4352_ (.B(_1165_),
    .C(_1166_),
    .A(_1148_),
    .Y(_1168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4353_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1165_),
    .A2(_1166_),
    .Y(_1169_),
    .B1(_1148_));
 sg13g2_or3_1 _4354_ (.A(_1147_),
    .B(_1167_),
    .C(_1169_),
    .X(_1170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4355_ (.B1(_1147_),
    .VDD(VPWR),
    .Y(_1171_),
    .VSS(VGND),
    .A1(_1167_),
    .A2(_1169_));
 sg13g2_and3_1 _4356_ (.X(_1172_),
    .A(_1136_),
    .B(_1170_),
    .C(_1171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4357_ (.B(_1170_),
    .C(_1171_),
    .A(_1136_),
    .Y(_1173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4358_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1170_),
    .A2(_1171_),
    .Y(_1174_),
    .B1(_1136_));
 sg13g2_or3_1 _4359_ (.A(_1102_),
    .B(_1172_),
    .C(_1174_),
    .X(_1175_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4360_ (.B1(_1102_),
    .VDD(VPWR),
    .Y(_1176_),
    .VSS(VGND),
    .A1(_1172_),
    .A2(_1174_));
 sg13g2_o21ai_1 _4361_ (.B1(_1129_),
    .VDD(VPWR),
    .Y(_1177_),
    .VSS(VGND),
    .A1(_1068_),
    .A2(_1130_));
 sg13g2_nand3_1 _4362_ (.B(_1176_),
    .C(_1177_),
    .A(_1175_),
    .Y(_1178_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4363_ (.A2(_1176_),
    .A1(_1175_),
    .B1(_1177_),
    .X(_1179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4364_ (.Y(_1180_),
    .A(_1178_),
    .B(_1179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4365_ (.A(_1133_),
    .B(_1134_),
    .C(_1178_),
    .D(_1179_),
    .X(_1181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4366_ (.B(_1180_),
    .A(_1135_),
    .X(_0136_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4367_ (.B1(_1178_),
    .VDD(VPWR),
    .Y(_1182_),
    .VSS(VGND),
    .A1(_1135_),
    .A2(_1180_));
 sg13g2_o21ai_1 _4368_ (.B1(_1173_),
    .VDD(VPWR),
    .Y(_1183_),
    .VSS(VGND),
    .A1(_1102_),
    .A2(_1174_));
 sg13g2_o21ai_1 _4369_ (.B1(_1145_),
    .VDD(VPWR),
    .Y(_1184_),
    .VSS(VGND),
    .A1(_1100_),
    .A2(_1146_));
 sg13g2_o21ai_1 _4370_ (.B1(_1168_),
    .VDD(VPWR),
    .Y(_1185_),
    .VSS(VGND),
    .A1(_1147_),
    .A2(_1169_));
 sg13g2_nor2_1 _4371_ (.A(_1140_),
    .B(_1143_),
    .Y(_1186_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4372_ (.B1(_1152_),
    .VDD(VPWR),
    .Y(_1187_),
    .VSS(VGND),
    .A1(_1149_),
    .A2(_1153_));
 sg13g2_nand2_1 _4373_ (.Y(_1188_),
    .A(net885),
    .B(net1022),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4374_ (.Y(_1189_),
    .A(net881),
    .B(net815),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4375_ (.Y(_1190_),
    .A(net881),
    .B(net817),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4376_ (.B(_1190_),
    .A(_1139_),
    .X(_1191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4377_ (.Y(_1192_),
    .B(_1191_),
    .A_N(_1188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4378_ (.Y(_1193_),
    .A(_1188_),
    .B(_1191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4379_ (.Y(_1194_),
    .A(_1187_),
    .B(_1193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4380_ (.A(_1186_),
    .B(_1194_),
    .Y(_1195_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4381_ (.Y(_1196_),
    .A(_1186_),
    .B(_1194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4382_ (.B1(_1163_),
    .VDD(VPWR),
    .Y(_1197_),
    .VSS(VGND),
    .A1(_1154_),
    .A2(_1164_));
 sg13g2_nand2_1 _4383_ (.Y(_1198_),
    .A(net879),
    .B(\DP_4.matrix[41] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4384_ (.Y(_1199_),
    .A(net821),
    .B(net873),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4385_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1200_),
    .B(_1199_),
    .A(_1150_));
 sg13g2_and2_1 _4386_ (.A(_1150_),
    .B(_1199_),
    .X(_1201_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4387_ (.Y(_1202_),
    .A(_1150_),
    .B(_1199_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4388_ (.Y(_1203_),
    .A(_1198_),
    .B(_1202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4389_ (.B1(_1158_),
    .VDD(VPWR),
    .Y(_1204_),
    .VSS(VGND),
    .A1(_1156_),
    .A2(_1159_));
 sg13g2_nand2_1 _4390_ (.Y(_1205_),
    .A(net823),
    .B(net1027),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4391_ (.A(net826),
    .B(net824),
    .C(net870),
    .D(net1026),
    .X(_1206_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4392_ (.Y(_1207_),
    .B1(net1027),
    .B2(net826),
    .A2(net870),
    .A1(net823),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4393_ (.A(_1206_),
    .B(_1207_),
    .Y(_1208_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4394_ (.Y(_1209_),
    .A(_1204_),
    .B(_1208_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4395_ (.Y(_1210_),
    .A(_1204_),
    .B(_1208_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4396_ (.B(_1210_),
    .A(_1203_),
    .X(_1211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4397_ (.Y(_1212_),
    .A(_1197_),
    .B(_1211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4398_ (.Y(_1213_),
    .A(_1197_),
    .B(_1211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4399_ (.B(_1213_),
    .A(_1196_),
    .X(_1214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4400_ (.Y(_1215_),
    .A(_1185_),
    .B(_1214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4401_ (.Y(_1216_),
    .A(_1185_),
    .B(_1214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4402_ (.Y(_1217_),
    .B(_1184_),
    .A_N(_1216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4403_ (.Y(_1218_),
    .A(_1184_),
    .B(_1216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4404_ (.A(_1183_),
    .B(_1218_),
    .Y(_1219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4405_ (.Y(_1220_),
    .A(_1183_),
    .B(_1218_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _4406_ (.A(_1219_),
    .B_N(_1220_),
    .Y(_1221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4407_ (.B(_1221_),
    .A(_1182_),
    .X(_0137_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4408_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1187_),
    .A2(_1193_),
    .Y(_1222_),
    .B1(_1195_));
 sg13g2_o21ai_1 _4409_ (.B1(_1212_),
    .VDD(VPWR),
    .Y(_1223_),
    .VSS(VGND),
    .A1(_1196_),
    .A2(_1213_));
 sg13g2_o21ai_1 _4410_ (.B1(_1192_),
    .VDD(VPWR),
    .Y(_1224_),
    .VSS(VGND),
    .A1(_1139_),
    .A2(_1190_));
 sg13g2_o21ai_1 _4411_ (.B1(_1200_),
    .VDD(VPWR),
    .Y(_1225_),
    .VSS(VGND),
    .A1(_1198_),
    .A2(_1201_));
 sg13g2_nand2_1 _4412_ (.Y(_1226_),
    .A(net883),
    .B(net1022),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4413_ (.Y(_1227_),
    .A(net879),
    .B(net815),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4414_ (.Y(_1228_),
    .A(net879),
    .B(net816),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4415_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1229_),
    .B(_1227_),
    .A(_1190_));
 sg13g2_xnor2_1 _4416_ (.Y(_1230_),
    .A(_1189_),
    .B(_1228_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4417_ (.B(_1230_),
    .A(_1226_),
    .X(_1231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4418_ (.Y(_1232_),
    .A(_1225_),
    .B(_1231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4419_ (.A(_1232_),
    .B_N(_1224_),
    .Y(_1233_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4420_ (.B(_1232_),
    .A(_1224_),
    .X(_1234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4421_ (.B1(_1209_),
    .VDD(VPWR),
    .Y(_1235_),
    .VSS(VGND),
    .A1(_1203_),
    .A2(_1210_));
 sg13g2_a21oi_1 _4422_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net828),
    .A2(net870),
    .Y(_1236_),
    .B1(_1205_));
 sg13g2_nand2_1 _4423_ (.Y(_1237_),
    .A(net877),
    .B(net818),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4424_ (.Y(_1238_),
    .A(net819),
    .B(net870),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4425_ (.A(net821),
    .B(net819),
    .C(net873),
    .D(net870),
    .X(_1239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4426_ (.Y(_1240_),
    .B1(net870),
    .B2(net821),
    .A2(net874),
    .A1(net819),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4427_ (.A(_1237_),
    .B(_1239_),
    .C(_1240_),
    .Y(_1241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4428_ (.B1(_1237_),
    .VDD(VPWR),
    .Y(_1242_),
    .VSS(VGND),
    .A1(_1239_),
    .A2(_1240_));
 sg13g2_nor2b_1 _4429_ (.A(_1241_),
    .B_N(_1242_),
    .Y(_1243_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4430_ (.Y(_1244_),
    .A(_1236_),
    .B(_1243_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4431_ (.Y(_1245_),
    .B(_1235_),
    .A_N(_1244_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4432_ (.B(_1244_),
    .A(_1235_),
    .X(_1246_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4433_ (.B(_1246_),
    .A(_1234_),
    .X(_1247_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4434_ (.Y(_1248_),
    .A(_1223_),
    .B(_1247_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4435_ (.B(_1247_),
    .A(_1223_),
    .X(_1249_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4436_ (.Y(_1250_),
    .B(_1249_),
    .A_N(_1222_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4437_ (.B(_1249_),
    .A(_1222_),
    .X(_1251_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4438_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1215_),
    .A2(_1217_),
    .Y(_1252_),
    .B1(_1251_));
 sg13g2_nand3_1 _4439_ (.B(_1217_),
    .C(_1251_),
    .A(_1215_),
    .Y(_1253_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4440_ (.Y(_1254_),
    .B(_1253_),
    .A_N(_1252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4441_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1178_),
    .A2(_1220_),
    .Y(_1255_),
    .B1(_1219_));
 sg13g2_a21oi_2 _4442_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_1255_),
    .Y(_1256_),
    .A2(_1221_),
    .A1(_1181_));
 sg13g2_nor2_1 _4443_ (.A(_1254_),
    .B(_1256_),
    .Y(_1257_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4444_ (.B(_1256_),
    .A(_1254_),
    .X(_0128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4445_ (.A2(_1231_),
    .A1(_1225_),
    .B1(_1233_),
    .X(_1258_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4446_ (.B1(_1245_),
    .VDD(VPWR),
    .Y(_1259_),
    .VSS(VGND),
    .A1(_1234_),
    .A2(_1246_));
 sg13g2_a21o_1 _4447_ (.A2(_1243_),
    .A1(_1236_),
    .B1(_1206_),
    .X(_1260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4448_ (.Y(_1261_),
    .A(net818),
    .B(net873),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4449_ (.Y(_1262_),
    .A(net821),
    .B(net1026),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4450_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1263_),
    .B(_1262_),
    .A(_1238_));
 sg13g2_xnor2_1 _4451_ (.Y(_1264_),
    .A(_1238_),
    .B(_1262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4452_ (.B(_1264_),
    .A(_1261_),
    .X(_1265_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4453_ (.Y(_1266_),
    .A(_1260_),
    .B(_1265_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4454_ (.B1(_1229_),
    .VDD(VPWR),
    .Y(_1267_),
    .VSS(VGND),
    .A1(_1226_),
    .A2(_1230_));
 sg13g2_or2_1 _4455_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1268_),
    .B(_1241_),
    .A(_1239_));
 sg13g2_nand2_1 _4456_ (.Y(_1269_),
    .A(net881),
    .B(net1022),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4457_ (.Y(_1270_),
    .A(net877),
    .B(net815),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4458_ (.Y(_1271_),
    .A(net877),
    .B(net816),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4459_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1272_),
    .B(_1270_),
    .A(_1228_));
 sg13g2_xnor2_1 _4460_ (.Y(_1273_),
    .A(_1227_),
    .B(_1271_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4461_ (.B(_1273_),
    .A(_1269_),
    .X(_1274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4462_ (.Y(_1275_),
    .A(_1268_),
    .B(_1274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4463_ (.A(_1275_),
    .B_N(_1267_),
    .Y(_1276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4464_ (.B(_1275_),
    .A(_1267_),
    .X(_1277_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4465_ (.A(_1266_),
    .B(_1277_),
    .Y(_1278_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4466_ (.B(_1277_),
    .A(_1266_),
    .X(_1279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4467_ (.Y(_1280_),
    .A(_1259_),
    .B(_1279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4468_ (.A(_1280_),
    .B_N(_1258_),
    .Y(_1281_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4469_ (.B(_1280_),
    .A(_1258_),
    .X(_1282_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4470_ (.B(_1250_),
    .C(_1282_),
    .A(_1248_),
    .Y(_1283_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4471_ (.VDD(VPWR),
    .Y(_1284_),
    .A(_1283_),
    .VSS(VGND));
 sg13g2_a21oi_1 _4472_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1248_),
    .A2(_1250_),
    .Y(_1285_),
    .B1(_1282_));
 sg13g2_nor2_1 _4473_ (.A(_1284_),
    .B(_1285_),
    .Y(_1286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4474_ (.A(_1252_),
    .B(_1257_),
    .Y(_1287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4475_ (.Y(_0129_),
    .A(_1286_),
    .B(_1287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4476_ (.A2(_1274_),
    .A1(_1268_),
    .B1(_1276_),
    .X(_1288_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4477_ (.Y(_1289_),
    .B1(net1026),
    .B2(net819),
    .A2(net871),
    .A1(net818),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4478_ (.Y(_1290_),
    .A(net818),
    .B(net1027),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4479_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1291_),
    .B(_1290_),
    .A(_1238_));
 sg13g2_nand2b_1 _4480_ (.Y(_1292_),
    .B(_1291_),
    .A_N(_1289_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4481_ (.B1(_1272_),
    .VDD(VPWR),
    .Y(_1293_),
    .VSS(VGND),
    .A1(_1269_),
    .A2(_1273_));
 sg13g2_o21ai_1 _4482_ (.B1(_1263_),
    .VDD(VPWR),
    .Y(_1294_),
    .VSS(VGND),
    .A1(_1261_),
    .A2(_1264_));
 sg13g2_nand2_1 _4483_ (.Y(_1295_),
    .A(net879),
    .B(net1022),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4484_ (.Y(_1296_),
    .A(net873),
    .B(net814),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4485_ (.Y(_1297_),
    .A(net873),
    .B(net816),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4486_ (.B(_1297_),
    .A(_1270_),
    .X(_1298_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4487_ (.Y(_1299_),
    .B(_1298_),
    .A_N(_1295_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4488_ (.Y(_1300_),
    .A(_1295_),
    .B(_1298_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4489_ (.Y(_1301_),
    .A(_1294_),
    .B(_1300_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4490_ (.A(_1301_),
    .B_N(_1293_),
    .Y(_1302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4491_ (.B(_1301_),
    .A(_1293_),
    .X(_1303_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4492_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1304_),
    .B(_1303_),
    .A(_1292_));
 sg13g2_xor2_1 _4493_ (.B(_1303_),
    .A(_1292_),
    .X(_1305_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4494_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1260_),
    .A2(_1265_),
    .Y(_1306_),
    .B1(_1278_));
 sg13g2_nor2b_1 _4495_ (.A(_1306_),
    .B_N(_1305_),
    .Y(_1307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4496_ (.B(_1306_),
    .A(_1305_),
    .X(_1308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4497_ (.A(_1308_),
    .B_N(_1288_),
    .Y(_1309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4498_ (.B(_1308_),
    .A(_1288_),
    .X(_1310_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4499_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1259_),
    .A2(_1279_),
    .Y(_1311_),
    .B1(_1281_));
 sg13g2_nor2_1 _4500_ (.A(_1310_),
    .B(_1311_),
    .Y(_1312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4501_ (.B(_1311_),
    .A(_1310_),
    .X(_1313_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4502_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1252_),
    .A2(_1283_),
    .Y(_1314_),
    .B1(_1285_));
 sg13g2_a21oi_1 _4503_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1253_),
    .A2(_1283_),
    .Y(_1315_),
    .B1(_1285_));
 sg13g2_a21oi_2 _4504_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_1315_),
    .Y(_1316_),
    .A2(_1314_),
    .A1(_1256_));
 sg13g2_xor2_1 _4505_ (.B(_1316_),
    .A(_1313_),
    .X(_0130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4506_ (.A2(_1300_),
    .A1(_1294_),
    .B1(_1302_),
    .X(_1317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4507_ (.B1(_1299_),
    .VDD(VPWR),
    .Y(_1318_),
    .VSS(VGND),
    .A1(_1270_),
    .A2(_1297_));
 sg13g2_nand2_1 _4508_ (.Y(_1319_),
    .A(net877),
    .B(net1022),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4509_ (.Y(_1320_),
    .A(net870),
    .B(net814),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4510_ (.Y(_1321_),
    .A(net816),
    .B(net871),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4511_ (.B(_1321_),
    .A(_1296_),
    .X(_1322_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4512_ (.Y(_1323_),
    .B(_1322_),
    .A_N(_1319_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4513_ (.Y(_1324_),
    .A(_1319_),
    .B(_1322_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4514_ (.A(_1291_),
    .B_N(_1324_),
    .Y(_1325_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4515_ (.Y(_1326_),
    .A(_1291_),
    .B(_1324_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4516_ (.Y(_1327_),
    .A(_1318_),
    .B(_1326_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4517_ (.A(_1290_),
    .B(_1327_),
    .Y(_1328_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4518_ (.B(_1327_),
    .A(_1290_),
    .X(_1329_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4519_ (.Y(_1330_),
    .B(_1329_),
    .A_N(_1304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4520_ (.Y(_1331_),
    .A(_1304_),
    .B(_1329_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4521_ (.Y(_1332_),
    .A(_1317_),
    .B(_1331_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4522_ (.B(_1331_),
    .A(_1317_),
    .X(_1333_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4523_ (.B1(_1333_),
    .VDD(VPWR),
    .Y(_1334_),
    .VSS(VGND),
    .A1(_1307_),
    .A2(_1309_));
 sg13g2_or3_1 _4524_ (.A(_1307_),
    .B(_1309_),
    .C(_1333_),
    .X(_1335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4525_ (.A(_1334_),
    .B(_1335_),
    .X(_1336_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4526_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1313_),
    .A2(_1316_),
    .Y(_1337_),
    .B1(_1312_));
 sg13g2_xnor2_1 _4527_ (.Y(_0131_),
    .A(_1336_),
    .B(_1337_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4528_ (.A(_1313_),
    .B(_1336_),
    .X(_1338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4529_ (.Y(_1339_),
    .A(_1312_),
    .B(_1335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4530_ (.Y(_1340_),
    .A(_1334_),
    .B(_1339_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4531_ (.A2(_1338_),
    .A1(_1316_),
    .B1(_1340_),
    .X(_1341_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4532_ (.A(_1330_),
    .B(_1332_),
    .X(_1342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4533_ (.A2(_1326_),
    .A1(_1318_),
    .B1(_1325_),
    .X(_1343_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4534_ (.Y(_1344_),
    .A(net873),
    .B(net1022),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4535_ (.Y(_1345_),
    .A(net814),
    .B(net1027),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4536_ (.Y(_1346_),
    .A(net816),
    .B(net1027),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4537_ (.B(_1346_),
    .A(_1320_),
    .X(_1347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4538_ (.Y(_1348_),
    .B(_1347_),
    .A_N(_1344_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4539_ (.Y(_1349_),
    .A(_1344_),
    .B(_1347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4540_ (.B1(_1323_),
    .VDD(VPWR),
    .Y(_1350_),
    .VSS(VGND),
    .A1(_1296_),
    .A2(_1321_));
 sg13g2_nand2_1 _4541_ (.Y(_1351_),
    .A(_1349_),
    .B(_1350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4542_ (.B(_1350_),
    .A(_1349_),
    .X(_1352_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4543_ (.Y(_1353_),
    .A(_1328_),
    .B(_1352_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4544_ (.A(_1353_),
    .B_N(_1343_),
    .Y(_1354_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4545_ (.B(_1353_),
    .A(_1343_),
    .X(_1355_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4546_ (.A(_1342_),
    .B(_1355_),
    .Y(_1356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4547_ (.B(_1355_),
    .A(_1342_),
    .X(_1357_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4548_ (.B(_1357_),
    .A(_1341_),
    .X(_0132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4549_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1341_),
    .A2(_1357_),
    .Y(_1358_),
    .B1(_1356_));
 sg13g2_a21oi_1 _4550_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1328_),
    .A2(_1352_),
    .Y(_1359_),
    .B1(_1354_));
 sg13g2_o21ai_1 _4551_ (.B1(_1348_),
    .VDD(VPWR),
    .Y(_1360_),
    .VSS(VGND),
    .A1(_1320_),
    .A2(_1346_));
 sg13g2_nand2_1 _4552_ (.Y(_1361_),
    .A(net870),
    .B(\DP_4.matrix[44] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4553_ (.Y(_1362_),
    .A(_1345_),
    .B(_1361_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4554_ (.Y(_1363_),
    .A(_1360_),
    .B(_1362_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4555_ (.Y(_1364_),
    .A(_1351_),
    .B(_1363_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4556_ (.Y(_1365_),
    .A(_1359_),
    .B(_1364_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4557_ (.Y(_0133_),
    .A(_1358_),
    .B(_1365_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4558_ (.A(net903),
    .B(net847),
    .X(_0084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _4559_ (.X(_1366_),
    .A(net901),
    .B(net843),
    .C(_0084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4560_ (.Y(_1367_),
    .B1(net843),
    .B2(net903),
    .A2(net901),
    .A1(net847),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4561_ (.A(_1366_),
    .B(_1367_),
    .Y(_0085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4562_ (.Y(_1368_),
    .A(net903),
    .B(net841),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4563_ (.A(net847),
    .B(net901),
    .C(net843),
    .D(net899),
    .X(_1369_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4564_ (.Y(_1370_),
    .B1(net899),
    .B2(net847),
    .A2(net843),
    .A1(net901),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4565_ (.A(_1368_),
    .B(_1369_),
    .C(_1370_),
    .Y(_1371_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4566_ (.B1(_1368_),
    .VDD(VPWR),
    .Y(_1372_),
    .VSS(VGND),
    .A1(_1369_),
    .A2(_1370_));
 sg13g2_nor2b_1 _4567_ (.A(_1371_),
    .B_N(_1372_),
    .Y(_1373_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4568_ (.Y(_1374_),
    .A(_1366_),
    .B(_1373_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4569_ (.B(_1373_),
    .A(_1366_),
    .X(_0086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4570_ (.Y(_1375_),
    .A(net903),
    .B(net839),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4571_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1376_),
    .B(_1371_),
    .A(_1369_));
 sg13g2_nand2_1 _4572_ (.Y(_1377_),
    .A(net901),
    .B(net841),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4573_ (.A(net847),
    .B(net843),
    .C(net899),
    .D(net897),
    .X(_1378_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4574_ (.B(net844),
    .C(net899),
    .A(net847),
    .Y(_1379_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net897));
 sg13g2_a22oi_1 _4575_ (.Y(_1380_),
    .B1(net897),
    .B2(net848),
    .A2(net899),
    .A1(net843),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4576_ (.A(_1377_),
    .B(_1378_),
    .C(_1380_),
    .Y(_1381_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4577_ (.B1(_1377_),
    .VDD(VPWR),
    .Y(_1382_),
    .VSS(VGND),
    .A1(_1378_),
    .A2(_1380_));
 sg13g2_nor2b_1 _4578_ (.A(_1381_),
    .B_N(_1382_),
    .Y(_1383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4579_ (.Y(_1384_),
    .A(_1376_),
    .B(_1383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4580_ (.Y(_1385_),
    .A(_1376_),
    .B(_1383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4581_ (.B(_1385_),
    .A(_1375_),
    .X(_1386_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4582_ (.Y(_1387_),
    .B(_1386_),
    .A_N(_1374_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4583_ (.Y(_0087_),
    .A(_1374_),
    .B(_1386_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4584_ (.Y(_1388_),
    .B1(net837),
    .B2(net903),
    .A2(net839),
    .A1(net901),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4585_ (.Y(_1389_),
    .A(net902),
    .B(net837),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4586_ (.A(net903),
    .B(net902),
    .C(net839),
    .D(net837),
    .X(_1390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4587_ (.A(_1388_),
    .B(_1390_),
    .Y(_1391_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4588_ (.VDD(VPWR),
    .Y(_1392_),
    .A(_1391_),
    .VSS(VGND));
 sg13g2_o21ai_1 _4589_ (.B1(_1379_),
    .VDD(VPWR),
    .Y(_1393_),
    .VSS(VGND),
    .A1(_1377_),
    .A2(_1380_));
 sg13g2_nand2_1 _4590_ (.Y(_1394_),
    .A(net899),
    .B(net841),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4591_ (.A(net848),
    .B(net844),
    .C(net897),
    .D(net895),
    .X(_1395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4592_ (.B(net844),
    .C(net897),
    .A(net848),
    .Y(_1396_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net895));
 sg13g2_a22oi_1 _4593_ (.Y(_1397_),
    .B1(net895),
    .B2(net848),
    .A2(net897),
    .A1(net844),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4594_ (.A(_1394_),
    .B(_1395_),
    .C(_1397_),
    .X(_1398_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4595_ (.B1(_1394_),
    .VDD(VPWR),
    .Y(_1399_),
    .VSS(VGND),
    .A1(_1395_),
    .A2(_1397_));
 sg13g2_nand3_1 _4596_ (.B(_1398_),
    .C(_1399_),
    .A(_1393_),
    .Y(_1400_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4597_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1398_),
    .A2(_1399_),
    .Y(_1401_),
    .B1(_1393_));
 sg13g2_a21o_1 _4598_ (.A2(_1399_),
    .A1(_1398_),
    .B1(_1393_),
    .X(_1402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4599_ (.Y(_1403_),
    .A(_1400_),
    .B(_1402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4600_ (.Y(_1404_),
    .A(_1392_),
    .B(_1403_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4601_ (.B1(_1384_),
    .VDD(VPWR),
    .Y(_1405_),
    .VSS(VGND),
    .A1(_1375_),
    .A2(_1385_));
 sg13g2_nor2b_2 _4602_ (.A(_1404_),
    .B_N(_1405_),
    .Y(_1406_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4603_ (.B(_1405_),
    .A(_1404_),
    .X(_1407_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4604_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1408_),
    .B(_1407_),
    .A(_1387_));
 sg13g2_xor2_1 _4605_ (.B(_1407_),
    .A(_1387_),
    .X(_0088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4606_ (.B1(_1400_),
    .VDD(VPWR),
    .Y(_1409_),
    .VSS(VGND),
    .A1(_1392_),
    .A2(_1401_));
 sg13g2_nand2_1 _4607_ (.Y(_1410_),
    .A(net904),
    .B(net836),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4608_ (.Y(_1411_),
    .A(net900),
    .B(net837),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4609_ (.Y(_1412_),
    .A(net900),
    .B(net839),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4610_ (.B(_1412_),
    .A(_1389_),
    .X(_1413_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4611_ (.Y(_1414_),
    .B(_1413_),
    .A_N(_1410_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4612_ (.B(_1413_),
    .A(_1410_),
    .X(_1415_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4613_ (.B1(_1396_),
    .VDD(VPWR),
    .Y(_1416_),
    .VSS(VGND),
    .A1(_1394_),
    .A2(_1397_));
 sg13g2_nand2_1 _4614_ (.Y(_1417_),
    .A(net841),
    .B(net898),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4615_ (.A(net850),
    .B(net846),
    .C(net895),
    .D(net894),
    .X(_1418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4616_ (.B(net846),
    .C(net895),
    .A(net850),
    .Y(_1419_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net894));
 sg13g2_a22oi_1 _4617_ (.Y(_1420_),
    .B1(net894),
    .B2(net850),
    .A2(net895),
    .A1(net846),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4618_ (.A(_1417_),
    .B(_1418_),
    .C(_1420_),
    .X(_1421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4619_ (.B1(_1417_),
    .VDD(VPWR),
    .Y(_1422_),
    .VSS(VGND),
    .A1(_1418_),
    .A2(_1420_));
 sg13g2_and3_1 _4620_ (.X(_1423_),
    .A(_1416_),
    .B(_1421_),
    .C(_1422_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4621_ (.B(_1421_),
    .C(_1422_),
    .A(_1416_),
    .Y(_1424_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4622_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1421_),
    .A2(_1422_),
    .Y(_1425_),
    .B1(_1416_));
 sg13g2_or3_1 _4623_ (.A(_1415_),
    .B(_1423_),
    .C(_1425_),
    .X(_1426_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4624_ (.B1(_1415_),
    .VDD(VPWR),
    .Y(_1427_),
    .VSS(VGND),
    .A1(_1423_),
    .A2(_1425_));
 sg13g2_nand3_1 _4625_ (.B(_1426_),
    .C(_1427_),
    .A(_1409_),
    .Y(_1428_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4626_ (.A2(_1427_),
    .A1(_1426_),
    .B1(_1409_),
    .X(_1429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4627_ (.B(_1428_),
    .C(_1429_),
    .A(_1390_),
    .Y(_1430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4628_ (.A2(_1429_),
    .A1(_1428_),
    .B1(_1390_),
    .X(_1431_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4629_ (.A(_1430_),
    .B(_1431_),
    .X(_1432_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4630_ (.B(_1430_),
    .C(_1431_),
    .A(_1406_),
    .Y(_1433_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4631_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1430_),
    .A2(_1431_),
    .Y(_1434_),
    .B1(_1406_));
 sg13g2_xor2_1 _4632_ (.B(_1432_),
    .A(_1406_),
    .X(_1435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4633_ (.Y(_0138_),
    .A(_1408_),
    .B(_1435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4634_ (.Y(_1436_),
    .A(_1428_),
    .B(_1430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4635_ (.B1(_1414_),
    .VDD(VPWR),
    .Y(_1437_),
    .VSS(VGND),
    .A1(_1389_),
    .A2(_1412_));
 sg13g2_nand2_1 _4636_ (.Y(_1438_),
    .A(net904),
    .B(net835),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4637_ (.Y(_1439_),
    .B(_1437_),
    .A_N(_1438_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4638_ (.B(_1438_),
    .A(_1437_),
    .X(_1440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4639_ (.B1(_1424_),
    .VDD(VPWR),
    .Y(_1441_),
    .VSS(VGND),
    .A1(_1415_),
    .A2(_1425_));
 sg13g2_nand2_1 _4640_ (.Y(_1442_),
    .A(net902),
    .B(\DP_4.matrix[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4641_ (.Y(_1443_),
    .A(net898),
    .B(net837),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4642_ (.Y(_1444_),
    .A(net898),
    .B(net840),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4643_ (.B(_1444_),
    .A(_1411_),
    .X(_1445_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4644_ (.Y(_1446_),
    .B(_1445_),
    .A_N(_1442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4645_ (.Y(_1447_),
    .A(_1442_),
    .B(_1445_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4646_ (.B1(_1419_),
    .VDD(VPWR),
    .Y(_1448_),
    .VSS(VGND),
    .A1(_1417_),
    .A2(_1420_));
 sg13g2_nand2_1 _4647_ (.Y(_1449_),
    .A(net841),
    .B(net896),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4648_ (.A(net849),
    .B(net846),
    .C(net894),
    .D(net892),
    .X(_1450_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4649_ (.B(net845),
    .C(net893),
    .A(net849),
    .Y(_1451_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net892));
 sg13g2_a22oi_1 _4650_ (.Y(_1452_),
    .B1(net892),
    .B2(net849),
    .A2(net893),
    .A1(net846),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4651_ (.A(_1449_),
    .B(_1450_),
    .C(_1452_),
    .X(_1453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4652_ (.B1(_1449_),
    .VDD(VPWR),
    .Y(_1454_),
    .VSS(VGND),
    .A1(_1450_),
    .A2(_1452_));
 sg13g2_and3_1 _4653_ (.X(_1455_),
    .A(_1448_),
    .B(_1453_),
    .C(_1454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4654_ (.B(_1453_),
    .C(_1454_),
    .A(_1448_),
    .Y(_1456_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4655_ (.A2(_1454_),
    .A1(_1453_),
    .B1(_1448_),
    .X(_1457_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4656_ (.B(_1456_),
    .C(_1457_),
    .A(_1447_),
    .Y(_1458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4657_ (.A2(_1457_),
    .A1(_1456_),
    .B1(_1447_),
    .X(_1459_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4658_ (.B(_1458_),
    .C(_1459_),
    .A(_1441_),
    .Y(_1460_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4659_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1458_),
    .A2(_1459_),
    .Y(_1461_),
    .B1(_1441_));
 sg13g2_a21o_1 _4660_ (.A2(_1459_),
    .A1(_1458_),
    .B1(_1441_),
    .X(_1462_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4661_ (.Y(_1463_),
    .A(_1460_),
    .B(_1462_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4662_ (.Y(_1464_),
    .A(_1440_),
    .B(_1463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4663_ (.A(_1464_),
    .B_N(_1436_),
    .Y(_1465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4664_ (.Y(_1466_),
    .A(_1436_),
    .B(_1464_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4665_ (.B1(_1433_),
    .VDD(VPWR),
    .Y(_1467_),
    .VSS(VGND),
    .A1(_1408_),
    .A2(_1434_));
 sg13g2_xor2_1 _4666_ (.B(_1467_),
    .A(_1466_),
    .X(_0145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4667_ (.B1(_1460_),
    .VDD(VPWR),
    .Y(_1468_),
    .VSS(VGND),
    .A1(_1440_),
    .A2(_1461_));
 sg13g2_o21ai_1 _4668_ (.B1(_1446_),
    .VDD(VPWR),
    .Y(_1469_),
    .VSS(VGND),
    .A1(_1411_),
    .A2(_1444_));
 sg13g2_a22oi_1 _4669_ (.Y(_1470_),
    .B1(net832),
    .B2(net904),
    .A2(net834),
    .A1(net902),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4670_ (.B(\DP_3.matrix[1] ),
    .C(net834),
    .A(net904),
    .Y(_1471_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net832));
 sg13g2_nor2b_1 _4671_ (.A(_1470_),
    .B_N(_1471_),
    .Y(_1472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4672_ (.Y(_1473_),
    .A(_1469_),
    .B(_1472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4673_ (.Y(_1474_),
    .A(_1469_),
    .B(_1472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4674_ (.A2(_1457_),
    .A1(_1447_),
    .B1(_1455_),
    .X(_1475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4675_ (.Y(_1476_),
    .A(net900),
    .B(net836),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4676_ (.Y(_1477_),
    .A(net896),
    .B(net838),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4677_ (.Y(_1478_),
    .A(net840),
    .B(net896),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4678_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1479_),
    .B(_1477_),
    .A(_1444_));
 sg13g2_and2_1 _4679_ (.A(_1443_),
    .B(_1478_),
    .X(_1480_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4680_ (.Y(_1481_),
    .A(_1443_),
    .B(_1478_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4681_ (.Y(_1482_),
    .A(_1476_),
    .B(_1481_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4682_ (.B1(_1451_),
    .VDD(VPWR),
    .Y(_1483_),
    .VSS(VGND),
    .A1(_1449_),
    .A2(_1452_));
 sg13g2_nand2_1 _4683_ (.Y(_1484_),
    .A(net841),
    .B(net893),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4684_ (.A(net849),
    .B(net845),
    .C(net892),
    .D(net890),
    .X(_1485_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4685_ (.B(net845),
    .C(net891),
    .A(net849),
    .Y(_1486_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net890));
 sg13g2_a22oi_1 _4686_ (.Y(_1487_),
    .B1(net890),
    .B2(net849),
    .A2(net891),
    .A1(net845),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4687_ (.A(_1484_),
    .B(_1485_),
    .C(_1487_),
    .X(_1488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4688_ (.B1(_1484_),
    .VDD(VPWR),
    .Y(_1489_),
    .VSS(VGND),
    .A1(_1485_),
    .A2(_1487_));
 sg13g2_and3_1 _4689_ (.X(_1490_),
    .A(_1483_),
    .B(_1488_),
    .C(_1489_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4690_ (.B(_1488_),
    .C(_1489_),
    .A(_1483_),
    .Y(_1491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4691_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1488_),
    .A2(_1489_),
    .Y(_1492_),
    .B1(_1483_));
 sg13g2_or3_1 _4692_ (.A(_1482_),
    .B(_1490_),
    .C(_1492_),
    .X(_1493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4693_ (.B1(_1482_),
    .VDD(VPWR),
    .Y(_1494_),
    .VSS(VGND),
    .A1(_1490_),
    .A2(_1492_));
 sg13g2_and3_1 _4694_ (.X(_1495_),
    .A(_1475_),
    .B(_1493_),
    .C(_1494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4695_ (.B(_1493_),
    .C(_1494_),
    .A(_1475_),
    .Y(_1496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4696_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1493_),
    .A2(_1494_),
    .Y(_1497_),
    .B1(_1475_));
 sg13g2_or3_1 _4697_ (.A(_1474_),
    .B(_1495_),
    .C(_1497_),
    .X(_1498_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4698_ (.B1(_1474_),
    .VDD(VPWR),
    .Y(_1499_),
    .VSS(VGND),
    .A1(_1495_),
    .A2(_1497_));
 sg13g2_nand3_1 _4699_ (.B(_1498_),
    .C(_1499_),
    .A(_1468_),
    .Y(_1500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4700_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1498_),
    .A2(_1499_),
    .Y(_1501_),
    .B1(_1468_));
 sg13g2_a21o_1 _4701_ (.A2(_1499_),
    .A1(_1498_),
    .B1(_1468_),
    .X(_1502_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4702_ (.Y(_1503_),
    .A(_1500_),
    .B(_1502_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4703_ (.B(_1503_),
    .A(_1439_),
    .X(_1504_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _4704_ (.A2(_1467_),
    .A1(_1466_),
    .B1(_1465_),
    .X(_1505_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4705_ (.Y(_1506_),
    .A(_1504_),
    .B(_1505_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4706_ (.B(_1505_),
    .A(_1504_),
    .X(_0146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4707_ (.B1(_1496_),
    .VDD(VPWR),
    .Y(_1507_),
    .VSS(VGND),
    .A1(_1474_),
    .A2(_1497_));
 sg13g2_o21ai_1 _4708_ (.B1(_1479_),
    .VDD(VPWR),
    .Y(_1508_),
    .VSS(VGND),
    .A1(_1476_),
    .A2(_1480_));
 sg13g2_nand2_1 _4709_ (.Y(_1509_),
    .A(net904),
    .B(net1023),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4710_ (.Y(_1510_),
    .A(net900),
    .B(net832),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4711_ (.A(net902),
    .B(net900),
    .C(net834),
    .D(net832),
    .X(_1511_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4712_ (.Y(_1512_),
    .B1(net832),
    .B2(net902),
    .A2(net834),
    .A1(net900),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4713_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1513_),
    .B(_1512_),
    .A(_1511_));
 sg13g2_nor2_1 _4714_ (.A(_1509_),
    .B(_1513_),
    .Y(_1514_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4715_ (.B(_1513_),
    .A(_1509_),
    .X(_1515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4716_ (.Y(_1516_),
    .A(_1508_),
    .B(_1515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4717_ (.Y(_1517_),
    .A(_1508_),
    .B(_1515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4718_ (.Y(_1518_),
    .A(_1471_),
    .B(_1517_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4719_ (.B1(_1491_),
    .VDD(VPWR),
    .Y(_1519_),
    .VSS(VGND),
    .A1(_1482_),
    .A2(_1492_));
 sg13g2_nand2_1 _4720_ (.Y(_1520_),
    .A(net898),
    .B(net836),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4721_ (.Y(_1521_),
    .A(net838),
    .B(net893),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4722_ (.Y(_1522_),
    .A(net839),
    .B(net894),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4723_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1523_),
    .B(_1521_),
    .A(_1478_));
 sg13g2_xnor2_1 _4724_ (.Y(_1524_),
    .A(_1477_),
    .B(_1522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4725_ (.Y(_1525_),
    .A(_1520_),
    .B(_1524_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4726_ (.B1(_1486_),
    .VDD(VPWR),
    .Y(_1526_),
    .VSS(VGND),
    .A1(_1484_),
    .A2(_1487_));
 sg13g2_nand2_1 _4727_ (.Y(_1527_),
    .A(net842),
    .B(net891),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4728_ (.A(net850),
    .B(net845),
    .C(net888),
    .D(net1028),
    .X(_1528_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4729_ (.B(net845),
    .C(net888),
    .A(net849),
    .Y(_1529_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net1028));
 sg13g2_a22oi_1 _4730_ (.Y(_1530_),
    .B1(net1028),
    .B2(net849),
    .A2(net888),
    .A1(net845),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4731_ (.A(_1527_),
    .B(_1528_),
    .C(_1530_),
    .X(_1531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4732_ (.B1(_1527_),
    .VDD(VPWR),
    .Y(_1532_),
    .VSS(VGND),
    .A1(_1528_),
    .A2(_1530_));
 sg13g2_and3_1 _4733_ (.X(_1533_),
    .A(_1526_),
    .B(_1531_),
    .C(_1532_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4734_ (.B(_1531_),
    .C(_1532_),
    .A(_1526_),
    .Y(_1534_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4735_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1531_),
    .A2(_1532_),
    .Y(_1535_),
    .B1(_1526_));
 sg13g2_or3_1 _4736_ (.A(_1525_),
    .B(_1533_),
    .C(_1535_),
    .X(_1536_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4737_ (.B1(_1525_),
    .VDD(VPWR),
    .Y(_1537_),
    .VSS(VGND),
    .A1(_1533_),
    .A2(_1535_));
 sg13g2_and3_1 _4738_ (.X(_1538_),
    .A(_1519_),
    .B(_1536_),
    .C(_1537_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4739_ (.B(_1536_),
    .C(_1537_),
    .A(_1519_),
    .Y(_1539_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4740_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1536_),
    .A2(_1537_),
    .Y(_1540_),
    .B1(_1519_));
 sg13g2_or3_1 _4741_ (.A(_1518_),
    .B(_1538_),
    .C(_1540_),
    .X(_1541_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4742_ (.B1(_1518_),
    .VDD(VPWR),
    .Y(_1542_),
    .VSS(VGND),
    .A1(_1538_),
    .A2(_1540_));
 sg13g2_and3_1 _4743_ (.X(_1543_),
    .A(_1507_),
    .B(_1541_),
    .C(_1542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4744_ (.B(_1541_),
    .C(_1542_),
    .A(_1507_),
    .Y(_1544_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4745_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1541_),
    .A2(_1542_),
    .Y(_1545_),
    .B1(_1507_));
 sg13g2_or3_1 _4746_ (.A(_1473_),
    .B(_1543_),
    .C(_1545_),
    .X(_1546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4747_ (.B1(_1473_),
    .VDD(VPWR),
    .Y(_1547_),
    .VSS(VGND),
    .A1(_1543_),
    .A2(_1545_));
 sg13g2_o21ai_1 _4748_ (.B1(_1500_),
    .VDD(VPWR),
    .Y(_1548_),
    .VSS(VGND),
    .A1(_1439_),
    .A2(_1501_));
 sg13g2_nand3_1 _4749_ (.B(_1547_),
    .C(_1548_),
    .A(_1546_),
    .Y(_1549_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4750_ (.A2(_1547_),
    .A1(_1546_),
    .B1(_1548_),
    .X(_1550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4751_ (.Y(_1551_),
    .A(_1549_),
    .B(_1550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4752_ (.A(_1504_),
    .B(_1505_),
    .C(_1549_),
    .D(_1550_),
    .X(_1552_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4753_ (.B(_1551_),
    .A(_1506_),
    .X(_0147_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4754_ (.B1(_1549_),
    .VDD(VPWR),
    .Y(_1553_),
    .VSS(VGND),
    .A1(_1506_),
    .A2(_1551_));
 sg13g2_o21ai_1 _4755_ (.B1(_1544_),
    .VDD(VPWR),
    .Y(_1554_),
    .VSS(VGND),
    .A1(_1473_),
    .A2(_1545_));
 sg13g2_o21ai_1 _4756_ (.B1(_1516_),
    .VDD(VPWR),
    .Y(_1555_),
    .VSS(VGND),
    .A1(_1471_),
    .A2(_1517_));
 sg13g2_o21ai_1 _4757_ (.B1(_1539_),
    .VDD(VPWR),
    .Y(_1556_),
    .VSS(VGND),
    .A1(_1518_),
    .A2(_1540_));
 sg13g2_nor2_1 _4758_ (.A(_1511_),
    .B(_1514_),
    .Y(_1557_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4759_ (.B1(_1523_),
    .VDD(VPWR),
    .Y(_1558_),
    .VSS(VGND),
    .A1(_1520_),
    .A2(_1524_));
 sg13g2_nand2_1 _4760_ (.Y(_1559_),
    .A(net902),
    .B(net1023),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4761_ (.Y(_1560_),
    .A(net898),
    .B(net832),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4762_ (.Y(_1561_),
    .A(net898),
    .B(net834),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4763_ (.B(_1561_),
    .A(_1510_),
    .X(_1562_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4764_ (.Y(_1563_),
    .B(_1562_),
    .A_N(_1559_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4765_ (.Y(_1564_),
    .A(_1559_),
    .B(_1562_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4766_ (.Y(_1565_),
    .A(_1558_),
    .B(_1564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4767_ (.A(_1557_),
    .B(_1565_),
    .Y(_1566_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4768_ (.Y(_1567_),
    .A(_1557_),
    .B(_1565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4769_ (.B1(_1534_),
    .VDD(VPWR),
    .Y(_1568_),
    .VSS(VGND),
    .A1(_1525_),
    .A2(_1535_));
 sg13g2_nand2_1 _4770_ (.Y(_1569_),
    .A(net896),
    .B(net836),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4771_ (.Y(_1570_),
    .A(net839),
    .B(net891),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4772_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1571_),
    .B(_1570_),
    .A(_1521_));
 sg13g2_and2_1 _4773_ (.A(_1521_),
    .B(_1570_),
    .X(_1572_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4774_ (.Y(_1573_),
    .A(_1521_),
    .B(_1570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4775_ (.Y(_1574_),
    .A(_1569_),
    .B(_1573_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4776_ (.B1(_1529_),
    .VDD(VPWR),
    .Y(_1575_),
    .VSS(VGND),
    .A1(_1527_),
    .A2(_1530_));
 sg13g2_nand2_1 _4777_ (.Y(_1576_),
    .A(net842),
    .B(net1029),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4778_ (.A(net845),
    .B(net842),
    .C(net888),
    .D(net1029),
    .X(_1577_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4779_ (.Y(_1578_),
    .B1(net1029),
    .B2(net846),
    .A2(net888),
    .A1(net842),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4780_ (.A(_1577_),
    .B(_1578_),
    .Y(_1579_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4781_ (.Y(_1580_),
    .A(_1575_),
    .B(_1579_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4782_ (.Y(_1581_),
    .A(_1575_),
    .B(_1579_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4783_ (.B(_1581_),
    .A(_1574_),
    .X(_1582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4784_ (.Y(_1583_),
    .A(_1568_),
    .B(_1582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4785_ (.Y(_1584_),
    .A(_1568_),
    .B(_1582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4786_ (.B(_1584_),
    .A(_1567_),
    .X(_1585_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4787_ (.Y(_1586_),
    .A(_1556_),
    .B(_1585_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4788_ (.Y(_1587_),
    .A(_1556_),
    .B(_1585_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4789_ (.Y(_1588_),
    .B(_1555_),
    .A_N(_1587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4790_ (.Y(_1589_),
    .A(_1555_),
    .B(_1587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4791_ (.A(_1554_),
    .B(_1589_),
    .Y(_1590_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4792_ (.Y(_1591_),
    .A(_1554_),
    .B(_1589_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4793_ (.A(_1590_),
    .B_N(_1591_),
    .Y(_1592_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4794_ (.B(_1592_),
    .A(_1553_),
    .X(_0148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4795_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1558_),
    .A2(_1564_),
    .Y(_1593_),
    .B1(_1566_));
 sg13g2_o21ai_1 _4796_ (.B1(_1583_),
    .VDD(VPWR),
    .Y(_1594_),
    .VSS(VGND),
    .A1(_1567_),
    .A2(_1584_));
 sg13g2_o21ai_1 _4797_ (.B1(_1563_),
    .VDD(VPWR),
    .Y(_1595_),
    .VSS(VGND),
    .A1(_1510_),
    .A2(_1561_));
 sg13g2_o21ai_1 _4798_ (.B1(_1571_),
    .VDD(VPWR),
    .Y(_1596_),
    .VSS(VGND),
    .A1(_1569_),
    .A2(_1572_));
 sg13g2_nand2_1 _4799_ (.Y(_1597_),
    .A(net900),
    .B(net1023),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4800_ (.Y(_1598_),
    .A(net896),
    .B(net833),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4801_ (.Y(_1599_),
    .A(net896),
    .B(net835),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4802_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1600_),
    .B(_1598_),
    .A(_1561_));
 sg13g2_xnor2_1 _4803_ (.Y(_1601_),
    .A(_1560_),
    .B(_1599_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4804_ (.B(_1601_),
    .A(_1597_),
    .X(_1602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4805_ (.Y(_1603_),
    .A(_1596_),
    .B(_1602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4806_ (.A(_1603_),
    .B_N(_1595_),
    .Y(_1604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4807_ (.B(_1603_),
    .A(_1595_),
    .X(_1605_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4808_ (.B1(_1580_),
    .VDD(VPWR),
    .Y(_1606_),
    .VSS(VGND),
    .A1(_1574_),
    .A2(_1581_));
 sg13g2_a21oi_1 _4809_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net846),
    .A2(net888),
    .Y(_1607_),
    .B1(_1576_));
 sg13g2_nand2_1 _4810_ (.Y(_1608_),
    .A(net893),
    .B(net836),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4811_ (.Y(_1609_),
    .A(net838),
    .B(net889),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4812_ (.A(net840),
    .B(net837),
    .C(net891),
    .D(net888),
    .X(_1610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4813_ (.Y(_1611_),
    .B1(net888),
    .B2(net840),
    .A2(net891),
    .A1(net838),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4814_ (.A(_1608_),
    .B(_1610_),
    .C(_1611_),
    .Y(_1612_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4815_ (.B1(_1608_),
    .VDD(VPWR),
    .Y(_1613_),
    .VSS(VGND),
    .A1(_1610_),
    .A2(_1611_));
 sg13g2_nor2b_1 _4816_ (.A(_1612_),
    .B_N(_1613_),
    .Y(_1614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4817_ (.Y(_1615_),
    .A(_1607_),
    .B(_1614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4818_ (.Y(_1616_),
    .B(_1606_),
    .A_N(_1615_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4819_ (.B(_1615_),
    .A(_1606_),
    .X(_1617_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4820_ (.B(_1617_),
    .A(_1605_),
    .X(_1618_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4821_ (.Y(_1619_),
    .A(_1594_),
    .B(_1618_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4822_ (.B(_1618_),
    .A(_1594_),
    .X(_1620_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4823_ (.Y(_1621_),
    .B(_1620_),
    .A_N(_1593_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4824_ (.B(_1620_),
    .A(_1593_),
    .X(_1622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4825_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1586_),
    .A2(_1588_),
    .Y(_1623_),
    .B1(_1622_));
 sg13g2_nand3_1 _4826_ (.B(_1588_),
    .C(_1622_),
    .A(_1586_),
    .Y(_1624_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4827_ (.Y(_1625_),
    .B(_1624_),
    .A_N(_1623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4828_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1549_),
    .A2(_1591_),
    .Y(_1626_),
    .B1(_1590_));
 sg13g2_a21oi_2 _4829_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_1626_),
    .Y(_1627_),
    .A2(_1592_),
    .A1(_1552_));
 sg13g2_nor2_1 _4830_ (.A(_1625_),
    .B(_1627_),
    .Y(_1628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4831_ (.B(_1627_),
    .A(_1625_),
    .X(_0139_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4832_ (.A2(_1602_),
    .A1(_1596_),
    .B1(_1604_),
    .X(_1629_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4833_ (.B1(_1616_),
    .VDD(VPWR),
    .Y(_1630_),
    .VSS(VGND),
    .A1(_1605_),
    .A2(_1617_));
 sg13g2_a21o_2 _4834_ (.A2(_1614_),
    .A1(_1607_),
    .B1(_1577_),
    .X(_1631_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4835_ (.Y(_1632_),
    .A(net836),
    .B(net891),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4836_ (.Y(_1633_),
    .A(net840),
    .B(net1028),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4837_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1634_),
    .B(_1633_),
    .A(_1609_));
 sg13g2_xnor2_1 _4838_ (.Y(_1635_),
    .A(_1609_),
    .B(_1633_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4839_ (.B(_1635_),
    .A(_1632_),
    .X(_1636_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4840_ (.Y(_1637_),
    .A(_1631_),
    .B(_1636_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4841_ (.B1(_1600_),
    .VDD(VPWR),
    .Y(_1638_),
    .VSS(VGND),
    .A1(_1597_),
    .A2(_1601_));
 sg13g2_or2_1 _4842_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1639_),
    .B(_1612_),
    .A(_1610_));
 sg13g2_nand2_1 _4843_ (.Y(_1640_),
    .A(net898),
    .B(net1023),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4844_ (.Y(_1641_),
    .A(net893),
    .B(net834),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4845_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1642_),
    .B(_1641_),
    .A(_1598_));
 sg13g2_xnor2_1 _4846_ (.Y(_1643_),
    .A(_1598_),
    .B(_1641_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4847_ (.B(_1643_),
    .A(_1640_),
    .X(_1644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4848_ (.Y(_1645_),
    .A(_1639_),
    .B(_1644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4849_ (.A(_1645_),
    .B_N(_1638_),
    .Y(_1646_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4850_ (.B(_1645_),
    .A(_1638_),
    .X(_1647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4851_ (.A(_1637_),
    .B(_1647_),
    .Y(_1648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4852_ (.B(_1647_),
    .A(_1637_),
    .X(_1649_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4853_ (.Y(_1650_),
    .A(_1630_),
    .B(_1649_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4854_ (.A(_1650_),
    .B_N(_1629_),
    .Y(_1651_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4855_ (.B(_1650_),
    .A(_1629_),
    .X(_1652_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4856_ (.B(_1621_),
    .C(_1652_),
    .A(_1619_),
    .Y(_1653_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4857_ (.VDD(VPWR),
    .Y(_1654_),
    .A(_1653_),
    .VSS(VGND));
 sg13g2_a21oi_1 _4858_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1619_),
    .A2(_1621_),
    .Y(_1655_),
    .B1(_1652_));
 sg13g2_nor2_1 _4859_ (.A(_1654_),
    .B(_1655_),
    .Y(_1656_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4860_ (.A(_1623_),
    .B(_1628_),
    .Y(_1657_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4861_ (.Y(_0140_),
    .A(_1656_),
    .B(_1657_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4862_ (.A2(_1644_),
    .A1(_1639_),
    .B1(_1646_),
    .X(_1658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4863_ (.Y(_1659_),
    .B1(net1028),
    .B2(net838),
    .A2(net889),
    .A1(\DP_4.matrix[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4864_ (.Y(_1660_),
    .A(\DP_4.matrix[5] ),
    .B(net1028),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4865_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1661_),
    .B(_1660_),
    .A(_1609_));
 sg13g2_nand2b_1 _4866_ (.Y(_1662_),
    .B(_1661_),
    .A_N(_1659_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4867_ (.B1(_1642_),
    .VDD(VPWR),
    .Y(_1663_),
    .VSS(VGND),
    .A1(_1640_),
    .A2(_1643_));
 sg13g2_o21ai_1 _4868_ (.B1(_1634_),
    .VDD(VPWR),
    .Y(_1664_),
    .VSS(VGND),
    .A1(_1632_),
    .A2(_1635_));
 sg13g2_nand2_1 _4869_ (.Y(_1665_),
    .A(net896),
    .B(net1023),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4870_ (.Y(_1666_),
    .A(net891),
    .B(net833),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4871_ (.A(_1641_),
    .B(_1666_),
    .Y(_1667_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4872_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1668_),
    .B(_1666_),
    .A(_1641_));
 sg13g2_a22oi_1 _4873_ (.Y(_1669_),
    .B1(net833),
    .B2(net893),
    .A2(net834),
    .A1(\DP_3.matrix[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4874_ (.A(_1667_),
    .B(_1669_),
    .Y(_1670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4875_ (.Y(_1671_),
    .A(_1665_),
    .B(_1670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4876_ (.Y(_1672_),
    .A(_1664_),
    .B(_1671_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4877_ (.A(_1672_),
    .B_N(_1663_),
    .Y(_1673_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4878_ (.B(_1672_),
    .A(_1663_),
    .X(_1674_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4879_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1675_),
    .B(_1674_),
    .A(_1662_));
 sg13g2_xor2_1 _4880_ (.B(_1674_),
    .A(_1662_),
    .X(_1676_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4881_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1631_),
    .A2(_1636_),
    .Y(_1677_),
    .B1(_1648_));
 sg13g2_nor2b_1 _4882_ (.A(_1677_),
    .B_N(_1676_),
    .Y(_1678_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4883_ (.B(_1677_),
    .A(_1676_),
    .X(_1679_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4884_ (.A(_1679_),
    .B_N(_1658_),
    .Y(_1680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4885_ (.B(_1679_),
    .A(_1658_),
    .X(_1681_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4886_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1630_),
    .A2(_1649_),
    .Y(_1682_),
    .B1(_1651_));
 sg13g2_nor2_1 _4887_ (.A(_1681_),
    .B(_1682_),
    .Y(_1683_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4888_ (.B(_1682_),
    .A(_1681_),
    .X(_1684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4889_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1623_),
    .A2(_1653_),
    .Y(_1685_),
    .B1(_1655_));
 sg13g2_a21oi_1 _4890_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1624_),
    .A2(_1653_),
    .Y(_1686_),
    .B1(_1655_));
 sg13g2_a21oi_2 _4891_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_1686_),
    .Y(_1687_),
    .A2(_1685_),
    .A1(_1627_));
 sg13g2_xor2_1 _4892_ (.B(_1687_),
    .A(_1684_),
    .X(_0141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4893_ (.A2(_1671_),
    .A1(_1664_),
    .B1(_1673_),
    .X(_1688_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4894_ (.B1(_1668_),
    .VDD(VPWR),
    .Y(_1689_),
    .VSS(VGND),
    .A1(_1665_),
    .A2(_1669_));
 sg13g2_nand2_1 _4895_ (.Y(_1690_),
    .A(net893),
    .B(net1023),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4896_ (.Y(_1691_),
    .A(net889),
    .B(net833),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4897_ (.Y(_1692_),
    .A(net835),
    .B(net889),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4898_ (.B(_1692_),
    .A(_1666_),
    .X(_1693_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4899_ (.Y(_1694_),
    .B(_1693_),
    .A_N(_1690_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4900_ (.Y(_1695_),
    .A(_1690_),
    .B(_1693_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4901_ (.A(_1661_),
    .B_N(_1695_),
    .Y(_1696_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4902_ (.Y(_1697_),
    .A(_1661_),
    .B(_1695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4903_ (.Y(_1698_),
    .A(_1689_),
    .B(_1697_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4904_ (.A(_1660_),
    .B(_1698_),
    .Y(_1699_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4905_ (.B(_1698_),
    .A(_1660_),
    .X(_1700_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4906_ (.Y(_1701_),
    .B(_1700_),
    .A_N(_1675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4907_ (.Y(_1702_),
    .A(_1675_),
    .B(_1700_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4908_ (.Y(_1703_),
    .A(_1688_),
    .B(_1702_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4909_ (.B(_1702_),
    .A(_1688_),
    .X(_1704_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4910_ (.B1(_1704_),
    .VDD(VPWR),
    .Y(_1705_),
    .VSS(VGND),
    .A1(_1678_),
    .A2(_1680_));
 sg13g2_or3_1 _4911_ (.A(_1678_),
    .B(_1680_),
    .C(_1704_),
    .X(_1706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4912_ (.A(_1705_),
    .B(_1706_),
    .X(_1707_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4913_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1684_),
    .A2(_1687_),
    .Y(_1708_),
    .B1(_1683_));
 sg13g2_xnor2_1 _4914_ (.Y(_0142_),
    .A(_1707_),
    .B(_1708_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4915_ (.A(_1684_),
    .B(_1707_),
    .X(_1709_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4916_ (.Y(_1710_),
    .A(_1683_),
    .B(_1706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4917_ (.Y(_1711_),
    .A(_1705_),
    .B(_1710_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4918_ (.A2(_1709_),
    .A1(_1687_),
    .B1(_1711_),
    .X(_1712_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4919_ (.A(_1701_),
    .B(_1703_),
    .X(_1713_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4920_ (.A2(_1697_),
    .A1(_1689_),
    .B1(_1696_),
    .X(_1714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4921_ (.B1(_1694_),
    .VDD(VPWR),
    .Y(_1715_),
    .VSS(VGND),
    .A1(_1666_),
    .A2(_1692_));
 sg13g2_nand2_1 _4922_ (.Y(_1716_),
    .A(net892),
    .B(\DP_4.matrix[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4923_ (.Y(_1717_),
    .A(net833),
    .B(net1029),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4924_ (.Y(_1718_),
    .A(net834),
    .B(net1029),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4925_ (.B(_1718_),
    .A(_1691_),
    .X(_1719_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4926_ (.Y(_1720_),
    .B(_1719_),
    .A_N(_1716_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4927_ (.Y(_1721_),
    .A(_1716_),
    .B(_1719_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4928_ (.Y(_1722_),
    .A(_1715_),
    .B(_1721_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4929_ (.B(_1721_),
    .A(_1715_),
    .X(_1723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4930_ (.Y(_1724_),
    .A(_1699_),
    .B(_1723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4931_ (.A(_1724_),
    .B_N(_1714_),
    .Y(_1725_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4932_ (.B(_1724_),
    .A(_1714_),
    .X(_1726_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4933_ (.A(_1713_),
    .B(_1726_),
    .Y(_1727_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4934_ (.B(_1726_),
    .A(_1713_),
    .X(_1728_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4935_ (.B(_1728_),
    .A(_1712_),
    .X(_0143_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4936_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1712_),
    .A2(_1728_),
    .Y(_1729_),
    .B1(_1727_));
 sg13g2_a21oi_1 _4937_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1699_),
    .A2(_1723_),
    .Y(_1730_),
    .B1(_1725_));
 sg13g2_o21ai_1 _4938_ (.B1(_1720_),
    .VDD(VPWR),
    .Y(_1731_),
    .VSS(VGND),
    .A1(_1691_),
    .A2(_1718_));
 sg13g2_nand2_1 _4939_ (.Y(_1732_),
    .A(net889),
    .B(\DP_4.matrix[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4940_ (.Y(_1733_),
    .A(_1717_),
    .B(_1732_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4941_ (.Y(_1734_),
    .A(_1731_),
    .B(_1733_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4942_ (.Y(_1735_),
    .A(_1722_),
    .B(_1734_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4943_ (.Y(_1736_),
    .A(_1730_),
    .B(_1735_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4944_ (.Y(_0144_),
    .A(_1729_),
    .B(_1736_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4945_ (.A(net869),
    .B(net282),
    .X(_0089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _4946_ (.X(_1737_),
    .A(net867),
    .B(net810),
    .C(_0089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4947_ (.Y(_1738_),
    .B1(net809),
    .B2(net869),
    .A2(net293),
    .A1(net812),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4948_ (.A(_1737_),
    .B(net294),
    .Y(_0090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4949_ (.Y(_1739_),
    .A(net869),
    .B(net805),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4950_ (.A(net812),
    .B(net867),
    .C(net809),
    .D(net865),
    .X(_1740_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4951_ (.Y(_1741_),
    .B1(net865),
    .B2(net812),
    .A2(net809),
    .A1(net867),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4952_ (.A(_1739_),
    .B(_1740_),
    .C(_1741_),
    .Y(_1742_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4953_ (.B1(_1739_),
    .VDD(VPWR),
    .Y(_1743_),
    .VSS(VGND),
    .A1(_1740_),
    .A2(_1741_));
 sg13g2_nor2b_1 _4954_ (.A(_1742_),
    .B_N(_1743_),
    .Y(_1744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4955_ (.Y(_1745_),
    .A(_1737_),
    .B(_1744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4956_ (.B(_1744_),
    .A(_1737_),
    .X(_0091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4957_ (.Y(_1746_),
    .A(net868),
    .B(net803),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4958_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1747_),
    .B(_1742_),
    .A(_1740_));
 sg13g2_nand2_1 _4959_ (.Y(_1748_),
    .A(net867),
    .B(net805),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4960_ (.A(net812),
    .B(net809),
    .C(net863),
    .D(net861),
    .X(_1749_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4961_ (.B(net809),
    .C(net864),
    .A(net812),
    .Y(_1750_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net860));
 sg13g2_a22oi_1 _4962_ (.Y(_1751_),
    .B1(net860),
    .B2(net812),
    .A2(net864),
    .A1(net809),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4963_ (.A(_1748_),
    .B(_1749_),
    .C(_1751_),
    .Y(_1752_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4964_ (.B1(_1748_),
    .VDD(VPWR),
    .Y(_1753_),
    .VSS(VGND),
    .A1(_1749_),
    .A2(_1751_));
 sg13g2_nor2b_1 _4965_ (.A(_1752_),
    .B_N(_1753_),
    .Y(_1754_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4966_ (.Y(_1755_),
    .A(_1747_),
    .B(_1754_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4967_ (.Y(_1756_),
    .A(_1747_),
    .B(_1754_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4968_ (.B(_1756_),
    .A(_1746_),
    .X(_1757_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4969_ (.Y(_1758_),
    .B(_1757_),
    .A_N(_1745_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4970_ (.Y(_0092_),
    .A(_1745_),
    .B(_1757_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4971_ (.Y(_1759_),
    .B1(net800),
    .B2(net869),
    .A2(net802),
    .A1(net867),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4972_ (.Y(_1760_),
    .A(net866),
    .B(net800),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4973_ (.A(net868),
    .B(net866),
    .C(net802),
    .D(net800),
    .X(_1761_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4974_ (.A(_1759_),
    .B(_1761_),
    .Y(_1762_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4975_ (.VDD(VPWR),
    .Y(_1763_),
    .A(_1762_),
    .VSS(VGND));
 sg13g2_o21ai_1 _4976_ (.B1(_1750_),
    .VDD(VPWR),
    .Y(_1764_),
    .VSS(VGND),
    .A1(_1748_),
    .A2(_1751_));
 sg13g2_nand2_1 _4977_ (.Y(_1765_),
    .A(net864),
    .B(net804),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4978_ (.A(net811),
    .B(net808),
    .C(net861),
    .D(net859),
    .X(_1766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4979_ (.B(net808),
    .C(net861),
    .A(net812),
    .Y(_1767_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net859));
 sg13g2_a22oi_1 _4980_ (.Y(_1768_),
    .B1(net859),
    .B2(net811),
    .A2(net861),
    .A1(net808),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4981_ (.A(_1765_),
    .B(_1766_),
    .C(_1768_),
    .X(_1769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4982_ (.B1(_1765_),
    .VDD(VPWR),
    .Y(_1770_),
    .VSS(VGND),
    .A1(_1766_),
    .A2(_1768_));
 sg13g2_nand3_1 _4983_ (.B(_1769_),
    .C(_1770_),
    .A(_1764_),
    .Y(_1771_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4984_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1769_),
    .A2(_1770_),
    .Y(_1772_),
    .B1(_1764_));
 sg13g2_a21o_1 _4985_ (.A2(_1770_),
    .A1(_1769_),
    .B1(_1764_),
    .X(_1773_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4986_ (.Y(_1774_),
    .A(_1771_),
    .B(_1773_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4987_ (.Y(_1775_),
    .A(_1763_),
    .B(_1774_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4988_ (.B1(_1755_),
    .VDD(VPWR),
    .Y(_1776_),
    .VSS(VGND),
    .A1(_1746_),
    .A2(_1756_));
 sg13g2_nor2b_2 _4989_ (.A(_1775_),
    .B_N(_1776_),
    .Y(_1777_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4990_ (.B(_1776_),
    .A(_1775_),
    .X(_1778_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4991_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1779_),
    .B(_1778_),
    .A(_1758_));
 sg13g2_xor2_1 _4992_ (.B(_1778_),
    .A(_1758_),
    .X(_0093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4993_ (.B1(_1771_),
    .VDD(VPWR),
    .Y(_1780_),
    .VSS(VGND),
    .A1(_1763_),
    .A2(_1772_));
 sg13g2_nand2_1 _4994_ (.Y(_1781_),
    .A(net868),
    .B(net798),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4995_ (.Y(_1782_),
    .A(net863),
    .B(net800),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4996_ (.Y(_1783_),
    .A(net863),
    .B(net802),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4997_ (.B(_1783_),
    .A(_1760_),
    .X(_1784_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4998_ (.Y(_1785_),
    .B(_1784_),
    .A_N(_1781_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4999_ (.B(_1784_),
    .A(_1781_),
    .X(_1786_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5000_ (.B1(_1767_),
    .VDD(VPWR),
    .Y(_1787_),
    .VSS(VGND),
    .A1(_1765_),
    .A2(_1768_));
 sg13g2_nand2_1 _5001_ (.Y(_1788_),
    .A(net804),
    .B(net861),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _5002_ (.A(net811),
    .B(net808),
    .C(net858),
    .D(net857),
    .X(_1789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _5003_ (.B(net808),
    .C(net858),
    .A(net811),
    .Y(_1790_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net857));
 sg13g2_a22oi_1 _5004_ (.Y(_1791_),
    .B1(net857),
    .B2(net811),
    .A2(net859),
    .A1(net808),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _5005_ (.A(_1788_),
    .B(_1789_),
    .C(_1791_),
    .X(_1792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5006_ (.B1(_1788_),
    .VDD(VPWR),
    .Y(_1793_),
    .VSS(VGND),
    .A1(_1789_),
    .A2(_1791_));
 sg13g2_and3_1 _5007_ (.X(_1794_),
    .A(_1787_),
    .B(_1792_),
    .C(_1793_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5008_ (.B(_1792_),
    .C(_1793_),
    .A(_1787_),
    .Y(_1795_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5009_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1792_),
    .A2(_1793_),
    .Y(_1796_),
    .B1(_1787_));
 sg13g2_or3_1 _5010_ (.A(_1786_),
    .B(_1794_),
    .C(_1796_),
    .X(_1797_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5011_ (.B1(_1786_),
    .VDD(VPWR),
    .Y(_1798_),
    .VSS(VGND),
    .A1(_1794_),
    .A2(_1796_));
 sg13g2_nand3_1 _5012_ (.B(_1797_),
    .C(_1798_),
    .A(_1780_),
    .Y(_1799_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5013_ (.A2(_1798_),
    .A1(_1797_),
    .B1(_1780_),
    .X(_1800_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5014_ (.B(_1799_),
    .C(_1800_),
    .A(_1761_),
    .Y(_1801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5015_ (.A2(_1800_),
    .A1(_1799_),
    .B1(_1761_),
    .X(_1802_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5016_ (.A(_1801_),
    .B(_1802_),
    .X(_1803_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5017_ (.B(_1801_),
    .C(_1802_),
    .A(_1777_),
    .Y(_1804_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5018_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1801_),
    .A2(_1802_),
    .Y(_1805_),
    .B1(_1777_));
 sg13g2_xor2_1 _5019_ (.B(_1803_),
    .A(_1777_),
    .X(_1806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5020_ (.Y(_0149_),
    .A(_1779_),
    .B(_1806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5021_ (.Y(_1807_),
    .A(_1799_),
    .B(_1801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5022_ (.B1(_1785_),
    .VDD(VPWR),
    .Y(_1808_),
    .VSS(VGND),
    .A1(_1760_),
    .A2(_1783_));
 sg13g2_nand2_1 _5023_ (.Y(_1809_),
    .A(net868),
    .B(net795),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5024_ (.Y(_1810_),
    .B(_1808_),
    .A_N(_1809_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5025_ (.B(_1809_),
    .A(_1808_),
    .X(_1811_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5026_ (.B1(_1795_),
    .VDD(VPWR),
    .Y(_1812_),
    .VSS(VGND),
    .A1(_1786_),
    .A2(_1796_));
 sg13g2_nand2_1 _5027_ (.Y(_1813_),
    .A(net866),
    .B(net798),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5028_ (.Y(_1814_),
    .A(net860),
    .B(net800),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5029_ (.Y(_1815_),
    .A(net860),
    .B(net802),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5030_ (.B(_1815_),
    .A(_1782_),
    .X(_1816_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5031_ (.Y(_1817_),
    .B(_1816_),
    .A_N(_1813_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5032_ (.Y(_1818_),
    .A(_1813_),
    .B(_1816_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5033_ (.B1(_1790_),
    .VDD(VPWR),
    .Y(_1819_),
    .VSS(VGND),
    .A1(_1788_),
    .A2(_1791_));
 sg13g2_nand2_1 _5034_ (.Y(_1820_),
    .A(net804),
    .B(net859),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _5035_ (.A(net811),
    .B(net806),
    .C(net856),
    .D(net855),
    .X(_1821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _5036_ (.B(net806),
    .C(net856),
    .A(net811),
    .Y(_1822_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net855));
 sg13g2_a22oi_1 _5037_ (.Y(_1823_),
    .B1(net855),
    .B2(net811),
    .A2(net857),
    .A1(net806),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _5038_ (.A(_1820_),
    .B(_1821_),
    .C(_1823_),
    .X(_1824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5039_ (.B1(_1820_),
    .VDD(VPWR),
    .Y(_1825_),
    .VSS(VGND),
    .A1(_1821_),
    .A2(_1823_));
 sg13g2_and3_1 _5040_ (.X(_1826_),
    .A(_1819_),
    .B(_1824_),
    .C(_1825_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5041_ (.B(_1824_),
    .C(_1825_),
    .A(_1819_),
    .Y(_1827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5042_ (.A2(_1825_),
    .A1(_1824_),
    .B1(_1819_),
    .X(_1828_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5043_ (.B(_1827_),
    .C(_1828_),
    .A(_1818_),
    .Y(_1829_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5044_ (.A2(_1828_),
    .A1(_1827_),
    .B1(_1818_),
    .X(_1830_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5045_ (.B(_1829_),
    .C(_1830_),
    .A(_1812_),
    .Y(_1831_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5046_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1829_),
    .A2(_1830_),
    .Y(_1832_),
    .B1(_1812_));
 sg13g2_a21o_1 _5047_ (.A2(_1830_),
    .A1(_1829_),
    .B1(_1812_),
    .X(_1833_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5048_ (.Y(_1834_),
    .A(_1831_),
    .B(_1833_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5049_ (.Y(_1835_),
    .A(_1811_),
    .B(_1834_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5050_ (.A(_1835_),
    .B_N(_1807_),
    .Y(_1836_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5051_ (.Y(_1837_),
    .A(_1807_),
    .B(_1835_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5052_ (.B1(_1804_),
    .VDD(VPWR),
    .Y(_1838_),
    .VSS(VGND),
    .A1(_1779_),
    .A2(_1805_));
 sg13g2_xor2_1 _5053_ (.B(_1838_),
    .A(_1837_),
    .X(_0156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5054_ (.B1(_1831_),
    .VDD(VPWR),
    .Y(_1839_),
    .VSS(VGND),
    .A1(_1811_),
    .A2(_1832_));
 sg13g2_o21ai_1 _5055_ (.B1(_1817_),
    .VDD(VPWR),
    .Y(_1840_),
    .VSS(VGND),
    .A1(_1782_),
    .A2(_1815_));
 sg13g2_a22oi_1 _5056_ (.Y(_1841_),
    .B1(net792),
    .B2(net868),
    .A2(net795),
    .A1(net866),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _5057_ (.B(net866),
    .C(net795),
    .A(net868),
    .Y(_1842_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net792));
 sg13g2_nor2b_1 _5058_ (.A(_1841_),
    .B_N(_1842_),
    .Y(_1843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5059_ (.Y(_1844_),
    .A(_1840_),
    .B(_1843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5060_ (.Y(_1845_),
    .A(_1840_),
    .B(_1843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5061_ (.A2(_1828_),
    .A1(_1818_),
    .B1(_1826_),
    .X(_1846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5062_ (.Y(_1847_),
    .A(net863),
    .B(net798),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5063_ (.Y(_1848_),
    .A(net858),
    .B(net800),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5064_ (.Y(_1849_),
    .A(net802),
    .B(net858),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5065_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1850_),
    .B(_1848_),
    .A(_1815_));
 sg13g2_and2_1 _5066_ (.A(_1814_),
    .B(_1849_),
    .X(_1851_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5067_ (.Y(_1852_),
    .A(_1814_),
    .B(_1849_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5068_ (.Y(_1853_),
    .A(_1847_),
    .B(_1852_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5069_ (.B1(_1822_),
    .VDD(VPWR),
    .Y(_1854_),
    .VSS(VGND),
    .A1(_1820_),
    .A2(_1823_));
 sg13g2_nand2_1 _5070_ (.Y(_1855_),
    .A(net804),
    .B(net856),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _5071_ (.A(net813),
    .B(net806),
    .C(net855),
    .D(net853),
    .X(_1856_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _5072_ (.B(net806),
    .C(net855),
    .A(net813),
    .Y(_1857_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net853));
 sg13g2_a22oi_1 _5073_ (.Y(_1858_),
    .B1(net853),
    .B2(net813),
    .A2(net855),
    .A1(net806),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _5074_ (.A(_1855_),
    .B(_1856_),
    .C(_1858_),
    .X(_1859_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5075_ (.B1(_1855_),
    .VDD(VPWR),
    .Y(_1860_),
    .VSS(VGND),
    .A1(_1856_),
    .A2(_1858_));
 sg13g2_and3_1 _5076_ (.X(_1861_),
    .A(_1854_),
    .B(_1859_),
    .C(_1860_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5077_ (.B(_1859_),
    .C(_1860_),
    .A(_1854_),
    .Y(_1862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5078_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1859_),
    .A2(_1860_),
    .Y(_1863_),
    .B1(_1854_));
 sg13g2_or3_1 _5079_ (.A(_1853_),
    .B(_1861_),
    .C(_1863_),
    .X(_1864_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5080_ (.B1(_1853_),
    .VDD(VPWR),
    .Y(_1865_),
    .VSS(VGND),
    .A1(_1861_),
    .A2(_1863_));
 sg13g2_and3_1 _5081_ (.X(_1866_),
    .A(_1846_),
    .B(_1864_),
    .C(_1865_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5082_ (.B(_1864_),
    .C(_1865_),
    .A(_1846_),
    .Y(_1867_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5083_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1864_),
    .A2(_1865_),
    .Y(_1868_),
    .B1(_1846_));
 sg13g2_or3_1 _5084_ (.A(_1845_),
    .B(_1866_),
    .C(_1868_),
    .X(_1869_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5085_ (.B1(_1845_),
    .VDD(VPWR),
    .Y(_1870_),
    .VSS(VGND),
    .A1(_1866_),
    .A2(_1868_));
 sg13g2_nand3_1 _5086_ (.B(_1869_),
    .C(_1870_),
    .A(_1839_),
    .Y(_1871_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5087_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1869_),
    .A2(_1870_),
    .Y(_1872_),
    .B1(_1839_));
 sg13g2_a21o_1 _5088_ (.A2(_1870_),
    .A1(_1869_),
    .B1(_1839_),
    .X(_1873_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5089_ (.Y(_1874_),
    .A(_1871_),
    .B(_1873_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5090_ (.B(_1874_),
    .A(_1810_),
    .X(_1875_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _5091_ (.A2(_1838_),
    .A1(_1837_),
    .B1(_1836_),
    .X(_1876_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5092_ (.Y(_1877_),
    .A(_1875_),
    .B(_1876_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5093_ (.B(_1876_),
    .A(_1875_),
    .X(_0157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5094_ (.B1(_1867_),
    .VDD(VPWR),
    .Y(_1878_),
    .VSS(VGND),
    .A1(_1845_),
    .A2(_1868_));
 sg13g2_o21ai_1 _5095_ (.B1(_1850_),
    .VDD(VPWR),
    .Y(_1879_),
    .VSS(VGND),
    .A1(_1847_),
    .A2(_1851_));
 sg13g2_nand2_1 _5096_ (.Y(_1880_),
    .A(net868),
    .B(net1021),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5097_ (.Y(_1881_),
    .A(net863),
    .B(net792),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _5098_ (.A(net866),
    .B(net863),
    .C(net795),
    .D(net792),
    .X(_1882_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5099_ (.Y(_1883_),
    .B1(net792),
    .B2(net866),
    .A2(net795),
    .A1(net863),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5100_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1884_),
    .B(_1883_),
    .A(_1882_));
 sg13g2_nor2_1 _5101_ (.A(_1880_),
    .B(_1884_),
    .Y(_1885_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5102_ (.B(_1884_),
    .A(_1880_),
    .X(_1886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5103_ (.Y(_1887_),
    .A(_1879_),
    .B(_1886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5104_ (.Y(_1888_),
    .A(_1879_),
    .B(_1886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5105_ (.Y(_1889_),
    .A(_1842_),
    .B(_1888_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5106_ (.B1(_1862_),
    .VDD(VPWR),
    .Y(_1890_),
    .VSS(VGND),
    .A1(_1853_),
    .A2(_1863_));
 sg13g2_nand2_1 _5107_ (.Y(_1891_),
    .A(net860),
    .B(net798),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _5108_ (.Y(_1892_),
    .A(net800),
    .B(net856),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5109_ (.Y(_1893_),
    .A(net802),
    .B(net856),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5110_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1894_),
    .B(_1892_),
    .A(_1849_));
 sg13g2_xnor2_1 _5111_ (.Y(_1895_),
    .A(_1848_),
    .B(_1893_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5112_ (.Y(_1896_),
    .A(_1891_),
    .B(_1895_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5113_ (.B1(_1857_),
    .VDD(VPWR),
    .Y(_1897_),
    .VSS(VGND),
    .A1(_1855_),
    .A2(_1858_));
 sg13g2_nand2_1 _5114_ (.Y(_1898_),
    .A(net804),
    .B(net854),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _5115_ (.A(net813),
    .B(net807),
    .C(net851),
    .D(net1024),
    .X(_1899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _5116_ (.B(net806),
    .C(net851),
    .A(net813),
    .Y(_1900_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net1024));
 sg13g2_a22oi_1 _5117_ (.Y(_1901_),
    .B1(net1025),
    .B2(net813),
    .A2(net853),
    .A1(net807),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _5118_ (.A(_1898_),
    .B(_1899_),
    .C(_1901_),
    .X(_1902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5119_ (.B1(_1898_),
    .VDD(VPWR),
    .Y(_1903_),
    .VSS(VGND),
    .A1(_1899_),
    .A2(_1901_));
 sg13g2_and3_1 _5120_ (.X(_1904_),
    .A(_1897_),
    .B(_1902_),
    .C(_1903_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5121_ (.B(_1902_),
    .C(_1903_),
    .A(_1897_),
    .Y(_1905_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5122_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1902_),
    .A2(_1903_),
    .Y(_1906_),
    .B1(_1897_));
 sg13g2_or3_1 _5123_ (.A(_1896_),
    .B(_1904_),
    .C(_1906_),
    .X(_1907_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5124_ (.B1(_1896_),
    .VDD(VPWR),
    .Y(_1908_),
    .VSS(VGND),
    .A1(_1904_),
    .A2(_1906_));
 sg13g2_and3_1 _5125_ (.X(_1909_),
    .A(_1890_),
    .B(_1907_),
    .C(_1908_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5126_ (.B(_1907_),
    .C(_1908_),
    .A(_1890_),
    .Y(_1910_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5127_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1907_),
    .A2(_1908_),
    .Y(_1911_),
    .B1(_1890_));
 sg13g2_or3_1 _5128_ (.A(_1889_),
    .B(_1909_),
    .C(_1911_),
    .X(_1912_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5129_ (.B1(_1889_),
    .VDD(VPWR),
    .Y(_1913_),
    .VSS(VGND),
    .A1(_1909_),
    .A2(_1911_));
 sg13g2_and3_1 _5130_ (.X(_1914_),
    .A(_1878_),
    .B(_1912_),
    .C(_1913_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5131_ (.B(_1912_),
    .C(_1913_),
    .A(_1878_),
    .Y(_1915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5132_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1912_),
    .A2(_1913_),
    .Y(_1916_),
    .B1(_1878_));
 sg13g2_or3_1 _5133_ (.A(_1844_),
    .B(_1914_),
    .C(_1916_),
    .X(_1917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5134_ (.B1(_1844_),
    .VDD(VPWR),
    .Y(_1918_),
    .VSS(VGND),
    .A1(_1914_),
    .A2(_1916_));
 sg13g2_o21ai_1 _5135_ (.B1(_1871_),
    .VDD(VPWR),
    .Y(_1919_),
    .VSS(VGND),
    .A1(_1810_),
    .A2(_1872_));
 sg13g2_nand3_1 _5136_ (.B(_1918_),
    .C(_1919_),
    .A(_1917_),
    .Y(_1920_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5137_ (.A2(_1918_),
    .A1(_1917_),
    .B1(_1919_),
    .X(_1921_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5138_ (.Y(_1922_),
    .A(_1920_),
    .B(_1921_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _5139_ (.A(_1875_),
    .B(_1876_),
    .C(_1920_),
    .D(_1921_),
    .X(_1923_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5140_ (.B(_1922_),
    .A(_1877_),
    .X(_0158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5141_ (.B1(_1920_),
    .VDD(VPWR),
    .Y(_1924_),
    .VSS(VGND),
    .A1(_1877_),
    .A2(_1922_));
 sg13g2_o21ai_1 _5142_ (.B1(_1915_),
    .VDD(VPWR),
    .Y(_1925_),
    .VSS(VGND),
    .A1(_1844_),
    .A2(_1916_));
 sg13g2_o21ai_1 _5143_ (.B1(_1887_),
    .VDD(VPWR),
    .Y(_1926_),
    .VSS(VGND),
    .A1(_1842_),
    .A2(_1888_));
 sg13g2_o21ai_1 _5144_ (.B1(_1910_),
    .VDD(VPWR),
    .Y(_1927_),
    .VSS(VGND),
    .A1(_1889_),
    .A2(_1911_));
 sg13g2_nor2_1 _5145_ (.A(_1882_),
    .B(_1885_),
    .Y(_1928_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5146_ (.B1(_1894_),
    .VDD(VPWR),
    .Y(_1929_),
    .VSS(VGND),
    .A1(_1891_),
    .A2(_1895_));
 sg13g2_nand2_1 _5147_ (.Y(_1930_),
    .A(net866),
    .B(net1021),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5148_ (.Y(_1931_),
    .A(net860),
    .B(net793),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5149_ (.Y(_1932_),
    .A(net860),
    .B(net795),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5150_ (.B(_1932_),
    .A(_1881_),
    .X(_1933_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5151_ (.Y(_1934_),
    .B(_1933_),
    .A_N(_1930_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5152_ (.Y(_1935_),
    .A(_1930_),
    .B(_1933_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5153_ (.Y(_1936_),
    .A(_1929_),
    .B(_1935_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5154_ (.A(_1928_),
    .B(_1936_),
    .Y(_1937_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5155_ (.Y(_1938_),
    .A(_1928_),
    .B(_1936_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5156_ (.B1(_1905_),
    .VDD(VPWR),
    .Y(_1939_),
    .VSS(VGND),
    .A1(_1896_),
    .A2(_1906_));
 sg13g2_nand2_1 _5157_ (.Y(_1940_),
    .A(net858),
    .B(net798),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5158_ (.Y(_1941_),
    .A(net802),
    .B(net854),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5159_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1942_),
    .B(_1941_),
    .A(_1892_));
 sg13g2_and2_1 _5160_ (.A(_1892_),
    .B(_1941_),
    .X(_1943_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5161_ (.Y(_1944_),
    .A(_1892_),
    .B(_1941_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5162_ (.Y(_1945_),
    .A(_1940_),
    .B(_1944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5163_ (.B1(_1900_),
    .VDD(VPWR),
    .Y(_1946_),
    .VSS(VGND),
    .A1(_1898_),
    .A2(_1901_));
 sg13g2_nand2_1 _5164_ (.Y(_1947_),
    .A(net804),
    .B(net1025),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _5165_ (.A(net807),
    .B(net804),
    .C(net851),
    .D(net1025),
    .X(_1948_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5166_ (.Y(_1949_),
    .B1(net1025),
    .B2(net806),
    .A2(net851),
    .A1(net804),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5167_ (.A(_1948_),
    .B(_1949_),
    .Y(_1950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5168_ (.Y(_1951_),
    .A(_1946_),
    .B(_1950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5169_ (.Y(_1952_),
    .A(_1946_),
    .B(_1950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5170_ (.B(_1952_),
    .A(_1945_),
    .X(_1953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5171_ (.Y(_1954_),
    .A(_1939_),
    .B(_1953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5172_ (.Y(_1955_),
    .A(_1939_),
    .B(_1953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5173_ (.B(_1955_),
    .A(_1938_),
    .X(_1956_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5174_ (.Y(_1957_),
    .A(_1927_),
    .B(_1956_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5175_ (.Y(_1958_),
    .A(_1927_),
    .B(_1956_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5176_ (.Y(_1959_),
    .B(_1926_),
    .A_N(_1958_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5177_ (.Y(_1960_),
    .A(_1926_),
    .B(_1958_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5178_ (.A(_1925_),
    .B(_1960_),
    .Y(_1961_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5179_ (.Y(_1962_),
    .A(_1925_),
    .B(_1960_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5180_ (.A(_1961_),
    .B_N(_1962_),
    .Y(_1963_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5181_ (.B(_1963_),
    .A(_1924_),
    .X(_0159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5182_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1929_),
    .A2(_1935_),
    .Y(_1964_),
    .B1(_1937_));
 sg13g2_o21ai_1 _5183_ (.B1(_1954_),
    .VDD(VPWR),
    .Y(_1965_),
    .VSS(VGND),
    .A1(_1938_),
    .A2(_1955_));
 sg13g2_o21ai_1 _5184_ (.B1(_1934_),
    .VDD(VPWR),
    .Y(_1966_),
    .VSS(VGND),
    .A1(_1881_),
    .A2(_1932_));
 sg13g2_o21ai_1 _5185_ (.B1(_1942_),
    .VDD(VPWR),
    .Y(_1967_),
    .VSS(VGND),
    .A1(_1940_),
    .A2(_1943_));
 sg13g2_nand2_1 _5186_ (.Y(_1968_),
    .A(net863),
    .B(net1021),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5187_ (.Y(_1969_),
    .A(net858),
    .B(net793),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5188_ (.Y(_1970_),
    .A(net858),
    .B(net795),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5189_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1971_),
    .B(_1969_),
    .A(_1932_));
 sg13g2_xnor2_1 _5190_ (.Y(_1972_),
    .A(_1931_),
    .B(_1970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5191_ (.B(_1972_),
    .A(_1968_),
    .X(_1973_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5192_ (.Y(_1974_),
    .A(_1967_),
    .B(_1973_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5193_ (.A(_1974_),
    .B_N(_1966_),
    .Y(_1975_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5194_ (.B(_1974_),
    .A(_1966_),
    .X(_1976_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5195_ (.B1(_1951_),
    .VDD(VPWR),
    .Y(_1977_),
    .VSS(VGND),
    .A1(_1945_),
    .A2(_1952_));
 sg13g2_a21oi_1 _5196_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net807),
    .A2(net851),
    .Y(_1978_),
    .B1(_1947_));
 sg13g2_nand2_1 _5197_ (.Y(_1979_),
    .A(net857),
    .B(net798),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5198_ (.Y(_1980_),
    .A(net800),
    .B(net852),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _5199_ (.A(net802),
    .B(net801),
    .C(net854),
    .D(net851),
    .X(_1981_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5200_ (.Y(_1982_),
    .B1(net851),
    .B2(net803),
    .A2(net854),
    .A1(net801),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5201_ (.A(_1979_),
    .B(_1981_),
    .C(_1982_),
    .Y(_1983_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5202_ (.B1(_1979_),
    .VDD(VPWR),
    .Y(_1984_),
    .VSS(VGND),
    .A1(_1981_),
    .A2(_1982_));
 sg13g2_nor2b_1 _5203_ (.A(_1983_),
    .B_N(_1984_),
    .Y(_1985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5204_ (.Y(_1986_),
    .A(_1978_),
    .B(_1985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5205_ (.Y(_1987_),
    .B(_1977_),
    .A_N(_1986_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5206_ (.B(_1986_),
    .A(_1977_),
    .X(_1988_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5207_ (.B(_1988_),
    .A(_1976_),
    .X(_1989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5208_ (.Y(_1990_),
    .A(_1965_),
    .B(_1989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5209_ (.B(_1989_),
    .A(_1965_),
    .X(_1991_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5210_ (.Y(_1992_),
    .B(_1991_),
    .A_N(_1964_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5211_ (.B(_1991_),
    .A(_1964_),
    .X(_1993_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5212_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1957_),
    .A2(_1959_),
    .Y(_1994_),
    .B1(_1993_));
 sg13g2_nand3_1 _5213_ (.B(_1959_),
    .C(_1993_),
    .A(_1957_),
    .Y(_1995_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5214_ (.Y(_1996_),
    .B(_1995_),
    .A_N(_1994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5215_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1920_),
    .A2(_1962_),
    .Y(_1997_),
    .B1(_1961_));
 sg13g2_a21oi_2 _5216_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_1997_),
    .Y(_1998_),
    .A2(_1963_),
    .A1(_1923_));
 sg13g2_nor2_1 _5217_ (.A(_1996_),
    .B(_1998_),
    .Y(_1999_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5218_ (.B(_1998_),
    .A(_1996_),
    .X(_0150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5219_ (.A2(_1973_),
    .A1(_1967_),
    .B1(_1975_),
    .X(_2000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5220_ (.B1(_1987_),
    .VDD(VPWR),
    .Y(_2001_),
    .VSS(VGND),
    .A1(_1976_),
    .A2(_1988_));
 sg13g2_a21o_2 _5221_ (.A2(_1985_),
    .A1(_1978_),
    .B1(_1948_),
    .X(_2002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5222_ (.Y(_2003_),
    .A(net798),
    .B(net854),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5223_ (.Y(_2004_),
    .A(net803),
    .B(net1024),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5224_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2005_),
    .B(_2004_),
    .A(_1980_));
 sg13g2_xnor2_1 _5225_ (.Y(_2006_),
    .A(_1980_),
    .B(_2004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5226_ (.B(_2006_),
    .A(_2003_),
    .X(_2007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5227_ (.A(_2002_),
    .B(_2007_),
    .X(_2008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5228_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2009_),
    .B(_2007_),
    .A(_2002_));
 sg13g2_xnor2_1 _5229_ (.Y(_2010_),
    .A(_2002_),
    .B(_2007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5230_ (.B1(_1971_),
    .VDD(VPWR),
    .Y(_2011_),
    .VSS(VGND),
    .A1(_1968_),
    .A2(_1972_));
 sg13g2_or2_1 _5231_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2012_),
    .B(_1983_),
    .A(_1981_));
 sg13g2_nand2_1 _5232_ (.Y(_2013_),
    .A(net860),
    .B(net1021),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5233_ (.Y(_2014_),
    .A(net856),
    .B(net795),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5234_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2015_),
    .B(_2014_),
    .A(_1969_));
 sg13g2_xnor2_1 _5235_ (.Y(_2016_),
    .A(_1969_),
    .B(_2014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5236_ (.B(_2016_),
    .A(_2013_),
    .X(_2017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5237_ (.Y(_2018_),
    .A(_2012_),
    .B(_2017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5238_ (.A(_2018_),
    .B_N(_2011_),
    .Y(_2019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5239_ (.Y(_2020_),
    .A(_2011_),
    .B(_2018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5240_ (.Y(_2021_),
    .A(_2010_),
    .B(_2020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5241_ (.Y(_2022_),
    .A(_2001_),
    .B(_2021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5242_ (.A(_2022_),
    .B_N(_2000_),
    .Y(_2023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5243_ (.B(_2022_),
    .A(_2000_),
    .X(_2024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5244_ (.B(_1992_),
    .C(_2024_),
    .A(_1990_),
    .Y(_2025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5245_ (.VDD(VPWR),
    .Y(_2026_),
    .A(_2025_),
    .VSS(VGND));
 sg13g2_a21oi_1 _5246_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1990_),
    .A2(_1992_),
    .Y(_2027_),
    .B1(_2024_));
 sg13g2_nor2_1 _5247_ (.A(_2026_),
    .B(_2027_),
    .Y(_2028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5248_ (.A(_1994_),
    .B(_1999_),
    .Y(_2029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5249_ (.Y(_0151_),
    .A(_2028_),
    .B(_2029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5250_ (.A2(_2017_),
    .A1(_2012_),
    .B1(_2019_),
    .X(_2030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5251_ (.Y(_2031_),
    .B1(net1024),
    .B2(net801),
    .A2(net852),
    .A1(net798),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _5252_ (.Y(_2032_),
    .A(net799),
    .B(net1024),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5253_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2033_),
    .B(_2032_),
    .A(_1980_));
 sg13g2_nand2b_1 _5254_ (.Y(_2034_),
    .B(_2033_),
    .A_N(_2031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5255_ (.B1(_2015_),
    .VDD(VPWR),
    .Y(_2035_),
    .VSS(VGND),
    .A1(_2013_),
    .A2(_2016_));
 sg13g2_o21ai_1 _5256_ (.B1(_2005_),
    .VDD(VPWR),
    .Y(_2036_),
    .VSS(VGND),
    .A1(_2003_),
    .A2(_2006_));
 sg13g2_nand2_1 _5257_ (.Y(_2037_),
    .A(net858),
    .B(net1021),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5258_ (.Y(_2038_),
    .A(net854),
    .B(net792),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _5259_ (.A(net856),
    .B(net854),
    .C(net796),
    .D(net793),
    .X(_2039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5260_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2040_),
    .B(_2038_),
    .A(_2014_));
 sg13g2_a22oi_1 _5261_ (.Y(_2041_),
    .B1(net793),
    .B2(net857),
    .A2(net796),
    .A1(net855),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5262_ (.A(_2039_),
    .B(_2041_),
    .Y(_2042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5263_ (.Y(_2043_),
    .A(_2037_),
    .B(_2042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5264_ (.Y(_2044_),
    .A(_2036_),
    .B(_2043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5265_ (.A(_2044_),
    .B_N(_2035_),
    .Y(_2045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5266_ (.B(_2044_),
    .A(_2035_),
    .X(_2046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5267_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2047_),
    .B(_2046_),
    .A(_2034_));
 sg13g2_xor2_1 _5268_ (.B(_2046_),
    .A(_2034_),
    .X(_2048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5269_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2009_),
    .A2(_2020_),
    .Y(_2049_),
    .B1(_2008_));
 sg13g2_nor2b_1 _5270_ (.A(_2049_),
    .B_N(_2048_),
    .Y(_2050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5271_ (.B(_2049_),
    .A(_2048_),
    .X(_2051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5272_ (.A(_2051_),
    .B_N(_2030_),
    .Y(_2052_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5273_ (.B(_2051_),
    .A(_2030_),
    .X(_2053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5274_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2001_),
    .A2(_2021_),
    .Y(_2054_),
    .B1(_2023_));
 sg13g2_nor2_1 _5275_ (.A(_2053_),
    .B(_2054_),
    .Y(_2055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5276_ (.B(_2054_),
    .A(_2053_),
    .X(_2056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5277_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1994_),
    .A2(_2025_),
    .Y(_2057_),
    .B1(_2027_));
 sg13g2_a21oi_1 _5278_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1995_),
    .A2(_2025_),
    .Y(_2058_),
    .B1(_2027_));
 sg13g2_a21oi_2 _5279_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_2058_),
    .Y(_2059_),
    .A2(_2057_),
    .A1(_1998_));
 sg13g2_xor2_1 _5280_ (.B(_2059_),
    .A(_2056_),
    .X(_0152_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5281_ (.A2(_2043_),
    .A1(_2036_),
    .B1(_2045_),
    .X(_2060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5282_ (.B1(_2040_),
    .VDD(VPWR),
    .Y(_2061_),
    .VSS(VGND),
    .A1(_2037_),
    .A2(_2041_));
 sg13g2_nand2_1 _5283_ (.Y(_2062_),
    .A(net856),
    .B(net1021),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5284_ (.Y(_2063_),
    .A(net851),
    .B(net792),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5285_ (.Y(_2064_),
    .A(net796),
    .B(net852),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5286_ (.B(_2064_),
    .A(_2038_),
    .X(_2065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5287_ (.Y(_2066_),
    .B(_2065_),
    .A_N(_2062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5288_ (.Y(_2067_),
    .A(_2062_),
    .B(_2065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5289_ (.A(_2033_),
    .B_N(_2067_),
    .Y(_2068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5290_ (.Y(_2069_),
    .A(_2033_),
    .B(_2067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5291_ (.Y(_2070_),
    .A(_2061_),
    .B(_2069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5292_ (.A(_2032_),
    .B(_2070_),
    .Y(_2071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5293_ (.Y(_2072_),
    .A(_2032_),
    .B(_2070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5294_ (.A(_2047_),
    .B(_2072_),
    .Y(_2073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5295_ (.B(_2072_),
    .A(_2047_),
    .X(_2074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5296_ (.B(_2074_),
    .A(_2060_),
    .X(_2075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5297_ (.B1(_2075_),
    .VDD(VPWR),
    .Y(_2076_),
    .VSS(VGND),
    .A1(_2050_),
    .A2(_2052_));
 sg13g2_or3_1 _5298_ (.A(_2050_),
    .B(_2052_),
    .C(_2075_),
    .X(_2077_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5299_ (.A(_2076_),
    .B(_2077_),
    .X(_2078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5300_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2056_),
    .A2(_2059_),
    .Y(_2079_),
    .B1(_2055_));
 sg13g2_xnor2_1 _5301_ (.Y(_0153_),
    .A(_2078_),
    .B(_2079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5302_ (.Y(_2080_),
    .A(_2056_),
    .B(_2078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5303_ (.VDD(VPWR),
    .Y(_2081_),
    .A(_2080_),
    .VSS(VGND));
 sg13g2_o21ai_1 _5304_ (.B1(_2076_),
    .VDD(VPWR),
    .Y(_2082_),
    .VSS(VGND),
    .A1(_2053_),
    .A2(_2054_));
 sg13g2_a22oi_1 _5305_ (.Y(_2083_),
    .B1(_2082_),
    .B2(_2077_),
    .A2(_2081_),
    .A1(_2059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5306_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2060_),
    .A2(_2074_),
    .Y(_2084_),
    .B1(_2073_));
 sg13g2_a21o_1 _5307_ (.A2(_2069_),
    .A1(_2061_),
    .B1(_2068_),
    .X(_2085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5308_ (.B1(_2066_),
    .VDD(VPWR),
    .Y(_2086_),
    .VSS(VGND),
    .A1(_2038_),
    .A2(_2064_));
 sg13g2_nand2_1 _5309_ (.Y(_2087_),
    .A(net854),
    .B(net1021),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5310_ (.Y(_2088_),
    .A(net792),
    .B(net1024),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5311_ (.Y(_2089_),
    .A(net796),
    .B(net1024),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5312_ (.B(_2089_),
    .A(_2063_),
    .X(_2090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5313_ (.Y(_2091_),
    .B(_2090_),
    .A_N(_2087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5314_ (.Y(_2092_),
    .A(_2087_),
    .B(_2090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5315_ (.Y(_2093_),
    .A(_2086_),
    .B(_2092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5316_ (.B(_2092_),
    .A(_2086_),
    .X(_2094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5317_ (.Y(_2095_),
    .A(_2071_),
    .B(_2094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5318_ (.A(_2095_),
    .B_N(_2085_),
    .Y(_2096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5319_ (.B(_2095_),
    .A(_2085_),
    .X(_2097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5320_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2098_),
    .B(_2097_),
    .A(_2084_));
 sg13g2_xor2_1 _5321_ (.B(_2097_),
    .A(_2084_),
    .X(_2099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5322_ (.VDD(VPWR),
    .Y(_2100_),
    .A(_2099_),
    .VSS(VGND));
 sg13g2_xnor2_1 _5323_ (.Y(_0154_),
    .A(_2083_),
    .B(_2099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5324_ (.B1(_2098_),
    .VDD(VPWR),
    .Y(_2101_),
    .VSS(VGND),
    .A1(_2083_),
    .A2(_2100_));
 sg13g2_a21oi_1 _5325_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2071_),
    .A2(_2094_),
    .Y(_2102_),
    .B1(_2096_));
 sg13g2_o21ai_1 _5326_ (.B1(_2091_),
    .VDD(VPWR),
    .Y(_2103_),
    .VSS(VGND),
    .A1(_2063_),
    .A2(_2089_));
 sg13g2_nand2_1 _5327_ (.Y(_2104_),
    .A(net852),
    .B(net1021),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5328_ (.B(_2104_),
    .A(_2088_),
    .X(_2105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5329_ (.Y(_2106_),
    .A(_2103_),
    .B(_2105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5330_ (.Y(_2107_),
    .A(_2093_),
    .B(_2106_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5331_ (.Y(_2108_),
    .A(_2102_),
    .B(_2107_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5332_ (.Y(_0155_),
    .A(_2101_),
    .B(_2108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5333_ (.Y(_2109_),
    .A(net356),
    .B(net286),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5334_ (.Y(_2110_),
    .A(\mac1.sum_lvl2_ff[20] ),
    .B(\mac1.sum_lvl2_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5335_ (.A(\mac1.sum_lvl2_ff[20] ),
    .B(\mac1.sum_lvl2_ff[1] ),
    .Y(_2111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5336_ (.B(\mac1.sum_lvl2_ff[1] ),
    .A(\mac1.sum_lvl2_ff[20] ),
    .X(_2112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5337_ (.Y(_0007_),
    .A(_2109_),
    .B(_2112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5338_ (.B1(_2110_),
    .VDD(VPWR),
    .Y(_2113_),
    .VSS(VGND),
    .A1(_2109_),
    .A2(_2111_));
 sg13g2_and2_1 _5339_ (.A(\mac1.sum_lvl2_ff[21] ),
    .B(\mac1.sum_lvl2_ff[2] ),
    .X(_2114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5340_ (.B(net380),
    .A(\mac1.sum_lvl2_ff[21] ),
    .X(_2115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5341_ (.B(net381),
    .A(_2113_),
    .X(_0008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5342_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2113_),
    .A2(_2115_),
    .Y(_2116_),
    .B1(_2114_));
 sg13g2_nand2_1 _5343_ (.Y(_2117_),
    .A(\mac1.sum_lvl2_ff[22] ),
    .B(net370),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5344_ (.Y(_2118_),
    .A(\mac1.sum_lvl2_ff[22] ),
    .B(net370),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5345_ (.B(net371),
    .A(_2116_),
    .X(_0009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5346_ (.B1(_2117_),
    .VDD(VPWR),
    .Y(_2119_),
    .VSS(VGND),
    .A1(_2116_),
    .A2(_2118_));
 sg13g2_and2_1 _5347_ (.A(\mac1.sum_lvl2_ff[23] ),
    .B(\mac1.sum_lvl2_ff[4] ),
    .X(_2120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5348_ (.B(net512),
    .A(\mac1.sum_lvl2_ff[23] ),
    .X(_2121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5349_ (.B(net513),
    .A(_2119_),
    .X(_0010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5350_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2119_),
    .A2(_2121_),
    .Y(_2122_),
    .B1(_2120_));
 sg13g2_nor2_1 _5351_ (.A(net505),
    .B(\mac1.sum_lvl2_ff[5] ),
    .Y(_2123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5352_ (.B(\mac1.sum_lvl2_ff[5] ),
    .A(net505),
    .X(_2124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5353_ (.Y(_0011_),
    .A(_2122_),
    .B(net506),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5354_ (.A(\mac1.sum_lvl2_ff[25] ),
    .B(net508),
    .X(_2125_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5355_ (.Y(_2126_),
    .A(\mac1.sum_lvl2_ff[25] ),
    .B(net508),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5356_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2121_),
    .C1(_2120_),
    .B1(_2119_),
    .A1(\mac1.sum_lvl2_ff[24] ),
    .Y(_2127_),
    .A2(\mac1.sum_lvl2_ff[5] ));
 sg13g2_nor3_1 _5357_ (.A(_2123_),
    .B(net509),
    .C(_2127_),
    .Y(_2128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5358_ (.B1(net509),
    .VDD(VPWR),
    .Y(_2129_),
    .VSS(VGND),
    .A1(_2123_),
    .A2(_2127_));
 sg13g2_nor2b_2 _5359_ (.A(_2128_),
    .B_N(net510),
    .Y(_0012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5360_ (.Y(_2130_),
    .A(\mac1.sum_lvl2_ff[26] ),
    .B(\mac1.sum_lvl2_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5361_ (.B(net529),
    .A(\mac1.sum_lvl2_ff[26] ),
    .X(_2131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5362_ (.B1(net530),
    .VDD(VPWR),
    .Y(_2132_),
    .VSS(VGND),
    .A1(_2125_),
    .A2(_2128_));
 sg13g2_or3_1 _5363_ (.A(_2125_),
    .B(_2128_),
    .C(net530),
    .X(_2133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5364_ (.A(_2132_),
    .B(net531),
    .X(_0013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5365_ (.Y(_2134_),
    .A(\mac1.sum_lvl2_ff[27] ),
    .B(net375),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5366_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2130_),
    .A2(_2132_),
    .Y(_2135_),
    .B1(net376));
 sg13g2_nand3_1 _5367_ (.B(_2132_),
    .C(net376),
    .A(_2130_),
    .Y(_2136_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5368_ (.A(net377),
    .B_N(_2136_),
    .Y(_0014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5369_ (.A2(net375),
    .A1(\mac1.sum_lvl2_ff[27] ),
    .B1(net377),
    .X(_2137_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5370_ (.A(\mac1.sum_lvl2_ff[28] ),
    .B(net434),
    .X(_2138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5371_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2139_),
    .B(net434),
    .A(\mac1.sum_lvl2_ff[28] ));
 sg13g2_nand2b_1 _5372_ (.Y(_2140_),
    .B(net435),
    .A_N(_2138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5373_ (.Y(_0015_),
    .A(_2137_),
    .B(net436),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5374_ (.Y(_2141_),
    .A(\mac1.sum_lvl2_ff[29] ),
    .B(\mac1.sum_lvl2_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5375_ (.B(\mac1.sum_lvl2_ff[10] ),
    .A(\mac1.sum_lvl2_ff[29] ),
    .X(_2142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5376_ (.VDD(VPWR),
    .Y(_2143_),
    .A(_2142_),
    .VSS(VGND));
 sg13g2_a21o_2 _5377_ (.A2(_2139_),
    .A1(_2137_),
    .B1(_2138_),
    .X(_2144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5378_ (.Y(_2145_),
    .A(_2142_),
    .B(_2144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5379_ (.Y(_0001_),
    .A(_2143_),
    .B(_2144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5380_ (.A(\mac1.sum_lvl2_ff[30] ),
    .B(\mac1.sum_lvl2_ff[11] ),
    .Y(_2146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5381_ (.Y(_2147_),
    .A(\mac1.sum_lvl2_ff[30] ),
    .B(\mac1.sum_lvl2_ff[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5382_ (.Y(_2148_),
    .A(_2141_),
    .B(_2145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5383_ (.Y(_0002_),
    .A(_2147_),
    .B(_2148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5384_ (.Y(_2149_),
    .A(net546),
    .B(net481),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5385_ (.A(\mac1.sum_lvl2_ff[31] ),
    .B(\mac1.sum_lvl2_ff[12] ),
    .Y(_2150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5386_ (.B(net481),
    .A(\mac1.sum_lvl2_ff[31] ),
    .X(_2151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5387_ (.A(_2141_),
    .B(_2146_),
    .Y(_2152_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5388_ (.A(_2143_),
    .B(_2147_),
    .Y(_2153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5389_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2153_),
    .C1(_2152_),
    .B1(_2144_),
    .A1(\mac1.sum_lvl2_ff[30] ),
    .Y(_2154_),
    .A2(\mac1.sum_lvl2_ff[11] ));
 sg13g2_xnor2_1 _5390_ (.Y(_0003_),
    .A(net482),
    .B(_2154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5391_ (.B1(_2149_),
    .VDD(VPWR),
    .Y(_2155_),
    .VSS(VGND),
    .A1(_2150_),
    .A2(_2154_));
 sg13g2_and2_1 _5392_ (.A(\mac1.sum_lvl2_ff[32] ),
    .B(\mac1.sum_lvl2_ff[13] ),
    .X(_2156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5393_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2157_),
    .B(\mac1.sum_lvl2_ff[13] ),
    .A(\mac1.sum_lvl2_ff[32] ));
 sg13g2_nand2b_1 _5394_ (.Y(_2158_),
    .B(_2157_),
    .A_N(_2156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5395_ (.Y(_0004_),
    .A(_2155_),
    .B(_2158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5396_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2155_),
    .A2(_2157_),
    .Y(_2159_),
    .B1(_2156_));
 sg13g2_nand2_1 _5397_ (.Y(_2160_),
    .A(\mac1.sum_lvl2_ff[33] ),
    .B(\mac1.sum_lvl2_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5398_ (.A(\mac1.sum_lvl2_ff[33] ),
    .B(\mac1.sum_lvl2_ff[14] ),
    .Y(_2161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5399_ (.B(net460),
    .A(\mac1.sum_lvl2_ff[33] ),
    .X(_2162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5400_ (.Y(_0005_),
    .A(_2159_),
    .B(net461),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5401_ (.B1(_2160_),
    .VDD(VPWR),
    .Y(_2163_),
    .VSS(VGND),
    .A1(_2159_),
    .A2(_2161_));
 sg13g2_xnor2_1 _5402_ (.Y(_2164_),
    .A(\mac1.sum_lvl2_ff[34] ),
    .B(net390),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5403_ (.Y(_0006_),
    .A(_2163_),
    .B(net391),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5404_ (.B(net286),
    .A(\mac1.sum_lvl2_ff[19] ),
    .X(_0000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5405_ (.Y(_2165_),
    .A(net288),
    .B(net265),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5406_ (.Y(_2166_),
    .A(\mac1.sum_lvl3_ff[21] ),
    .B(\mac1.sum_lvl3_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5407_ (.A(\mac1.sum_lvl3_ff[21] ),
    .B(\mac1.sum_lvl3_ff[1] ),
    .Y(_2167_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5408_ (.B(\mac1.sum_lvl3_ff[1] ),
    .A(\mac1.sum_lvl3_ff[21] ),
    .X(_2168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5409_ (.Y(_0023_),
    .A(_2165_),
    .B(_2168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5410_ (.B1(_2166_),
    .VDD(VPWR),
    .Y(_2169_),
    .VSS(VGND),
    .A1(_2165_),
    .A2(_2167_));
 sg13g2_and2_1 _5411_ (.A(\mac1.sum_lvl3_ff[22] ),
    .B(\mac1.sum_lvl3_ff[2] ),
    .X(_2170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5412_ (.B(net454),
    .A(\mac1.sum_lvl3_ff[22] ),
    .X(_2171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5413_ (.B(net455),
    .A(_2169_),
    .X(_0024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5414_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2169_),
    .A2(_2171_),
    .Y(_2172_),
    .B1(_2170_));
 sg13g2_nand2_1 _5415_ (.Y(_2173_),
    .A(net361),
    .B(\mac1.sum_lvl3_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5416_ (.Y(_2174_),
    .A(net361),
    .B(\mac1.sum_lvl3_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5417_ (.B(net362),
    .A(_2172_),
    .X(_0025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5418_ (.B1(_2173_),
    .VDD(VPWR),
    .Y(_2175_),
    .VSS(VGND),
    .A1(_2172_),
    .A2(_2174_));
 sg13g2_and2_1 _5419_ (.A(net406),
    .B(\mac1.sum_lvl3_ff[4] ),
    .X(_2176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5420_ (.B(\mac1.sum_lvl3_ff[4] ),
    .A(net406),
    .X(_2177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5421_ (.B(net407),
    .A(_2175_),
    .X(_0026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5422_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2175_),
    .A2(_2177_),
    .Y(_2178_),
    .B1(_2176_));
 sg13g2_nor2_1 _5423_ (.A(\mac1.sum_lvl3_ff[25] ),
    .B(net320),
    .Y(_2179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5424_ (.B(net320),
    .A(\mac1.sum_lvl3_ff[25] ),
    .X(_2180_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5425_ (.Y(_0027_),
    .A(_2178_),
    .B(net321),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5426_ (.A(net533),
    .B(net501),
    .X(_2181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5427_ (.Y(_2182_),
    .A(\mac1.sum_lvl3_ff[26] ),
    .B(net501),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5428_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2177_),
    .C1(_2176_),
    .B1(_2175_),
    .A1(\mac1.sum_lvl3_ff[25] ),
    .Y(_2183_),
    .A2(net320));
 sg13g2_nor3_1 _5429_ (.A(_2179_),
    .B(net502),
    .C(_2183_),
    .Y(_2184_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5430_ (.B1(net502),
    .VDD(VPWR),
    .Y(_2185_),
    .VSS(VGND),
    .A1(_2179_),
    .A2(_2183_));
 sg13g2_nor2b_1 _5431_ (.A(_2184_),
    .B_N(net503),
    .Y(_0028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5432_ (.Y(_2186_),
    .A(net419),
    .B(\mac1.sum_lvl3_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5433_ (.B(\mac1.sum_lvl3_ff[7] ),
    .A(net419),
    .X(_2187_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5434_ (.B1(_2187_),
    .VDD(VPWR),
    .Y(_2188_),
    .VSS(VGND),
    .A1(_2181_),
    .A2(_2184_));
 sg13g2_or3_1 _5435_ (.A(_2181_),
    .B(_2184_),
    .C(_2187_),
    .X(_2189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5436_ (.A(_2188_),
    .B(_2189_),
    .X(_0029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5437_ (.A(\mac1.sum_lvl3_ff[28] ),
    .B(\mac1.sum_lvl3_ff[8] ),
    .X(_2190_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5438_ (.Y(_2191_),
    .A(\mac1.sum_lvl3_ff[28] ),
    .B(\mac1.sum_lvl3_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5439_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net420),
    .A2(_2188_),
    .Y(_2192_),
    .B1(_2191_));
 sg13g2_nand3_1 _5440_ (.B(_2188_),
    .C(_2191_),
    .A(net420),
    .Y(_2193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5441_ (.A(_2192_),
    .B_N(net421),
    .Y(_0030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5442_ (.A(_2190_),
    .B(_2192_),
    .Y(_2194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5443_ (.Y(_2195_),
    .A(net358),
    .B(\mac1.sum_lvl3_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5444_ (.B(\mac1.sum_lvl3_ff[9] ),
    .A(net358),
    .X(_2196_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5445_ (.B1(_2196_),
    .VDD(VPWR),
    .Y(_2197_),
    .VSS(VGND),
    .A1(_2190_),
    .A2(_2192_));
 sg13g2_xnor2_1 _5446_ (.Y(_0031_),
    .A(_2194_),
    .B(net359),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5447_ (.Y(_2198_),
    .A(_2195_),
    .B(_2197_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5448_ (.Y(_2199_),
    .A(net348),
    .B(net364),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5449_ (.B(\mac1.sum_lvl3_ff[10] ),
    .A(net348),
    .X(_2200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5450_ (.Y(_2201_),
    .A(_2198_),
    .B(net349),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5451_ (.B(net349),
    .A(_2198_),
    .X(_0017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5452_ (.A(\mac1.sum_lvl3_ff[31] ),
    .B(\mac1.sum_lvl3_ff[11] ),
    .Y(_2202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5453_ (.Y(_2203_),
    .A(\mac1.sum_lvl3_ff[31] ),
    .B(\mac1.sum_lvl3_ff[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5454_ (.Y(_2204_),
    .B(_2203_),
    .A_N(_2202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5455_ (.Y(_2205_),
    .A(_2199_),
    .B(_2201_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5456_ (.Y(_0018_),
    .A(_2204_),
    .B(_2205_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5457_ (.Y(_2206_),
    .A(\mac1.sum_lvl3_ff[32] ),
    .B(\mac1.sum_lvl3_ff[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5458_ (.B(\mac1.sum_lvl3_ff[12] ),
    .A(\mac1.sum_lvl3_ff[32] ),
    .X(_2207_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5459_ (.B1(_2203_),
    .VDD(VPWR),
    .Y(_2208_),
    .VSS(VGND),
    .A1(_2199_),
    .A2(_2202_));
 sg13g2_nand3b_1 _5460_ (.B(_2203_),
    .C(_2200_),
    .Y(_2209_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_2202_));
 sg13g2_a21oi_1 _5461_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2195_),
    .A2(_2197_),
    .Y(_2210_),
    .B1(_2209_));
 sg13g2_o21ai_1 _5462_ (.B1(_2207_),
    .VDD(VPWR),
    .Y(_2211_),
    .VSS(VGND),
    .A1(_2208_),
    .A2(_2210_));
 sg13g2_or3_1 _5463_ (.A(_2207_),
    .B(_2208_),
    .C(_2210_),
    .X(_2212_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5464_ (.A(_2211_),
    .B(_2212_),
    .X(_0019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5465_ (.Y(_2213_),
    .A(_2206_),
    .B(_2211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5466_ (.Y(_2214_),
    .A(\mac1.sum_lvl3_ff[33] ),
    .B(\mac1.sum_lvl3_ff[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5467_ (.Y(_2215_),
    .A(\mac1.sum_lvl3_ff[33] ),
    .B(net367),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5468_ (.Y(_0020_),
    .A(_2213_),
    .B(net368),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5469_ (.Y(_2216_),
    .A(\mac1.sum_lvl3_ff[34] ),
    .B(\mac1.sum_lvl3_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5470_ (.A(\mac1.sum_lvl3_ff[34] ),
    .B(\mac1.sum_lvl3_ff[14] ),
    .Y(_2217_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5471_ (.B(net477),
    .A(\mac1.sum_lvl3_ff[34] ),
    .X(_2218_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5472_ (.B(_2211_),
    .C(_2214_),
    .A(_2206_),
    .Y(_2219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5473_ (.B1(_2219_),
    .VDD(VPWR),
    .Y(_2220_),
    .VSS(VGND),
    .A1(\mac1.sum_lvl3_ff[33] ),
    .A2(net367));
 sg13g2_xnor2_1 _5474_ (.Y(_0021_),
    .A(net478),
    .B(_2220_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5475_ (.B1(_2216_),
    .VDD(VPWR),
    .Y(_2221_),
    .VSS(VGND),
    .A1(_2217_),
    .A2(_2220_));
 sg13g2_xnor2_1 _5476_ (.Y(_2222_),
    .A(\mac1.sum_lvl3_ff[35] ),
    .B(net438),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5477_ (.Y(_0022_),
    .A(_2221_),
    .B(net439),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5478_ (.B(net265),
    .A(\mac1.sum_lvl3_ff[20] ),
    .X(_0016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5479_ (.Y(_2223_),
    .A(net284),
    .B(net267),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5480_ (.Y(_2224_),
    .A(\mac2.sum_lvl2_ff[20] ),
    .B(\mac2.sum_lvl2_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5481_ (.A(\mac2.sum_lvl2_ff[20] ),
    .B(\mac2.sum_lvl2_ff[1] ),
    .Y(_2225_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5482_ (.B(\mac2.sum_lvl2_ff[1] ),
    .A(\mac2.sum_lvl2_ff[20] ),
    .X(_2226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5483_ (.Y(_0039_),
    .A(_2223_),
    .B(_2226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5484_ (.B1(_2224_),
    .VDD(VPWR),
    .Y(_2227_),
    .VSS(VGND),
    .A1(_2223_),
    .A2(_2225_));
 sg13g2_and2_1 _5485_ (.A(\mac2.sum_lvl2_ff[21] ),
    .B(net305),
    .X(_2228_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5486_ (.B(net305),
    .A(\mac2.sum_lvl2_ff[21] ),
    .X(_2229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5487_ (.B(net306),
    .A(_2227_),
    .X(_0040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5488_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2227_),
    .A2(net306),
    .Y(_2230_),
    .B1(_2228_));
 sg13g2_nand2_1 _5489_ (.Y(_2231_),
    .A(\mac2.sum_lvl2_ff[22] ),
    .B(net353),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5490_ (.Y(_2232_),
    .A(\mac2.sum_lvl2_ff[22] ),
    .B(net353),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5491_ (.B(net354),
    .A(_2230_),
    .X(_0041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5492_ (.B1(_2231_),
    .VDD(VPWR),
    .Y(_2233_),
    .VSS(VGND),
    .A1(_2230_),
    .A2(_2232_));
 sg13g2_and2_1 _5493_ (.A(\mac2.sum_lvl2_ff[23] ),
    .B(\mac2.sum_lvl2_ff[4] ),
    .X(_2234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5494_ (.B(net451),
    .A(\mac2.sum_lvl2_ff[23] ),
    .X(_2235_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5495_ (.B(net452),
    .A(_2233_),
    .X(_0042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5496_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2233_),
    .A2(_2235_),
    .Y(_2236_),
    .B1(_2234_));
 sg13g2_nor2_1 _5497_ (.A(net387),
    .B(\mac2.sum_lvl2_ff[5] ),
    .Y(_2237_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5498_ (.B(\mac2.sum_lvl2_ff[5] ),
    .A(net387),
    .X(_2238_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5499_ (.Y(_0043_),
    .A(_2236_),
    .B(net388),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5500_ (.A(\mac2.sum_lvl2_ff[25] ),
    .B(\mac2.sum_lvl2_ff[6] ),
    .X(_2239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5501_ (.Y(_2240_),
    .A(\mac2.sum_lvl2_ff[25] ),
    .B(net517),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5502_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2235_),
    .C1(_2234_),
    .B1(_2233_),
    .A1(net387),
    .Y(_2241_),
    .A2(\mac2.sum_lvl2_ff[5] ));
 sg13g2_nor3_1 _5503_ (.A(_2237_),
    .B(net518),
    .C(_2241_),
    .Y(_2242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5504_ (.B1(net518),
    .VDD(VPWR),
    .Y(_2243_),
    .VSS(VGND),
    .A1(_2237_),
    .A2(_2241_));
 sg13g2_nor2b_2 _5505_ (.A(_2242_),
    .B_N(net519),
    .Y(_0044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5506_ (.Y(_2244_),
    .A(\mac2.sum_lvl2_ff[26] ),
    .B(\mac2.sum_lvl2_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5507_ (.B(\mac2.sum_lvl2_ff[7] ),
    .A(\mac2.sum_lvl2_ff[26] ),
    .X(_2245_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5508_ (.B1(_2245_),
    .VDD(VPWR),
    .Y(_2246_),
    .VSS(VGND),
    .A1(_2239_),
    .A2(_2242_));
 sg13g2_or3_1 _5509_ (.A(_2239_),
    .B(_2242_),
    .C(_2245_),
    .X(_2247_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5510_ (.A(_2246_),
    .B(_2247_),
    .X(_0045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5511_ (.Y(_2248_),
    .A(\mac2.sum_lvl2_ff[27] ),
    .B(net490),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5512_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2244_),
    .A2(_2246_),
    .Y(_2249_),
    .B1(net491));
 sg13g2_nand3_1 _5513_ (.B(_2246_),
    .C(net491),
    .A(_2244_),
    .Y(_2250_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _5514_ (.A(net492),
    .B_N(_2250_),
    .Y(_0046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5515_ (.A2(net490),
    .A1(\mac2.sum_lvl2_ff[27] ),
    .B1(_2249_),
    .X(_2251_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5516_ (.A(\mac2.sum_lvl2_ff[28] ),
    .B(\mac2.sum_lvl2_ff[9] ),
    .X(_2252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5517_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2253_),
    .B(net545),
    .A(\mac2.sum_lvl2_ff[28] ));
 sg13g2_nand2b_1 _5518_ (.Y(_2254_),
    .B(_2253_),
    .A_N(_2252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5519_ (.Y(_0047_),
    .A(_2251_),
    .B(_2254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5520_ (.Y(_2255_),
    .A(\mac2.sum_lvl2_ff[29] ),
    .B(\mac2.sum_lvl2_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5521_ (.B(\mac2.sum_lvl2_ff[10] ),
    .A(\mac2.sum_lvl2_ff[29] ),
    .X(_2256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5522_ (.VDD(VPWR),
    .Y(_2257_),
    .A(_2256_),
    .VSS(VGND));
 sg13g2_a21o_2 _5523_ (.A2(_2253_),
    .A1(_2251_),
    .B1(_2252_),
    .X(_2258_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5524_ (.Y(_2259_),
    .A(_2256_),
    .B(_2258_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5525_ (.Y(_0033_),
    .A(_2257_),
    .B(_2258_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5526_ (.A(\mac2.sum_lvl2_ff[30] ),
    .B(\mac2.sum_lvl2_ff[11] ),
    .Y(_2260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5527_ (.Y(_2261_),
    .A(\mac2.sum_lvl2_ff[30] ),
    .B(\mac2.sum_lvl2_ff[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5528_ (.Y(_2262_),
    .A(_2255_),
    .B(_2259_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5529_ (.Y(_0034_),
    .A(_2261_),
    .B(_2262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5530_ (.Y(_2263_),
    .A(\mac2.sum_lvl2_ff[31] ),
    .B(\mac2.sum_lvl2_ff[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5531_ (.A(\mac2.sum_lvl2_ff[31] ),
    .B(\mac2.sum_lvl2_ff[12] ),
    .Y(_2264_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5532_ (.B(\mac2.sum_lvl2_ff[12] ),
    .A(\mac2.sum_lvl2_ff[31] ),
    .X(_2265_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5533_ (.A(_2255_),
    .B(_2260_),
    .Y(_2266_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5534_ (.A(_2257_),
    .B(_2261_),
    .Y(_2267_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5535_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2267_),
    .C1(_2266_),
    .B1(_2258_),
    .A1(\mac2.sum_lvl2_ff[30] ),
    .Y(_2268_),
    .A2(\mac2.sum_lvl2_ff[11] ));
 sg13g2_xnor2_1 _5536_ (.Y(_0035_),
    .A(_2265_),
    .B(_2268_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5537_ (.B1(_2263_),
    .VDD(VPWR),
    .Y(_2269_),
    .VSS(VGND),
    .A1(_2264_),
    .A2(_2268_));
 sg13g2_and2_1 _5538_ (.A(\mac2.sum_lvl2_ff[32] ),
    .B(\mac2.sum_lvl2_ff[13] ),
    .X(_2270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5539_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2271_),
    .B(\mac2.sum_lvl2_ff[13] ),
    .A(\mac2.sum_lvl2_ff[32] ));
 sg13g2_nand2b_1 _5540_ (.Y(_2272_),
    .B(_2271_),
    .A_N(_2270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5541_ (.Y(_0036_),
    .A(_2269_),
    .B(_2272_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5542_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2269_),
    .A2(_2271_),
    .Y(_2273_),
    .B1(_2270_));
 sg13g2_nand2_1 _5543_ (.Y(_2274_),
    .A(\mac2.sum_lvl2_ff[33] ),
    .B(\mac2.sum_lvl2_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5544_ (.A(\mac2.sum_lvl2_ff[33] ),
    .B(\mac2.sum_lvl2_ff[14] ),
    .Y(_2275_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5545_ (.B(net542),
    .A(\mac2.sum_lvl2_ff[33] ),
    .X(_2276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5546_ (.Y(_0037_),
    .A(_2273_),
    .B(net543),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5547_ (.B1(_2274_),
    .VDD(VPWR),
    .Y(_2277_),
    .VSS(VGND),
    .A1(_2273_),
    .A2(_2275_));
 sg13g2_xnor2_1 _5548_ (.Y(_2278_),
    .A(\mac2.sum_lvl2_ff[34] ),
    .B(net527),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5549_ (.Y(_0038_),
    .A(_2277_),
    .B(net528),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5550_ (.B(net267),
    .A(\mac2.sum_lvl2_ff[19] ),
    .X(_0032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5551_ (.Y(_2279_),
    .A(net449),
    .B(net290),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5552_ (.Y(_2280_),
    .A(\mac2.sum_lvl3_ff[21] ),
    .B(\mac2.sum_lvl3_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5553_ (.A(\mac2.sum_lvl3_ff[21] ),
    .B(\mac2.sum_lvl3_ff[1] ),
    .Y(_2281_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5554_ (.B(\mac2.sum_lvl3_ff[1] ),
    .A(\mac2.sum_lvl3_ff[21] ),
    .X(_2282_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5555_ (.Y(_0055_),
    .A(_2279_),
    .B(_2282_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5556_ (.B1(_2280_),
    .VDD(VPWR),
    .Y(_2283_),
    .VSS(VGND),
    .A1(_2279_),
    .A2(_2281_));
 sg13g2_and2_1 _5557_ (.A(net473),
    .B(\mac2.sum_lvl3_ff[2] ),
    .X(_2284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5558_ (.B(\mac2.sum_lvl3_ff[2] ),
    .A(net473),
    .X(_2285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5559_ (.B(net474),
    .A(_2283_),
    .X(_0056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5560_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2283_),
    .A2(_2285_),
    .Y(_2286_),
    .B1(_2284_));
 sg13g2_nand2_1 _5561_ (.Y(_2287_),
    .A(\mac2.sum_lvl3_ff[23] ),
    .B(\mac2.sum_lvl3_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5562_ (.Y(_2288_),
    .A(\mac2.sum_lvl3_ff[23] ),
    .B(net484),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5563_ (.B(net485),
    .A(_2286_),
    .X(_0057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5564_ (.B1(_2287_),
    .VDD(VPWR),
    .Y(_2289_),
    .VSS(VGND),
    .A1(_2286_),
    .A2(_2288_));
 sg13g2_and2_1 _5565_ (.A(\mac2.sum_lvl3_ff[24] ),
    .B(net457),
    .X(_2290_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5566_ (.B(net457),
    .A(\mac2.sum_lvl3_ff[24] ),
    .X(_2291_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5567_ (.B(net458),
    .A(_2289_),
    .X(_0058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5568_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2289_),
    .A2(_2291_),
    .Y(_2292_),
    .B1(_2290_));
 sg13g2_nor2_1 _5569_ (.A(\mac2.sum_lvl3_ff[25] ),
    .B(net396),
    .Y(_2293_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5570_ (.B(net396),
    .A(\mac2.sum_lvl3_ff[25] ),
    .X(_2294_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5571_ (.Y(_0059_),
    .A(_2292_),
    .B(net397),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5572_ (.A(\mac2.sum_lvl3_ff[26] ),
    .B(net463),
    .X(_2295_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5573_ (.Y(_2296_),
    .A(\mac2.sum_lvl3_ff[26] ),
    .B(net463),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5574_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2291_),
    .C1(_2290_),
    .B1(_2289_),
    .A1(\mac2.sum_lvl3_ff[25] ),
    .Y(_2297_),
    .A2(net396));
 sg13g2_nor3_1 _5575_ (.A(_2293_),
    .B(net464),
    .C(_2297_),
    .Y(_2298_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5576_ (.B1(net464),
    .VDD(VPWR),
    .Y(_2299_),
    .VSS(VGND),
    .A1(_2293_),
    .A2(_2297_));
 sg13g2_nor2b_1 _5577_ (.A(_2298_),
    .B_N(net465),
    .Y(_0060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5578_ (.Y(_2300_),
    .A(\mac2.sum_lvl3_ff[27] ),
    .B(\mac2.sum_lvl3_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5579_ (.B(net537),
    .A(\mac2.sum_lvl3_ff[27] ),
    .X(_2301_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5580_ (.B1(net538),
    .VDD(VPWR),
    .Y(_2302_),
    .VSS(VGND),
    .A1(_2295_),
    .A2(_2298_));
 sg13g2_or3_1 _5581_ (.A(_2295_),
    .B(_2298_),
    .C(net538),
    .X(_2303_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5582_ (.A(net539),
    .B(_2303_),
    .X(_0061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5583_ (.Y(_2304_),
    .A(\mac2.sum_lvl3_ff[28] ),
    .B(net423),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5584_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2300_),
    .A2(_2302_),
    .Y(_2305_),
    .B1(net424));
 sg13g2_nand3_1 _5585_ (.B(_2302_),
    .C(net424),
    .A(_2300_),
    .Y(_2306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5586_ (.A(net425),
    .B_N(_2306_),
    .Y(_0062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5587_ (.A2(net423),
    .A1(net429),
    .B1(net425),
    .X(_2307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5588_ (.A(\mac2.sum_lvl3_ff[29] ),
    .B(\mac2.sum_lvl3_ff[9] ),
    .X(_2308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5589_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2309_),
    .B(\mac2.sum_lvl3_ff[9] ),
    .A(\mac2.sum_lvl3_ff[29] ));
 sg13g2_nand2b_1 _5590_ (.Y(_2310_),
    .B(_2309_),
    .A_N(_2308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5591_ (.Y(_0063_),
    .A(_2307_),
    .B(_2310_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5592_ (.Y(_2311_),
    .A(net336),
    .B(\mac2.sum_lvl3_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5593_ (.B(net444),
    .A(net336),
    .X(_2312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5594_ (.VDD(VPWR),
    .Y(_2313_),
    .A(_2312_),
    .VSS(VGND));
 sg13g2_a21o_2 _5595_ (.A2(_2309_),
    .A1(_2307_),
    .B1(_2308_),
    .X(_2314_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5596_ (.Y(_2315_),
    .A(_2312_),
    .B(_2314_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5597_ (.Y(_0049_),
    .A(_2313_),
    .B(_2314_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5598_ (.A(\mac2.sum_lvl3_ff[31] ),
    .B(\mac2.sum_lvl3_ff[11] ),
    .Y(_2316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5599_ (.Y(_2317_),
    .A(\mac2.sum_lvl3_ff[31] ),
    .B(\mac2.sum_lvl3_ff[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5600_ (.Y(_2318_),
    .A(net337),
    .B(_2315_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5601_ (.Y(_0050_),
    .A(_2317_),
    .B(net338),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5602_ (.Y(_2319_),
    .A(\mac2.sum_lvl3_ff[32] ),
    .B(net310),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5603_ (.A(\mac2.sum_lvl3_ff[32] ),
    .B(net310),
    .Y(_2320_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5604_ (.B(net310),
    .A(\mac2.sum_lvl3_ff[32] ),
    .X(_2321_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5605_ (.A(_2311_),
    .B(_2316_),
    .Y(_2322_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5606_ (.A(_2313_),
    .B(_2317_),
    .Y(_2323_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5607_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2323_),
    .C1(_2322_),
    .B1(_2314_),
    .A1(\mac2.sum_lvl3_ff[31] ),
    .Y(_2324_),
    .A2(\mac2.sum_lvl3_ff[11] ));
 sg13g2_xnor2_1 _5608_ (.Y(_0051_),
    .A(net311),
    .B(_2324_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5609_ (.B1(_2319_),
    .VDD(VPWR),
    .Y(_2325_),
    .VSS(VGND),
    .A1(_2320_),
    .A2(_2324_));
 sg13g2_and2_1 _5610_ (.A(\mac2.sum_lvl3_ff[33] ),
    .B(net467),
    .X(_2326_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5611_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2327_),
    .B(net467),
    .A(\mac2.sum_lvl3_ff[33] ));
 sg13g2_nand2b_1 _5612_ (.Y(_2328_),
    .B(net468),
    .A_N(_2326_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5613_ (.Y(_0052_),
    .A(_2325_),
    .B(net469),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5614_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2325_),
    .A2(_2327_),
    .Y(_2329_),
    .B1(_2326_));
 sg13g2_nand2_1 _5615_ (.Y(_2330_),
    .A(\mac2.sum_lvl3_ff[34] ),
    .B(net328),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5616_ (.A(\mac2.sum_lvl3_ff[34] ),
    .B(net328),
    .Y(_2331_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5617_ (.B(net328),
    .A(\mac2.sum_lvl3_ff[34] ),
    .X(_2332_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5618_ (.Y(_0053_),
    .A(_2329_),
    .B(net329),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5619_ (.B1(_2330_),
    .VDD(VPWR),
    .Y(_2333_),
    .VSS(VGND),
    .A1(_2329_),
    .A2(_2331_));
 sg13g2_xnor2_1 _5620_ (.Y(_2334_),
    .A(\mac2.sum_lvl3_ff[35] ),
    .B(net343),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5621_ (.Y(_0054_),
    .A(_2333_),
    .B(net344),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5622_ (.B(net290),
    .A(\mac2.sum_lvl3_ff[20] ),
    .X(_0048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5623_ (.Y(_2335_),
    .A(\mac1.total_sum[0] ),
    .B(\mac2.total_sum[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5624_ (.Y(_2336_),
    .A(\mac1.total_sum[1] ),
    .B(\mac2.total_sum[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5625_ (.A(\mac1.total_sum[1] ),
    .B(\mac2.total_sum[1] ),
    .Y(_2337_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5626_ (.B(\mac2.total_sum[1] ),
    .A(\mac1.total_sum[1] ),
    .X(_2338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5627_ (.Y(net26),
    .A(_2335_),
    .B(_2338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5628_ (.B1(_2336_),
    .VDD(VPWR),
    .Y(_2339_),
    .VSS(VGND),
    .A1(_2335_),
    .A2(_2337_));
 sg13g2_and2_1 _5629_ (.A(\mac1.total_sum[2] ),
    .B(\mac2.total_sum[2] ),
    .X(_2340_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5630_ (.B(\mac2.total_sum[2] ),
    .A(\mac1.total_sum[2] ),
    .X(_2341_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5631_ (.B(_2341_),
    .A(_2339_),
    .X(net27),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5632_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2339_),
    .A2(_2341_),
    .Y(_2342_),
    .B1(_2340_));
 sg13g2_nand2_1 _5633_ (.Y(_2343_),
    .A(\mac1.total_sum[3] ),
    .B(\mac2.total_sum[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5634_ (.Y(_2344_),
    .A(\mac1.total_sum[3] ),
    .B(\mac2.total_sum[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5635_ (.B(_2344_),
    .A(_2342_),
    .X(net28),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5636_ (.B1(_2343_),
    .VDD(VPWR),
    .Y(_2345_),
    .VSS(VGND),
    .A1(_2342_),
    .A2(_2344_));
 sg13g2_and2_1 _5637_ (.A(\mac1.total_sum[4] ),
    .B(\mac2.total_sum[4] ),
    .X(_2346_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5638_ (.B(\mac2.total_sum[4] ),
    .A(\mac1.total_sum[4] ),
    .X(_2347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5639_ (.B(_2347_),
    .A(_2345_),
    .X(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5640_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2345_),
    .A2(_2347_),
    .Y(_2348_),
    .B1(_2346_));
 sg13g2_nor2_1 _5641_ (.A(\mac1.total_sum[5] ),
    .B(\mac2.total_sum[5] ),
    .Y(_2349_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5642_ (.B(\mac2.total_sum[5] ),
    .A(\mac1.total_sum[5] ),
    .X(_2350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5643_ (.Y(net30),
    .A(_2348_),
    .B(_2350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5644_ (.A(\mac1.total_sum[6] ),
    .B(\mac2.total_sum[6] ),
    .X(_2351_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5645_ (.Y(_2352_),
    .A(\mac1.total_sum[6] ),
    .B(\mac2.total_sum[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5646_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2347_),
    .C1(_2346_),
    .B1(_2345_),
    .A1(\mac1.total_sum[5] ),
    .Y(_2353_),
    .A2(\mac2.total_sum[5] ));
 sg13g2_nor3_1 _5647_ (.A(_2349_),
    .B(_2352_),
    .C(_2353_),
    .Y(_2354_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5648_ (.B1(_2352_),
    .VDD(VPWR),
    .Y(_2355_),
    .VSS(VGND),
    .A1(_2349_),
    .A2(_2353_));
 sg13g2_nor2b_1 _5649_ (.A(_2354_),
    .B_N(_2355_),
    .Y(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5650_ (.Y(_2356_),
    .A(\mac1.total_sum[7] ),
    .B(\mac2.total_sum[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5651_ (.B(\mac2.total_sum[7] ),
    .A(\mac1.total_sum[7] ),
    .X(_2357_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5652_ (.B1(_2357_),
    .VDD(VPWR),
    .Y(_2358_),
    .VSS(VGND),
    .A1(_2351_),
    .A2(_2354_));
 sg13g2_or3_1 _5653_ (.A(_2351_),
    .B(_2354_),
    .C(_2357_),
    .X(_2359_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5654_ (.A(_2358_),
    .B(_2359_),
    .X(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5655_ (.Y(_2360_),
    .A(\mac1.total_sum[8] ),
    .B(\mac2.total_sum[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5656_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2356_),
    .A2(_2358_),
    .Y(_2361_),
    .B1(_2360_));
 sg13g2_nand3_1 _5657_ (.B(_2358_),
    .C(_2360_),
    .A(_2356_),
    .Y(_2362_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5658_ (.A(_2361_),
    .B_N(_2362_),
    .Y(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5659_ (.A2(\mac2.total_sum[8] ),
    .A1(\mac1.total_sum[8] ),
    .B1(_2361_),
    .X(_2363_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5660_ (.A(\mac1.total_sum[9] ),
    .B(\mac2.total_sum[9] ),
    .X(_2364_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5661_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2365_),
    .B(\mac2.total_sum[9] ),
    .A(\mac1.total_sum[9] ));
 sg13g2_nand2b_1 _5662_ (.Y(_2366_),
    .B(_2365_),
    .A_N(_2364_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5663_ (.Y(net18),
    .A(_2363_),
    .B(_2366_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5664_ (.Y(_2367_),
    .A(\mac1.total_sum[10] ),
    .B(\mac2.total_sum[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5665_ (.B(\mac2.total_sum[10] ),
    .A(\mac1.total_sum[10] ),
    .X(_2368_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5666_ (.VDD(VPWR),
    .Y(_2369_),
    .A(_2368_),
    .VSS(VGND));
 sg13g2_a21o_2 _5667_ (.A2(_2365_),
    .A1(_2363_),
    .B1(_2364_),
    .X(_2370_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5668_ (.Y(_2371_),
    .A(_2368_),
    .B(_2370_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5669_ (.Y(net19),
    .A(_2369_),
    .B(_2370_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5670_ (.A(\mac1.total_sum[11] ),
    .B(\mac2.total_sum[11] ),
    .Y(_2372_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5671_ (.Y(_2373_),
    .A(\mac1.total_sum[11] ),
    .B(\mac2.total_sum[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5672_ (.Y(_2374_),
    .A(_2367_),
    .B(_2371_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5673_ (.Y(net20),
    .A(_2373_),
    .B(_2374_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5674_ (.Y(_2375_),
    .A(\mac1.total_sum[12] ),
    .B(\mac2.total_sum[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5675_ (.A(\mac1.total_sum[12] ),
    .B(\mac2.total_sum[12] ),
    .Y(_2376_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5676_ (.B(\mac2.total_sum[12] ),
    .A(\mac1.total_sum[12] ),
    .X(_2377_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5677_ (.A(_2367_),
    .B(_2372_),
    .Y(_2378_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5678_ (.A(_2369_),
    .B(_2373_),
    .Y(_2379_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5679_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2379_),
    .C1(_2378_),
    .B1(_2370_),
    .A1(\mac1.total_sum[11] ),
    .Y(_2380_),
    .A2(\mac2.total_sum[11] ));
 sg13g2_xnor2_1 _5680_ (.Y(net21),
    .A(_2377_),
    .B(_2380_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5681_ (.B1(_2375_),
    .VDD(VPWR),
    .Y(_2381_),
    .VSS(VGND),
    .A1(_2376_),
    .A2(_2380_));
 sg13g2_and2_1 _5682_ (.A(\mac1.total_sum[13] ),
    .B(\mac2.total_sum[13] ),
    .X(_2382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5683_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2383_),
    .B(\mac2.total_sum[13] ),
    .A(\mac1.total_sum[13] ));
 sg13g2_nand2b_1 _5684_ (.Y(_2384_),
    .B(_2383_),
    .A_N(_2382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5685_ (.Y(net22),
    .A(_2381_),
    .B(_2384_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5686_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2381_),
    .A2(_2383_),
    .Y(_2385_),
    .B1(_2382_));
 sg13g2_nand2_1 _5687_ (.Y(_2386_),
    .A(\mac1.total_sum[14] ),
    .B(\mac2.total_sum[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5688_ (.A(\mac1.total_sum[14] ),
    .B(\mac2.total_sum[14] ),
    .Y(_2387_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5689_ (.B(\mac2.total_sum[14] ),
    .A(\mac1.total_sum[14] ),
    .X(_2388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5690_ (.Y(net23),
    .A(_2385_),
    .B(_2388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5691_ (.B1(_2386_),
    .VDD(VPWR),
    .Y(_2389_),
    .VSS(VGND),
    .A1(_2385_),
    .A2(_2387_));
 sg13g2_xnor2_1 _5692_ (.Y(_2390_),
    .A(\mac1.total_sum[15] ),
    .B(\mac2.total_sum[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5693_ (.Y(net24),
    .A(_2389_),
    .B(_2390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5694_ (.B(\mac2.total_sum[0] ),
    .A(\mac1.total_sum[0] ),
    .X(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _5695_ (.A(\DP_1.I_range.out_data[4] ),
    .B(_2602_),
    .C(\DP_1.Q_range.out_data[4] ),
    .D(\DP_1.Q_range.out_data[6] ),
    .X(_2391_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _5696_ (.A(\DP_1.I_range.out_data[2] ),
    .B(\DP_1.Q_range.out_data[2] ),
    .C(\DP_1.I_range.out_data[6] ),
    .D(_2601_),
    .X(_2392_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _5697_ (.A(net443),
    .B(_2600_),
    .C(_2391_),
    .D(_2392_),
    .Y(_2393_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _5698_ (.A(\DP_1.I_range.out_data[3] ),
    .B(_2600_),
    .C(\DP_1.I_range.out_data[2] ),
    .D(_2601_),
    .X(_2394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _5699_ (.A(\DP_1.Q_range.out_data[2] ),
    .B(\DP_1.I_range.out_data[6] ),
    .C(_2391_),
    .D(_2394_),
    .X(_2395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5700_ (.A(\DP_1.Q_range.out_data[2] ),
    .B_N(\DP_1.I_range.out_data[2] ),
    .Y(_2396_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5701_ (.Y(_2397_),
    .A(\DP_1.I_range.out_data[3] ),
    .B(\DP_1.Q_range.out_data[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5702_ (.Y(_2398_),
    .A(_2396_),
    .B(_2397_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5703_ (.Y(_2399_),
    .A(\DP_1.I_range.out_data[2] ),
    .B(\DP_1.Q_range.out_data[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5704_ (.B(\DP_1.Q_range.out_data[2] ),
    .A(\DP_1.I_range.out_data[2] ),
    .X(_2400_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5705_ (.B1(net784),
    .VDD(VPWR),
    .Y(_2401_),
    .VSS(VGND),
    .A1(net1037),
    .A2(net789));
 sg13g2_inv_1 _5706_ (.VDD(VPWR),
    .Y(_2402_),
    .A(_2401_),
    .VSS(VGND));
 sg13g2_o21ai_1 _5707_ (.B1(_2402_),
    .VDD(VPWR),
    .Y(_2403_),
    .VSS(VGND),
    .A1(net403),
    .A2(net791));
 sg13g2_and2_1 _5708_ (.A(net772),
    .B(_2403_),
    .X(_2404_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5709_ (.A(_2397_),
    .B(net790),
    .X(_2405_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5710_ (.A2(_2395_),
    .A1(net1037),
    .B1(_2404_),
    .X(_2406_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5711_ (.A(\DP_1.matrix[43] ),
    .B(net791),
    .Y(_2407_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5712_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2605_),
    .A2(net791),
    .Y(_2408_),
    .B1(_2407_));
 sg13g2_a22oi_1 _5713_ (.Y(_2409_),
    .B1(_2408_),
    .B2(net783),
    .A2(net780),
    .A1(net966),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5714_ (.A0(net1009),
    .A1(\DP_1.matrix[41] ),
    .S(net788),
    .X(_2410_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5715_ (.Y(_2411_),
    .B1(_2410_),
    .B2(net783),
    .A2(net780),
    .A1(net327),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5716_ (.A0(net1013),
    .A1(net998),
    .S(net788),
    .X(_2412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5717_ (.Y(_2413_),
    .B1(_2412_),
    .B2(net784),
    .A2(net780),
    .A1(net977),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5718_ (.A0(net1003),
    .A1(net1019),
    .S(net790),
    .X(_2414_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5719_ (.Y(_2415_),
    .B1(_2414_),
    .B2(net782),
    .A2(net781),
    .A1(net273),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5720_ (.A(net1018),
    .B(net789),
    .Y(_2416_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5721_ (.Y(_2417_),
    .A(net983),
    .B(net790),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5722_ (.B1(net782),
    .VDD(VPWR),
    .Y(_2418_),
    .VSS(VGND),
    .A1(net1002),
    .A2(net790));
 sg13g2_a22oi_1 _5723_ (.Y(_2419_),
    .B1(_2417_),
    .B2(_2418_),
    .A2(_2416_),
    .A1(net782),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5724_ (.Y(_2420_),
    .B(_2419_),
    .A_N(_2415_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5725_ (.A0(net1015),
    .A1(net1000),
    .S(net789),
    .X(_2421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5726_ (.Y(_2422_),
    .B1(_2421_),
    .B2(net782),
    .A2(net781),
    .A1(net980),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5727_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2423_),
    .B(_2422_),
    .A(_2420_));
 sg13g2_or2_1 _5728_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2424_),
    .B(_2423_),
    .A(_2413_));
 sg13g2_mux2_1 _5729_ (.A0(net1011),
    .A1(net996),
    .S(net788),
    .X(_2425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5730_ (.Y(_2426_),
    .B1(_2425_),
    .B2(net783),
    .A2(net780),
    .A1(net974),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5731_ (.A(_2424_),
    .B(_2426_),
    .Y(_2427_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5732_ (.A(_2411_),
    .B(_2424_),
    .C(_2426_),
    .Y(_2428_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5733_ (.A0(net1007),
    .A1(\DP_1.matrix[42] ),
    .S(net788),
    .X(_2429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5734_ (.Y(_2430_),
    .B1(_2429_),
    .B2(net783),
    .A2(net780),
    .A1(net315),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5735_ (.A(_2430_),
    .B_N(_2428_),
    .Y(_2431_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5736_ (.Y(_2432_),
    .B(_2431_),
    .A_N(_2409_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5737_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net773),
    .A2(_2432_),
    .Y(_2433_),
    .B1(_2406_));
 sg13g2_a21oi_1 _5738_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2404_),
    .A2(_2432_),
    .Y(_0160_),
    .B1(_2433_));
 sg13g2_o21ai_1 _5739_ (.B1(net783),
    .VDD(VPWR),
    .Y(_2434_),
    .VSS(VGND),
    .A1(net1032),
    .A2(net789));
 sg13g2_inv_1 _5740_ (.VDD(VPWR),
    .Y(_2435_),
    .A(_2434_),
    .VSS(VGND));
 sg13g2_o21ai_1 _5741_ (.B1(_2435_),
    .VDD(VPWR),
    .Y(_2436_),
    .VSS(VGND),
    .A1(net384),
    .A2(net791));
 sg13g2_and2_1 _5742_ (.A(net773),
    .B(_2436_),
    .X(_2437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5743_ (.A2(_2395_),
    .A1(net1032),
    .B1(_2437_),
    .X(_2438_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5744_ (.A(\DP_2.matrix[43] ),
    .B(net790),
    .Y(_2439_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5745_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2606_),
    .A2(net791),
    .Y(_2440_),
    .B1(_2439_));
 sg13g2_a22oi_1 _5746_ (.Y(_2441_),
    .B1(_2440_),
    .B2(net783),
    .A2(net780),
    .A1(net906),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5747_ (.A0(net949),
    .A1(net930),
    .S(net788),
    .X(_2442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5748_ (.Y(_2443_),
    .B1(_2442_),
    .B2(net784),
    .A2(net780),
    .A1(net910),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5749_ (.A0(net952),
    .A1(net934),
    .S(net788),
    .X(_2444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5750_ (.Y(_2445_),
    .B1(_2444_),
    .B2(net783),
    .A2(net780),
    .A1(net279),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5751_ (.A0(net943),
    .A1(net960),
    .S(net790),
    .X(_2446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5752_ (.Y(_2447_),
    .B1(_2446_),
    .B2(net782),
    .A2(net781),
    .A1(net924),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5753_ (.A(net956),
    .B(net789),
    .Y(_2448_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5754_ (.Y(_2449_),
    .A(net272),
    .B(net790),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5755_ (.B1(net782),
    .VDD(VPWR),
    .Y(_2450_),
    .VSS(VGND),
    .A1(net940),
    .A2(net790));
 sg13g2_a22oi_1 _5756_ (.Y(_2451_),
    .B1(_2449_),
    .B2(_2450_),
    .A2(_2448_),
    .A1(net782),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5757_ (.Y(_2452_),
    .B(_2451_),
    .A_N(_2447_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5758_ (.A0(net954),
    .A1(net936),
    .S(net789),
    .X(_2453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5759_ (.Y(_2454_),
    .B1(_2453_),
    .B2(net782),
    .A2(net781),
    .A1(\DP_2.matrix[74] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5760_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2455_),
    .B(_2454_),
    .A(_2452_));
 sg13g2_or2_1 _5761_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2456_),
    .B(_2455_),
    .A(_2445_));
 sg13g2_nand2_1 _5762_ (.Y(_2457_),
    .A(net269),
    .B(net781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5763_ (.A(\DP_2.matrix[40] ),
    .B(net791),
    .Y(_2458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5764_ (.B1(net783),
    .VDD(VPWR),
    .Y(_2459_),
    .VSS(VGND),
    .A1(net951),
    .A2(net788));
 sg13g2_o21ai_1 _5765_ (.B1(_2457_),
    .VDD(VPWR),
    .Y(_2460_),
    .VSS(VGND),
    .A1(_2458_),
    .A2(_2459_));
 sg13g2_nor2b_1 _5766_ (.A(_2456_),
    .B_N(_2460_),
    .Y(_2461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5767_ (.A(_2443_),
    .B_N(_2461_),
    .Y(_2462_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5768_ (.A0(net948),
    .A1(\DP_2.matrix[42] ),
    .S(net788),
    .X(_2463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5769_ (.Y(_2464_),
    .B1(_2463_),
    .B2(net784),
    .A2(net781),
    .A1(net908),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5770_ (.A(_2464_),
    .B_N(_2462_),
    .Y(_2465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5771_ (.Y(_2466_),
    .B(_2465_),
    .A_N(_2441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5772_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net773),
    .A2(_2466_),
    .Y(_2467_),
    .B1(_2438_));
 sg13g2_a21oi_1 _5773_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2437_),
    .A2(_2466_),
    .Y(_0163_),
    .B1(_2467_));
 sg13g2_nor2b_1 _5774_ (.A(\DP_3.I_range.out_data[3] ),
    .B_N(\DP_3.Q_range.out_data[3] ),
    .Y(_2468_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5775_ (.B(\DP_3.Q_range.out_data[3] ),
    .A(\DP_3.I_range.out_data[3] ),
    .X(_2469_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5776_ (.Y(_2470_),
    .B(\DP_3.I_range.out_data[2] ),
    .A_N(\DP_3.Q_range.out_data[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5777_ (.Y(_2471_),
    .A(_2469_),
    .B(_2470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5778_ (.Y(_2472_),
    .A(\DP_3.I_range.out_data[2] ),
    .B(\DP_3.Q_range.out_data[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5779_ (.B(\DP_3.Q_range.out_data[2] ),
    .A(\DP_3.I_range.out_data[2] ),
    .X(_2473_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5780_ (.B1(net778),
    .VDD(VPWR),
    .Y(_2474_),
    .VSS(VGND),
    .A1(net1028),
    .A2(net785));
 sg13g2_a21oi_1 _5781_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2607_),
    .A2(net785),
    .Y(_2475_),
    .B1(_2474_));
 sg13g2_nor4_1 _5782_ (.A(\DP_3.Q_range.out_data[2] ),
    .B(_2604_),
    .C(\DP_3.Q_range.out_data[4] ),
    .D(\DP_3.Q_range.out_data[6] ),
    .Y(_2476_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _5783_ (.A(\DP_3.I_range.out_data[6] ),
    .B(\DP_3.I_range.out_data[2] ),
    .C(_2603_),
    .D(\DP_3.I_range.out_data[4] ),
    .Y(_2477_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _5784_ (.X(_2478_),
    .A(_2468_),
    .B(_2476_),
    .C(_2477_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5785_ (.B(_2476_),
    .C(_2477_),
    .A(_2468_),
    .Y(_2479_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5786_ (.Y(_2480_),
    .A(net1028),
    .B(net767),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5787_ (.B1(_2480_),
    .VDD(VPWR),
    .Y(_2481_),
    .VSS(VGND),
    .A1(_2475_),
    .A2(net767));
 sg13g2_nor2_1 _5788_ (.A(_2469_),
    .B(net785),
    .Y(_2482_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5789_ (.Y(_2483_),
    .A(\DP_3.matrix[77] ),
    .B(net775),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5790_ (.A(net876),
    .B(_2472_),
    .Y(_2484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5791_ (.B1(net778),
    .VDD(VPWR),
    .Y(_2485_),
    .VSS(VGND),
    .A1(net894),
    .A2(net785));
 sg13g2_o21ai_1 _5792_ (.B1(_2483_),
    .VDD(VPWR),
    .Y(_2486_),
    .VSS(VGND),
    .A1(_2484_),
    .A2(_2485_));
 sg13g2_mux2_1 _5793_ (.A0(net880),
    .A1(net897),
    .S(net786),
    .X(_2487_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5794_ (.Y(_2488_),
    .B1(_2487_),
    .B2(net777),
    .A2(net775),
    .A1(net862),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5795_ (.Y(_2489_),
    .A(net869),
    .B(net775),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5796_ (.A(net886),
    .B(net786),
    .Y(_2490_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5797_ (.B1(net777),
    .VDD(VPWR),
    .Y(_2491_),
    .VSS(VGND),
    .A1(net903),
    .A2(net785));
 sg13g2_o21ai_1 _5798_ (.B1(_2489_),
    .VDD(VPWR),
    .Y(_2492_),
    .VSS(VGND),
    .A1(_2490_),
    .A2(_2491_));
 sg13g2_nand2_1 _5799_ (.Y(_2493_),
    .A(_2469_),
    .B(net786),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5800_ (.Y(_2494_),
    .B1(net786),
    .B2(net867),
    .A2(net777),
    .A1(net885),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5801_ (.A(net901),
    .B(_2493_),
    .Y(_2495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5802_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2493_),
    .A2(_2494_),
    .Y(_2496_),
    .B1(_2495_));
 sg13g2_and2_1 _5803_ (.A(_2492_),
    .B(_2496_),
    .X(_2497_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5804_ (.A0(net882),
    .A1(net899),
    .S(net786),
    .X(_2498_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5805_ (.Y(_2499_),
    .B1(_2498_),
    .B2(net777),
    .A2(net775),
    .A1(net865),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5806_ (.A(_2499_),
    .B_N(_2497_),
    .Y(_2500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5807_ (.Y(_2501_),
    .B(_2500_),
    .A_N(_2488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5808_ (.A0(net878),
    .A1(net895),
    .S(net787),
    .X(_2502_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5809_ (.Y(_2503_),
    .B1(_2502_),
    .B2(net777),
    .A2(net775),
    .A1(net274),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _5810_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2504_),
    .B(_2503_),
    .A(_2501_));
 sg13g2_nand2b_1 _5811_ (.Y(_2505_),
    .B(_2486_),
    .A_N(_2504_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5812_ (.Y(_2506_),
    .A(net280),
    .B(net775),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5813_ (.A(net875),
    .B(_2472_),
    .Y(_2507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5814_ (.B1(net778),
    .VDD(VPWR),
    .Y(_2508_),
    .VSS(VGND),
    .A1(net892),
    .A2(net785));
 sg13g2_o21ai_1 _5815_ (.B1(_2506_),
    .VDD(VPWR),
    .Y(_2509_),
    .VSS(VGND),
    .A1(_2507_),
    .A2(_2508_));
 sg13g2_nor2b_1 _5816_ (.A(_2505_),
    .B_N(_2509_),
    .Y(_2510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5817_ (.A0(net872),
    .A1(net890),
    .S(net787),
    .X(_2511_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5818_ (.Y(_2512_),
    .B1(_2511_),
    .B2(net778),
    .A2(net776),
    .A1(net275),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5819_ (.Y(_2513_),
    .B(_2510_),
    .A_N(_2512_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5820_ (.Y(_2514_),
    .A(net770),
    .B(_2513_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5821_ (.A0(_2475_),
    .A1(_2481_),
    .S(_2514_),
    .X(_0166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5822_ (.A0(\DP_4.matrix[44] ),
    .A1(net1023),
    .S(net787),
    .X(_2515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5823_ (.A(net778),
    .B(_2515_),
    .X(_2516_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5824_ (.Y(_2517_),
    .A(net1023),
    .B(net767),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5825_ (.B1(_2517_),
    .VDD(VPWR),
    .Y(_2518_),
    .VSS(VGND),
    .A1(net767),
    .A2(_2516_));
 sg13g2_nand2_1 _5826_ (.Y(_2519_),
    .A(net799),
    .B(net776),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5827_ (.A(net818),
    .B(net787),
    .Y(_2520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5828_ (.B1(net779),
    .VDD(VPWR),
    .Y(_2521_),
    .VSS(VGND),
    .A1(net836),
    .A2(net785));
 sg13g2_o21ai_1 _5829_ (.B1(_2519_),
    .VDD(VPWR),
    .Y(_2522_),
    .VSS(VGND),
    .A1(_2520_),
    .A2(_2521_));
 sg13g2_mux2_1 _5830_ (.A0(net822),
    .A1(net839),
    .S(net787),
    .X(_2523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5831_ (.Y(_2524_),
    .B1(_2523_),
    .B2(net779),
    .A2(net776),
    .A1(net374),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5832_ (.A0(net831),
    .A1(net847),
    .S(net786),
    .X(_2525_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5833_ (.Y(_2526_),
    .B1(_2525_),
    .B2(net777),
    .A2(net775),
    .A1(net282),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5834_ (.Y(_2527_),
    .B1(net786),
    .B2(net810),
    .A2(net777),
    .A1(net825),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5835_ (.A(net843),
    .B(_2493_),
    .Y(_2528_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5836_ (.A2(_2527_),
    .A1(_2493_),
    .B1(_2528_),
    .X(_2529_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5837_ (.A(_2526_),
    .B(_2529_),
    .Y(_2530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5838_ (.A0(net823),
    .A1(net841),
    .S(net786),
    .X(_2531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5839_ (.Y(_2532_),
    .B1(_2531_),
    .B2(net777),
    .A2(net775),
    .A1(net805),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5840_ (.A(_2526_),
    .B(_2529_),
    .C(_2532_),
    .Y(_2533_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5841_ (.Y(_2534_),
    .B(_2533_),
    .A_N(_2524_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5842_ (.Y(_2535_),
    .A(net276),
    .B(net776),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5843_ (.A(net820),
    .B(net787),
    .Y(_2536_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5844_ (.B1(net778),
    .VDD(VPWR),
    .Y(_2537_),
    .VSS(VGND),
    .A1(net837),
    .A2(net785));
 sg13g2_o21ai_1 _5845_ (.B1(_2535_),
    .VDD(VPWR),
    .Y(_2538_),
    .VSS(VGND),
    .A1(_2536_),
    .A2(_2537_));
 sg13g2_nand2b_1 _5846_ (.Y(_2539_),
    .B(_2538_),
    .A_N(_2534_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5847_ (.Y(_2540_),
    .B(_2522_),
    .A_N(_2539_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5848_ (.Y(_2541_),
    .A(net797),
    .B(net776),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5849_ (.A(net817),
    .B(net787),
    .Y(_2542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5850_ (.B1(net778),
    .VDD(VPWR),
    .Y(_2543_),
    .VSS(VGND),
    .A1(net835),
    .A2(_2473_));
 sg13g2_o21ai_1 _5851_ (.B1(_2541_),
    .VDD(VPWR),
    .Y(_2544_),
    .VSS(VGND),
    .A1(_2542_),
    .A2(_2543_));
 sg13g2_nor2b_1 _5852_ (.A(_2540_),
    .B_N(_2544_),
    .Y(_2545_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5853_ (.A0(\DP_4.matrix[43] ),
    .A1(net832),
    .S(_2472_),
    .X(_2546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5854_ (.Y(_2547_),
    .B1(_2546_),
    .B2(net778),
    .A2(net776),
    .A1(net794),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5855_ (.Y(_2548_),
    .B(_2545_),
    .A_N(_2547_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5856_ (.Y(_2549_),
    .A(net770),
    .B(_2548_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5857_ (.A0(_2516_),
    .A1(_2518_),
    .S(_2549_),
    .X(_0169_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5858_ (.Y(_0172_),
    .A(net1019),
    .B(_2395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5859_ (.A(net1018),
    .B(net771),
    .Y(_2550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5860_ (.B(_2419_),
    .A(_2415_),
    .X(_2551_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5861_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net771),
    .A2(_2551_),
    .Y(_0173_),
    .B1(_2550_));
 sg13g2_nor2_1 _5862_ (.A(net1015),
    .B(net771),
    .Y(_2552_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5863_ (.Y(_2553_),
    .A(_2420_),
    .B(_2422_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5864_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net771),
    .A2(_2553_),
    .Y(_0174_),
    .B1(_2552_));
 sg13g2_nor2_1 _5865_ (.A(net1013),
    .B(net774),
    .Y(_2554_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5866_ (.Y(_2555_),
    .A(_2413_),
    .B(_2423_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5867_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net774),
    .A2(_2555_),
    .Y(_0175_),
    .B1(_2554_));
 sg13g2_nor2_1 _5868_ (.A(net1011),
    .B(net772),
    .Y(_2556_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5869_ (.Y(_2557_),
    .A(_2424_),
    .B(_2426_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5870_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net772),
    .A2(_2557_),
    .Y(_0176_),
    .B1(_2556_));
 sg13g2_xnor2_1 _5871_ (.Y(_2558_),
    .A(_2411_),
    .B(_2427_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5872_ (.A0(_2558_),
    .A1(net1010),
    .S(_2395_),
    .X(_0177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5873_ (.Y(_2559_),
    .A(_2428_),
    .B(_2430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5874_ (.A0(_2559_),
    .A1(net1008),
    .S(_2395_),
    .X(_0178_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5875_ (.Y(_2560_),
    .B(_2409_),
    .A_N(_2431_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5876_ (.B(_2432_),
    .C(_2560_),
    .A(net773),
    .Y(_2561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5877_ (.B1(_2561_),
    .VDD(VPWR),
    .Y(_0179_),
    .VSS(VGND),
    .A1(_2605_),
    .A2(net773));
 sg13g2_xnor2_1 _5878_ (.Y(_0196_),
    .A(net960),
    .B(_2395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5879_ (.A(net956),
    .B(net771),
    .Y(_2562_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5880_ (.B(_2451_),
    .A(_2447_),
    .X(_2563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5881_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net771),
    .A2(_2563_),
    .Y(_0197_),
    .B1(_2562_));
 sg13g2_nor2_1 _5882_ (.A(net954),
    .B(net771),
    .Y(_2564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5883_ (.Y(_2565_),
    .A(_2452_),
    .B(_2454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5884_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net771),
    .A2(_2565_),
    .Y(_0198_),
    .B1(_2564_));
 sg13g2_nor2_1 _5885_ (.A(net952),
    .B(net772),
    .Y(_2566_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5886_ (.Y(_2567_),
    .A(_2445_),
    .B(_2455_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5887_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net772),
    .A2(_2567_),
    .Y(_0199_),
    .B1(_2566_));
 sg13g2_nor2_1 _5888_ (.A(net951),
    .B(net772),
    .Y(_2568_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5889_ (.B(_2460_),
    .A(_2456_),
    .X(_2569_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5890_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net772),
    .A2(_2569_),
    .Y(_0200_),
    .B1(_2568_));
 sg13g2_xnor2_1 _5891_ (.Y(_2570_),
    .A(_2443_),
    .B(_2461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5892_ (.A0(_2570_),
    .A1(net949),
    .S(_2395_),
    .X(_0201_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5893_ (.Y(_2571_),
    .A(_2462_),
    .B(_2464_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5894_ (.A0(_2571_),
    .A1(net948),
    .S(_2395_),
    .X(_0202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5895_ (.Y(_2572_),
    .B(_2441_),
    .A_N(_2465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5896_ (.B(_2466_),
    .C(_2572_),
    .A(net772),
    .Y(_2573_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5897_ (.B1(_2573_),
    .VDD(VPWR),
    .Y(_0203_),
    .VSS(VGND),
    .A1(_2606_),
    .A2(net773));
 sg13g2_xnor2_1 _5898_ (.Y(_0220_),
    .A(net903),
    .B(net767),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5899_ (.A(net901),
    .B(net768),
    .Y(_2574_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5900_ (.Y(_2575_),
    .A(_2492_),
    .B(_2496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5901_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net768),
    .A2(_2575_),
    .Y(_0221_),
    .B1(_2574_));
 sg13g2_nor2_1 _5902_ (.A(net899),
    .B(net768),
    .Y(_2576_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5903_ (.B(_2499_),
    .A(_2497_),
    .X(_2577_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5904_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net768),
    .A2(_2577_),
    .Y(_0222_),
    .B1(_2576_));
 sg13g2_nor2_1 _5905_ (.A(net897),
    .B(net768),
    .Y(_2578_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5906_ (.B(_2500_),
    .A(_2488_),
    .X(_2579_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5907_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net768),
    .A2(_2579_),
    .Y(_0223_),
    .B1(_2578_));
 sg13g2_nor2_1 _5908_ (.A(net895),
    .B(net769),
    .Y(_2580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5909_ (.Y(_2581_),
    .A(_2501_),
    .B(_2503_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5910_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net769),
    .A2(_2581_),
    .Y(_0224_),
    .B1(_2580_));
 sg13g2_xnor2_1 _5911_ (.Y(_2582_),
    .A(_2486_),
    .B(_2504_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5912_ (.A0(_2582_),
    .A1(net894),
    .S(_2479_),
    .X(_0225_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5913_ (.A(net892),
    .B(net770),
    .Y(_2583_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5914_ (.B(_2509_),
    .A(_2505_),
    .X(_2584_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5915_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net770),
    .A2(_2584_),
    .Y(_0226_),
    .B1(_2583_));
 sg13g2_nand2_1 _5916_ (.Y(_2585_),
    .A(net890),
    .B(_2479_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5917_ (.A(_2510_),
    .B_N(_2512_),
    .Y(_2586_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5918_ (.B1(net325),
    .VDD(VPWR),
    .Y(_0227_),
    .VSS(VGND),
    .A1(_2514_),
    .A2(_2586_));
 sg13g2_xnor2_1 _5919_ (.Y(_0244_),
    .A(net847),
    .B(net767),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5920_ (.A(net843),
    .B(net768),
    .Y(_2587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5921_ (.Y(_2588_),
    .A(_2526_),
    .B(_2529_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5922_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net768),
    .A2(_2588_),
    .Y(_0245_),
    .B1(_2587_));
 sg13g2_nor2_1 _5923_ (.A(net841),
    .B(net769),
    .Y(_2589_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5924_ (.B(_2532_),
    .A(_2530_),
    .X(_2590_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5925_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net769),
    .A2(_2590_),
    .Y(_0246_),
    .B1(_2589_));
 sg13g2_nor2_1 _5926_ (.A(net839),
    .B(net769),
    .Y(_2591_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5927_ (.B(_2533_),
    .A(_2524_),
    .X(_2592_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5928_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net769),
    .A2(_2592_),
    .Y(_0247_),
    .B1(_2591_));
 sg13g2_nor2_1 _5929_ (.A(net837),
    .B(net770),
    .Y(_2593_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5930_ (.B(_2538_),
    .A(_2534_),
    .X(_2594_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5931_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2478_),
    .A2(_2594_),
    .Y(_0248_),
    .B1(_2593_));
 sg13g2_xnor2_1 _5932_ (.Y(_2595_),
    .A(_2522_),
    .B(_2539_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5933_ (.A0(_2595_),
    .A1(net836),
    .S(net767),
    .X(_0249_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5934_ (.A(net835),
    .B(net770),
    .Y(_2596_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5935_ (.B(_2544_),
    .A(_2540_),
    .X(_2597_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5936_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net770),
    .A2(_2597_),
    .Y(_0250_),
    .B1(_2596_));
 sg13g2_nand2_1 _5937_ (.Y(_2598_),
    .A(net832),
    .B(net767),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5938_ (.A(_2545_),
    .B_N(_2547_),
    .Y(_2599_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5939_ (.B1(_2598_),
    .VDD(VPWR),
    .Y(_0251_),
    .VSS(VGND),
    .A1(_2549_),
    .A2(_2599_));
 sg13g2_buf_1 _5940_ (.A(net1036),
    .X(_0161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5941_ (.A(net1033),
    .X(_0162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5942_ (.A(net1031),
    .X(_0164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5943_ (.A(net271),
    .X(_0165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5944_ (.A(net1026),
    .X(_0167_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5945_ (.A(net1024),
    .X(_0168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5946_ (.A(net1022),
    .X(_0170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5947_ (.A(net270),
    .X(_0171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5948_ (.A(net1004),
    .X(_0180_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5949_ (.A(net1001),
    .X(_0181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5950_ (.A(net999),
    .X(_0182_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5951_ (.A(net997),
    .X(_0183_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5952_ (.A(net994),
    .X(_0184_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5953_ (.A(net992),
    .X(_0185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5954_ (.A(net990),
    .X(_0186_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5955_ (.A(net278),
    .X(_0187_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5956_ (.A(net273),
    .X(_0188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5957_ (.A(net983),
    .X(_0189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5958_ (.A(net980),
    .X(_0190_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5959_ (.A(net977),
    .X(_0191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5960_ (.A(net974),
    .X(_0192_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5961_ (.A(net971),
    .X(_0193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5962_ (.A(net968),
    .X(_0194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5963_ (.A(net966),
    .X(_0195_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5964_ (.A(net942),
    .X(_0204_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5965_ (.A(net938),
    .X(_0205_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5966_ (.A(net935),
    .X(_0206_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5967_ (.A(net933),
    .X(_0207_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5968_ (.A(net931),
    .X(_0208_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5969_ (.A(net929),
    .X(_0209_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5970_ (.A(net928),
    .X(_0210_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5971_ (.A(net281),
    .X(_0211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5972_ (.A(net924),
    .X(_0212_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5973_ (.A(net272),
    .X(_0213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5974_ (.A(net916),
    .X(_0214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5975_ (.A(net279),
    .X(_0215_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5976_ (.A(net269),
    .X(_0216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5977_ (.A(net910),
    .X(_0217_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5978_ (.A(net908),
    .X(_0218_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5979_ (.A(net906),
    .X(_0219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5980_ (.A(net886),
    .X(_0228_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5981_ (.A(net884),
    .X(_0229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5982_ (.A(net882),
    .X(_0230_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5983_ (.A(net880),
    .X(_0231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5984_ (.A(net878),
    .X(_0232_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5985_ (.A(net876),
    .X(_0233_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5986_ (.A(net873),
    .X(_0234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5987_ (.A(net872),
    .X(_0235_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5988_ (.A(net868),
    .X(_0236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5989_ (.A(net867),
    .X(_0237_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5990_ (.A(net864),
    .X(_0238_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5991_ (.A(net862),
    .X(_0239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5992_ (.A(net274),
    .X(_0240_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5993_ (.A(net277),
    .X(_0241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5994_ (.A(net280),
    .X(_0242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5995_ (.A(net275),
    .X(_0243_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5996_ (.A(net829),
    .X(_0252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5997_ (.A(net826),
    .X(_0253_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5998_ (.A(net823),
    .X(_0254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _5999_ (.A(net821),
    .X(_0255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _6000_ (.A(net819),
    .X(_0256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _6001_ (.A(net818),
    .X(_0257_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _6002_ (.A(net816),
    .X(_0258_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _6003_ (.A(net815),
    .X(_0259_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _6004_ (.A(net813),
    .X(_0260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _6005_ (.A(net810),
    .X(_0261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _6006_ (.A(net805),
    .X(_0262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _6007_ (.A(net803),
    .X(_0263_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _6008_ (.A(net276),
    .X(_0264_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _6009_ (.A(net799),
    .X(_0265_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _6010_ (.A(net797),
    .X(_0266_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _6011_ (.A(net794),
    .X(_0267_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbpq_2 _6012_ (.RESET_B(net1056),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net9),
    .Q(\DP_3.Q_range.out_data[2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6013_ (.RESET_B(net1056),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net10),
    .Q(\DP_3.Q_range.out_data[3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6014_ (.RESET_B(net1056),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net11),
    .Q(\DP_3.Q_range.out_data[4] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6015_ (.RESET_B(net1056),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\DP_3.Q_range.data_plus_4[6] ),
    .Q(\DP_3.Q_range.out_data[5] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6016_ (.RESET_B(net1056),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net12),
    .Q(\DP_3.Q_range.out_data[6] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6017_ (.RESET_B(net1066),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0069_),
    .Q(\mac1.products_ff[0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6018_ (.RESET_B(net1070),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0070_),
    .Q(\mac1.products_ff[1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6019_ (.RESET_B(net1072),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0071_),
    .Q(\mac1.products_ff[2] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6020_ (.RESET_B(net1092),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0072_),
    .Q(\mac1.products_ff[3] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6021_ (.RESET_B(net1092),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0073_),
    .Q(\mac1.products_ff[4] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6022_ (.RESET_B(net1092),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0105_),
    .Q(\mac1.products_ff[5] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6023_ (.RESET_B(net1097),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0112_),
    .Q(\mac1.products_ff[6] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6024_ (.RESET_B(net1097),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0113_),
    .Q(\mac1.products_ff[7] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6025_ (.RESET_B(net1098),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0114_),
    .Q(\mac1.products_ff[8] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6026_ (.RESET_B(net1098),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0115_),
    .Q(\mac1.products_ff[9] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6027_ (.RESET_B(net1098),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0106_),
    .Q(\mac1.products_ff[10] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6028_ (.RESET_B(net1098),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0107_),
    .Q(\mac1.products_ff[11] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6029_ (.RESET_B(net1110),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0108_),
    .Q(\mac1.products_ff[12] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6030_ (.RESET_B(net1111),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0109_),
    .Q(\mac1.products_ff[13] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6031_ (.RESET_B(net1111),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0110_),
    .Q(\mac1.products_ff[14] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6032_ (.RESET_B(net1125),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0111_),
    .Q(\mac1.products_ff[15] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6033_ (.RESET_B(net1066),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0074_),
    .Q(\mac1.products_ff[68] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6034_ (.RESET_B(net1070),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net433),
    .Q(\mac1.products_ff[69] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6035_ (.RESET_B(net1072),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0076_),
    .Q(\mac1.products_ff[70] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6036_ (.RESET_B(net1092),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0077_),
    .Q(\mac1.products_ff[71] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6037_ (.RESET_B(net1097),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0078_),
    .Q(\mac1.products_ff[72] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6038_ (.RESET_B(net1096),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0116_),
    .Q(\mac1.products_ff[73] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6039_ (.RESET_B(net1096),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0123_),
    .Q(\mac1.products_ff[74] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6040_ (.RESET_B(net1108),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0124_),
    .Q(\mac1.products_ff[75] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6041_ (.RESET_B(net1117),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0125_),
    .Q(\mac1.products_ff[76] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6042_ (.RESET_B(net1113),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0126_),
    .Q(\mac1.products_ff[77] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6043_ (.RESET_B(net1113),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0117_),
    .Q(\mac1.products_ff[78] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6044_ (.RESET_B(net1113),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0118_),
    .Q(\mac1.products_ff[79] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6045_ (.RESET_B(net1115),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0119_),
    .Q(\mac1.products_ff[80] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6046_ (.RESET_B(net1114),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0120_),
    .Q(\mac1.products_ff[81] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6047_ (.RESET_B(net1114),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0121_),
    .Q(\mac1.products_ff[82] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6048_ (.RESET_B(net1116),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0122_),
    .Q(\mac1.products_ff[83] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6049_ (.RESET_B(net1093),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0160_),
    .Q(\DP_1.matrix[8] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _6050_ (.RESET_B(net1111),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0161_),
    .Q(\DP_1.matrix[44] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6051_ (.RESET_B(net1068),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0162_),
    .Q(\DP_1.matrix[80] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _6052_ (.RESET_B(net1093),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0163_),
    .Q(\DP_2.matrix[8] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _6053_ (.RESET_B(net1111),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0164_),
    .Q(\DP_2.matrix[44] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6054_ (.RESET_B(net1068),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0165_),
    .Q(\DP_2.matrix[80] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6055_ (.RESET_B(net1101),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0166_),
    .Q(\DP_3.matrix[8] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6056_ (.RESET_B(net1124),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0167_),
    .Q(\DP_3.matrix[44] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6057_ (.RESET_B(net1062),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0168_),
    .Q(\DP_3.matrix[80] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6058_ (.RESET_B(net1101),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0169_),
    .Q(\DP_4.matrix[8] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6059_ (.RESET_B(net1105),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0170_),
    .Q(\DP_4.matrix[44] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6060_ (.RESET_B(net1062),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0171_),
    .Q(\DP_4.matrix[80] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6061_ (.RESET_B(net1073),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0172_),
    .Q(\DP_1.matrix[0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _6062_ (.RESET_B(net1070),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0173_),
    .Q(\DP_1.matrix[1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6063_ (.RESET_B(net1072),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0174_),
    .Q(\DP_1.matrix[2] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6064_ (.RESET_B(net1075),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0175_),
    .Q(\DP_1.matrix[3] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6065_ (.RESET_B(net1075),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0176_),
    .Q(\DP_1.matrix[4] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6066_ (.RESET_B(net1093),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0177_),
    .Q(\DP_1.matrix[5] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _6067_ (.RESET_B(net1093),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0178_),
    .Q(\DP_1.matrix[6] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _6068_ (.RESET_B(net1094),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0179_),
    .Q(\DP_1.matrix[7] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6069_ (.RESET_B(net1108),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0180_),
    .Q(\DP_1.matrix[36] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6070_ (.RESET_B(net1108),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0181_),
    .Q(\DP_1.matrix[37] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6071_ (.RESET_B(net1108),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0182_),
    .Q(\DP_1.matrix[38] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6072_ (.RESET_B(net1118),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0183_),
    .Q(\DP_1.matrix[39] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6073_ (.RESET_B(net1108),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0184_),
    .Q(\DP_1.matrix[40] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _6074_ (.RESET_B(net1111),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0185_),
    .Q(\DP_1.matrix[41] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6075_ (.RESET_B(net1041),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0064_),
    .Q(\mac1.products_ff[136] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _6076_ (.RESET_B(net1111),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0186_),
    .Q(\DP_1.matrix[42] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _6077_ (.RESET_B(net1110),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0187_),
    .Q(\DP_1.matrix[43] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6078_ (.RESET_B(net1049),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0065_),
    .Q(\mac1.products_ff[137] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _6079_ (.RESET_B(net1071),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0188_),
    .Q(\DP_1.matrix[72] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6080_ (.RESET_B(net1071),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0189_),
    .Q(\DP_1.matrix[73] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6081_ (.RESET_B(net1050),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0066_),
    .Q(\mac1.products_ff[138] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6082_ (.RESET_B(net1071),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0190_),
    .Q(\DP_1.matrix[74] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6083_ (.RESET_B(net1067),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0191_),
    .Q(\DP_1.matrix[75] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6084_ (.RESET_B(net1050),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0067_),
    .Q(\mac1.products_ff[139] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6085_ (.RESET_B(net1067),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0192_),
    .Q(\DP_1.matrix[76] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6086_ (.RESET_B(net1067),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0193_),
    .Q(\DP_1.matrix[77] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6087_ (.RESET_B(net1064),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0068_),
    .Q(\mac1.products_ff[140] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _6088_ (.RESET_B(net1073),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0194_),
    .Q(\DP_1.matrix[78] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6089_ (.RESET_B(net1073),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0195_),
    .Q(\DP_1.matrix[79] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6090_ (.RESET_B(net1041),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0094_),
    .Q(\mac1.products_ff[141] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _6091_ (.RESET_B(net1073),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0196_),
    .Q(\DP_2.matrix[0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6092_ (.RESET_B(net1075),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0197_),
    .Q(\DP_2.matrix[1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6093_ (.RESET_B(net1064),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0101_),
    .Q(\mac1.products_ff[142] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _6094_ (.RESET_B(net1076),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net394),
    .Q(\DP_2.matrix[2] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6095_ (.RESET_B(net1072),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0199_),
    .Q(\DP_2.matrix[3] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6096_ (.RESET_B(net1042),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0102_),
    .Q(\mac1.products_ff[143] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6097_ (.RESET_B(net1093),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0200_),
    .Q(\DP_2.matrix[4] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _6098_ (.RESET_B(net1093),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0201_),
    .Q(\DP_2.matrix[5] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6099_ (.RESET_B(net1042),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0103_),
    .Q(\mac1.products_ff[144] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6100_ (.RESET_B(net1093),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0202_),
    .Q(\DP_2.matrix[6] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _6101_ (.RESET_B(net1094),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0203_),
    .Q(\DP_2.matrix[7] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6102_ (.RESET_B(net1047),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0104_),
    .Q(\mac1.products_ff[145] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _6103_ (.RESET_B(net1113),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0204_),
    .Q(\DP_2.matrix[36] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _6104_ (.RESET_B(net1113),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0205_),
    .Q(\DP_2.matrix[37] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6105_ (.RESET_B(net1044),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0095_),
    .Q(\mac1.products_ff[146] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6106_ (.RESET_B(net1109),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0206_),
    .Q(\DP_2.matrix[38] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6107_ (.RESET_B(net1098),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0207_),
    .Q(\DP_2.matrix[39] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6108_ (.RESET_B(net1046),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0096_),
    .Q(\mac1.products_ff[147] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _6109_ (.RESET_B(net1108),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0208_),
    .Q(\DP_2.matrix[40] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6110_ (.RESET_B(net1110),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0209_),
    .Q(\DP_2.matrix[41] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6111_ (.RESET_B(net1051),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0097_),
    .Q(\mac1.products_ff[148] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6112_ (.RESET_B(net1110),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0210_),
    .Q(\DP_2.matrix[42] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _6113_ (.RESET_B(net1110),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0211_),
    .Q(\DP_2.matrix[43] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6114_ (.RESET_B(net1068),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0098_),
    .Q(\mac1.products_ff[149] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6115_ (.RESET_B(net1067),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0212_),
    .Q(\DP_2.matrix[72] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6116_ (.RESET_B(net1069),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0213_),
    .Q(\DP_2.matrix[73] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6117_ (.RESET_B(net1068),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0099_),
    .Q(\mac1.products_ff[150] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6118_ (.RESET_B(net1065),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0214_),
    .Q(\DP_2.matrix[74] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6119_ (.RESET_B(net1071),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0215_),
    .Q(\DP_2.matrix[75] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6120_ (.RESET_B(net1074),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0100_),
    .Q(\mac1.products_ff[151] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6121_ (.RESET_B(net1067),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0216_),
    .Q(\DP_2.matrix[76] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6122_ (.RESET_B(net1073),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0217_),
    .Q(\DP_2.matrix[77] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6123_ (.RESET_B(net1067),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net210),
    .Q(\mac1.sum_lvl1_ff[0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6124_ (.RESET_B(net1073),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0218_),
    .Q(\DP_2.matrix[78] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6125_ (.RESET_B(net1073),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0219_),
    .Q(\DP_2.matrix[79] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6126_ (.RESET_B(net1070),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net182),
    .Q(\mac1.sum_lvl1_ff[1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _6127_ (.RESET_B(net1081),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0220_),
    .Q(\DP_3.matrix[0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6128_ (.RESET_B(net1088),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0221_),
    .Q(\DP_3.matrix[1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6129_ (.RESET_B(net1072),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net186),
    .Q(\mac1.sum_lvl1_ff[2] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6130_ (.RESET_B(net1088),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0222_),
    .Q(\DP_3.matrix[2] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6131_ (.RESET_B(net1088),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0223_),
    .Q(\DP_3.matrix[3] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6132_ (.RESET_B(net1092),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net127),
    .Q(\mac1.sum_lvl1_ff[3] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6133_ (.RESET_B(net1087),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0224_),
    .Q(\DP_3.matrix[4] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6134_ (.RESET_B(net1089),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net417),
    .Q(\DP_3.matrix[5] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6135_ (.RESET_B(net1092),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net147),
    .Q(\mac1.sum_lvl1_ff[4] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _6136_ (.RESET_B(net1089),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0226_),
    .Q(\DP_3.matrix[6] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6137_ (.RESET_B(net1101),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0227_),
    .Q(\DP_3.matrix[7] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6138_ (.RESET_B(net1097),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net80),
    .Q(\mac1.sum_lvl1_ff[5] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6139_ (.RESET_B(net1106),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0228_),
    .Q(\DP_3.matrix[36] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6140_ (.RESET_B(net1122),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0229_),
    .Q(\DP_3.matrix[37] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6141_ (.RESET_B(net1096),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net144),
    .Q(\mac1.sum_lvl1_ff[6] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _6142_ (.RESET_B(net1106),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0230_),
    .Q(\DP_3.matrix[38] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6143_ (.RESET_B(net1124),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0231_),
    .Q(\DP_3.matrix[39] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6144_ (.RESET_B(net1096),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net88),
    .Q(\mac1.sum_lvl1_ff[7] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _6145_ (.RESET_B(net1106),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0232_),
    .Q(\DP_3.matrix[40] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6146_ (.RESET_B(net1122),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0233_),
    .Q(\DP_3.matrix[41] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6147_ (.RESET_B(net1096),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net116),
    .Q(\mac1.sum_lvl1_ff[8] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6148_ (.RESET_B(net1123),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0234_),
    .Q(\DP_3.matrix[42] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6149_ (.RESET_B(net1123),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0235_),
    .Q(\DP_3.matrix[43] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6150_ (.RESET_B(net1098),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net168),
    .Q(\mac1.sum_lvl1_ff[9] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6151_ (.RESET_B(net1081),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0236_),
    .Q(\DP_3.matrix[72] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6152_ (.RESET_B(net1081),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0237_),
    .Q(\DP_3.matrix[73] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6153_ (.RESET_B(net1110),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net142),
    .Q(\mac1.sum_lvl1_ff[10] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6154_ (.RESET_B(net1081),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0238_),
    .Q(\DP_3.matrix[74] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6155_ (.RESET_B(net1082),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0239_),
    .Q(\DP_3.matrix[75] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6156_ (.RESET_B(net1112),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net70),
    .Q(\mac1.sum_lvl1_ff[11] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6157_ (.RESET_B(net1087),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0240_),
    .Q(\DP_3.matrix[76] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6158_ (.RESET_B(net1081),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0241_),
    .Q(\DP_3.matrix[77] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6159_ (.RESET_B(net1111),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net175),
    .Q(\mac1.sum_lvl1_ff[12] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _6160_ (.RESET_B(net1081),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0242_),
    .Q(\DP_3.matrix[78] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6161_ (.RESET_B(net1087),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0243_),
    .Q(\DP_3.matrix[79] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6162_ (.RESET_B(net1116),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net213),
    .Q(\mac1.sum_lvl1_ff[13] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _6163_ (.RESET_B(net1087),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0244_),
    .Q(\DP_4.matrix[0] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6164_ (.RESET_B(net1087),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0245_),
    .Q(\DP_4.matrix[1] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6165_ (.RESET_B(net1125),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net260),
    .Q(\mac1.sum_lvl1_ff[14] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6166_ (.RESET_B(net1087),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0246_),
    .Q(\DP_4.matrix[2] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6167_ (.RESET_B(net1087),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0247_),
    .Q(\DP_4.matrix[3] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6168_ (.RESET_B(net1125),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net231),
    .Q(\mac1.sum_lvl1_ff[15] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6169_ (.RESET_B(net1089),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net415),
    .Q(\DP_4.matrix[4] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6170_ (.RESET_B(net1089),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0249_),
    .Q(\DP_4.matrix[5] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6171_ (.RESET_B(net1101),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0250_),
    .Q(\DP_4.matrix[6] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6172_ (.RESET_B(net1101),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0251_),
    .Q(\DP_4.matrix[7] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6173_ (.RESET_B(net1106),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0252_),
    .Q(\DP_4.matrix[36] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6174_ (.RESET_B(net1121),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0253_),
    .Q(\DP_4.matrix[37] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_1 _6175_ (.RESET_B(net1122),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0254_),
    .Q(\DP_4.matrix[38] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6176_ (.RESET_B(net1106),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0255_),
    .Q(\DP_4.matrix[39] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6177_ (.RESET_B(net1122),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0256_),
    .Q(\DP_4.matrix[40] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6178_ (.RESET_B(net1106),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0257_),
    .Q(\DP_4.matrix[41] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6179_ (.RESET_B(net1123),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0258_),
    .Q(\DP_4.matrix[42] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6180_ (.RESET_B(net1106),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0259_),
    .Q(\DP_4.matrix[43] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6181_ (.RESET_B(net1081),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0260_),
    .Q(\DP_4.matrix[72] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6182_ (.RESET_B(net1082),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0261_),
    .Q(\DP_4.matrix[73] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6183_ (.RESET_B(net1082),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0262_),
    .Q(\DP_4.matrix[74] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6184_ (.RESET_B(net1081),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0263_),
    .Q(\DP_4.matrix[75] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6185_ (.RESET_B(net1087),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0264_),
    .Q(\DP_4.matrix[76] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6186_ (.RESET_B(net1088),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0265_),
    .Q(\DP_4.matrix[77] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6187_ (.RESET_B(net1082),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0266_),
    .Q(\DP_4.matrix[78] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6188_ (.RESET_B(net1088),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0267_),
    .Q(\DP_4.matrix[79] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6189_ (.RESET_B(net1066),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net181),
    .Q(\mac1.sum_lvl1_ff[36] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6190_ (.RESET_B(net1070),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net199),
    .Q(\mac1.sum_lvl1_ff[37] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6191_ (.RESET_B(net1072),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net202),
    .Q(\mac1.sum_lvl1_ff[38] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6192_ (.RESET_B(net1095),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net228),
    .Q(\mac1.sum_lvl1_ff[39] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6193_ (.RESET_B(net1097),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net248),
    .Q(\mac1.sum_lvl1_ff[40] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6194_ (.RESET_B(net1096),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net251),
    .Q(\mac1.sum_lvl1_ff[41] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6195_ (.RESET_B(net1109),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net91),
    .Q(\mac1.sum_lvl1_ff[42] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6196_ (.RESET_B(net1108),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net221),
    .Q(\mac1.sum_lvl1_ff[43] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6197_ (.RESET_B(net1117),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net224),
    .Q(\mac1.sum_lvl1_ff[44] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6198_ (.RESET_B(net1113),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net219),
    .Q(\mac1.sum_lvl1_ff[45] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6199_ (.RESET_B(net1115),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net206),
    .Q(\mac1.sum_lvl1_ff[46] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6200_ (.RESET_B(net1115),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net170),
    .Q(\mac1.sum_lvl1_ff[47] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6201_ (.RESET_B(net1114),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net162),
    .Q(\mac1.sum_lvl1_ff[48] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6202_ (.RESET_B(net1114),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net78),
    .Q(\mac1.sum_lvl1_ff[49] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6203_ (.RESET_B(net1114),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net141),
    .Q(\mac1.sum_lvl1_ff[50] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6204_ (.RESET_B(net1114),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net258),
    .Q(\mac1.sum_lvl1_ff[51] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6205_ (.RESET_B(net1070),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net66),
    .Q(\mac1.sum_lvl2_ff[0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6206_ (.RESET_B(net1070),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net148),
    .Q(\mac1.sum_lvl2_ff[1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6207_ (.RESET_B(net1092),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net130),
    .Q(\mac1.sum_lvl2_ff[2] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6208_ (.RESET_B(net1095),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net120),
    .Q(\mac1.sum_lvl2_ff[3] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6209_ (.RESET_B(net1097),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net118),
    .Q(\mac1.sum_lvl2_ff[4] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6210_ (.RESET_B(net1097),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net140),
    .Q(\mac1.sum_lvl2_ff[5] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6211_ (.RESET_B(net1096),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net76),
    .Q(\mac1.sum_lvl2_ff[6] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6212_ (.RESET_B(net1109),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net92),
    .Q(\mac1.sum_lvl2_ff[7] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6213_ (.RESET_B(net1109),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net50),
    .Q(\mac1.sum_lvl2_ff[8] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6214_ (.RESET_B(net1110),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net246),
    .Q(\mac1.sum_lvl2_ff[9] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6215_ (.RESET_B(net1112),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net113),
    .Q(\mac1.sum_lvl2_ff[10] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6216_ (.RESET_B(net1111),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net77),
    .Q(\mac1.sum_lvl2_ff[11] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6217_ (.RESET_B(net1116),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net95),
    .Q(\mac1.sum_lvl2_ff[12] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6218_ (.RESET_B(net1116),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net58),
    .Q(\mac1.sum_lvl2_ff[13] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6219_ (.RESET_B(net1128),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net133),
    .Q(\mac1.sum_lvl2_ff[14] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6220_ (.RESET_B(net1128),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net169),
    .Q(\mac1.sum_lvl2_ff[15] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6221_ (.RESET_B(net1066),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net146),
    .Q(\mac1.sum_lvl2_ff[19] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6222_ (.RESET_B(net1070),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net149),
    .Q(\mac1.sum_lvl2_ff[20] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6223_ (.RESET_B(net1092),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net106),
    .Q(\mac1.sum_lvl2_ff[21] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6224_ (.RESET_B(net1095),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net171),
    .Q(\mac1.sum_lvl2_ff[22] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6225_ (.RESET_B(net1097),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net143),
    .Q(\mac1.sum_lvl2_ff[23] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _6226_ (.RESET_B(net1096),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net174),
    .Q(\mac1.sum_lvl2_ff[24] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6227_ (.RESET_B(net1109),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net178),
    .Q(\mac1.sum_lvl2_ff[25] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _6228_ (.RESET_B(net1108),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net184),
    .Q(\mac1.sum_lvl2_ff[26] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _6229_ (.RESET_B(net1113),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net159),
    .Q(\mac1.sum_lvl2_ff[27] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _6230_ (.RESET_B(net1113),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net135),
    .Q(\mac1.sum_lvl2_ff[28] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _6231_ (.RESET_B(net1115),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net209),
    .Q(\mac1.sum_lvl2_ff[29] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _6232_ (.RESET_B(net1115),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net241),
    .Q(\mac1.sum_lvl2_ff[30] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _6233_ (.RESET_B(net1114),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net190),
    .Q(\mac1.sum_lvl2_ff[31] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6234_ (.RESET_B(net1114),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net55),
    .Q(\mac1.sum_lvl2_ff[32] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _6235_ (.RESET_B(net1115),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net218),
    .Q(\mac1.sum_lvl2_ff[33] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6236_ (.RESET_B(net1128),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net102),
    .Q(\mac1.sum_lvl2_ff[34] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6237_ (.RESET_B(net1041),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net200),
    .Q(\mac1.sum_lvl2_ff[38] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6238_ (.RESET_B(net1049),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net259),
    .Q(\mac1.sum_lvl2_ff[39] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _6239_ (.RESET_B(net1065),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net256),
    .Q(\mac1.sum_lvl2_ff[40] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6240_ (.RESET_B(net1050),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net93),
    .Q(\mac1.sum_lvl2_ff[41] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6241_ (.RESET_B(net1066),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net249),
    .Q(\mac1.sum_lvl2_ff[42] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6242_ (.RESET_B(net1041),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net158),
    .Q(\mac1.sum_lvl2_ff[43] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6243_ (.RESET_B(net1066),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net203),
    .Q(\mac1.sum_lvl2_ff[44] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6244_ (.RESET_B(net1041),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net165),
    .Q(\mac1.sum_lvl2_ff[45] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6245_ (.RESET_B(net1042),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net177),
    .Q(\mac1.sum_lvl2_ff[46] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6246_ (.RESET_B(net1047),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net83),
    .Q(\mac1.sum_lvl2_ff[47] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6247_ (.RESET_B(net1046),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net205),
    .Q(\mac1.sum_lvl2_ff[48] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6248_ (.RESET_B(net1046),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net167),
    .Q(\mac1.sum_lvl2_ff[49] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6249_ (.RESET_B(net1051),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net180),
    .Q(\mac1.sum_lvl2_ff[50] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6250_ (.RESET_B(net1068),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net134),
    .Q(\mac1.sum_lvl2_ff[51] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6251_ (.RESET_B(net1074),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net254),
    .Q(\mac1.sum_lvl2_ff[52] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6252_ (.RESET_B(net1075),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net136),
    .Q(\mac1.sum_lvl2_ff[53] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6253_ (.RESET_B(net1083),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net242),
    .Q(\mac2.sum_lvl2_ff[38] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6254_ (.RESET_B(net1084),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net87),
    .Q(\mac2.sum_lvl2_ff[39] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6255_ (.RESET_B(net1078),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net150),
    .Q(\mac2.sum_lvl2_ff[40] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6256_ (.RESET_B(net1078),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net124),
    .Q(\mac2.sum_lvl2_ff[41] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6257_ (.RESET_B(net1077),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net229),
    .Q(\mac2.sum_lvl2_ff[42] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6258_ (.RESET_B(net1077),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net208),
    .Q(\mac2.sum_lvl2_ff[43] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6259_ (.RESET_B(net1061),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net195),
    .Q(\mac2.sum_lvl2_ff[44] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6260_ (.RESET_B(net1061),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net132),
    .Q(\mac2.sum_lvl2_ff[45] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6261_ (.RESET_B(net1061),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net117),
    .Q(\mac2.sum_lvl2_ff[46] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6262_ (.RESET_B(net1060),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net154),
    .Q(\mac2.sum_lvl2_ff[47] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6263_ (.RESET_B(net1055),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net112),
    .Q(\mac2.sum_lvl2_ff[48] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6264_ (.RESET_B(net1054),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net115),
    .Q(\mac2.sum_lvl2_ff[49] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6265_ (.RESET_B(net1055),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net255),
    .Q(\mac2.sum_lvl2_ff[50] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6266_ (.RESET_B(net1059),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net194),
    .Q(\mac2.sum_lvl2_ff[51] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6267_ (.RESET_B(net1058),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net264),
    .Q(\mac2.sum_lvl2_ff[52] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6268_ (.RESET_B(net1057),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net235),
    .Q(\mac2.sum_lvl2_ff[53] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6269_ (.RESET_B(net1041),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net155),
    .Q(\mac1.sum_lvl1_ff[72] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _6270_ (.RESET_B(net1049),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net67),
    .Q(\mac1.sum_lvl1_ff[73] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _6271_ (.RESET_B(net1064),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net193),
    .Q(\mac1.sum_lvl1_ff[74] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6272_ (.RESET_B(net1049),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net262),
    .Q(\mac1.sum_lvl1_ff[75] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _6273_ (.RESET_B(net1064),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net57),
    .Q(\mac1.sum_lvl1_ff[76] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6274_ (.RESET_B(net1041),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net204),
    .Q(\mac1.sum_lvl1_ff[77] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6275_ (.RESET_B(net1064),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net152),
    .Q(\mac1.sum_lvl1_ff[78] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6276_ (.RESET_B(net1042),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net145),
    .Q(\mac1.sum_lvl1_ff[79] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6277_ (.RESET_B(net1041),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net201),
    .Q(\mac1.sum_lvl1_ff[80] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6278_ (.RESET_B(net1047),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net119),
    .Q(\mac1.sum_lvl1_ff[81] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6279_ (.RESET_B(net1045),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net250),
    .Q(\mac1.sum_lvl1_ff[82] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6280_ (.RESET_B(net1046),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net166),
    .Q(\mac1.sum_lvl1_ff[83] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6281_ (.RESET_B(net1051),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net238),
    .Q(\mac1.sum_lvl1_ff[84] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6282_ (.RESET_B(net1068),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net212),
    .Q(\mac1.sum_lvl1_ff[85] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6283_ (.RESET_B(net1074),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net103),
    .Q(\mac1.sum_lvl1_ff[86] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6284_ (.RESET_B(net1073),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net211),
    .Q(\mac1.sum_lvl1_ff[87] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6285_ (.RESET_B(net1079),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net74),
    .Q(\mac2.sum_lvl1_ff[72] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6286_ (.RESET_B(net1079),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net71),
    .Q(\mac2.sum_lvl1_ff[73] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6287_ (.RESET_B(net1078),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net164),
    .Q(\mac2.sum_lvl1_ff[74] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6288_ (.RESET_B(net1078),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net54),
    .Q(\mac2.sum_lvl1_ff[75] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6289_ (.RESET_B(net1080),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net65),
    .Q(\mac2.sum_lvl1_ff[76] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6290_ (.RESET_B(net1062),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net191),
    .Q(\mac2.sum_lvl1_ff[77] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6291_ (.RESET_B(net1061),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net139),
    .Q(\mac2.sum_lvl1_ff[78] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6292_ (.RESET_B(net1060),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net232),
    .Q(\mac2.sum_lvl1_ff[79] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6293_ (.RESET_B(net1060),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net187),
    .Q(\mac2.sum_lvl1_ff[80] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6294_ (.RESET_B(net1060),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net198),
    .Q(\mac2.sum_lvl1_ff[81] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6295_ (.RESET_B(net1052),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net215),
    .Q(\mac2.sum_lvl1_ff[82] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6296_ (.RESET_B(net1053),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net261),
    .Q(\mac2.sum_lvl1_ff[83] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6297_ (.RESET_B(net1052),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net253),
    .Q(\mac2.sum_lvl1_ff[84] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6298_ (.RESET_B(net1058),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net105),
    .Q(\mac2.sum_lvl1_ff[85] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6299_ (.RESET_B(net1057),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net173),
    .Q(\mac2.sum_lvl1_ff[86] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6300_ (.RESET_B(net1057),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net257),
    .Q(\mac2.sum_lvl1_ff[87] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6301_ (.RESET_B(net1049),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net107),
    .Q(\mac1.sum_lvl3_ff[20] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6302_ (.RESET_B(net1050),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net100),
    .Q(\mac1.sum_lvl3_ff[21] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6303_ (.RESET_B(net1066),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net72),
    .Q(\mac1.sum_lvl3_ff[22] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6304_ (.RESET_B(net1050),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net89),
    .Q(\mac1.sum_lvl3_ff[23] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6305_ (.RESET_B(net1050),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net263),
    .Q(\mac1.sum_lvl3_ff[24] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6306_ (.RESET_B(net1049),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net68),
    .Q(\mac1.sum_lvl3_ff[25] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _6307_ (.RESET_B(net1067),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net217),
    .Q(\mac1.sum_lvl3_ff[26] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6308_ (.RESET_B(net1050),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net86),
    .Q(\mac1.sum_lvl3_ff[27] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6309_ (.RESET_B(net1049),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net90),
    .Q(\mac1.sum_lvl3_ff[28] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6310_ (.RESET_B(net1051),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net79),
    .Q(\mac1.sum_lvl3_ff[29] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6311_ (.RESET_B(net1047),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net156),
    .Q(\mac1.sum_lvl3_ff[30] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6312_ (.RESET_B(net1046),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net84),
    .Q(\mac1.sum_lvl3_ff[31] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6313_ (.RESET_B(net1068),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net46),
    .Q(\mac1.sum_lvl3_ff[32] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _6314_ (.RESET_B(net1069),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net99),
    .Q(\mac1.sum_lvl3_ff[33] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6315_ (.RESET_B(net1074),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net81),
    .Q(\mac1.sum_lvl3_ff[34] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6316_ (.RESET_B(net1093),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net185),
    .Q(\mac1.sum_lvl3_ff[35] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6317_ (.RESET_B(net1049),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net287),
    .Q(\mac1.sum_lvl3_ff[0] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _6318_ (.RESET_B(net1064),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net357),
    .Q(\mac1.sum_lvl3_ff[1] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6319_ (.RESET_B(net1065),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net382),
    .Q(\mac1.sum_lvl3_ff[2] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _6320_ (.RESET_B(net1076),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net372),
    .Q(\mac1.sum_lvl3_ff[3] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _6321_ (.RESET_B(net1064),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net514),
    .Q(\mac1.sum_lvl3_ff[4] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _6322_ (.RESET_B(net1064),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net507),
    .Q(\mac1.sum_lvl3_ff[5] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _6323_ (.RESET_B(net1066),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net511),
    .Q(\mac1.sum_lvl3_ff[6] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _6324_ (.RESET_B(net1109),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net532),
    .Q(\mac1.sum_lvl3_ff[7] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _6325_ (.RESET_B(net1109),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net378),
    .Q(\mac1.sum_lvl3_ff[8] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _6326_ (.RESET_B(net1110),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net437),
    .Q(\mac1.sum_lvl3_ff[9] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6327_ (.RESET_B(net1046),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0001_),
    .Q(\mac1.sum_lvl3_ff[10] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6328_ (.RESET_B(net1046),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0002_),
    .Q(\mac1.sum_lvl3_ff[11] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _6329_ (.RESET_B(net1075),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net483),
    .Q(\mac1.sum_lvl3_ff[12] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6330_ (.RESET_B(net1068),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0004_),
    .Q(\mac1.sum_lvl3_ff[13] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6331_ (.RESET_B(net1075),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net462),
    .Q(\mac1.sum_lvl3_ff[14] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6332_ (.RESET_B(net1094),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net392),
    .Q(\mac1.sum_lvl3_ff[15] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6333_ (.RESET_B(net1083),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net131),
    .Q(\mac2.sum_lvl3_ff[20] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6334_ (.RESET_B(net1083),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net230),
    .Q(\mac2.sum_lvl3_ff[21] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6335_ (.RESET_B(net1083),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net214),
    .Q(\mac2.sum_lvl3_ff[22] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6336_ (.RESET_B(net1083),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net137),
    .Q(\mac2.sum_lvl3_ff[23] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6337_ (.RESET_B(net1078),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net44),
    .Q(\mac2.sum_lvl3_ff[24] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6338_ (.RESET_B(net1077),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net94),
    .Q(\mac2.sum_lvl3_ff[25] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6339_ (.RESET_B(net1077),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net122),
    .Q(\mac2.sum_lvl3_ff[26] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6340_ (.RESET_B(net1061),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net128),
    .Q(\mac2.sum_lvl3_ff[27] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6341_ (.RESET_B(net1051),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net247),
    .Q(\mac2.sum_lvl3_ff[28] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6342_ (.RESET_B(net1060),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net160),
    .Q(\mac2.sum_lvl3_ff[29] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6343_ (.RESET_B(net1054),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net69),
    .Q(\mac2.sum_lvl3_ff[30] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6344_ (.RESET_B(net1054),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net110),
    .Q(\mac2.sum_lvl3_ff[31] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6345_ (.RESET_B(net1055),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net129),
    .Q(\mac2.sum_lvl3_ff[32] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6346_ (.RESET_B(net1059),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net236),
    .Q(\mac2.sum_lvl3_ff[33] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6347_ (.RESET_B(net1059),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net60),
    .Q(\mac2.sum_lvl3_ff[34] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6348_ (.RESET_B(net1059),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net227),
    .Q(\mac2.sum_lvl3_ff[35] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6349_ (.RESET_B(net1039),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net266),
    .Q(\mac1.total_sum[0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6350_ (.RESET_B(net1040),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net289),
    .Q(\mac1.total_sum[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6351_ (.RESET_B(net1039),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net456),
    .Q(\mac1.total_sum[2] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6352_ (.RESET_B(net1039),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net363),
    .Q(\mac1.total_sum[3] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6353_ (.RESET_B(net1039),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net408),
    .Q(\mac1.total_sum[4] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6354_ (.RESET_B(net1040),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net322),
    .Q(\mac1.total_sum[5] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6355_ (.RESET_B(net1040),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net504),
    .Q(\mac1.total_sum[6] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6356_ (.RESET_B(net1040),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0029_),
    .Q(\mac1.total_sum[7] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6357_ (.RESET_B(net1040),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net422),
    .Q(\mac1.total_sum[8] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6358_ (.RESET_B(net1044),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net360),
    .Q(\mac1.total_sum[9] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6359_ (.RESET_B(net1044),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net350),
    .Q(\mac1.total_sum[10] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6360_ (.RESET_B(net1044),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net365),
    .Q(\mac1.total_sum[11] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6361_ (.RESET_B(net1045),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0019_),
    .Q(\mac1.total_sum[12] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6362_ (.RESET_B(net1045),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net369),
    .Q(\mac1.total_sum[13] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6363_ (.RESET_B(net1045),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net479),
    .Q(\mac1.total_sum[14] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6364_ (.RESET_B(net1046),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net440),
    .Q(\mac1.total_sum[15] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6365_ (.RESET_B(net1078),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0084_),
    .Q(\mac2.products_ff[0] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6366_ (.RESET_B(net1083),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0085_),
    .Q(\mac2.products_ff[1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6367_ (.RESET_B(net1086),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0086_),
    .Q(\mac2.products_ff[2] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6368_ (.RESET_B(net1085),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0087_),
    .Q(\mac2.products_ff[3] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6369_ (.RESET_B(net1099),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0088_),
    .Q(\mac2.products_ff[4] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6370_ (.RESET_B(net1099),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0138_),
    .Q(\mac2.products_ff[5] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6371_ (.RESET_B(net1100),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0145_),
    .Q(\mac2.products_ff[6] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6372_ (.RESET_B(net1102),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0146_),
    .Q(\mac2.products_ff[7] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6373_ (.RESET_B(net1102),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0147_),
    .Q(\mac2.products_ff[8] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6374_ (.RESET_B(net1102),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0148_),
    .Q(\mac2.products_ff[9] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6375_ (.RESET_B(net1104),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0139_),
    .Q(\mac2.products_ff[10] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6376_ (.RESET_B(net1104),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0140_),
    .Q(\mac2.products_ff[11] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6377_ (.RESET_B(net1105),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0141_),
    .Q(\mac2.products_ff[12] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6378_ (.RESET_B(net1105),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0142_),
    .Q(\mac2.products_ff[13] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6379_ (.RESET_B(net1105),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0143_),
    .Q(\mac2.products_ff[14] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6380_ (.RESET_B(net1105),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0144_),
    .Q(\mac2.products_ff[15] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6381_ (.RESET_B(net1079),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0079_),
    .Q(\mac2.products_ff[68] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6382_ (.RESET_B(net1084),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net402),
    .Q(\mac2.products_ff[69] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6383_ (.RESET_B(net1085),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0081_),
    .Q(\mac2.products_ff[70] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6384_ (.RESET_B(net1099),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0082_),
    .Q(\mac2.products_ff[71] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6385_ (.RESET_B(net1100),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0083_),
    .Q(\mac2.products_ff[72] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6386_ (.RESET_B(net1102),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0127_),
    .Q(\mac2.products_ff[73] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6387_ (.RESET_B(net1103),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0134_),
    .Q(\mac2.products_ff[74] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6388_ (.RESET_B(net1119),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0135_),
    .Q(\mac2.products_ff[75] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6389_ (.RESET_B(net1119),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0136_),
    .Q(\mac2.products_ff[76] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6390_ (.RESET_B(net1119),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0137_),
    .Q(\mac2.products_ff[77] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6391_ (.RESET_B(net1121),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0128_),
    .Q(\mac2.products_ff[78] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6392_ (.RESET_B(net1125),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0129_),
    .Q(\mac2.products_ff[79] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6393_ (.RESET_B(net1126),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0130_),
    .Q(\mac2.products_ff[80] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6394_ (.RESET_B(net1126),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0131_),
    .Q(\mac2.products_ff[81] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6395_ (.RESET_B(net1127),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0132_),
    .Q(\mac2.products_ff[82] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6396_ (.RESET_B(net1126),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0133_),
    .Q(\mac2.products_ff[83] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6397_ (.RESET_B(net1079),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net283),
    .Q(\mac2.products_ff[136] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6398_ (.RESET_B(net1080),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net295),
    .Q(\mac2.products_ff[137] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6399_ (.RESET_B(net1080),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0091_),
    .Q(\mac2.products_ff[138] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6400_ (.RESET_B(net1077),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0092_),
    .Q(\mac2.products_ff[139] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6401_ (.RESET_B(net1077),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0093_),
    .Q(\mac2.products_ff[140] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6402_ (.RESET_B(net1062),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0149_),
    .Q(\mac2.products_ff[141] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6403_ (.RESET_B(net1061),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0156_),
    .Q(\mac2.products_ff[142] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6404_ (.RESET_B(net1060),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0157_),
    .Q(\mac2.products_ff[143] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6405_ (.RESET_B(net1060),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0158_),
    .Q(\mac2.products_ff[144] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6406_ (.RESET_B(net1060),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0159_),
    .Q(\mac2.products_ff[145] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6407_ (.RESET_B(net1054),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0150_),
    .Q(\mac2.products_ff[146] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6408_ (.RESET_B(net1052),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0151_),
    .Q(\mac2.products_ff[147] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6409_ (.RESET_B(net1056),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0152_),
    .Q(\mac2.products_ff[148] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6410_ (.RESET_B(net1058),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0153_),
    .Q(\mac2.products_ff[149] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6411_ (.RESET_B(net1057),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0154_),
    .Q(\mac2.products_ff[150] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6412_ (.RESET_B(net1057),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0155_),
    .Q(\mac2.products_ff[151] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6413_ (.RESET_B(net1084),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net176),
    .Q(\mac2.sum_lvl1_ff[0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6414_ (.RESET_B(net1084),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net51),
    .Q(\mac2.sum_lvl1_ff[1] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6415_ (.RESET_B(net1085),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net138),
    .Q(\mac2.sum_lvl1_ff[2] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6416_ (.RESET_B(net1099),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net183),
    .Q(\mac2.sum_lvl1_ff[3] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6417_ (.RESET_B(net1100),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net240),
    .Q(\mac2.sum_lvl1_ff[4] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6418_ (.RESET_B(net1100),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net111),
    .Q(\mac2.sum_lvl1_ff[5] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6419_ (.RESET_B(net1102),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net96),
    .Q(\mac2.sum_lvl1_ff[6] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6420_ (.RESET_B(net1104),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net234),
    .Q(\mac2.sum_lvl1_ff[7] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6421_ (.RESET_B(net1103),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net104),
    .Q(\mac2.sum_lvl1_ff[8] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6422_ (.RESET_B(net1103),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net245),
    .Q(\mac2.sum_lvl1_ff[9] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6423_ (.RESET_B(net1119),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net48),
    .Q(\mac2.sum_lvl1_ff[10] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6424_ (.RESET_B(net1120),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net97),
    .Q(\mac2.sum_lvl1_ff[11] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6425_ (.RESET_B(net1105),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net62),
    .Q(\mac2.sum_lvl1_ff[12] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6426_ (.RESET_B(net1105),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net75),
    .Q(\mac2.sum_lvl1_ff[13] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6427_ (.RESET_B(net1105),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net125),
    .Q(\mac2.sum_lvl1_ff[14] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6428_ (.RESET_B(net1122),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net47),
    .Q(\mac2.sum_lvl1_ff[15] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6429_ (.RESET_B(net1084),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net114),
    .Q(\mac2.sum_lvl1_ff[36] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6430_ (.RESET_B(net1083),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net207),
    .Q(\mac2.sum_lvl1_ff[37] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6431_ (.RESET_B(net1085),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net163),
    .Q(\mac2.sum_lvl1_ff[38] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6432_ (.RESET_B(net1099),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net197),
    .Q(\mac2.sum_lvl1_ff[39] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6433_ (.RESET_B(net1100),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net126),
    .Q(\mac2.sum_lvl1_ff[40] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6434_ (.RESET_B(net1102),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net233),
    .Q(\mac2.sum_lvl1_ff[41] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6435_ (.RESET_B(net1103),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net172),
    .Q(\mac2.sum_lvl1_ff[42] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6436_ (.RESET_B(net1120),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net196),
    .Q(\mac2.sum_lvl1_ff[43] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6437_ (.RESET_B(net1120),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net98),
    .Q(\mac2.sum_lvl1_ff[44] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6438_ (.RESET_B(net1119),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net225),
    .Q(\mac2.sum_lvl1_ff[45] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6439_ (.RESET_B(net1125),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net188),
    .Q(\mac2.sum_lvl1_ff[46] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6440_ (.RESET_B(net1125),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net223),
    .Q(\mac2.sum_lvl1_ff[47] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6441_ (.RESET_B(net1126),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net244),
    .Q(\mac2.sum_lvl1_ff[48] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6442_ (.RESET_B(net1126),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net222),
    .Q(\mac2.sum_lvl1_ff[49] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6443_ (.RESET_B(net1127),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net64),
    .Q(\mac2.sum_lvl1_ff[50] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6444_ (.RESET_B(net1126),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net151),
    .Q(\mac2.sum_lvl1_ff[51] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6445_ (.RESET_B(net1053),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1),
    .Q(\DP_1.I_range.out_data[2] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6446_ (.RESET_B(net1053),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2),
    .Q(\DP_1.I_range.out_data[3] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6447_ (.RESET_B(net1052),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3),
    .Q(\DP_1.I_range.out_data[4] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6448_ (.RESET_B(net1053),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\DP_1.I_range.data_plus_4[6] ),
    .Q(\DP_1.I_range.out_data[5] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6449_ (.RESET_B(net1053),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net4),
    .Q(\DP_1.I_range.out_data[6] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6450_ (.RESET_B(net1084),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net59),
    .Q(\mac2.sum_lvl2_ff[0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6451_ (.RESET_B(net1086),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net101),
    .Q(\mac2.sum_lvl2_ff[1] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6452_ (.RESET_B(net1099),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net161),
    .Q(\mac2.sum_lvl2_ff[2] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6453_ (.RESET_B(net1099),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net157),
    .Q(\mac2.sum_lvl2_ff[3] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6454_ (.RESET_B(net1100),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net85),
    .Q(\mac2.sum_lvl2_ff[4] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6455_ (.RESET_B(net1102),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net109),
    .Q(\mac2.sum_lvl2_ff[5] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6456_ (.RESET_B(net1104),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net153),
    .Q(\mac2.sum_lvl2_ff[6] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6457_ (.RESET_B(net1103),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net61),
    .Q(\mac2.sum_lvl2_ff[7] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6458_ (.RESET_B(net1103),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net45),
    .Q(\mac2.sum_lvl2_ff[8] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6459_ (.RESET_B(net1103),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net189),
    .Q(\mac2.sum_lvl2_ff[9] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6460_ (.RESET_B(net1119),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net52),
    .Q(\mac2.sum_lvl2_ff[10] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6461_ (.RESET_B(net1119),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net56),
    .Q(\mac2.sum_lvl2_ff[11] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6462_ (.RESET_B(net1122),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net41),
    .Q(\mac2.sum_lvl2_ff[12] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6463_ (.RESET_B(net1123),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net42),
    .Q(\mac2.sum_lvl2_ff[13] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6464_ (.RESET_B(net1122),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net43),
    .Q(\mac2.sum_lvl2_ff[14] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6465_ (.RESET_B(net1122),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net220),
    .Q(\mac2.sum_lvl2_ff[15] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6466_ (.RESET_B(net1084),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net49),
    .Q(\mac2.sum_lvl2_ff[19] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6467_ (.RESET_B(net1085),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net192),
    .Q(\mac2.sum_lvl2_ff[20] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6468_ (.RESET_B(net1099),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net63),
    .Q(\mac2.sum_lvl2_ff[21] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6469_ (.RESET_B(net1100),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net73),
    .Q(\mac2.sum_lvl2_ff[22] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6470_ (.RESET_B(net1102),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net53),
    .Q(\mac2.sum_lvl2_ff[23] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _6471_ (.RESET_B(net1103),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net252),
    .Q(\mac2.sum_lvl2_ff[24] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _6472_ (.RESET_B(net1119),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net226),
    .Q(\mac2.sum_lvl2_ff[25] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _6473_ (.RESET_B(net1121),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net237),
    .Q(\mac2.sum_lvl2_ff[26] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _6474_ (.RESET_B(net1121),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net239),
    .Q(\mac2.sum_lvl2_ff[27] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6475_ (.RESET_B(net1121),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net216),
    .Q(\mac2.sum_lvl2_ff[28] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _6476_ (.RESET_B(net1125),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net121),
    .Q(\mac2.sum_lvl2_ff[29] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _6477_ (.RESET_B(net1125),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net82),
    .Q(\mac2.sum_lvl2_ff[30] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _6478_ (.RESET_B(net1126),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net108),
    .Q(\mac2.sum_lvl2_ff[31] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6479_ (.RESET_B(net1127),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net123),
    .Q(\mac2.sum_lvl2_ff[32] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _6480_ (.RESET_B(net1127),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net243),
    .Q(\mac2.sum_lvl2_ff[33] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6481_ (.RESET_B(net1126),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net179),
    .Q(\mac2.sum_lvl2_ff[34] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6482_ (.RESET_B(net1083),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net268),
    .Q(\mac2.sum_lvl3_ff[0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6483_ (.RESET_B(net1085),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net285),
    .Q(\mac2.sum_lvl3_ff[1] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6484_ (.RESET_B(net1085),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net307),
    .Q(\mac2.sum_lvl3_ff[2] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6485_ (.RESET_B(net1085),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net355),
    .Q(\mac2.sum_lvl3_ff[3] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6486_ (.RESET_B(net1078),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net453),
    .Q(\mac2.sum_lvl3_ff[4] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6487_ (.RESET_B(net1078),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net389),
    .Q(\mac2.sum_lvl3_ff[5] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6488_ (.RESET_B(net1077),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net520),
    .Q(\mac2.sum_lvl3_ff[6] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6489_ (.RESET_B(net1077),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0045_),
    .Q(\mac2.sum_lvl3_ff[7] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6490_ (.RESET_B(net1051),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net493),
    .Q(\mac2.sum_lvl3_ff[8] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6491_ (.RESET_B(net1061),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0047_),
    .Q(\mac2.sum_lvl3_ff[9] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6492_ (.RESET_B(net1054),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0033_),
    .Q(\mac2.sum_lvl3_ff[10] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6493_ (.RESET_B(net1054),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0034_),
    .Q(\mac2.sum_lvl3_ff[11] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6494_ (.RESET_B(net1054),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0035_),
    .Q(\mac2.sum_lvl3_ff[12] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6495_ (.RESET_B(net1059),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0036_),
    .Q(\mac2.sum_lvl3_ff[13] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _6496_ (.RESET_B(net1059),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0037_),
    .Q(\mac2.sum_lvl3_ff[14] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6497_ (.RESET_B(net1059),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0038_),
    .Q(\mac2.sum_lvl3_ff[15] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6498_ (.RESET_B(net1039),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net291),
    .Q(\mac2.total_sum[0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6499_ (.RESET_B(net1039),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net450),
    .Q(\mac2.total_sum[1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6500_ (.RESET_B(net1039),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net475),
    .Q(\mac2.total_sum[2] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6501_ (.RESET_B(net1039),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net486),
    .Q(\mac2.total_sum[3] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6502_ (.RESET_B(net1040),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net459),
    .Q(\mac2.total_sum[4] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6503_ (.RESET_B(net1043),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net398),
    .Q(\mac2.total_sum[5] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6504_ (.RESET_B(net1043),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net466),
    .Q(\mac2.total_sum[6] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6505_ (.RESET_B(net1040),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net540),
    .Q(\mac2.total_sum[7] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6506_ (.RESET_B(net1044),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net426),
    .Q(\mac2.total_sum[8] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6507_ (.RESET_B(net1044),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net430),
    .Q(\mac2.total_sum[9] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6508_ (.RESET_B(net1044),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net445),
    .Q(\mac2.total_sum[10] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6509_ (.RESET_B(net1044),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net339),
    .Q(\mac2.total_sum[11] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6510_ (.RESET_B(net1045),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net312),
    .Q(\mac2.total_sum[12] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6511_ (.RESET_B(net1045),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net470),
    .Q(\mac2.total_sum[13] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6512_ (.RESET_B(net1045),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net330),
    .Q(\mac2.total_sum[14] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6513_ (.RESET_B(net1054),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net345),
    .Q(\mac2.total_sum[15] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _6514_ (.RESET_B(net1053),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net5),
    .Q(\DP_1.Q_range.out_data[2] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _6515_ (.RESET_B(net1052),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net6),
    .Q(\DP_1.Q_range.out_data[3] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6516_ (.RESET_B(net1052),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net7),
    .Q(\DP_1.Q_range.out_data[4] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6517_ (.RESET_B(net1052),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\DP_1.Q_range.data_plus_4[6] ),
    .Q(\DP_1.Q_range.out_data[5] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6518_ (.RESET_B(net1052),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net8),
    .Q(\DP_1.Q_range.out_data[6] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _6519_ (.RESET_B(net1056),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net13),
    .Q(\DP_3.I_range.out_data[2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6520_ (.RESET_B(net1056),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net14),
    .Q(\DP_3.I_range.out_data[3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6521_ (.RESET_B(net1057),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net15),
    .Q(\DP_3.I_range.out_data[4] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6522_ (.RESET_B(net1057),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\DP_3.I_range.data_plus_4[6] ),
    .Q(\DP_3.I_range.out_data[5] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6523_ (.RESET_B(net1057),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net16),
    .Q(\DP_3.I_range.out_data[6] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_tiehi heichips25_template_34 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net34));
 sg13g2_tiehi heichips25_template_35 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net35));
 sg13g2_tiehi heichips25_template_36 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net36));
 sg13g2_tiehi heichips25_template_37 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net37));
 sg13g2_tiehi heichips25_template_38 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net38));
 sg13g2_tiehi heichips25_template_39 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net39));
 sg13g2_tiehi heichips25_template_40 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net40));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout767 (.A(_2479_),
    .X(net767),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout768 (.A(net769),
    .X(net768),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout769 (.A(net770),
    .X(net769),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout770 (.A(_2478_),
    .X(net770),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout771 (.A(net774),
    .X(net771),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout772 (.A(net774),
    .X(net772),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout773 (.A(net774),
    .X(net773),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout774 (.A(_2393_),
    .X(net774),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout775 (.A(_2482_),
    .X(net775),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout776 (.A(_2482_),
    .X(net776),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout777 (.A(net779),
    .X(net777),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout778 (.A(net779),
    .X(net778),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout779 (.A(_2471_),
    .X(net779),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout780 (.A(net781),
    .X(net780),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout781 (.A(_2405_),
    .X(net781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout782 (.A(net784),
    .X(net782),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout783 (.A(net784),
    .X(net783),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout784 (.A(_2398_),
    .X(net784),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout785 (.A(_2473_),
    .X(net785),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout786 (.A(net787),
    .X(net786),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout787 (.A(_2472_),
    .X(net787),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout788 (.A(net789),
    .X(net788),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout789 (.A(_2400_),
    .X(net789),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout790 (.A(_2399_),
    .X(net790),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout791 (.A(_2399_),
    .X(net791),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout792 (.A(net794),
    .X(net792),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout793 (.A(net794),
    .X(net793),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout794 (.A(net302),
    .X(net794),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout795 (.A(net797),
    .X(net795),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout796 (.A(net797),
    .X(net796),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout797 (.A(net352),
    .X(net797),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout798 (.A(net799),
    .X(net798),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout799 (.A(net297),
    .X(net799),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout800 (.A(net801),
    .X(net800),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout801 (.A(\DP_4.matrix[76] ),
    .X(net801),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout802 (.A(net803),
    .X(net802),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout803 (.A(net374),
    .X(net803),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout804 (.A(net805),
    .X(net804),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout805 (.A(net308),
    .X(net805),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout806 (.A(net808),
    .X(net806),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout807 (.A(net808),
    .X(net807),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout808 (.A(net809),
    .X(net808),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout809 (.A(net810),
    .X(net809),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout810 (.A(net301),
    .X(net810),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout811 (.A(net812),
    .X(net811),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout812 (.A(net813),
    .X(net812),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout813 (.A(net282),
    .X(net813),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout814 (.A(net815),
    .X(net814),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout815 (.A(net342),
    .X(net815),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout816 (.A(net817),
    .X(net816),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout817 (.A(net500),
    .X(net817),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout818 (.A(net379),
    .X(net818),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout819 (.A(net820),
    .X(net819),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout820 (.A(net496),
    .X(net820),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout821 (.A(net822),
    .X(net821),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout822 (.A(net497),
    .X(net822),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout823 (.A(net319),
    .X(net823),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout824 (.A(\DP_4.matrix[38] ),
    .X(net824),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout825 (.A(net828),
    .X(net825),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout826 (.A(net828),
    .X(net826),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout827 (.A(net828),
    .X(net827),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout828 (.A(net400),
    .X(net828),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout829 (.A(net830),
    .X(net829),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout830 (.A(net373),
    .X(net830),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout831 (.A(net373),
    .X(net831),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout832 (.A(net366),
    .X(net832),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout833 (.A(\DP_4.matrix[7] ),
    .X(net833),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout834 (.A(net835),
    .X(net834),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout835 (.A(net386),
    .X(net835),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout836 (.A(net480),
    .X(net836),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout837 (.A(net414),
    .X(net837),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout838 (.A(\DP_4.matrix[4] ),
    .X(net838),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout839 (.A(net409),
    .X(net839),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout840 (.A(\DP_4.matrix[3] ),
    .X(net840),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout841 (.A(net410),
    .X(net841),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout842 (.A(\DP_4.matrix[2] ),
    .X(net842),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout843 (.A(net404),
    .X(net843),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout844 (.A(\DP_4.matrix[1] ),
    .X(net844),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout845 (.A(net846),
    .X(net845),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout846 (.A(\DP_4.matrix[1] ),
    .X(net846),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout847 (.A(net316),
    .X(net847),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout848 (.A(\DP_4.matrix[0] ),
    .X(net848),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout849 (.A(net850),
    .X(net849),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout850 (.A(\DP_4.matrix[0] ),
    .X(net850),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout851 (.A(net853),
    .X(net851),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout852 (.A(net853),
    .X(net852),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout853 (.A(\DP_3.matrix[79] ),
    .X(net853),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout854 (.A(net855),
    .X(net854),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout855 (.A(\DP_3.matrix[78] ),
    .X(net855),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout856 (.A(net857),
    .X(net856),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout857 (.A(\DP_3.matrix[77] ),
    .X(net857),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout858 (.A(net859),
    .X(net858),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout859 (.A(\DP_3.matrix[76] ),
    .X(net859),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout860 (.A(net862),
    .X(net860),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout861 (.A(net862),
    .X(net861),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout862 (.A(net351),
    .X(net862),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout863 (.A(net865),
    .X(net863),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout864 (.A(net865),
    .X(net864),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout865 (.A(net521),
    .X(net865),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout866 (.A(net867),
    .X(net866),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout867 (.A(net293),
    .X(net867),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout868 (.A(net869),
    .X(net868),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout869 (.A(net489),
    .X(net869),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout870 (.A(net871),
    .X(net870),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout871 (.A(net872),
    .X(net871),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout872 (.A(net299),
    .X(net872),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout873 (.A(net874),
    .X(net873),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout874 (.A(net875),
    .X(net874),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout875 (.A(\DP_3.matrix[42] ),
    .X(net875),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout876 (.A(net340),
    .X(net876),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout877 (.A(\DP_3.matrix[41] ),
    .X(net877),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout878 (.A(net326),
    .X(net878),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout879 (.A(\DP_3.matrix[40] ),
    .X(net879),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout880 (.A(net334),
    .X(net880),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout881 (.A(\DP_3.matrix[39] ),
    .X(net881),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout882 (.A(net331),
    .X(net882),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout883 (.A(\DP_3.matrix[38] ),
    .X(net883),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout884 (.A(net885),
    .X(net884),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout885 (.A(net516),
    .X(net885),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout886 (.A(net323),
    .X(net886),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout887 (.A(\DP_3.matrix[36] ),
    .X(net887),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout888 (.A(net890),
    .X(net888),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout889 (.A(net890),
    .X(net889),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout890 (.A(net324),
    .X(net890),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout891 (.A(net892),
    .X(net891),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout892 (.A(net428),
    .X(net892),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout893 (.A(net894),
    .X(net893),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout894 (.A(net416),
    .X(net894),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout895 (.A(net385),
    .X(net895),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout896 (.A(\DP_3.matrix[4] ),
    .X(net896),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout897 (.A(net898),
    .X(net897),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout898 (.A(net525),
    .X(net898),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout899 (.A(net476),
    .X(net899),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout900 (.A(\DP_3.matrix[2] ),
    .X(net900),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout901 (.A(net902),
    .X(net901),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout902 (.A(net427),
    .X(net902),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout903 (.A(net332),
    .X(net903),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout904 (.A(\DP_3.matrix[0] ),
    .X(net904),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout905 (.A(net906),
    .X(net905),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout906 (.A(net298),
    .X(net906),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout907 (.A(net908),
    .X(net907),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout908 (.A(net300),
    .X(net908),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout909 (.A(net910),
    .X(net909),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout910 (.A(net347),
    .X(net910),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout911 (.A(net912),
    .X(net911),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout912 (.A(\DP_2.matrix[76] ),
    .X(net912),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout913 (.A(net914),
    .X(net913),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout914 (.A(\DP_2.matrix[75] ),
    .X(net914),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout915 (.A(net916),
    .X(net915),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout916 (.A(net413),
    .X(net916),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout917 (.A(net919),
    .X(net917),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout918 (.A(net919),
    .X(net918),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout919 (.A(net920),
    .X(net919),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout920 (.A(\DP_2.matrix[73] ),
    .X(net920),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout921 (.A(net923),
    .X(net921),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout922 (.A(net923),
    .X(net922),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout923 (.A(net924),
    .X(net923),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout924 (.A(net333),
    .X(net924),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout925 (.A(net926),
    .X(net925),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout926 (.A(\DP_2.matrix[43] ),
    .X(net926),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout927 (.A(net928),
    .X(net927),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout928 (.A(net412),
    .X(net928),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout929 (.A(net930),
    .X(net929),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout930 (.A(net494),
    .X(net930),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout931 (.A(net932),
    .X(net931),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout932 (.A(net534),
    .X(net932),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout933 (.A(net934),
    .X(net933),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout934 (.A(net499),
    .X(net934),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout935 (.A(net936),
    .X(net935),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout936 (.A(net488),
    .X(net936),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout937 (.A(net938),
    .X(net937),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout938 (.A(net939),
    .X(net938),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout939 (.A(net431),
    .X(net939),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout940 (.A(net431),
    .X(net940),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout941 (.A(net942),
    .X(net941),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout942 (.A(net405),
    .X(net942),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout943 (.A(net405),
    .X(net943),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout944 (.A(\DP_2.matrix[7] ),
    .X(net944),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout945 (.A(\DP_2.matrix[7] ),
    .X(net945),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout946 (.A(net948),
    .X(net946),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout947 (.A(net948),
    .X(net947),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout948 (.A(net411),
    .X(net948),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout949 (.A(net472),
    .X(net949),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout950 (.A(net951),
    .X(net950),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout951 (.A(net418),
    .X(net951),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout952 (.A(net399),
    .X(net952),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout953 (.A(\DP_2.matrix[3] ),
    .X(net953),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout954 (.A(net393),
    .X(net954),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout955 (.A(\DP_2.matrix[2] ),
    .X(net955),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout956 (.A(net959),
    .X(net956),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout957 (.A(net959),
    .X(net957),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout958 (.A(net959),
    .X(net958),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout959 (.A(net523),
    .X(net959),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout960 (.A(net341),
    .X(net960),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout961 (.A(net962),
    .X(net961),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout962 (.A(net963),
    .X(net962),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout963 (.A(\DP_2.matrix[0] ),
    .X(net963),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout964 (.A(net965),
    .X(net964),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout965 (.A(net966),
    .X(net965),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout966 (.A(net304),
    .X(net966),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout967 (.A(net968),
    .X(net967),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout968 (.A(net315),
    .X(net968),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout969 (.A(net970),
    .X(net969),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout970 (.A(net971),
    .X(net970),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout971 (.A(net327),
    .X(net971),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout972 (.A(net973),
    .X(net972),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout973 (.A(net974),
    .X(net973),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout974 (.A(net318),
    .X(net974),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout975 (.A(net977),
    .X(net975),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout976 (.A(net977),
    .X(net976),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout977 (.A(net303),
    .X(net977),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout978 (.A(net980),
    .X(net978),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout979 (.A(net980),
    .X(net979),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout980 (.A(net309),
    .X(net980),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout981 (.A(net983),
    .X(net981),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout982 (.A(net983),
    .X(net982),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout983 (.A(net296),
    .X(net983),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout984 (.A(net985),
    .X(net984),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout985 (.A(net273),
    .X(net985),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout986 (.A(net987),
    .X(net986),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout987 (.A(net988),
    .X(net987),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout988 (.A(\DP_1.matrix[43] ),
    .X(net988),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout989 (.A(net990),
    .X(net989),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout990 (.A(net346),
    .X(net990),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout991 (.A(net992),
    .X(net991),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout992 (.A(net993),
    .X(net992),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout993 (.A(net544),
    .X(net993),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout994 (.A(net996),
    .X(net994),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout995 (.A(net996),
    .X(net995),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout996 (.A(net487),
    .X(net996),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout997 (.A(net998),
    .X(net997),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout998 (.A(net498),
    .X(net998),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout999 (.A(net1000),
    .X(net999),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1000 (.A(net495),
    .X(net1000),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1001 (.A(net1002),
    .X(net1001),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1002 (.A(net515),
    .X(net1002),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1003 (.A(net395),
    .X(net1003),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1004 (.A(net395),
    .X(net1004),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1005 (.A(net1006),
    .X(net1005),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1006 (.A(net447),
    .X(net1006),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1007 (.A(net1008),
    .X(net1007),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1008 (.A(net446),
    .X(net1008),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1009 (.A(net1010),
    .X(net1009),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1010 (.A(net448),
    .X(net1010),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1011 (.A(net1012),
    .X(net1011),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1012 (.A(net526),
    .X(net1012),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1013 (.A(net1014),
    .X(net1013),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1014 (.A(net524),
    .X(net1014),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1015 (.A(net471),
    .X(net1015),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1016 (.A(\DP_1.matrix[2] ),
    .X(net1016),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1017 (.A(net1018),
    .X(net1017),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1018 (.A(net441),
    .X(net1018),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1019 (.A(net335),
    .X(net1019),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1020 (.A(\DP_1.matrix[0] ),
    .X(net1020),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1021 (.A(\DP_4.matrix[80] ),
    .X(net1021),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1022 (.A(net383),
    .X(net1022),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1023 (.A(net541),
    .X(net1023),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1024 (.A(net317),
    .X(net1024),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1025 (.A(\DP_3.matrix[80] ),
    .X(net1025),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1026 (.A(net313),
    .X(net1026),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1027 (.A(\DP_3.matrix[44] ),
    .X(net1027),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1028 (.A(net536),
    .X(net1028),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1029 (.A(\DP_3.matrix[8] ),
    .X(net1029),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1030 (.A(\DP_2.matrix[80] ),
    .X(net1030),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1031 (.A(net384),
    .X(net1031),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1032 (.A(net535),
    .X(net1032),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1033 (.A(net314),
    .X(net1033),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1034 (.A(\DP_1.matrix[80] ),
    .X(net1034),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1035 (.A(net1036),
    .X(net1035),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1036 (.A(net403),
    .X(net1036),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1037 (.A(net522),
    .X(net1037),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1038 (.A(\DP_1.matrix[8] ),
    .X(net1038),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1039 (.A(net1040),
    .X(net1039),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1040 (.A(net1043),
    .X(net1040),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1041 (.A(net1043),
    .X(net1041),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1042 (.A(net1043),
    .X(net1042),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1043 (.A(net1048),
    .X(net1043),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1044 (.A(net1048),
    .X(net1044),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1045 (.A(net1048),
    .X(net1045),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1046 (.A(net1047),
    .X(net1046),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1047 (.A(net1048),
    .X(net1047),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1048 (.A(net1063),
    .X(net1048),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1049 (.A(net1050),
    .X(net1049),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1050 (.A(net1051),
    .X(net1050),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1051 (.A(net1063),
    .X(net1051),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1052 (.A(net1053),
    .X(net1052),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1053 (.A(net1055),
    .X(net1053),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1054 (.A(net1055),
    .X(net1054),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1055 (.A(net1063),
    .X(net1055),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1056 (.A(net1058),
    .X(net1056),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1057 (.A(net1058),
    .X(net1057),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1058 (.A(net1059),
    .X(net1058),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1059 (.A(net1063),
    .X(net1059),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1060 (.A(net1061),
    .X(net1060),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1061 (.A(net1062),
    .X(net1061),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1062 (.A(net1063),
    .X(net1062),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1063 (.A(net1091),
    .X(net1063),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1064 (.A(net1065),
    .X(net1064),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1065 (.A(net1069),
    .X(net1065),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1066 (.A(net1067),
    .X(net1066),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1067 (.A(net1069),
    .X(net1067),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1068 (.A(net1069),
    .X(net1068),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1069 (.A(net1091),
    .X(net1069),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1070 (.A(net1072),
    .X(net1070),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1071 (.A(net1072),
    .X(net1071),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1072 (.A(net1076),
    .X(net1072),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1073 (.A(net1075),
    .X(net1073),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1074 (.A(net1075),
    .X(net1074),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1075 (.A(net1076),
    .X(net1075),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1076 (.A(net1091),
    .X(net1076),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1077 (.A(net1080),
    .X(net1077),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1078 (.A(net1080),
    .X(net1078),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1079 (.A(net1080),
    .X(net1079),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1080 (.A(net1090),
    .X(net1080),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1081 (.A(net1090),
    .X(net1081),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1082 (.A(net1090),
    .X(net1082),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1083 (.A(net1086),
    .X(net1083),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1084 (.A(net1086),
    .X(net1084),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1085 (.A(net1086),
    .X(net1085),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1086 (.A(net1090),
    .X(net1086),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1087 (.A(net1088),
    .X(net1087),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1088 (.A(net1089),
    .X(net1088),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1089 (.A(net1090),
    .X(net1089),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1090 (.A(net1091),
    .X(net1090),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1091 (.A(rst_n),
    .X(net1091),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1092 (.A(net1095),
    .X(net1092),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1093 (.A(net1094),
    .X(net1093),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1094 (.A(net1095),
    .X(net1094),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1095 (.A(net1107),
    .X(net1095),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1096 (.A(net1098),
    .X(net1096),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1097 (.A(net1098),
    .X(net1097),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1098 (.A(net1107),
    .X(net1098),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1099 (.A(net1101),
    .X(net1099),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1100 (.A(net1101),
    .X(net1100),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1101 (.A(net1107),
    .X(net1101),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1102 (.A(net1104),
    .X(net1102),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1103 (.A(net1104),
    .X(net1103),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1104 (.A(net1107),
    .X(net1104),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1105 (.A(net1106),
    .X(net1105),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1106 (.A(net1107),
    .X(net1106),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1107 (.A(rst_n),
    .X(net1107),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1108 (.A(net1109),
    .X(net1108),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1109 (.A(net1118),
    .X(net1109),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1110 (.A(net1112),
    .X(net1110),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1111 (.A(net1112),
    .X(net1111),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1112 (.A(net1118),
    .X(net1112),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1113 (.A(net1117),
    .X(net1113),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1114 (.A(net1115),
    .X(net1114),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1115 (.A(net1116),
    .X(net1115),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1116 (.A(net1117),
    .X(net1116),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1117 (.A(net1118),
    .X(net1117),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1118 (.A(net1129),
    .X(net1118),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1119 (.A(net1120),
    .X(net1119),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1120 (.A(net1121),
    .X(net1120),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1121 (.A(net1129),
    .X(net1121),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1122 (.A(net1124),
    .X(net1122),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1123 (.A(net1124),
    .X(net1123),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1124 (.A(net1129),
    .X(net1124),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1125 (.A(net1128),
    .X(net1125),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1126 (.A(net1127),
    .X(net1126),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1127 (.A(net1128),
    .X(net1127),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1128 (.A(net1129),
    .X(net1128),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1129 (.A(rst_n),
    .X(net1129),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input14 (.A(uio_in[5]),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input16 (.A(uio_in[7]),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uio_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uio_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uio_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uio_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uo_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uo_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uo_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output30 (.A(net30),
    .X(uo_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output31 (.A(net31),
    .X(uo_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output32 (.A(net32),
    .X(uo_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tiehi heichips25_template_33 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net33));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_2_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_3_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_5_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_6_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_7_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_8_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_9_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_10_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_11_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_12_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_13_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_14_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_15_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_16_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_17_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_18_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_19_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_20_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_21_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_22_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_23_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_24_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_25_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_26_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_27_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_28_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_29_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_30_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_31_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_32_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_33_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_34_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_35_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_36_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_37_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_39_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_40_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_41_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_42_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_43_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_44_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_45_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_46_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_47_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_48_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_49_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_50_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_51_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_52_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_53_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_54_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_55_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_56_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_57_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_58_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_59_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_60_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_61_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_62_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_63_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_64_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_65_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_66_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_67_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload0 (.A(clknet_4_1_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload1 (.A(clknet_4_2_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload2 (.A(clknet_4_3_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload3 (.A(clknet_4_5_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload4 (.A(clknet_4_6_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload5 (.A(clknet_4_7_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload6 (.A(clknet_4_9_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload7 (.A(clknet_4_10_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload8 (.A(clknet_4_11_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload9 (.A(clknet_4_13_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload10 (.A(clknet_4_14_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload11 (.A(clknet_4_15_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload12 (.A(clknet_leaf_65_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload13 (.VDD(VPWR),
    .A(clknet_leaf_28_clk),
    .VSS(VGND));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_44_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload15 (.A(clknet_leaf_57_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_50_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload17 (.VDD(VPWR),
    .A(clknet_leaf_48_clk),
    .VSS(VGND));
 sg13g2_inv_2 clkload18 (.A(clknet_leaf_31_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_32_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload20 (.VDD(VPWR),
    .A(clknet_leaf_35_clk),
    .VSS(VGND));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_37_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd3_1 hold1 (.A(\mac2.sum_lvl1_ff[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold2 (.A(\mac2.sum_lvl1_ff[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold3 (.A(\mac2.sum_lvl1_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold4 (.A(\mac2.sum_lvl2_ff[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold5 (.A(\mac2.sum_lvl1_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold6 (.A(\mac1.sum_lvl2_ff[50] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold7 (.A(\mac2.products_ff[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold8 (.A(\mac2.products_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold9 (.A(\mac2.sum_lvl1_ff[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold10 (.A(\mac1.sum_lvl1_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold11 (.A(\mac2.products_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold12 (.A(\mac2.sum_lvl1_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold13 (.A(\mac2.sum_lvl1_ff[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold14 (.A(\mac2.products_ff[139] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold15 (.A(\mac1.sum_lvl1_ff[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold16 (.A(\mac2.sum_lvl1_ff[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold17 (.A(\mac1.products_ff[140] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold18 (.A(\mac1.sum_lvl1_ff[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold19 (.A(\mac2.sum_lvl1_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold20 (.A(\mac2.sum_lvl2_ff[52] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold21 (.A(\mac2.sum_lvl1_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold22 (.A(\mac2.products_ff[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold23 (.A(\mac2.sum_lvl1_ff[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold24 (.A(\mac2.products_ff[82] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold25 (.A(\mac2.products_ff[140] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold26 (.A(\mac1.sum_lvl1_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold27 (.A(\mac1.products_ff[137] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold28 (.A(\mac1.sum_lvl2_ff[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold29 (.A(\mac2.sum_lvl2_ff[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold30 (.A(\mac1.products_ff[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold31 (.A(\mac2.products_ff[137] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold32 (.A(\mac1.sum_lvl2_ff[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold33 (.A(\mac2.sum_lvl1_ff[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold34 (.A(\mac2.products_ff[136] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold35 (.A(\mac2.products_ff[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold36 (.A(\mac1.sum_lvl1_ff[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold37 (.A(\mac1.sum_lvl1_ff[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold38 (.A(\mac1.products_ff[81] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold39 (.A(\mac1.sum_lvl2_ff[47] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold40 (.A(\mac1.products_ff[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold41 (.A(\mac1.sum_lvl2_ff[52] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold42 (.A(\mac2.sum_lvl1_ff[47] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold43 (.A(\mac1.sum_lvl1_ff[81] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold44 (.A(\mac1.sum_lvl2_ff[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold45 (.A(\mac2.sum_lvl1_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold46 (.A(\mac1.sum_lvl2_ff[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold47 (.A(\mac2.sum_lvl1_ff[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold48 (.A(\mac1.products_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold49 (.A(\mac1.sum_lvl2_ff[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold50 (.A(\mac1.sum_lvl2_ff[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold51 (.A(\mac1.products_ff[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold52 (.A(\mac1.sum_lvl1_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold53 (.A(\mac1.sum_lvl1_ff[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold54 (.A(\mac2.sum_lvl2_ff[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold55 (.A(\mac1.sum_lvl1_ff[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold56 (.A(\mac2.products_ff[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold57 (.A(\mac2.products_ff[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold58 (.A(\mac2.products_ff[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold59 (.A(\mac1.sum_lvl2_ff[51] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold60 (.A(\mac1.sum_lvl2_ff[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold61 (.A(\mac2.sum_lvl1_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold62 (.A(\mac1.sum_lvl1_ff[51] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold63 (.A(\mac1.products_ff[150] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold64 (.A(\mac2.products_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold65 (.A(\mac2.products_ff[149] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold66 (.A(\mac1.sum_lvl1_ff[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold67 (.A(\mac1.sum_lvl2_ff[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold68 (.A(\mac2.sum_lvl1_ff[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold69 (.A(\mac2.sum_lvl1_ff[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold70 (.A(\mac2.sum_lvl2_ff[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold71 (.A(\mac2.products_ff[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold72 (.A(\mac2.sum_lvl1_ff[82] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold73 (.A(\mac1.sum_lvl1_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold74 (.A(\mac2.products_ff[68] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold75 (.A(\mac2.sum_lvl1_ff[83] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold76 (.A(\mac1.products_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold77 (.A(\mac2.sum_lvl1_ff[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold78 (.A(\mac1.sum_lvl1_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold79 (.A(\mac1.products_ff[145] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold80 (.A(\mac1.sum_lvl1_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold81 (.A(\mac2.sum_lvl1_ff[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold82 (.A(\mac2.sum_lvl2_ff[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold83 (.A(\mac2.sum_lvl1_ff[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold84 (.A(\mac2.sum_lvl1_ff[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold85 (.A(\mac2.products_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold86 (.A(\mac2.products_ff[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold87 (.A(\mac1.products_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold88 (.A(\mac2.sum_lvl2_ff[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold89 (.A(\mac2.sum_lvl2_ff[50] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold90 (.A(\mac1.sum_lvl1_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold91 (.A(\mac2.sum_lvl2_ff[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold92 (.A(\mac2.sum_lvl1_ff[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold93 (.A(\mac1.sum_lvl1_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold94 (.A(\mac1.sum_lvl1_ff[85] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold95 (.A(\mac1.sum_lvl1_ff[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold96 (.A(\mac1.sum_lvl1_ff[87] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold97 (.A(\mac2.sum_lvl2_ff[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold98 (.A(\mac2.products_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold99 (.A(\mac2.products_ff[142] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold100 (.A(\mac1.sum_lvl1_ff[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold101 (.A(\mac1.products_ff[82] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold102 (.A(\mac1.products_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold103 (.A(\mac1.sum_lvl1_ff[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold104 (.A(\mac1.products_ff[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold105 (.A(\mac1.products_ff[143] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold106 (.A(\mac1.sum_lvl1_ff[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold107 (.A(\mac1.products_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold108 (.A(\mac1.sum_lvl1_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold109 (.A(\mac1.sum_lvl1_ff[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold110 (.A(\mac2.sum_lvl1_ff[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold111 (.A(\mac2.products_ff[83] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold112 (.A(\mac1.products_ff[142] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold113 (.A(\mac2.sum_lvl1_ff[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold114 (.A(\mac2.sum_lvl1_ff[81] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold115 (.A(\mac1.products_ff[136] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold116 (.A(\mac1.sum_lvl2_ff[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold117 (.A(\mac2.sum_lvl1_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold118 (.A(\mac1.sum_lvl1_ff[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold119 (.A(\mac1.sum_lvl1_ff[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold120 (.A(\mac2.sum_lvl2_ff[47] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold121 (.A(\mac2.sum_lvl1_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold122 (.A(\mac1.products_ff[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold123 (.A(\mac2.products_ff[70] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold124 (.A(\mac2.products_ff[138] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold125 (.A(\mac1.sum_lvl1_ff[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold126 (.A(\mac1.products_ff[147] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold127 (.A(\mac1.sum_lvl1_ff[83] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold128 (.A(\mac1.products_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold129 (.A(\mac1.sum_lvl1_ff[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold130 (.A(\mac1.products_ff[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold131 (.A(\mac1.sum_lvl1_ff[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold132 (.A(\mac2.products_ff[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold133 (.A(\mac2.products_ff[150] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold134 (.A(\mac1.sum_lvl1_ff[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold135 (.A(\mac1.products_ff[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold136 (.A(\mac2.products_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold137 (.A(\mac1.sum_lvl1_ff[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold138 (.A(\mac1.sum_lvl1_ff[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold139 (.A(\mac2.sum_lvl1_ff[51] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold140 (.A(\mac1.sum_lvl1_ff[84] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold141 (.A(\mac1.products_ff[68] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold142 (.A(\mac1.products_ff[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold143 (.A(\mac2.products_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold144 (.A(\mac1.sum_lvl1_ff[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold145 (.A(\mac1.sum_lvl2_ff[53] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold146 (.A(\mac1.products_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold147 (.A(\mac2.products_ff[144] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold148 (.A(\mac2.products_ff[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold149 (.A(\mac2.sum_lvl1_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold150 (.A(\mac1.sum_lvl1_ff[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold151 (.A(\mac2.products_ff[141] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold152 (.A(\mac2.sum_lvl1_ff[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold153 (.A(\mac1.products_ff[138] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold154 (.A(\mac2.sum_lvl1_ff[85] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold155 (.A(\mac2.sum_lvl1_ff[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold156 (.A(\mac2.products_ff[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold157 (.A(\mac2.products_ff[71] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold158 (.A(\mac2.products_ff[145] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold159 (.A(\mac1.products_ff[69] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold160 (.A(\mac1.sum_lvl1_ff[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold161 (.A(\mac1.products_ff[144] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold162 (.A(\mac1.products_ff[70] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold163 (.A(\mac1.sum_lvl1_ff[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold164 (.A(\mac1.products_ff[141] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold165 (.A(\mac1.sum_lvl1_ff[82] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold166 (.A(\mac1.products_ff[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold167 (.A(\mac2.products_ff[69] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold168 (.A(\mac2.sum_lvl1_ff[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold169 (.A(\mac1.sum_lvl1_ff[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold170 (.A(\mac1.products_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold171 (.A(\mac1.products_ff[151] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold172 (.A(\mac1.products_ff[149] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold173 (.A(\mac1.products_ff[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold174 (.A(\mac2.sum_lvl2_ff[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold175 (.A(\mac2.products_ff[146] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold176 (.A(\mac2.sum_lvl1_ff[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold177 (.A(\mac1.sum_lvl2_ff[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold178 (.A(\mac1.sum_lvl1_ff[50] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold179 (.A(\mac1.products_ff[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold180 (.A(\mac2.sum_lvl1_ff[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold181 (.A(\mac1.products_ff[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold182 (.A(\mac2.products_ff[81] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold183 (.A(\mac2.products_ff[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold184 (.A(\mac1.products_ff[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold185 (.A(\mac2.products_ff[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold186 (.A(\mac2.sum_lvl1_ff[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold187 (.A(\mac2.sum_lvl2_ff[53] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold188 (.A(\mac1.products_ff[71] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold189 (.A(\mac2.sum_lvl1_ff[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold190 (.A(\mac2.sum_lvl2_ff[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold191 (.A(\mac1.products_ff[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold192 (.A(\mac2.products_ff[143] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold193 (.A(\mac2.products_ff[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold194 (.A(\mac2.products_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold195 (.A(\mac2.sum_lvl1_ff[87] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold196 (.A(\mac2.sum_lvl2_ff[51] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold197 (.A(\mac2.sum_lvl1_ff[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold198 (.A(\mac1.products_ff[148] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold199 (.A(\mac2.sum_lvl1_ff[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold200 (.A(\mac2.products_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold201 (.A(\mac1.sum_lvl1_ff[47] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold202 (.A(\mac2.sum_lvl1_ff[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold203 (.A(\mac2.sum_lvl1_ff[50] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold204 (.A(\mac2.products_ff[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold205 (.A(\mac2.products_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold206 (.A(\mac1.sum_lvl1_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold207 (.A(\mac2.sum_lvl2_ff[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold208 (.A(\mac1.products_ff[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold209 (.A(\mac1.sum_lvl1_ff[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold210 (.A(\mac1.products_ff[146] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold211 (.A(\mac1.products_ff[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold212 (.A(\mac2.sum_lvl1_ff[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold213 (.A(\mac2.products_ff[148] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold214 (.A(\mac1.sum_lvl1_ff[86] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold215 (.A(\mac2.sum_lvl1_ff[84] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold216 (.A(\mac1.sum_lvl1_ff[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold217 (.A(\mac2.products_ff[151] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold218 (.A(\mac1.products_ff[83] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold219 (.A(\mac1.sum_lvl1_ff[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold220 (.A(\mac1.products_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold221 (.A(\mac2.products_ff[147] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold222 (.A(\mac1.products_ff[139] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold223 (.A(\mac1.sum_lvl2_ff[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold224 (.A(\mac2.sum_lvl1_ff[86] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold225 (.A(\mac1.sum_lvl3_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0016_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold227 (.A(\mac2.sum_lvl2_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0032_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold229 (.A(\DP_2.matrix[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold230 (.A(\DP_4.matrix[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold231 (.A(\DP_2.matrix[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold232 (.A(\DP_2.matrix[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold233 (.A(\DP_1.matrix[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold234 (.A(\DP_3.matrix[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold235 (.A(\DP_3.matrix[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold236 (.A(\DP_4.matrix[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold237 (.A(\DP_3.matrix[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold238 (.A(\DP_1.matrix[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold239 (.A(\DP_2.matrix[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold240 (.A(\DP_3.matrix[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold241 (.A(\DP_2.matrix[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold242 (.A(\DP_4.matrix[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0089_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold244 (.A(\mac2.sum_lvl2_ff[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0039_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold246 (.A(\mac1.sum_lvl2_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0000_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold248 (.A(\mac1.sum_lvl3_ff[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0023_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold250 (.A(\mac2.sum_lvl3_ff[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0048_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold252 (.A(\DP_2.matrix[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold253 (.A(\DP_3.matrix[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold254 (.A(_1738_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0090_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold256 (.A(\DP_1.matrix[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold257 (.A(\DP_4.matrix[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold258 (.A(\DP_2.matrix[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold259 (.A(\DP_3.matrix[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold260 (.A(\DP_2.matrix[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold261 (.A(\DP_4.matrix[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold262 (.A(\DP_4.matrix[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold263 (.A(\DP_1.matrix[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold264 (.A(\DP_1.matrix[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold265 (.A(\mac2.sum_lvl2_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold266 (.A(_2229_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0040_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold268 (.A(\DP_4.matrix[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold269 (.A(\DP_1.matrix[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold270 (.A(\mac2.sum_lvl3_ff[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold271 (.A(_2321_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold272 (.A(_0051_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold273 (.A(\DP_3.matrix[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold274 (.A(\DP_1.matrix[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold275 (.A(\DP_1.matrix[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold276 (.A(\DP_4.matrix[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold277 (.A(\DP_3.matrix[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold278 (.A(\DP_1.matrix[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold279 (.A(\DP_4.matrix[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold280 (.A(\mac1.sum_lvl3_ff[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold281 (.A(_2180_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0027_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold283 (.A(\DP_3.matrix[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold284 (.A(\DP_3.matrix[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold285 (.A(_2585_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold286 (.A(\DP_3.matrix[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold287 (.A(\DP_1.matrix[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold288 (.A(\mac2.sum_lvl3_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold289 (.A(_2332_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0053_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold291 (.A(\DP_3.matrix[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold292 (.A(\DP_3.matrix[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold293 (.A(\DP_2.matrix[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold294 (.A(\DP_3.matrix[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold295 (.A(\DP_1.matrix[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold296 (.A(\mac2.sum_lvl3_ff[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold297 (.A(_2311_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold298 (.A(_2318_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold299 (.A(_0050_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold300 (.A(\DP_3.matrix[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold301 (.A(\DP_2.matrix[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold302 (.A(\DP_4.matrix[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold303 (.A(\mac2.sum_lvl3_ff[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold304 (.A(_2334_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0054_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold306 (.A(\DP_1.matrix[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold307 (.A(\DP_2.matrix[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold308 (.A(\mac1.sum_lvl3_ff[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold309 (.A(_2200_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold310 (.A(_0017_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold311 (.A(\DP_3.matrix[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold312 (.A(\DP_4.matrix[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold313 (.A(\mac2.sum_lvl2_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold314 (.A(_2232_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold315 (.A(_0041_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold316 (.A(\mac1.sum_lvl2_ff[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0007_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold318 (.A(\mac1.sum_lvl3_ff[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold319 (.A(_2196_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0031_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold321 (.A(\mac1.sum_lvl3_ff[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold322 (.A(_2174_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0025_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold324 (.A(\mac1.sum_lvl3_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold325 (.A(_0018_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold326 (.A(\DP_4.matrix[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold327 (.A(\mac1.sum_lvl3_ff[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold328 (.A(_2215_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold329 (.A(_0020_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold330 (.A(\mac1.sum_lvl2_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold331 (.A(_2118_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0009_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold333 (.A(\DP_4.matrix[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold334 (.A(\DP_4.matrix[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold335 (.A(\mac1.sum_lvl2_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold336 (.A(_2134_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold337 (.A(_2135_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold338 (.A(_0014_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold339 (.A(\DP_4.matrix[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold340 (.A(\mac1.sum_lvl2_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold341 (.A(_2115_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0008_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold343 (.A(\DP_4.matrix[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold344 (.A(\DP_2.matrix[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold345 (.A(\DP_3.matrix[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold346 (.A(\DP_4.matrix[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold347 (.A(\mac2.sum_lvl2_ff[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold348 (.A(_2238_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold349 (.A(_0043_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold350 (.A(\mac1.sum_lvl2_ff[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold351 (.A(_2164_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0006_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold353 (.A(\DP_2.matrix[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold354 (.A(_0198_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold355 (.A(\DP_1.matrix[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold356 (.A(\mac2.sum_lvl3_ff[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold357 (.A(_2294_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold358 (.A(_0059_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold359 (.A(\DP_2.matrix[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold360 (.A(\DP_4.matrix[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold361 (.A(_0996_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0080_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold363 (.A(\DP_1.matrix[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold364 (.A(\DP_4.matrix[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold365 (.A(\DP_2.matrix[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold366 (.A(\mac1.sum_lvl3_ff[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold367 (.A(_2177_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold368 (.A(_0026_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold369 (.A(\DP_4.matrix[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold370 (.A(\DP_4.matrix[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold371 (.A(\DP_2.matrix[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold372 (.A(\DP_2.matrix[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold373 (.A(\DP_2.matrix[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold374 (.A(\DP_4.matrix[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold375 (.A(_0248_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold376 (.A(\DP_3.matrix[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold377 (.A(_0225_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold378 (.A(\DP_2.matrix[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold379 (.A(\mac1.sum_lvl3_ff[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold380 (.A(_2186_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold381 (.A(_2193_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0030_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold383 (.A(\mac2.sum_lvl3_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold384 (.A(_2304_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold385 (.A(_2305_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold386 (.A(_0062_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold387 (.A(\DP_3.matrix[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold388 (.A(\DP_3.matrix[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold389 (.A(\mac2.sum_lvl3_ff[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold390 (.A(_0063_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold391 (.A(\DP_2.matrix[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold392 (.A(_0625_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold393 (.A(_0075_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold394 (.A(\mac1.sum_lvl2_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold395 (.A(_2139_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold396 (.A(_2140_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold397 (.A(_0015_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold398 (.A(\mac1.sum_lvl3_ff[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold399 (.A(_2222_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold400 (.A(_0022_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold401 (.A(\DP_1.matrix[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold402 (.A(_2981_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold403 (.A(\DP_1.I_range.out_data[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold404 (.A(\mac2.sum_lvl3_ff[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold405 (.A(_0049_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold406 (.A(\DP_1.matrix[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold407 (.A(\DP_1.matrix[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold408 (.A(\DP_1.matrix[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold409 (.A(\mac2.sum_lvl3_ff[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold410 (.A(_0055_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold411 (.A(\mac2.sum_lvl2_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold412 (.A(_2235_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold413 (.A(_0042_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold414 (.A(\mac1.sum_lvl3_ff[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold415 (.A(_2171_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold416 (.A(_0024_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold417 (.A(\mac2.sum_lvl3_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold418 (.A(_2291_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold419 (.A(_0058_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold420 (.A(\mac1.sum_lvl2_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold421 (.A(_2162_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold422 (.A(_0005_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold423 (.A(\mac2.sum_lvl3_ff[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold424 (.A(_2296_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold425 (.A(_2299_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold426 (.A(_0060_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold427 (.A(\mac2.sum_lvl3_ff[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold428 (.A(_2327_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold429 (.A(_2328_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold430 (.A(_0052_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold431 (.A(\DP_1.matrix[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold432 (.A(\DP_2.matrix[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold433 (.A(\mac2.sum_lvl3_ff[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold434 (.A(_2285_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold435 (.A(_0056_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold436 (.A(\DP_3.matrix[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold437 (.A(\mac1.sum_lvl3_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold438 (.A(_2218_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold439 (.A(_0021_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold440 (.A(\DP_4.matrix[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold441 (.A(\mac1.sum_lvl2_ff[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold442 (.A(_2151_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold443 (.A(_0003_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold444 (.A(\mac2.sum_lvl3_ff[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold445 (.A(_2288_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold446 (.A(_0057_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold447 (.A(\DP_1.matrix[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold448 (.A(\DP_2.matrix[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold449 (.A(\DP_3.matrix[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold450 (.A(\mac2.sum_lvl2_ff[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold451 (.A(_2248_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold452 (.A(_2249_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold453 (.A(_0046_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold454 (.A(\DP_2.matrix[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold455 (.A(\DP_1.matrix[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold456 (.A(\DP_4.matrix[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold457 (.A(\DP_4.matrix[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold458 (.A(\DP_1.matrix[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold459 (.A(\DP_2.matrix[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold460 (.A(\DP_4.matrix[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold461 (.A(\mac1.sum_lvl3_ff[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold462 (.A(_2182_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold463 (.A(_2185_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold464 (.A(_0028_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold465 (.A(\mac1.sum_lvl2_ff[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold466 (.A(_2124_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold467 (.A(_0011_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold468 (.A(\mac1.sum_lvl2_ff[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold469 (.A(_2126_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold470 (.A(_2129_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold471 (.A(_0012_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold472 (.A(\mac1.sum_lvl2_ff[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold473 (.A(_2121_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold474 (.A(_0010_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold475 (.A(\DP_1.matrix[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold476 (.A(\DP_3.matrix[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold477 (.A(\mac2.sum_lvl2_ff[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold478 (.A(_2240_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold479 (.A(_2243_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold480 (.A(_0044_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold481 (.A(\DP_3.matrix[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold482 (.A(\DP_1.matrix[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold483 (.A(\DP_2.matrix[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold484 (.A(\DP_1.matrix[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold485 (.A(\DP_3.matrix[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold486 (.A(\DP_1.matrix[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold487 (.A(\mac2.sum_lvl2_ff[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold488 (.A(_2278_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold489 (.A(\mac1.sum_lvl2_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold490 (.A(_2131_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold491 (.A(_2133_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold492 (.A(_0013_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold493 (.A(\mac1.sum_lvl3_ff[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold494 (.A(\DP_2.matrix[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold495 (.A(\DP_2.matrix[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold496 (.A(\DP_3.matrix[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold497 (.A(\mac2.sum_lvl3_ff[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold498 (.A(_2301_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold499 (.A(_2302_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold500 (.A(_0061_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold501 (.A(\DP_4.matrix[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold502 (.A(\mac2.sum_lvl2_ff[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold503 (.A(_2276_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold504 (.A(\DP_1.matrix[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold505 (.A(\mac2.sum_lvl2_ff[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold506 (.A(\mac1.sum_lvl2_ff[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net546));
 sg13g2_fill_1 FILLER_0_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_1027 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net33;
 assign uio_oe[1] = net34;
 assign uio_oe[2] = net35;
 assign uio_oe[3] = net36;
 assign uio_oe[4] = net37;
 assign uio_oe[5] = net38;
 assign uio_oe[6] = net39;
 assign uio_oe[7] = net40;
endmodule
