* NGSPICE file created from heichips25_template.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_2 abstract view
.subckt sg13g2_and3_2 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_2 abstract view
.subckt sg13g2_nor4_2 A B C Y VSS VDD D
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

.subckt heichips25_template VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
X_3155_ _2727_ _2717_ _2725_ _2745_ VPWR VGND sg13g2_a21o_1
X_3086_ _2677_ _2657_ _0068_ VPWR VGND sg13g2_xor2_1
X_3988_ _0777_ _0778_ _0780_ _0781_ VPWR VGND sg13g2_or3_1
XFILLER_23_667 VPWR VGND sg13g2_fill_2
X_5727_ DP_1.Q_range.out_data\[4\] DP_1.I_range.out_data\[5\] _2384_ VPWR VGND sg13g2_nor2b_1
X_5658_ mac2.total_sum\[1\] mac1.total_sum\[1\] _2331_ VPWR VGND sg13g2_xor2_1
X_5589_ net498 mac2.sum_lvl3_ff\[22\] _2277_ VPWR VGND sg13g2_xor2_1
X_4609_ _1373_ _1374_ _1375_ VPWR VGND sg13g2_nor2b_1
Xhold340 _0246_ VPWR VGND net380 sg13g2_dlygate4sd3_1
Xhold351 _0008_ VPWR VGND net391 sg13g2_dlygate4sd3_1
Xhold362 _2311_ VPWR VGND net402 sg13g2_dlygate4sd3_1
Xhold395 DP_3.matrix\[2\] VPWR VGND net435 sg13g2_dlygate4sd3_1
Xhold384 DP_1.matrix\[72\] VPWR VGND net424 sg13g2_dlygate4sd3_1
Xhold373 _0052_ VPWR VGND net413 sg13g2_dlygate4sd3_1
Xfanout820 net821 net820 VPWR VGND sg13g2_buf_8
Xfanout842 net329 net842 VPWR VGND sg13g2_buf_8
Xfanout831 net832 net831 VPWR VGND sg13g2_buf_1
Xfanout853 net405 net853 VPWR VGND sg13g2_buf_2
Xfanout875 net876 net875 VPWR VGND sg13g2_buf_8
Xfanout864 net865 net864 VPWR VGND sg13g2_buf_2
Xfanout897 net356 net897 VPWR VGND sg13g2_buf_8
Xfanout886 net887 net886 VPWR VGND sg13g2_buf_8
XFILLER_26_41 VPWR VGND sg13g2_fill_2
XFILLER_27_951 VPWR VGND sg13g2_decap_8
XFILLER_41_420 VPWR VGND sg13g2_fill_1
XFILLER_42_976 VPWR VGND sg13g2_decap_8
XFILLER_10_840 VPWR VGND sg13g2_decap_8
XFILLER_6_888 VPWR VGND sg13g2_decap_8
XFILLER_3_1007 VPWR VGND sg13g2_decap_8
XFILLER_37_726 VPWR VGND sg13g2_fill_1
XFILLER_18_973 VPWR VGND sg13g2_decap_8
X_4960_ _1713_ _1707_ _1715_ VPWR VGND sg13g2_xor2_1
XFILLER_45_792 VPWR VGND sg13g2_fill_2
X_4891_ _1649_ _1646_ _1648_ VPWR VGND sg13g2_nand2_1
X_3911_ _0703_ _0704_ _0698_ _0706_ VPWR VGND sg13g2_nand3_1
X_3842_ _0639_ net1022 net953 VPWR VGND sg13g2_nand2_1
X_6561_ net1067 VGND VPWR _0047_ mac2.sum_lvl3_ff\[9\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_3773_ _0577_ _0568_ _0576_ VPWR VGND sg13g2_xnor2_1
X_5512_ mac2.sum_lvl2_ff\[20\] mac2.sum_lvl2_ff\[1\] _2217_ VPWR VGND sg13g2_nor2_1
X_6492_ net1144 VGND VPWR net235 mac2.sum_lvl1_ff\[8\] clknet_leaf_41_clk sg13g2_dfrbpq_1
XFILLER_8_192 VPWR VGND sg13g2_fill_1
X_5443_ mac1.sum_lvl3_ff\[22\] net381 _2163_ VPWR VGND sg13g2_and2_1
X_5374_ VGND VPWR _2107_ _2109_ net390 _2106_ sg13g2_a21oi_2
X_4325_ _1103_ _1097_ _1102_ VPWR VGND sg13g2_xnor2_1
X_4256_ _1034_ _1031_ _1036_ VPWR VGND sg13g2_xor2_1
X_3207_ _2756_ VPWR _2796_ VGND _2754_ _2757_ sg13g2_o21ai_1
X_4187_ _0974_ _0949_ _0973_ VPWR VGND sg13g2_xnor2_1
X_3138_ _2727_ _2726_ _2717_ _2729_ VPWR VGND sg13g2_a21o_1
XFILLER_28_748 VPWR VGND sg13g2_fill_2
X_3069_ VPWR _2662_ _2661_ VGND sg13g2_inv_1
XFILLER_24_954 VPWR VGND sg13g2_decap_8
XFILLER_3_825 VPWR VGND sg13g2_decap_8
Xhold170 mac2.sum_lvl1_ff\[38\] VPWR VGND net210 sg13g2_dlygate4sd3_1
Xhold181 mac2.sum_lvl1_ff\[7\] VPWR VGND net221 sg13g2_dlygate4sd3_1
Xhold192 mac2.products_ff\[148\] VPWR VGND net232 sg13g2_dlygate4sd3_1
XFILLER_14_420 VPWR VGND sg13g2_fill_2
XFILLER_15_932 VPWR VGND sg13g2_decap_8
XFILLER_18_1015 VPWR VGND sg13g2_decap_8
XFILLER_14_475 VPWR VGND sg13g2_decap_4
XFILLER_14_486 VPWR VGND sg13g2_fill_1
XFILLER_5_173 VPWR VGND sg13g2_fill_2
X_5090_ _1834_ _1835_ _1836_ VPWR VGND sg13g2_nor2b_1
X_4110_ _0900_ _0880_ _0899_ VPWR VGND sg13g2_xnor2_1
X_4041_ _0833_ _0818_ _0832_ VPWR VGND sg13g2_nand2_1
X_5992_ _2620_ net863 net789 VPWR VGND sg13g2_nand2_1
X_4943_ _1697_ _1698_ _1699_ VPWR VGND sg13g2_and2_1
X_4874_ _1592_ VPWR _1632_ VGND _1589_ _1593_ sg13g2_o21ai_1
XFILLER_21_957 VPWR VGND sg13g2_decap_8
X_3825_ _0624_ _0616_ _0623_ VPWR VGND sg13g2_nand2_1
X_3756_ VGND VPWR _0508_ _0528_ _0561_ _0530_ sg13g2_a21oi_1
X_6544_ net1143 VGND VPWR net89 mac2.sum_lvl2_ff\[31\] clknet_leaf_42_clk sg13g2_dfrbpq_1
Xclkbuf_4_12_0_clk clknet_0_clk clknet_4_12_0_clk VPWR VGND sg13g2_buf_8
X_6475_ net1075 VGND VPWR _0157_ mac2.products_ff\[143\] clknet_leaf_22_clk sg13g2_dfrbpq_1
X_3687_ _0494_ _0484_ _0493_ VPWR VGND sg13g2_nand2b_1
X_5426_ _2151_ net466 _2149_ VPWR VGND sg13g2_nand2b_1
X_5357_ VGND VPWR _2064_ _2087_ _2095_ _2089_ sg13g2_a21oi_1
X_5288_ _1998_ VPWR _2029_ VGND _1996_ _1999_ sg13g2_o21ai_1
X_4308_ _1087_ _1057_ _1085_ VPWR VGND sg13g2_xnor2_1
X_4239_ _1015_ VPWR _1020_ VGND _1016_ _1018_ sg13g2_o21ai_1
XFILLER_15_228 VPWR VGND sg13g2_fill_1
XFILLER_24_740 VPWR VGND sg13g2_decap_8
XFILLER_12_913 VPWR VGND sg13g2_decap_8
XFILLER_24_751 VPWR VGND sg13g2_fill_2
XFILLER_8_906 VPWR VGND sg13g2_decap_8
XFILLER_48_1019 VPWR VGND sg13g2_decap_8
XFILLER_3_677 VPWR VGND sg13g2_fill_2
XFILLER_48_94 VPWR VGND sg13g2_fill_1
XFILLER_30_710 VPWR VGND sg13g2_fill_1
X_3610_ _0396_ _0416_ _0418_ _0419_ VPWR VGND sg13g2_or3_1
X_4590_ _1358_ net923 net863 _0084_ VPWR VGND sg13g2_and3_2
XFILLER_7_961 VPWR VGND sg13g2_decap_8
X_3541_ _0351_ _0347_ _0350_ VPWR VGND sg13g2_nand2_1
X_3472_ _0283_ _0282_ _0285_ VPWR VGND sg13g2_xor2_1
X_6260_ net1064 VGND VPWR net239 mac1.sum_lvl1_ff\[36\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_6191_ net1091 VGND VPWR _0211_ DP_2.matrix\[43\] clknet_leaf_65_clk sg13g2_dfrbpq_1
X_5211_ _1955_ _1918_ _1953_ VPWR VGND sg13g2_nand2_1
X_5142_ VGND VPWR _1887_ _1885_ _1842_ sg13g2_or2_1
XFILLER_29_0 VPWR VGND sg13g2_fill_1
XFILLER_29_309 VPWR VGND sg13g2_fill_1
X_5073_ _1817_ _1818_ _1812_ _1820_ VPWR VGND sg13g2_nand3_1
X_4024_ _0807_ _0815_ _0816_ VPWR VGND sg13g2_nor2_1
X_5975_ _2609_ _2489_ _2504_ VPWR VGND sg13g2_xnor2_1
X_4926_ _1661_ VPWR _1682_ VGND _1658_ _1662_ sg13g2_o21ai_1
X_4857_ _1580_ _1614_ _1578_ _1616_ VPWR VGND sg13g2_nand3_1
X_3808_ _0598_ VPWR _0610_ VGND _0570_ _0596_ sg13g2_o21ai_1
X_6527_ net1143 VGND VPWR net256 mac2.sum_lvl2_ff\[11\] clknet_leaf_42_clk sg13g2_dfrbpq_1
X_4788_ _1531_ VPWR _1548_ VGND _1510_ _1532_ sg13g2_o21ai_1
X_3739_ _0544_ net1032 net1053 VPWR VGND sg13g2_nand2_1
X_6458_ net1134 VGND VPWR _0134_ mac2.products_ff\[74\] clknet_leaf_44_clk sg13g2_dfrbpq_1
X_6389_ net1062 VGND VPWR net288 mac1.sum_lvl3_ff\[1\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_5409_ _2132_ _2130_ _2131_ _2137_ VPWR VGND sg13g2_a21o_2
XFILLER_47_139 VPWR VGND sg13g2_fill_2
XFILLER_28_353 VPWR VGND sg13g2_fill_1
XFILLER_44_868 VPWR VGND sg13g2_fill_2
XFILLER_11_220 VPWR VGND sg13g2_fill_1
XFILLER_12_754 VPWR VGND sg13g2_fill_2
XFILLER_7_257 VPWR VGND sg13g2_fill_2
XFILLER_4_964 VPWR VGND sg13g2_decap_8
XFILLER_19_386 VPWR VGND sg13g2_fill_1
X_5760_ _2417_ _2395_ net808 VPWR VGND sg13g2_nand2_1
X_5691_ mac2.total_sum\[8\] mac1.total_sum\[8\] _2354_ _2356_ VPWR VGND sg13g2_a21o_1
X_4711_ _1473_ _1435_ _1470_ VPWR VGND sg13g2_xnor2_1
X_4642_ _1406_ _1405_ _1402_ VPWR VGND sg13g2_nand2b_1
X_4573_ _1342_ _1336_ _1344_ VPWR VGND sg13g2_xor2_1
X_6312_ net1117 VGND VPWR net254 mac1.sum_lvl2_ff\[42\] clknet_leaf_54_clk sg13g2_dfrbpq_1
X_3524_ _0332_ _0331_ _0326_ _0335_ VPWR VGND sg13g2_a21o_1
X_6243_ net1126 VGND VPWR _0251_ DP_4.matrix\[7\] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_3455_ net1041 net1039 net974 net972 _0268_ VPWR VGND sg13g2_and4_1
X_3386_ _2931_ _2969_ _2970_ VPWR VGND sg13g2_nor2_1
X_6174_ net1067 VGND VPWR _0099_ mac1.products_ff\[150\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_5125_ _1869_ _1868_ _0157_ VPWR VGND sg13g2_xor2_1
X_5056_ _1803_ _1801_ _1802_ VPWR VGND sg13g2_nand2b_1
X_4007_ _0797_ _0796_ _0798_ _0800_ VPWR VGND sg13g2_a21o_1
XFILLER_25_345 VPWR VGND sg13g2_fill_2
X_5958_ VGND VPWR net783 _2598_ _0200_ _2597_ sg13g2_a21oi_1
XFILLER_25_389 VPWR VGND sg13g2_fill_1
XFILLER_41_838 VPWR VGND sg13g2_fill_1
X_4909_ _1665_ _1656_ _1666_ VPWR VGND sg13g2_nor2b_1
X_5889_ net806 VPWR _2543_ VGND DP_4.matrix\[73\] _2476_ sg13g2_o21ai_1
XFILLER_1_956 VPWR VGND sg13g2_decap_8
XFILLER_49_938 VPWR VGND sg13g2_decap_8
Xhold30 mac2.products_ff\[15\] VPWR VGND net70 sg13g2_dlygate4sd3_1
XFILLER_0_466 VPWR VGND sg13g2_decap_8
XFILLER_0_488 VPWR VGND sg13g2_fill_1
Xhold41 mac1.products_ff\[7\] VPWR VGND net81 sg13g2_dlygate4sd3_1
Xhold63 mac1.products_ff\[2\] VPWR VGND net103 sg13g2_dlygate4sd3_1
Xhold74 mac2.products_ff\[75\] VPWR VGND net114 sg13g2_dlygate4sd3_1
Xhold52 mac2.sum_lvl2_ff\[52\] VPWR VGND net92 sg13g2_dlygate4sd3_1
Xhold96 mac1.sum_lvl2_ff\[42\] VPWR VGND net136 sg13g2_dlygate4sd3_1
Xhold85 mac1.sum_lvl2_ff\[49\] VPWR VGND net125 sg13g2_dlygate4sd3_1
XFILLER_16_334 VPWR VGND sg13g2_fill_1
X_3240_ _2793_ VPWR _2828_ VGND _2790_ _2794_ sg13g2_o21ai_1
X_3171_ _2758_ _2759_ _2753_ _2761_ VPWR VGND sg13g2_nand3_1
Xfanout1050 net302 net1050 VPWR VGND sg13g2_buf_8
Xfanout1072 net1087 net1072 VPWR VGND sg13g2_buf_8
Xfanout1061 net1068 net1061 VPWR VGND sg13g2_buf_8
Xfanout1083 net1085 net1083 VPWR VGND sg13g2_buf_8
Xfanout1094 net1095 net1094 VPWR VGND sg13g2_buf_8
XFILLER_19_194 VPWR VGND sg13g2_decap_4
X_5812_ VPWR _2468_ _2467_ VGND sg13g2_inv_1
X_5743_ DP_1.Q_range.out_data\[2\] DP_1.I_range.out_data\[2\] _2400_ VPWR VGND sg13g2_nor2b_2
XFILLER_34_186 VPWR VGND sg13g2_fill_1
X_5674_ mac2.total_sum\[5\] mac1.total_sum\[5\] _2343_ VPWR VGND sg13g2_xor2_1
X_4625_ _1386_ _1387_ _1389_ _1390_ VPWR VGND sg13g2_or3_1
Xhold511 mac1.sum_lvl3_ff\[4\] VPWR VGND net551 sg13g2_dlygate4sd3_1
Xhold500 mac1.sum_lvl3_ff\[12\] VPWR VGND net540 sg13g2_dlygate4sd3_1
X_4556_ _1326_ _1327_ _1328_ VPWR VGND sg13g2_and2_1
X_3507_ _0316_ _0315_ _0318_ VPWR VGND sg13g2_xor2_1
X_4487_ _1261_ net901 net1043 VPWR VGND sg13g2_nand2_1
X_3438_ _3015_ _3008_ _0071_ VPWR VGND sg13g2_xor2_1
X_6226_ net1127 VGND VPWR _0234_ DP_3.matrix\[42\] clknet_leaf_45_clk sg13g2_dfrbpq_2
X_6157_ net1112 VGND VPWR _0188_ DP_1.matrix\[72\] clknet_leaf_58_clk sg13g2_dfrbpq_1
X_3369_ _2952_ _2953_ _2954_ VPWR VGND sg13g2_nor2_1
X_5108_ _1854_ _1847_ _1852_ _1853_ VPWR VGND sg13g2_and3_1
X_6088_ net1063 VGND VPWR _0069_ mac1.products_ff\[0\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_5039_ _1787_ _1780_ _1785_ _1786_ VPWR VGND sg13g2_and3_1
XFILLER_39_993 VPWR VGND sg13g2_decap_8
XFILLER_14_805 VPWR VGND sg13g2_decap_4
XFILLER_22_882 VPWR VGND sg13g2_fill_1
XFILLER_31_75 VPWR VGND sg13g2_fill_1
Xoutput31 net31 uo_out[6] VPWR VGND sg13g2_buf_1
Xoutput20 net20 uio_out[3] VPWR VGND sg13g2_buf_1
XFILLER_0_263 VPWR VGND sg13g2_decap_8
XFILLER_17_643 VPWR VGND sg13g2_fill_2
XFILLER_29_492 VPWR VGND sg13g2_fill_2
XFILLER_32_635 VPWR VGND sg13g2_fill_1
XFILLER_9_820 VPWR VGND sg13g2_decap_8
XFILLER_9_875 VPWR VGND sg13g2_decap_8
XFILLER_8_352 VPWR VGND sg13g2_fill_2
X_4410_ _1186_ _1179_ _1185_ VPWR VGND sg13g2_xnor2_1
X_5390_ net462 VPWR _2122_ VGND _2116_ _2120_ sg13g2_o21ai_1
X_4341_ _1095_ _1116_ _1118_ _1119_ VPWR VGND sg13g2_or3_1
X_4272_ _1050_ _1049_ _1011_ _1052_ VPWR VGND sg13g2_a21o_1
X_6011_ VPWR _0251_ _2632_ VGND sg13g2_inv_1
X_3223_ _2788_ VPWR _2812_ VGND _2808_ _2810_ sg13g2_o21ai_1
X_3154_ _2744_ _2739_ _2742_ VPWR VGND sg13g2_xnor2_1
XFILLER_11_0 VPWR VGND sg13g2_fill_1
X_3085_ VGND VPWR _2678_ _2677_ _2657_ sg13g2_or2_1
XFILLER_27_418 VPWR VGND sg13g2_decap_4
XFILLER_36_930 VPWR VGND sg13g2_decap_4
XFILLER_22_123 VPWR VGND sg13g2_decap_4
X_3987_ _0780_ net1057 net963 net1005 net959 VPWR VGND sg13g2_a22oi_1
X_5726_ mac2.total_sum\[0\] mac1.total_sum\[0\] net25 VPWR VGND sg13g2_xor2_1
XFILLER_22_178 VPWR VGND sg13g2_fill_1
X_5657_ mac1.total_sum\[1\] mac2.total_sum\[1\] _2330_ VPWR VGND sg13g2_nor2_1
X_5588_ mac2.sum_lvl3_ff\[22\] net498 _2276_ VPWR VGND sg13g2_and2_1
X_4608_ _1369_ VPWR _1374_ VGND _1370_ _1372_ sg13g2_o21ai_1
Xhold330 DP_4.matrix\[74\] VPWR VGND net370 sg13g2_dlygate4sd3_1
Xhold341 mac1.sum_lvl3_ff\[2\] VPWR VGND net381 sg13g2_dlygate4sd3_1
Xhold352 mac1.sum_lvl2_ff\[8\] VPWR VGND net392 sg13g2_dlygate4sd3_1
X_4539_ _1311_ net897 DP_4.matrix\[44\] VPWR VGND sg13g2_nand2_1
Xhold396 _0222_ VPWR VGND net436 sg13g2_dlygate4sd3_1
Xhold385 DP_1.matrix\[2\] VPWR VGND net425 sg13g2_dlygate4sd3_1
Xhold374 DP_2.matrix\[4\] VPWR VGND net414 sg13g2_dlygate4sd3_1
Xhold363 _0050_ VPWR VGND net403 sg13g2_dlygate4sd3_1
Xfanout821 DP_4.matrix\[75\] net821 VPWR VGND sg13g2_buf_2
Xfanout832 net376 net832 VPWR VGND sg13g2_buf_1
Xfanout810 _2396_ net810 VPWR VGND sg13g2_buf_8
Xfanout843 DP_4.matrix\[38\] net843 VPWR VGND sg13g2_buf_1
X_6209_ net1122 VGND VPWR net388 DP_3.matrix\[3\] clknet_leaf_35_clk sg13g2_dfrbpq_2
Xfanout876 DP_3.matrix\[77\] net876 VPWR VGND sg13g2_buf_8
Xfanout854 net855 net854 VPWR VGND sg13g2_buf_8
Xfanout865 net866 net865 VPWR VGND sg13g2_buf_2
Xfanout887 net888 net887 VPWR VGND sg13g2_buf_1
Xfanout898 DP_3.matrix\[40\] net898 VPWR VGND sg13g2_buf_8
XFILLER_26_462 VPWR VGND sg13g2_fill_2
XFILLER_42_911 VPWR VGND sg13g2_fill_2
XFILLER_22_690 VPWR VGND sg13g2_fill_2
XFILLER_10_896 VPWR VGND sg13g2_decap_8
XFILLER_6_867 VPWR VGND sg13g2_decap_8
XFILLER_1_550 VPWR VGND sg13g2_fill_2
XFILLER_18_952 VPWR VGND sg13g2_decap_8
X_4890_ VPWR _1648_ _1647_ VGND sg13g2_inv_1
X_3910_ _0705_ _0698_ _0703_ _0704_ VPWR VGND sg13g2_and3_1
XFILLER_17_484 VPWR VGND sg13g2_fill_1
X_3841_ _0638_ net953 net1024 net955 net1022 VPWR VGND sg13g2_a22oi_1
XFILLER_33_988 VPWR VGND sg13g2_decap_8
XFILLER_20_638 VPWR VGND sg13g2_fill_1
X_3772_ _0576_ _0540_ _0574_ VPWR VGND sg13g2_xnor2_1
X_6560_ net1073 VGND VPWR net520 mac2.sum_lvl3_ff\[8\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_5511_ _2216_ mac2.sum_lvl2_ff\[20\] mac2.sum_lvl2_ff\[1\] VPWR VGND sg13g2_nand2_1
X_6491_ net1141 VGND VPWR net160 mac2.sum_lvl1_ff\[7\] clknet_leaf_41_clk sg13g2_dfrbpq_1
X_5442_ _2159_ VPWR _2162_ VGND _2158_ _2160_ sg13g2_o21ai_1
X_5373_ net390 _2106_ _0008_ VPWR VGND sg13g2_xor2_1
X_4324_ _1102_ _1064_ _1099_ VPWR VGND sg13g2_xnor2_1
X_4255_ _1035_ _1034_ _1031_ VPWR VGND sg13g2_nand2b_1
X_3206_ _2795_ _2790_ _2794_ VPWR VGND sg13g2_xnor2_1
X_4186_ _0971_ _0965_ _0973_ VPWR VGND sg13g2_xor2_1
XFILLER_41_1014 VPWR VGND sg13g2_decap_8
X_3137_ _2726_ _2727_ _2717_ _2728_ VPWR VGND sg13g2_nand3_1
X_3068_ _2658_ _2660_ _2661_ VPWR VGND sg13g2_nor2_1
XFILLER_24_933 VPWR VGND sg13g2_decap_8
X_5709_ _2360_ _2365_ _2371_ VPWR VGND sg13g2_nor2_1
XFILLER_3_804 VPWR VGND sg13g2_decap_8
XFILLER_12_99 VPWR VGND sg13g2_fill_2
Xhold171 mac1.sum_lvl1_ff\[41\] VPWR VGND net211 sg13g2_dlygate4sd3_1
Xhold160 mac1.products_ff\[14\] VPWR VGND net200 sg13g2_dlygate4sd3_1
Xhold182 mac2.sum_lvl1_ff\[3\] VPWR VGND net222 sg13g2_dlygate4sd3_1
Xhold193 mac2.products_ff\[150\] VPWR VGND net233 sg13g2_dlygate4sd3_1
XFILLER_37_52 VPWR VGND sg13g2_fill_2
XFILLER_15_911 VPWR VGND sg13g2_decap_8
XFILLER_15_988 VPWR VGND sg13g2_decap_8
XFILLER_30_936 VPWR VGND sg13g2_fill_1
X_4040_ _0831_ _0824_ _0832_ VPWR VGND sg13g2_xor2_1
X_5991_ _2619_ _2541_ _2545_ VPWR VGND sg13g2_xnor2_1
X_4942_ _1671_ _1673_ _1696_ _1698_ VPWR VGND sg13g2_or3_1
X_4873_ _1631_ _1623_ _1628_ VPWR VGND sg13g2_xnor2_1
XFILLER_21_936 VPWR VGND sg13g2_decap_8
X_3824_ _0621_ _0622_ _0623_ VPWR VGND sg13g2_nor2b_1
XFILLER_20_479 VPWR VGND sg13g2_fill_1
X_6543_ net1136 VGND VPWR net111 mac2.sum_lvl2_ff\[30\] clknet_leaf_43_clk sg13g2_dfrbpq_1
X_3755_ _0558_ _0537_ _0560_ VPWR VGND sg13g2_xor2_1
X_3686_ _0493_ _0485_ _0492_ VPWR VGND sg13g2_xnor2_1
X_6474_ net1079 VGND VPWR _0156_ mac2.products_ff\[142\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_5425_ VGND VPWR _2150_ net465 mac1.sum_lvl2_ff\[32\] sg13g2_or2_1
X_5356_ _2091_ VPWR _2094_ VGND _2076_ _2093_ sg13g2_o21ai_1
X_5287_ _2008_ VPWR _2028_ VGND _2006_ _2009_ sg13g2_o21ai_1
X_4307_ _1085_ _1057_ _1086_ VPWR VGND sg13g2_nor2b_1
X_4238_ _1015_ _1016_ _1018_ _1019_ VPWR VGND sg13g2_or3_1
X_4169_ _0955_ _0956_ _0957_ VPWR VGND sg13g2_and2_1
XFILLER_43_527 VPWR VGND sg13g2_fill_1
XFILLER_12_969 VPWR VGND sg13g2_decap_8
XFILLER_11_468 VPWR VGND sg13g2_fill_1
XFILLER_47_822 VPWR VGND sg13g2_fill_2
XFILLER_19_502 VPWR VGND sg13g2_fill_1
XFILLER_19_557 VPWR VGND sg13g2_fill_2
XFILLER_46_354 VPWR VGND sg13g2_fill_2
XFILLER_15_752 VPWR VGND sg13g2_fill_2
XFILLER_15_785 VPWR VGND sg13g2_fill_2
XFILLER_15_796 VPWR VGND sg13g2_decap_8
XFILLER_31_1013 VPWR VGND sg13g2_decap_8
XFILLER_7_940 VPWR VGND sg13g2_decap_8
XFILLER_11_980 VPWR VGND sg13g2_decap_8
X_3540_ _0348_ _0349_ _0350_ VPWR VGND sg13g2_nor2b_1
XFILLER_6_472 VPWR VGND sg13g2_fill_2
X_5210_ _1918_ _1953_ _1954_ VPWR VGND sg13g2_nor2_1
X_3471_ _0282_ _0283_ _0284_ VPWR VGND sg13g2_nor2b_2
X_6190_ net1091 VGND VPWR _0210_ DP_2.matrix\[42\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_5141_ _1886_ net820 net875 VPWR VGND sg13g2_nand2_1
X_5072_ _1819_ _1812_ _1817_ _1818_ VPWR VGND sg13g2_and3_1
X_4023_ _0815_ _0808_ _0814_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_800 VPWR VGND sg13g2_fill_1
XFILLER_37_321 VPWR VGND sg13g2_fill_2
XFILLER_37_387 VPWR VGND sg13g2_fill_1
X_5974_ _2608_ VPWR _0222_ VGND net789 _2607_ sg13g2_o21ai_1
X_4925_ _1664_ _1657_ _1666_ _1681_ VPWR VGND sg13g2_a21o_1
X_4856_ VGND VPWR _1578_ _1580_ _1615_ _1614_ sg13g2_a21oi_1
X_3807_ VGND VPWR _0578_ _0601_ _0609_ _0603_ sg13g2_a21oi_1
X_6526_ net1143 VGND VPWR net257 mac2.sum_lvl2_ff\[10\] clknet_leaf_43_clk sg13g2_dfrbpq_1
X_4787_ _1508_ VPWR _1547_ VGND _1463_ _1509_ sg13g2_o21ai_1
X_3738_ _0512_ VPWR _0543_ VGND _0510_ _0513_ sg13g2_o21ai_1
X_3669_ _0476_ net1032 net966 VPWR VGND sg13g2_nand2_1
X_6457_ net1118 VGND VPWR _0127_ mac2.products_ff\[73\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_6388_ net1064 VGND VPWR net268 mac1.sum_lvl3_ff\[0\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_5408_ VPWR _2136_ _2135_ VGND sg13g2_inv_1
X_5339_ _2062_ _2054_ _2061_ _2078_ VPWR VGND sg13g2_a21o_1
Xclkbuf_leaf_67_clk clknet_4_0_0_clk clknet_leaf_67_clk VPWR VGND sg13g2_buf_8
XFILLER_44_825 VPWR VGND sg13g2_decap_8
XFILLER_29_877 VPWR VGND sg13g2_fill_1
XFILLER_29_888 VPWR VGND sg13g2_fill_1
XFILLER_44_836 VPWR VGND sg13g2_fill_1
XFILLER_28_376 VPWR VGND sg13g2_fill_1
XFILLER_31_519 VPWR VGND sg13g2_decap_8
XFILLER_7_247 VPWR VGND sg13g2_fill_1
XFILLER_12_799 VPWR VGND sg13g2_decap_8
XFILLER_4_943 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_58_clk clknet_4_10_0_clk clknet_leaf_58_clk VPWR VGND sg13g2_buf_8
Xclkbuf_4_11_0_clk clknet_0_clk clknet_4_11_0_clk VPWR VGND sg13g2_buf_8
XFILLER_35_836 VPWR VGND sg13g2_fill_2
X_5690_ _2354_ _2355_ net17 VPWR VGND sg13g2_nor2b_2
X_4710_ _1435_ _1470_ _1472_ VPWR VGND sg13g2_and2_1
X_4641_ _1404_ _1381_ _1405_ VPWR VGND sg13g2_xor2_1
X_4572_ _1343_ _1336_ _1342_ VPWR VGND sg13g2_nand2_1
X_6311_ net1071 VGND VPWR net157 mac1.sum_lvl2_ff\[41\] clknet_leaf_66_clk sg13g2_dfrbpq_1
X_3523_ _0331_ _0332_ _0326_ _0334_ VPWR VGND sg13g2_nand3_1
X_6242_ net1128 VGND VPWR net358 DP_4.matrix\[6\] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_3454_ _3031_ net1039 net972 VPWR VGND sg13g2_nand2_1
XFILLER_41_0 VPWR VGND sg13g2_fill_1
X_6173_ net1094 VGND VPWR net407 DP_2.matrix\[3\] clknet_leaf_61_clk sg13g2_dfrbpq_1
X_3385_ _2969_ _2960_ _2968_ VPWR VGND sg13g2_xnor2_1
X_5124_ _1870_ _1868_ _1869_ VPWR VGND sg13g2_nand2_1
X_5055_ _1802_ net889 net814 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_49_clk clknet_4_11_0_clk clknet_leaf_49_clk VPWR VGND sg13g2_buf_8
X_4006_ _0797_ _0798_ _0796_ _0799_ VPWR VGND sg13g2_nand3_1
X_5957_ _2598_ _2460_ _2462_ VPWR VGND sg13g2_xnor2_1
X_4908_ _1665_ _1657_ _1664_ VPWR VGND sg13g2_xnor2_1
X_5888_ _2542_ net847 net795 VPWR VGND sg13g2_nand2b_1
X_4839_ _1572_ VPWR _1598_ VGND _1566_ _1573_ sg13g2_o21ai_1
XFILLER_5_718 VPWR VGND sg13g2_fill_2
X_6509_ net1136 VGND VPWR net252 mac2.sum_lvl1_ff\[45\] clknet_leaf_50_clk sg13g2_dfrbpq_1
XFILLER_1_935 VPWR VGND sg13g2_decap_8
XFILLER_49_917 VPWR VGND sg13g2_decap_8
XFILLER_0_445 VPWR VGND sg13g2_fill_2
Xhold31 mac1.products_ff\[12\] VPWR VGND net71 sg13g2_dlygate4sd3_1
Xhold20 mac2.products_ff\[142\] VPWR VGND net60 sg13g2_dlygate4sd3_1
Xhold64 mac1.sum_lvl2_ff\[50\] VPWR VGND net104 sg13g2_dlygate4sd3_1
Xhold42 mac2.sum_lvl1_ff\[6\] VPWR VGND net82 sg13g2_dlygate4sd3_1
Xhold53 mac2.sum_lvl1_ff\[79\] VPWR VGND net93 sg13g2_dlygate4sd3_1
Xhold97 mac2.sum_lvl1_ff\[15\] VPWR VGND net137 sg13g2_dlygate4sd3_1
Xhold86 mac1.products_ff\[139\] VPWR VGND net126 sg13g2_dlygate4sd3_1
Xhold75 mac2.sum_lvl2_ff\[43\] VPWR VGND net115 sg13g2_dlygate4sd3_1
XFILLER_44_600 VPWR VGND sg13g2_fill_1
XFILLER_17_825 VPWR VGND sg13g2_fill_2
XFILLER_17_869 VPWR VGND sg13g2_decap_8
XFILLER_40_861 VPWR VGND sg13g2_decap_8
Xfanout1040 net336 net1040 VPWR VGND sg13g2_buf_8
XFILLER_6_1028 VPWR VGND sg13g2_fill_1
X_3170_ _2760_ _2753_ _2758_ _2759_ VPWR VGND sg13g2_and3_1
Xfanout1051 net386 net1051 VPWR VGND sg13g2_buf_8
Xfanout1062 net1064 net1062 VPWR VGND sg13g2_buf_8
Xfanout1073 net1074 net1073 VPWR VGND sg13g2_buf_8
Xfanout1095 net1108 net1095 VPWR VGND sg13g2_buf_8
Xfanout1084 net1085 net1084 VPWR VGND sg13g2_buf_8
X_5811_ _2464_ _2466_ _2467_ VPWR VGND sg13g2_nor2_1
XFILLER_35_699 VPWR VGND sg13g2_fill_2
X_5742_ _2399_ net418 net801 VPWR VGND sg13g2_nand2_1
X_5673_ mac1.total_sum\[5\] mac2.total_sum\[5\] _2342_ VPWR VGND sg13g2_nor2_1
X_4624_ _1389_ net916 net868 net918 net865 VPWR VGND sg13g2_a22oi_1
Xhold501 _2200_ VPWR VGND net541 sg13g2_dlygate4sd3_1
X_4555_ _1299_ _1301_ _1325_ _1327_ VPWR VGND sg13g2_or3_1
X_3506_ _0317_ _0315_ _0316_ VPWR VGND sg13g2_nand2b_1
Xhold512 mac2.sum_lvl2_ff\[14\] VPWR VGND net552 sg13g2_dlygate4sd3_1
X_4486_ VGND VPWR _1260_ _1233_ _1231_ sg13g2_or2_1
X_3437_ _3016_ _3008_ _3015_ VPWR VGND sg13g2_nand2_1
X_6225_ net1097 VGND VPWR net181 mac1.sum_lvl1_ff\[15\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_6156_ net1111 VGND VPWR _0103_ mac1.products_ff\[144\] clknet_leaf_54_clk sg13g2_dfrbpq_1
X_3368_ VGND VPWR _2922_ _2953_ _2920_ _2900_ sg13g2_a21oi_2
X_5107_ _1848_ VPWR _1853_ VGND _1849_ _1851_ sg13g2_o21ai_1
X_3299_ _2886_ _2876_ _2885_ VPWR VGND sg13g2_nand2b_1
Xheichips25_template_33 VPWR VGND uio_oe[0] sg13g2_tiehi
XFILLER_39_972 VPWR VGND sg13g2_decap_8
X_6087_ net1080 VGND VPWR DP_3.Q_range.data_plus_4\[6\] DP_3.Q_range.out_data\[5\]
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
X_5038_ _1781_ VPWR _1786_ VGND _1782_ _1784_ sg13g2_o21ai_1
XFILLER_41_625 VPWR VGND sg13g2_fill_1
XFILLER_40_102 VPWR VGND sg13g2_fill_1
XFILLER_40_146 VPWR VGND sg13g2_fill_1
Xoutput21 net21 uio_out[4] VPWR VGND sg13g2_buf_1
Xoutput32 net32 uo_out[7] VPWR VGND sg13g2_buf_1
XFILLER_29_482 VPWR VGND sg13g2_fill_1
XFILLER_16_121 VPWR VGND sg13g2_fill_2
XFILLER_45_986 VPWR VGND sg13g2_decap_8
XFILLER_44_496 VPWR VGND sg13g2_fill_2
XFILLER_9_854 VPWR VGND sg13g2_decap_8
X_4340_ VGND VPWR _1114_ _1115_ _1118_ _1096_ sg13g2_a21oi_1
X_4271_ _1049_ _1050_ _1011_ _1051_ VPWR VGND sg13g2_nand3_1
X_6010_ _2632_ _2573_ _2631_ net791 net853 VPWR VGND sg13g2_a22oi_1
X_3222_ _2788_ _2808_ _2810_ _2811_ VPWR VGND sg13g2_or3_1
X_3153_ _2743_ _2739_ _2742_ VPWR VGND sg13g2_nand2_1
XFILLER_48_780 VPWR VGND sg13g2_fill_1
X_3084_ _2675_ _2674_ _2677_ VPWR VGND sg13g2_xor2_1
XFILLER_22_102 VPWR VGND sg13g2_decap_8
XFILLER_10_308 VPWR VGND sg13g2_fill_2
X_3986_ net959 net1005 net963 _0779_ VPWR VGND net1057 sg13g2_nand4_1
X_5725_ net24 _2382_ _2383_ VPWR VGND sg13g2_xnor2_1
X_5656_ _2329_ mac1.total_sum\[1\] mac2.total_sum\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_11_1022 VPWR VGND sg13g2_decap_8
X_4607_ _1369_ _1370_ _1372_ _1373_ VPWR VGND sg13g2_nor3_1
Xhold320 _2286_ VPWR VGND net360 sg13g2_dlygate4sd3_1
X_5587_ _2272_ VPWR _2275_ VGND _2271_ _2273_ sg13g2_o21ai_1
Xhold331 DP_4.matrix\[4\] VPWR VGND net371 sg13g2_dlygate4sd3_1
Xhold353 _2127_ VPWR VGND net393 sg13g2_dlygate4sd3_1
Xhold342 _2164_ VPWR VGND net382 sg13g2_dlygate4sd3_1
X_4538_ _1289_ VPWR _1310_ VGND _1286_ _1290_ sg13g2_o21ai_1
Xfanout800 _2401_ net800 VPWR VGND sg13g2_buf_8
Xhold364 DP_2.matrix\[76\] VPWR VGND net404 sg13g2_dlygate4sd3_1
Xhold386 DP_2.matrix\[78\] VPWR VGND net426 sg13g2_dlygate4sd3_1
Xhold375 DP_2.matrix\[42\] VPWR VGND net415 sg13g2_dlygate4sd3_1
X_4469_ VGND VPWR _1207_ _1209_ _1244_ _1243_ sg13g2_a21oi_1
Xfanout811 net813 net811 VPWR VGND sg13g2_buf_8
Xfanout822 net823 net822 VPWR VGND sg13g2_buf_8
X_6208_ net1122 VGND VPWR net436 DP_3.matrix\[2\] clknet_leaf_35_clk sg13g2_dfrbpq_2
Xfanout833 net334 net833 VPWR VGND sg13g2_buf_8
Xhold397 mac2.sum_lvl3_ff\[35\] VPWR VGND net437 sg13g2_dlygate4sd3_1
Xfanout855 net357 net855 VPWR VGND sg13g2_buf_8
Xfanout866 net474 net866 VPWR VGND sg13g2_buf_8
Xfanout844 net846 net844 VPWR VGND sg13g2_buf_2
Xfanout877 net878 net877 VPWR VGND sg13g2_buf_2
X_6139_ net1094 VGND VPWR net397 DP_1.matrix\[4\] clknet_leaf_61_clk sg13g2_dfrbpq_1
XFILLER_19_909 VPWR VGND sg13g2_decap_8
Xfanout899 net337 net899 VPWR VGND sg13g2_buf_8
Xfanout888 net310 net888 VPWR VGND sg13g2_buf_2
XFILLER_26_43 VPWR VGND sg13g2_fill_1
XFILLER_27_986 VPWR VGND sg13g2_decap_8
XFILLER_14_658 VPWR VGND sg13g2_fill_1
XFILLER_10_875 VPWR VGND sg13g2_decap_8
XFILLER_6_846 VPWR VGND sg13g2_decap_8
XFILLER_18_931 VPWR VGND sg13g2_decap_8
XFILLER_45_783 VPWR VGND sg13g2_fill_1
XFILLER_17_474 VPWR VGND sg13g2_decap_4
XFILLER_45_794 VPWR VGND sg13g2_fill_1
X_3840_ _0077_ _0624_ _0636_ VPWR VGND sg13g2_xnor2_1
X_3771_ _0540_ _0574_ _0575_ VPWR VGND sg13g2_nor2b_1
XFILLER_34_1011 VPWR VGND sg13g2_decap_8
XFILLER_12_190 VPWR VGND sg13g2_decap_8
X_5510_ _2215_ net308 net271 VPWR VGND sg13g2_nand2_1
X_6490_ net1141 VGND VPWR net261 mac2.sum_lvl1_ff\[6\] clknet_leaf_44_clk sg13g2_dfrbpq_1
X_5441_ _0023_ _2158_ _2161_ VPWR VGND sg13g2_xnor2_1
X_5372_ net389 mac1.sum_lvl2_ff\[21\] _2108_ VPWR VGND sg13g2_xor2_1
X_4323_ _1064_ _1099_ _1101_ VPWR VGND sg13g2_and2_1
X_4254_ _1033_ _1010_ _1034_ VPWR VGND sg13g2_xor2_1
X_3205_ _2794_ _2747_ _2792_ VPWR VGND sg13g2_xnor2_1
X_4185_ _0972_ _0965_ _0971_ VPWR VGND sg13g2_nand2_1
X_3136_ _2724_ _2723_ _2718_ _2727_ VPWR VGND sg13g2_a21o_1
X_3067_ net1004 net1000 net934 net932 _2660_ VPWR VGND sg13g2_and4_1
XFILLER_24_912 VPWR VGND sg13g2_decap_8
XFILLER_24_989 VPWR VGND sg13g2_decap_8
X_3969_ _0762_ net947 net1022 net949 net1019 VPWR VGND sg13g2_a22oi_1
X_5708_ mac2.total_sum\[12\] mac1.total_sum\[12\] _2370_ VPWR VGND sg13g2_xor2_1
X_5639_ net531 VPWR _2317_ VGND _2314_ _2316_ sg13g2_o21ai_1
Xhold150 mac2.sum_lvl1_ff\[72\] VPWR VGND net190 sg13g2_dlygate4sd3_1
Xhold161 mac1.products_ff\[142\] VPWR VGND net201 sg13g2_dlygate4sd3_1
Xhold172 mac1.sum_lvl1_ff\[36\] VPWR VGND net212 sg13g2_dlygate4sd3_1
Xhold194 mac1.sum_lvl1_ff\[2\] VPWR VGND net234 sg13g2_dlygate4sd3_1
Xhold183 mac1.products_ff\[150\] VPWR VGND net223 sg13g2_dlygate4sd3_1
XFILLER_14_422 VPWR VGND sg13g2_fill_1
XFILLER_15_967 VPWR VGND sg13g2_decap_8
XFILLER_14_499 VPWR VGND sg13g2_fill_1
XFILLER_6_676 VPWR VGND sg13g2_fill_2
XFILLER_5_175 VPWR VGND sg13g2_fill_1
XFILLER_2_882 VPWR VGND sg13g2_decap_8
XFILLER_49_363 VPWR VGND sg13g2_fill_1
XFILLER_37_503 VPWR VGND sg13g2_decap_8
XFILLER_37_547 VPWR VGND sg13g2_fill_2
X_5990_ _0244_ net868 net793 VPWR VGND sg13g2_xnor2_1
X_4941_ _1696_ VPWR _1697_ VGND _1671_ _1673_ sg13g2_o21ai_1
X_4872_ VGND VPWR _1630_ _1628_ _1623_ sg13g2_or2_1
X_3823_ _0618_ VPWR _0622_ VGND _0619_ _0620_ sg13g2_o21ai_1
XFILLER_21_915 VPWR VGND sg13g2_decap_8
X_6542_ net1141 VGND VPWR net41 mac2.sum_lvl2_ff\[29\] clknet_leaf_43_clk sg13g2_dfrbpq_1
X_3754_ _0558_ _0537_ _0559_ VPWR VGND sg13g2_nor2b_1
X_3685_ _0490_ _0491_ _0492_ VPWR VGND sg13g2_nor2b_1
X_6473_ net1081 VGND VPWR _0149_ mac2.products_ff\[141\] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_5424_ mac1.sum_lvl2_ff\[32\] net465 _2149_ VPWR VGND sg13g2_and2_1
X_5355_ _0154_ _2076_ _2092_ VPWR VGND sg13g2_xnor2_1
XFILLER_0_819 VPWR VGND sg13g2_decap_8
X_5286_ _2027_ _2026_ _2024_ VPWR VGND sg13g2_nand2b_1
X_4306_ _1085_ _1061_ _1084_ VPWR VGND sg13g2_xnor2_1
X_4237_ _1018_ net898 net849 net900 net846 VPWR VGND sg13g2_a22oi_1
XFILLER_28_514 VPWR VGND sg13g2_fill_1
X_4168_ _0928_ _0930_ _0954_ _0956_ VPWR VGND sg13g2_or3_1
X_3119_ _2708_ _2707_ _2710_ VPWR VGND sg13g2_xor2_1
X_4099_ VGND VPWR _0889_ _0862_ _0860_ sg13g2_or2_1
XFILLER_24_720 VPWR VGND sg13g2_fill_2
XFILLER_23_241 VPWR VGND sg13g2_fill_1
XFILLER_24_786 VPWR VGND sg13g2_decap_4
XFILLER_12_948 VPWR VGND sg13g2_decap_8
XFILLER_20_992 VPWR VGND sg13g2_decap_8
XFILLER_2_167 VPWR VGND sg13g2_fill_2
XFILLER_24_1010 VPWR VGND sg13g2_decap_8
XFILLER_46_344 VPWR VGND sg13g2_fill_2
XFILLER_7_996 VPWR VGND sg13g2_decap_8
X_3470_ _3026_ VPWR _0283_ VGND _3017_ _3027_ sg13g2_o21ai_1
X_5140_ _1885_ net818 net876 VPWR VGND sg13g2_nand2_2
XFILLER_9_1015 VPWR VGND sg13g2_decap_8
X_5071_ _1813_ VPWR _1818_ VGND _1814_ _1816_ sg13g2_o21ai_1
X_4022_ _0814_ _0809_ _0812_ VPWR VGND sg13g2_xnor2_1
X_5973_ _2608_ net920 net789 VPWR VGND sg13g2_nand2_1
X_4924_ _1680_ _1677_ _0141_ VPWR VGND sg13g2_xor2_1
X_4855_ _1612_ _1585_ _1614_ VPWR VGND sg13g2_xor2_1
X_3806_ _0605_ VPWR _0608_ VGND _0590_ _0607_ sg13g2_o21ai_1
X_4786_ _1536_ VPWR _1546_ VGND _1465_ _1537_ sg13g2_o21ai_1
X_3737_ _0522_ VPWR _0542_ VGND _0520_ _0523_ sg13g2_o21ai_1
X_6525_ net1143 VGND VPWR net259 mac2.sum_lvl2_ff\[9\] clknet_leaf_42_clk sg13g2_dfrbpq_1
X_3668_ _0475_ net1037 net1053 VPWR VGND sg13g2_nand2_1
X_6456_ net1129 VGND VPWR _0083_ mac2.products_ff\[72\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_3599_ _0408_ net1058 net984 DP_1.matrix\[7\] net980 VPWR VGND sg13g2_a22oi_1
X_6387_ net1089 VGND VPWR net143 mac1.sum_lvl3_ff\[35\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_5407_ net478 net365 _2135_ VPWR VGND sg13g2_xor2_1
X_5338_ VGND VPWR _2053_ _2067_ _2077_ _2066_ sg13g2_a21oi_1
X_5269_ _2011_ _2005_ _2010_ VPWR VGND sg13g2_xnor2_1
XFILLER_16_506 VPWR VGND sg13g2_fill_2
XFILLER_16_528 VPWR VGND sg13g2_fill_1
XFILLER_12_756 VPWR VGND sg13g2_fill_1
XFILLER_15_1009 VPWR VGND sg13g2_decap_8
XFILLER_7_215 VPWR VGND sg13g2_decap_4
XFILLER_4_922 VPWR VGND sg13g2_decap_8
XFILLER_4_999 VPWR VGND sg13g2_decap_8
XFILLER_46_141 VPWR VGND sg13g2_fill_2
XFILLER_46_185 VPWR VGND sg13g2_fill_2
XFILLER_15_583 VPWR VGND sg13g2_fill_2
X_4640_ _1404_ net921 net860 VPWR VGND sg13g2_nand2_1
X_6310_ net1069 VGND VPWR net150 mac1.sum_lvl2_ff\[40\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_4571_ _1342_ _1337_ _1340_ VPWR VGND sg13g2_xnor2_1
X_3522_ _0333_ _0326_ _0331_ _0332_ VPWR VGND sg13g2_and3_1
X_6241_ net1126 VGND VPWR _0249_ DP_4.matrix\[5\] clknet_leaf_37_clk sg13g2_dfrbpq_2
X_3453_ _3030_ net972 net1040 net974 net1038 VPWR VGND sg13g2_a22oi_1
X_6172_ net1093 VGND VPWR _0198_ DP_2.matrix\[2\] clknet_leaf_61_clk sg13g2_dfrbpq_1
X_3384_ _2968_ _2932_ _2966_ VPWR VGND sg13g2_xnor2_1
XFILLER_34_0 VPWR VGND sg13g2_fill_2
X_5123_ _1831_ _1830_ _1829_ _1869_ VPWR VGND sg13g2_a21o_1
XFILLER_29_108 VPWR VGND sg13g2_fill_2
X_5054_ _1778_ VPWR _1801_ VGND _1753_ _1776_ sg13g2_o21ai_1
X_4005_ _0750_ VPWR _0798_ VGND _0689_ _0751_ sg13g2_o21ai_1
XFILLER_25_347 VPWR VGND sg13g2_fill_1
XFILLER_38_1009 VPWR VGND sg13g2_decap_8
X_5956_ net972 net783 _2597_ VPWR VGND sg13g2_nor2_1
XFILLER_41_829 VPWR VGND sg13g2_decap_4
X_4907_ _1664_ _1658_ _1663_ VPWR VGND sg13g2_xnor2_1
X_5887_ _2541_ _2538_ _2540_ VPWR VGND sg13g2_nand2_1
X_4838_ _1595_ _1587_ _1597_ VPWR VGND sg13g2_xor2_1
X_4769_ _1530_ _1511_ _1528_ _1529_ VPWR VGND sg13g2_and3_1
X_6508_ net1136 VGND VPWR net199 mac2.sum_lvl1_ff\[44\] clknet_leaf_49_clk sg13g2_dfrbpq_1
X_6439_ net1124 VGND VPWR _0087_ mac2.products_ff\[3\] clknet_leaf_32_clk sg13g2_dfrbpq_1
XFILLER_1_914 VPWR VGND sg13g2_decap_8
Xhold32 mac1.products_ff\[72\] VPWR VGND net72 sg13g2_dlygate4sd3_1
Xhold10 mac2.sum_lvl2_ff\[50\] VPWR VGND net50 sg13g2_dlygate4sd3_1
Xhold21 mac2.products_ff\[137\] VPWR VGND net61 sg13g2_dlygate4sd3_1
Xhold54 mac2.sum_lvl1_ff\[84\] VPWR VGND net94 sg13g2_dlygate4sd3_1
Xhold65 mac2.sum_lvl2_ff\[51\] VPWR VGND net105 sg13g2_dlygate4sd3_1
Xhold43 mac2.products_ff\[9\] VPWR VGND net83 sg13g2_dlygate4sd3_1
Xhold87 mac1.sum_lvl1_ff\[5\] VPWR VGND net127 sg13g2_dlygate4sd3_1
Xhold98 mac1.sum_lvl1_ff\[81\] VPWR VGND net138 sg13g2_dlygate4sd3_1
XFILLER_17_804 VPWR VGND sg13g2_decap_8
XFILLER_21_1013 VPWR VGND sg13g2_decap_8
Xhold76 mac2.sum_lvl2_ff\[38\] VPWR VGND net116 sg13g2_dlygate4sd3_1
XFILLER_17_848 VPWR VGND sg13g2_decap_8
XFILLER_29_686 VPWR VGND sg13g2_fill_2
XFILLER_28_196 VPWR VGND sg13g2_fill_2
XFILLER_43_177 VPWR VGND sg13g2_fill_2
XFILLER_3_262 VPWR VGND sg13g2_decap_4
XFILLER_6_1007 VPWR VGND sg13g2_decap_8
Xfanout1030 net1031 net1030 VPWR VGND sg13g2_buf_8
Xfanout1041 DP_1.matrix\[0\] net1041 VPWR VGND sg13g2_buf_1
Xfanout1063 net1064 net1063 VPWR VGND sg13g2_buf_8
XFILLER_0_980 VPWR VGND sg13g2_decap_8
Xfanout1052 DP_2.matrix\[44\] net1052 VPWR VGND sg13g2_buf_8
Xfanout1074 net1087 net1074 VPWR VGND sg13g2_buf_8
XFILLER_19_141 VPWR VGND sg13g2_decap_4
Xfanout1096 net1099 net1096 VPWR VGND sg13g2_buf_8
Xfanout1085 net1086 net1085 VPWR VGND sg13g2_buf_8
XFILLER_48_984 VPWR VGND sg13g2_decap_8
XFILLER_34_122 VPWR VGND sg13g2_fill_2
X_5810_ _2466_ net800 _2465_ net801 DP_2.matrix\[78\] VPWR VGND sg13g2_a22oi_1
XFILLER_22_306 VPWR VGND sg13g2_fill_2
X_5741_ _2395_ net809 _2398_ VPWR VGND sg13g2_nor2_1
X_5672_ VGND VPWR _2338_ _2340_ _2341_ _2339_ sg13g2_a21oi_1
X_4623_ net865 net918 net868 _1388_ VPWR VGND net916 sg13g2_nand4_1
Xhold502 DP_1.matrix\[77\] VPWR VGND net542 sg13g2_dlygate4sd3_1
X_4554_ _1325_ VPWR _1326_ VGND _1299_ _1301_ sg13g2_o21ai_1
X_3505_ _0316_ net1041 net970 VPWR VGND sg13g2_nand2_1
X_4485_ _1221_ VPWR _1259_ VGND _1218_ _1222_ sg13g2_o21ai_1
X_6224_ net1146 VGND VPWR _0233_ DP_3.matrix\[41\] clknet_leaf_45_clk sg13g2_dfrbpq_2
XFILLER_44_1013 VPWR VGND sg13g2_decap_8
X_3436_ _3013_ _3014_ _3015_ VPWR VGND sg13g2_nor2b_1
X_6155_ net1070 VGND VPWR _0187_ DP_1.matrix\[43\] clknet_leaf_3_clk sg13g2_dfrbpq_2
X_3367_ _2950_ _2929_ _2952_ VPWR VGND sg13g2_xor2_1
X_5106_ _1848_ _1849_ _1851_ _1852_ VPWR VGND sg13g2_or3_1
X_6086_ net1080 VGND VPWR net11 DP_3.Q_range.out_data\[4\] clknet_leaf_22_clk sg13g2_dfrbpq_1
X_5037_ _1781_ _1782_ _1784_ _1785_ VPWR VGND sg13g2_or3_1
X_3298_ _2885_ _2877_ _2884_ VPWR VGND sg13g2_xnor2_1
Xheichips25_template_34 VPWR VGND uio_oe[1] sg13g2_tiehi
XFILLER_26_656 VPWR VGND sg13g2_fill_1
X_5939_ VGND VPWR net787 _2586_ _0177_ _2585_ sg13g2_a21oi_1
Xclkbuf_4_10_0_clk clknet_0_clk clknet_4_10_0_clk VPWR VGND sg13g2_buf_8
Xoutput22 net22 uio_out[5] VPWR VGND sg13g2_buf_1
XFILLER_1_788 VPWR VGND sg13g2_decap_8
XFILLER_45_965 VPWR VGND sg13g2_decap_8
XFILLER_16_100 VPWR VGND sg13g2_fill_2
XFILLER_44_486 VPWR VGND sg13g2_fill_1
XFILLER_12_361 VPWR VGND sg13g2_fill_2
XFILLER_13_884 VPWR VGND sg13g2_decap_8
X_4270_ _1048_ _1047_ _1030_ _1050_ VPWR VGND sg13g2_a21o_1
X_3221_ VGND VPWR _2806_ _2807_ _2810_ _2789_ sg13g2_a21oi_1
X_3152_ _2740_ _2741_ _2742_ VPWR VGND sg13g2_nor2b_2
X_3083_ _2674_ _2675_ _2676_ VPWR VGND sg13g2_nor2b_2
XFILLER_23_615 VPWR VGND sg13g2_decap_8
XFILLER_36_987 VPWR VGND sg13g2_decap_8
XFILLER_23_626 VPWR VGND sg13g2_fill_1
X_3985_ net963 net959 net1005 net1056 _0778_ VPWR VGND sg13g2_and4_1
X_5724_ _2383_ mac1.total_sum\[15\] mac2.total_sum\[15\] VPWR VGND sg13g2_xnor2_1
X_5655_ _2328_ mac1.total_sum\[0\] mac2.total_sum\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_11_1001 VPWR VGND sg13g2_decap_8
X_4606_ _1372_ net918 net869 net920 net863 VPWR VGND sg13g2_a22oi_1
Xhold310 mac2.sum_lvl2_ff\[2\] VPWR VGND net350 sg13g2_dlygate4sd3_1
X_5586_ _0055_ _2271_ _2274_ VPWR VGND sg13g2_xnor2_1
Xhold332 _0248_ VPWR VGND net372 sg13g2_dlygate4sd3_1
Xhold343 _0024_ VPWR VGND net383 sg13g2_dlygate4sd3_1
Xhold321 _0059_ VPWR VGND net361 sg13g2_dlygate4sd3_1
X_4537_ _1292_ _1285_ _1294_ _1309_ VPWR VGND sg13g2_a21o_1
Xhold365 DP_4.matrix\[7\] VPWR VGND net405 sg13g2_dlygate4sd3_1
Xhold354 _2128_ VPWR VGND net394 sg13g2_dlygate4sd3_1
Xhold376 DP_2.matrix\[6\] VPWR VGND net416 sg13g2_dlygate4sd3_1
X_4468_ _1241_ _1214_ _1243_ VPWR VGND sg13g2_xor2_1
Xhold387 mac1.sum_lvl3_ff\[13\] VPWR VGND net427 sg13g2_dlygate4sd3_1
Xfanout812 net813 net812 VPWR VGND sg13g2_buf_1
Xfanout823 net370 net823 VPWR VGND sg13g2_buf_2
Xfanout801 _2398_ net801 VPWR VGND sg13g2_buf_8
X_6207_ net1114 VGND VPWR net74 mac1.sum_lvl1_ff\[9\] clknet_leaf_59_clk sg13g2_dfrbpq_1
X_3419_ VGND VPWR _2970_ _2993_ _3001_ _2995_ sg13g2_a21oi_1
Xhold398 _2327_ VPWR VGND net438 sg13g2_dlygate4sd3_1
Xfanout834 DP_4.matrix\[43\] net834 VPWR VGND sg13g2_buf_1
Xfanout856 net450 net856 VPWR VGND sg13g2_buf_8
Xfanout867 net868 net867 VPWR VGND sg13g2_buf_2
X_6138_ net1062 VGND VPWR _0066_ mac1.products_ff\[138\] clknet_leaf_67_clk sg13g2_dfrbpq_1
X_4399_ _1165_ VPWR _1175_ VGND _1094_ _1166_ sg13g2_o21ai_1
Xfanout845 DP_4.matrix\[37\] net845 VPWR VGND sg13g2_buf_1
Xfanout878 net879 net878 VPWR VGND sg13g2_buf_2
Xfanout889 net890 net889 VPWR VGND sg13g2_buf_8
X_6069_ net847 _0253_ VPWR VGND sg13g2_buf_1
XFILLER_39_781 VPWR VGND sg13g2_fill_2
XFILLER_26_464 VPWR VGND sg13g2_fill_1
XFILLER_27_965 VPWR VGND sg13g2_decap_8
XFILLER_26_497 VPWR VGND sg13g2_decap_4
XFILLER_41_489 VPWR VGND sg13g2_fill_1
XFILLER_10_854 VPWR VGND sg13g2_decap_8
XFILLER_22_692 VPWR VGND sg13g2_fill_1
XFILLER_21_191 VPWR VGND sg13g2_decap_4
XFILLER_42_98 VPWR VGND sg13g2_fill_2
XFILLER_18_910 VPWR VGND sg13g2_decap_8
XFILLER_18_987 VPWR VGND sg13g2_decap_8
XFILLER_20_629 VPWR VGND sg13g2_fill_1
X_3770_ _0574_ _0569_ _0572_ VPWR VGND sg13g2_xnor2_1
XFILLER_32_489 VPWR VGND sg13g2_fill_1
X_5440_ mac1.sum_lvl3_ff\[1\] mac1.sum_lvl3_ff\[21\] _2161_ VPWR VGND sg13g2_xor2_1
X_5371_ mac1.sum_lvl2_ff\[21\] net389 _2107_ VPWR VGND sg13g2_and2_1
XFILLER_5_891 VPWR VGND sg13g2_decap_8
X_4322_ VGND VPWR _1100_ _1098_ _1065_ sg13g2_or2_1
X_4253_ _1033_ net903 net840 VPWR VGND sg13g2_nand2_1
X_3204_ VGND VPWR _2793_ _2791_ _2748_ sg13g2_or2_1
X_4184_ _0971_ _0966_ _0969_ VPWR VGND sg13g2_xnor2_1
X_3135_ _2723_ _2724_ _2718_ _2726_ VPWR VGND sg13g2_nand3_1
X_3066_ _2659_ net1000 net932 VPWR VGND sg13g2_nand2_1
XFILLER_23_434 VPWR VGND sg13g2_fill_1
XFILLER_24_968 VPWR VGND sg13g2_decap_8
X_3968_ net1021 net1019 net949 net947 _0761_ VPWR VGND sg13g2_and4_1
XFILLER_10_117 VPWR VGND sg13g2_fill_1
X_5707_ mac1.total_sum\[12\] mac2.total_sum\[12\] _2369_ VPWR VGND sg13g2_nor2_1
X_3899_ _0694_ net1017 net954 VPWR VGND sg13g2_nand2_1
X_5638_ VGND VPWR _2301_ _2303_ _2316_ _2315_ sg13g2_a21oi_1
X_5569_ mac2.sum_lvl2_ff\[32\] mac2.sum_lvl2_ff\[13\] _2262_ VPWR VGND sg13g2_and2_1
XFILLER_3_839 VPWR VGND sg13g2_decap_8
Xhold151 mac2.sum_lvl1_ff\[44\] VPWR VGND net191 sg13g2_dlygate4sd3_1
Xhold140 mac2.sum_lvl1_ff\[42\] VPWR VGND net180 sg13g2_dlygate4sd3_1
Xhold162 mac2.sum_lvl1_ff\[85\] VPWR VGND net202 sg13g2_dlygate4sd3_1
Xhold173 mac1.sum_lvl2_ff\[51\] VPWR VGND net213 sg13g2_dlygate4sd3_1
Xhold184 mac2.products_ff\[79\] VPWR VGND net224 sg13g2_dlygate4sd3_1
Xhold195 mac2.products_ff\[8\] VPWR VGND net235 sg13g2_dlygate4sd3_1
XFILLER_19_729 VPWR VGND sg13g2_fill_1
XFILLER_15_946 VPWR VGND sg13g2_decap_8
XFILLER_2_861 VPWR VGND sg13g2_decap_8
X_4940_ _1695_ _1681_ _1696_ VPWR VGND sg13g2_xor2_1
X_4871_ _1623_ _1628_ _1629_ VPWR VGND sg13g2_and2_1
X_3822_ _0618_ _0619_ _0620_ _0621_ VPWR VGND sg13g2_nor3_1
X_6541_ net1137 VGND VPWR net55 mac2.sum_lvl2_ff\[28\] clknet_leaf_50_clk sg13g2_dfrbpq_1
XFILLER_9_460 VPWR VGND sg13g2_fill_2
X_3753_ _0556_ _0555_ _0558_ VPWR VGND sg13g2_xor2_1
X_3684_ _0486_ VPWR _0491_ VGND _0488_ _0489_ sg13g2_o21ai_1
X_6472_ net1081 VGND VPWR _0093_ mac2.products_ff\[140\] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_5423_ _2142_ VPWR _2148_ VGND _2143_ _2147_ sg13g2_o21ai_1
X_5354_ VPWR _2093_ _2092_ VGND sg13g2_inv_1
X_4305_ _1084_ _1081_ _1083_ VPWR VGND sg13g2_nand2_1
X_5285_ VGND VPWR _2026_ _2025_ _1973_ sg13g2_or2_1
X_4236_ net846 net900 net849 _1017_ VPWR VGND net898 sg13g2_nand4_1
X_4167_ _0954_ VPWR _0955_ VGND _0928_ _0930_ sg13g2_o21ai_1
X_3118_ _2709_ _2707_ VPWR VGND _2708_ sg13g2_nand2b_2
X_4098_ _0850_ VPWR _0888_ VGND _0847_ _0851_ sg13g2_o21ai_1
X_3049_ _2644_ _2636_ _2643_ VPWR VGND sg13g2_nand2_1
XFILLER_11_404 VPWR VGND sg13g2_fill_2
XFILLER_12_927 VPWR VGND sg13g2_decap_8
XFILLER_23_34 VPWR VGND sg13g2_fill_2
XFILLER_20_971 VPWR VGND sg13g2_decap_8
XFILLER_48_64 VPWR VGND sg13g2_fill_2
XFILLER_46_301 VPWR VGND sg13g2_fill_1
XFILLER_15_754 VPWR VGND sg13g2_fill_1
XFILLER_14_253 VPWR VGND sg13g2_fill_2
XFILLER_15_776 VPWR VGND sg13g2_fill_1
XFILLER_42_562 VPWR VGND sg13g2_fill_1
XFILLER_7_975 VPWR VGND sg13g2_decap_8
X_5070_ _1813_ _1814_ _1816_ _1817_ VPWR VGND sg13g2_or3_1
X_4021_ _0813_ _0812_ _0809_ VPWR VGND sg13g2_nand2b_1
XFILLER_38_813 VPWR VGND sg13g2_decap_8
X_5972_ _2503_ _2499_ _2607_ VPWR VGND sg13g2_xor2_1
X_4923_ _1680_ _1679_ _1648_ _1678_ _1619_ VPWR VGND sg13g2_a22oi_1
X_4854_ _1613_ _1612_ _1585_ VPWR VGND sg13g2_nand2b_1
X_3805_ _0110_ _0590_ _0606_ VPWR VGND sg13g2_xnor2_1
X_4785_ _1541_ VPWR _1545_ VGND _1498_ _1543_ sg13g2_o21ai_1
X_3736_ _0541_ _0540_ _0538_ VPWR VGND sg13g2_nand2b_1
X_6524_ net1143 VGND VPWR net247 mac2.sum_lvl2_ff\[8\] clknet_leaf_42_clk sg13g2_dfrbpq_1
X_3667_ _0449_ VPWR _0474_ VGND _0447_ _0450_ sg13g2_o21ai_1
X_6455_ net1120 VGND VPWR _0082_ mac2.products_ff\[71\] clknet_leaf_31_clk sg13g2_dfrbpq_1
XFILLER_47_1022 VPWR VGND sg13g2_decap_8
X_3598_ net979 net1025 net983 _0407_ VPWR VGND net1058 sg13g2_nand4_1
X_5406_ _2134_ net365 mac1.sum_lvl2_ff\[10\] VPWR VGND sg13g2_nand2_1
X_6386_ net1073 VGND VPWR net87 mac1.sum_lvl3_ff\[34\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_5337_ _2076_ _2075_ _2070_ _2074_ _2052_ VPWR VGND sg13g2_a22oi_1
X_5268_ _2009_ _2006_ _2010_ VPWR VGND sg13g2_xor2_1
X_4219_ _1001_ net900 net850 net902 net847 VPWR VGND sg13g2_a22oi_1
X_5199_ _1941_ _1942_ _1943_ VPWR VGND sg13g2_nor2_1
XFILLER_28_312 VPWR VGND sg13g2_fill_1
XFILLER_28_367 VPWR VGND sg13g2_fill_1
XFILLER_12_746 VPWR VGND sg13g2_fill_2
XFILLER_34_66 VPWR VGND sg13g2_fill_1
XFILLER_4_901 VPWR VGND sg13g2_decap_8
XFILLER_4_978 VPWR VGND sg13g2_decap_8
XFILLER_3_433 VPWR VGND sg13g2_fill_1
XFILLER_19_345 VPWR VGND sg13g2_fill_1
XFILLER_35_805 VPWR VGND sg13g2_fill_2
XFILLER_46_164 VPWR VGND sg13g2_fill_1
XFILLER_43_893 VPWR VGND sg13g2_fill_1
X_4570_ _1341_ _1340_ _1337_ VPWR VGND sg13g2_nand2b_1
X_3521_ _0327_ VPWR _0332_ VGND _0328_ _0330_ sg13g2_o21ai_1
X_6240_ net1126 VGND VPWR net372 DP_4.matrix\[4\] clknet_leaf_37_clk sg13g2_dfrbpq_1
X_3452_ _0072_ _3016_ _3028_ VPWR VGND sg13g2_xnor2_1
X_3383_ _2932_ _2966_ _2967_ VPWR VGND sg13g2_nor2b_1
X_6171_ net1067 VGND VPWR _0098_ mac1.products_ff\[149\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_5122_ _1867_ _1803_ _1868_ VPWR VGND sg13g2_xor2_1
X_5053_ _1800_ _1792_ _1794_ VPWR VGND sg13g2_nand2_1
X_4004_ _0723_ VPWR _0797_ VGND _0793_ _0795_ sg13g2_o21ai_1
XFILLER_38_687 VPWR VGND sg13g2_fill_2
X_5955_ VGND VPWR net783 _2596_ _0199_ _2595_ sg13g2_a21oi_1
X_4906_ _1660_ _1662_ _1663_ VPWR VGND sg13g2_nor2_1
X_5886_ _2539_ VPWR _2540_ VGND net869 net805 sg13g2_o21ai_1
X_4837_ _1595_ _1587_ _1596_ VPWR VGND sg13g2_nor2b_1
XFILLER_21_565 VPWR VGND sg13g2_fill_2
XFILLER_14_1021 VPWR VGND sg13g2_decap_8
X_4768_ _1517_ VPWR _1529_ VGND _1525_ _1527_ sg13g2_o21ai_1
X_6507_ net1136 VGND VPWR net114 mac2.sum_lvl1_ff\[43\] clknet_leaf_49_clk sg13g2_dfrbpq_1
X_3719_ _0525_ _0519_ _0524_ VPWR VGND sg13g2_xnor2_1
X_4699_ _1438_ VPWR _1461_ VGND _1403_ _1436_ sg13g2_o21ai_1
X_6438_ net1122 VGND VPWR _0086_ mac2.products_ff\[2\] clknet_leaf_26_clk sg13g2_dfrbpq_1
XFILLER_0_403 VPWR VGND sg13g2_fill_2
X_6369_ net1081 VGND VPWR net258 mac2.sum_lvl1_ff\[85\] clknet_leaf_21_clk sg13g2_dfrbpq_1
Xhold22 mac1.sum_lvl1_ff\[3\] VPWR VGND net62 sg13g2_dlygate4sd3_1
Xhold11 mac2.sum_lvl1_ff\[81\] VPWR VGND net51 sg13g2_dlygate4sd3_1
Xhold33 mac1.sum_lvl1_ff\[6\] VPWR VGND net73 sg13g2_dlygate4sd3_1
Xhold55 mac1.products_ff\[137\] VPWR VGND net95 sg13g2_dlygate4sd3_1
Xhold44 mac2.products_ff\[11\] VPWR VGND net84 sg13g2_dlygate4sd3_1
Xhold77 mac2.sum_lvl1_ff\[14\] VPWR VGND net117 sg13g2_dlygate4sd3_1
Xhold99 mac1.sum_lvl1_ff\[44\] VPWR VGND net139 sg13g2_dlygate4sd3_1
XFILLER_28_131 VPWR VGND sg13g2_fill_1
Xhold66 mac2.sum_lvl1_ff\[82\] VPWR VGND net106 sg13g2_dlygate4sd3_1
Xhold88 mac2.products_ff\[141\] VPWR VGND net128 sg13g2_dlygate4sd3_1
XFILLER_17_827 VPWR VGND sg13g2_fill_1
XFILLER_45_43 VPWR VGND sg13g2_fill_2
XFILLER_45_32 VPWR VGND sg13g2_fill_1
XFILLER_45_98 VPWR VGND sg13g2_fill_2
XFILLER_44_679 VPWR VGND sg13g2_fill_2
XFILLER_40_830 VPWR VGND sg13g2_fill_1
Xfanout1020 net493 net1020 VPWR VGND sg13g2_buf_2
Xfanout1031 DP_1.matrix\[5\] net1031 VPWR VGND sg13g2_buf_8
Xfanout1042 DP_4.matrix\[80\] net1042 VPWR VGND sg13g2_buf_8
Xfanout1064 net1068 net1064 VPWR VGND sg13g2_buf_8
Xfanout1053 net527 net1053 VPWR VGND sg13g2_buf_8
XFILLER_48_963 VPWR VGND sg13g2_decap_8
Xfanout1075 net1076 net1075 VPWR VGND sg13g2_buf_8
Xfanout1097 net1099 net1097 VPWR VGND sg13g2_buf_8
Xfanout1086 net1087 net1086 VPWR VGND sg13g2_buf_8
XFILLER_16_882 VPWR VGND sg13g2_decap_8
X_5740_ _2397_ DP_1.I_range.out_data\[2\] DP_1.Q_range.out_data\[2\] VPWR VGND sg13g2_xnor2_1
X_5671_ _2340_ _2338_ net29 VPWR VGND sg13g2_xor2_1
X_4622_ net868 net865 net918 net916 _1387_ VPWR VGND sg13g2_and4_1
X_4553_ _1323_ _1309_ _1325_ VPWR VGND sg13g2_xor2_1
Xhold503 DP_2.matrix\[73\] VPWR VGND net543 sg13g2_dlygate4sd3_1
X_3504_ _0292_ VPWR _0315_ VGND _3031_ _0290_ sg13g2_o21ai_1
X_4484_ _1258_ _1252_ _1257_ VPWR VGND sg13g2_xnor2_1
X_3435_ _3010_ VPWR _3014_ VGND _3011_ _3012_ sg13g2_o21ai_1
X_6223_ net1139 VGND VPWR _0232_ DP_3.matrix\[40\] clknet_leaf_45_clk sg13g2_dfrbpq_2
X_6154_ net1072 VGND VPWR _0186_ DP_1.matrix\[42\] clknet_leaf_3_clk sg13g2_dfrbpq_2
X_3366_ _2950_ _2929_ _2951_ VPWR VGND sg13g2_nor2b_1
X_5105_ _1851_ net870 net829 net873 net825 VPWR VGND sg13g2_a22oi_1
X_3297_ _2882_ _2883_ _2884_ VPWR VGND sg13g2_nor2b_1
X_6085_ net1080 VGND VPWR net10 DP_3.Q_range.out_data\[3\] clknet_leaf_22_clk sg13g2_dfrbpq_1
X_5036_ _1784_ net875 net828 net877 net824 VPWR VGND sg13g2_a22oi_1
Xheichips25_template_35 VPWR VGND uio_oe[2] sg13g2_tiehi
X_5938_ _2586_ _2408_ _2428_ VPWR VGND sg13g2_xnor2_1
X_5869_ net1050 net804 _2524_ VPWR VGND sg13g2_nor2_1
XFILLER_22_896 VPWR VGND sg13g2_decap_8
Xoutput23 net23 uio_out[6] VPWR VGND sg13g2_buf_1
XFILLER_1_767 VPWR VGND sg13g2_decap_8
XFILLER_0_277 VPWR VGND sg13g2_fill_2
XFILLER_29_451 VPWR VGND sg13g2_decap_4
XFILLER_16_123 VPWR VGND sg13g2_fill_1
XFILLER_17_668 VPWR VGND sg13g2_fill_1
XFILLER_13_863 VPWR VGND sg13g2_decap_8
XFILLER_9_834 VPWR VGND sg13g2_decap_8
XFILLER_8_344 VPWR VGND sg13g2_fill_2
XFILLER_40_693 VPWR VGND sg13g2_fill_2
XFILLER_9_889 VPWR VGND sg13g2_decap_8
XFILLER_28_1009 VPWR VGND sg13g2_decap_8
X_3220_ _2806_ _2807_ _2789_ _2809_ VPWR VGND sg13g2_nand3_1
X_3151_ net1000 net928 net1003 _2741_ VPWR VGND net927 sg13g2_nand4_1
X_3082_ _2654_ VPWR _2675_ VGND _2645_ _2655_ sg13g2_o21ai_1
X_3984_ _0777_ net956 net1009 VPWR VGND sg13g2_nand2_1
X_5723_ _2379_ VPWR _2382_ VGND _2378_ _2380_ sg13g2_o21ai_1
X_5654_ net325 mac2.sum_lvl3_ff\[20\] _0048_ VPWR VGND sg13g2_xor2_1
X_4605_ net866 net920 net869 _1371_ VPWR VGND net918 sg13g2_nand4_1
X_5585_ mac2.sum_lvl3_ff\[1\] mac2.sum_lvl3_ff\[21\] _2274_ VPWR VGND sg13g2_xor2_1
Xhold300 mac1.sum_lvl2_ff\[4\] VPWR VGND net340 sg13g2_dlygate4sd3_1
Xhold311 _2221_ VPWR VGND net351 sg13g2_dlygate4sd3_1
Xhold344 DP_4.matrix\[3\] VPWR VGND net384 sg13g2_dlygate4sd3_1
Xhold322 DP_1.matrix\[44\] VPWR VGND net362 sg13g2_dlygate4sd3_1
X_4536_ _1308_ _1305_ _0130_ VPWR VGND sg13g2_xor2_1
Xhold333 DP_4.matrix\[37\] VPWR VGND net373 sg13g2_dlygate4sd3_1
Xhold355 _0014_ VPWR VGND net395 sg13g2_dlygate4sd3_1
Xhold377 _0202_ VPWR VGND net417 sg13g2_dlygate4sd3_1
Xhold366 DP_2.matrix\[3\] VPWR VGND net406 sg13g2_dlygate4sd3_1
X_4467_ _1242_ _1241_ _1214_ VPWR VGND sg13g2_nand2b_1
Xfanout824 net826 net824 VPWR VGND sg13g2_buf_8
Xfanout813 net324 net813 VPWR VGND sg13g2_buf_2
Xfanout802 _2398_ net802 VPWR VGND sg13g2_buf_2
X_3418_ _2997_ VPWR _3000_ VGND _2982_ _2999_ sg13g2_o21ai_1
X_4398_ _1170_ VPWR _1174_ VGND _1127_ _1172_ sg13g2_o21ai_1
Xhold388 _2206_ VPWR VGND net428 sg13g2_dlygate4sd3_1
Xhold399 _0054_ VPWR VGND net439 sg13g2_dlygate4sd3_1
X_6206_ net1105 VGND VPWR net423 DP_3.matrix\[1\] clknet_leaf_35_clk sg13g2_dfrbpq_2
Xfanout857 net371 net857 VPWR VGND sg13g2_buf_8
X_6137_ net1094 VGND VPWR _0175_ DP_1.matrix\[3\] clknet_leaf_61_clk sg13g2_dfrbpq_2
X_3349_ _2914_ VPWR _2934_ VGND _2912_ _2915_ sg13g2_o21ai_1
Xfanout846 DP_4.matrix\[37\] net846 VPWR VGND sg13g2_buf_8
Xfanout835 net335 net835 VPWR VGND sg13g2_buf_8
Xfanout879 net353 net879 VPWR VGND sg13g2_buf_1
Xfanout868 net374 net868 VPWR VGND sg13g2_buf_8
X_6068_ net850 _0252_ VPWR VGND sg13g2_buf_1
XFILLER_26_421 VPWR VGND sg13g2_fill_2
XFILLER_27_944 VPWR VGND sg13g2_decap_8
X_5019_ _1768_ _1756_ _1767_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_432 VPWR VGND sg13g2_fill_1
XFILLER_10_833 VPWR VGND sg13g2_decap_8
XFILLER_42_88 VPWR VGND sg13g2_fill_2
XFILLER_1_520 VPWR VGND sg13g2_fill_2
XFILLER_18_966 VPWR VGND sg13g2_decap_8
XFILLER_45_774 VPWR VGND sg13g2_fill_1
XFILLER_33_936 VPWR VGND sg13g2_fill_2
XFILLER_8_185 VPWR VGND sg13g2_fill_2
X_5370_ _2103_ VPWR _2106_ VGND _2102_ _2104_ sg13g2_o21ai_1
XFILLER_5_870 VPWR VGND sg13g2_decap_8
X_4321_ _1099_ net840 net899 VPWR VGND sg13g2_nand2_1
X_4252_ _1032_ net903 net838 VPWR VGND sg13g2_nand2_1
X_3203_ _2792_ net934 net992 VPWR VGND sg13g2_nand2_1
X_4183_ _0970_ _0969_ _0966_ VPWR VGND sg13g2_nand2b_1
XFILLER_41_1028 VPWR VGND sg13g2_fill_1
X_3134_ _2725_ _2718_ _2723_ _2724_ VPWR VGND sg13g2_and3_1
X_3065_ _2658_ net932 net1004 net934 net1000 VPWR VGND sg13g2_a22oi_1
XFILLER_24_947 VPWR VGND sg13g2_decap_8
X_3967_ _0760_ net1019 net948 VPWR VGND sg13g2_nand2_1
X_5706_ _2368_ mac1.total_sum\[12\] mac2.total_sum\[12\] VPWR VGND sg13g2_nand2_1
XFILLER_32_991 VPWR VGND sg13g2_decap_8
X_3898_ _0693_ net1017 net952 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_30_clk clknet_4_12_0_clk clknet_leaf_30_clk VPWR VGND sg13g2_buf_8
X_5637_ _2309_ _2306_ _2315_ VPWR VGND _2308_ sg13g2_nand3b_1
XFILLER_3_818 VPWR VGND sg13g2_decap_8
X_5568_ _2255_ VPWR _2261_ VGND _2256_ _2260_ sg13g2_o21ai_1
Xhold130 mac1.sum_lvl2_ff\[38\] VPWR VGND net170 sg13g2_dlygate4sd3_1
Xhold152 mac1.products_ff\[149\] VPWR VGND net192 sg13g2_dlygate4sd3_1
X_4519_ _1292_ _1286_ _1291_ VPWR VGND sg13g2_xnor2_1
Xhold141 mac1.products_ff\[15\] VPWR VGND net181 sg13g2_dlygate4sd3_1
Xhold174 mac2.products_ff\[72\] VPWR VGND net214 sg13g2_dlygate4sd3_1
X_5499_ _2204_ net428 _2199_ _2208_ VPWR VGND sg13g2_nand3_1
Xhold163 mac2.sum_lvl1_ff\[39\] VPWR VGND net203 sg13g2_dlygate4sd3_1
Xhold185 mac2.products_ff\[12\] VPWR VGND net225 sg13g2_dlygate4sd3_1
Xhold196 mac2.products_ff\[146\] VPWR VGND net236 sg13g2_dlygate4sd3_1
XFILLER_2_1022 VPWR VGND sg13g2_decap_8
XFILLER_15_925 VPWR VGND sg13g2_decap_8
XFILLER_18_1008 VPWR VGND sg13g2_decap_8
XFILLER_42_788 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_21_clk clknet_4_5_0_clk clknet_leaf_21_clk VPWR VGND sg13g2_buf_8
XFILLER_2_840 VPWR VGND sg13g2_decap_8
XFILLER_1_361 VPWR VGND sg13g2_fill_2
X_4870_ _1627_ _1624_ _1628_ VPWR VGND sg13g2_xor2_1
X_3821_ _0620_ net1018 net962 net958 net1021 VPWR VGND sg13g2_a22oi_1
XFILLER_33_788 VPWR VGND sg13g2_fill_2
XFILLER_20_416 VPWR VGND sg13g2_fill_1
XFILLER_20_449 VPWR VGND sg13g2_fill_2
X_6540_ net1137 VGND VPWR net191 mac2.sum_lvl2_ff\[27\] clknet_leaf_43_clk sg13g2_dfrbpq_1
X_3752_ _0556_ _0555_ _0557_ VPWR VGND sg13g2_nor2b_1
Xclkbuf_leaf_12_clk clknet_4_6_0_clk clknet_leaf_12_clk VPWR VGND sg13g2_buf_8
XFILLER_9_494 VPWR VGND sg13g2_decap_8
X_3683_ _0486_ _0488_ _0489_ _0490_ VPWR VGND sg13g2_nor3_1
X_6471_ net1086 VGND VPWR _0092_ mac2.products_ff\[139\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_5422_ _0003_ net320 _2147_ VPWR VGND sg13g2_xnor2_1
X_5353_ _2090_ _2077_ _2092_ VPWR VGND sg13g2_xor2_1
X_4304_ _1080_ _1079_ _1062_ _1083_ VPWR VGND sg13g2_a21o_1
X_5284_ _2025_ net817 net1045 VPWR VGND sg13g2_nand2_1
X_4235_ net849 net846 net900 net898 _1016_ VPWR VGND sg13g2_and4_1
X_4166_ _0952_ _0938_ _0954_ VPWR VGND sg13g2_xor2_1
X_3117_ _2708_ net1004 net928 VPWR VGND sg13g2_nand2_1
X_4097_ _0887_ _0881_ _0886_ VPWR VGND sg13g2_xnor2_1
X_3048_ _2641_ _2642_ _2643_ VPWR VGND sg13g2_nor2b_1
XFILLER_24_722 VPWR VGND sg13g2_fill_1
XFILLER_12_906 VPWR VGND sg13g2_decap_8
X_4999_ _1749_ _1740_ _1747_ VPWR VGND sg13g2_xnor2_1
XFILLER_7_409 VPWR VGND sg13g2_fill_2
XFILLER_20_950 VPWR VGND sg13g2_decap_8
XFILLER_47_814 VPWR VGND sg13g2_fill_1
XFILLER_47_858 VPWR VGND sg13g2_fill_2
XFILLER_46_335 VPWR VGND sg13g2_fill_1
XFILLER_14_243 VPWR VGND sg13g2_fill_2
XFILLER_11_994 VPWR VGND sg13g2_decap_8
XFILLER_31_1027 VPWR VGND sg13g2_fill_2
XFILLER_7_954 VPWR VGND sg13g2_decap_8
XFILLER_6_486 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_1_clk clknet_4_0_0_clk clknet_leaf_1_clk VPWR VGND sg13g2_buf_8
X_4020_ _0811_ _0760_ _0812_ VPWR VGND sg13g2_xor2_1
XFILLER_25_508 VPWR VGND sg13g2_fill_2
X_5971_ _2606_ VPWR _0221_ VGND net789 _2605_ sg13g2_o21ai_1
XFILLER_45_390 VPWR VGND sg13g2_fill_2
X_4922_ _1679_ _1616_ _1646_ VPWR VGND sg13g2_nand2_1
X_4853_ _1610_ _1586_ _1612_ VPWR VGND sg13g2_xor2_1
X_3804_ VPWR _0607_ _0606_ VGND sg13g2_inv_1
X_4784_ _1543_ _1498_ _0147_ VPWR VGND sg13g2_xor2_1
X_3735_ VGND VPWR _0540_ _0539_ _0487_ sg13g2_or2_1
X_6523_ net1143 VGND VPWR net221 mac2.sum_lvl2_ff\[7\] clknet_leaf_42_clk sg13g2_dfrbpq_1
X_6454_ net1122 VGND VPWR _0081_ mac2.products_ff\[70\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_5405_ _0015_ _2130_ _2133_ VPWR VGND sg13g2_xnor2_1
X_3666_ _0441_ VPWR _0473_ VGND _0388_ _0439_ sg13g2_o21ai_1
XFILLER_47_1001 VPWR VGND sg13g2_decap_8
X_3597_ net984 net980 net1025 net1058 _0406_ VPWR VGND sg13g2_and4_1
X_6385_ net1074 VGND VPWR net213 mac1.sum_lvl3_ff\[33\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_5336_ _2069_ VPWR _2075_ VGND _2046_ _2047_ sg13g2_o21ai_1
X_5267_ _2009_ _1962_ _2007_ VPWR VGND sg13g2_xnor2_1
X_4218_ net846 net902 net850 _1000_ VPWR VGND net900 sg13g2_nand4_1
X_5198_ _1942_ net1045 net826 net871 net822 VPWR VGND sg13g2_a22oi_1
X_4149_ _0937_ _0934_ _0119_ VPWR VGND sg13g2_xor2_1
XFILLER_7_239 VPWR VGND sg13g2_fill_2
Xclkload0 clknet_4_1_0_clk clkload0/X VPWR VGND sg13g2_buf_8
XFILLER_4_957 VPWR VGND sg13g2_decap_8
XFILLER_46_110 VPWR VGND sg13g2_fill_2
XFILLER_46_143 VPWR VGND sg13g2_fill_1
X_3520_ _0327_ _0328_ _0330_ _0331_ VPWR VGND sg13g2_or3_1
X_3451_ _3029_ _3028_ _3016_ VPWR VGND sg13g2_nand2b_1
X_6170_ net1091 VGND VPWR _0197_ DP_2.matrix\[1\] clknet_leaf_62_clk sg13g2_dfrbpq_1
X_3382_ _2966_ _2961_ _2964_ VPWR VGND sg13g2_xnor2_1
X_5121_ _1867_ _1864_ _1866_ VPWR VGND sg13g2_nand2_1
X_5052_ _0149_ _1772_ _1799_ VPWR VGND sg13g2_xnor2_1
X_4003_ _0723_ _0793_ _0795_ _0796_ VPWR VGND sg13g2_or3_1
X_5954_ _2596_ _2448_ _2459_ VPWR VGND sg13g2_xnor2_1
XFILLER_34_850 VPWR VGND sg13g2_fill_2
XFILLER_34_872 VPWR VGND sg13g2_fill_2
X_4905_ _1662_ net852 DP_3.matrix\[5\] net855 net912 VPWR VGND sg13g2_a22oi_1
X_5885_ VGND VPWR _2635_ net805 _2539_ net795 sg13g2_a21oi_1
XFILLER_40_319 VPWR VGND sg13g2_fill_2
X_4836_ _1595_ _1588_ _1594_ VPWR VGND sg13g2_xnor2_1
XFILLER_14_1000 VPWR VGND sg13g2_decap_8
X_6506_ net1136 VGND VPWR net131 mac2.sum_lvl1_ff\[42\] clknet_leaf_43_clk sg13g2_dfrbpq_1
X_4767_ _1517_ _1525_ _1527_ _1528_ VPWR VGND sg13g2_or3_1
X_3718_ _0523_ _0520_ _0524_ VPWR VGND sg13g2_xor2_1
X_4698_ _1452_ VPWR _1460_ VGND _1432_ _1453_ sg13g2_o21ai_1
X_3649_ _0455_ _0456_ _0457_ VPWR VGND sg13g2_nor2_1
X_6437_ net1106 VGND VPWR _0085_ mac2.products_ff\[1\] clknet_leaf_26_clk sg13g2_dfrbpq_1
X_6368_ net1076 VGND VPWR net232 mac2.sum_lvl1_ff\[84\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_5319_ _2059_ _2058_ _2055_ VPWR VGND sg13g2_nand2b_1
XFILLER_1_949 VPWR VGND sg13g2_decap_8
X_6299_ net1110 VGND VPWR net260 mac1.sum_lvl2_ff\[26\] clknet_leaf_56_clk sg13g2_dfrbpq_1
XFILLER_0_459 VPWR VGND sg13g2_decap_8
Xhold12 mac1.sum_lvl1_ff\[42\] VPWR VGND net52 sg13g2_dlygate4sd3_1
Xhold23 mac1.products_ff\[79\] VPWR VGND net63 sg13g2_dlygate4sd3_1
Xhold56 mac1.products_ff\[3\] VPWR VGND net96 sg13g2_dlygate4sd3_1
Xhold34 mac1.products_ff\[9\] VPWR VGND net74 sg13g2_dlygate4sd3_1
Xhold45 mac2.sum_lvl2_ff\[45\] VPWR VGND net85 sg13g2_dlygate4sd3_1
Xhold67 mac1.products_ff\[0\] VPWR VGND net107 sg13g2_dlygate4sd3_1
Xhold89 mac1.sum_lvl2_ff\[40\] VPWR VGND net129 sg13g2_dlygate4sd3_1
Xhold78 mac2.sum_lvl2_ff\[49\] VPWR VGND net118 sg13g2_dlygate4sd3_1
XFILLER_29_688 VPWR VGND sg13g2_fill_1
XFILLER_28_198 VPWR VGND sg13g2_fill_1
XFILLER_29_699 VPWR VGND sg13g2_decap_8
XFILLER_43_124 VPWR VGND sg13g2_fill_1
XFILLER_43_179 VPWR VGND sg13g2_fill_1
Xfanout1010 net1012 net1010 VPWR VGND sg13g2_buf_8
Xfanout1021 net1022 net1021 VPWR VGND sg13g2_buf_8
Xfanout1032 net1033 net1032 VPWR VGND sg13g2_buf_8
Xfanout1054 net418 net1054 VPWR VGND sg13g2_buf_8
Xfanout1065 net1066 net1065 VPWR VGND sg13g2_buf_8
Xfanout1043 net344 net1043 VPWR VGND sg13g2_buf_8
XFILLER_48_942 VPWR VGND sg13g2_decap_8
Xfanout1087 net1148 net1087 VPWR VGND sg13g2_buf_8
Xfanout1076 net1080 net1076 VPWR VGND sg13g2_buf_8
Xfanout1098 net1099 net1098 VPWR VGND sg13g2_buf_8
XFILLER_19_165 VPWR VGND sg13g2_fill_2
XFILLER_47_485 VPWR VGND sg13g2_fill_2
XFILLER_34_124 VPWR VGND sg13g2_fill_1
XFILLER_16_850 VPWR VGND sg13g2_fill_2
XFILLER_16_861 VPWR VGND sg13g2_decap_8
X_5670_ mac2.total_sum\[4\] mac1.total_sum\[4\] _2340_ VPWR VGND sg13g2_xor2_1
X_4621_ _1386_ net920 net862 VPWR VGND sg13g2_nand2_1
X_4552_ _1324_ _1309_ _1323_ VPWR VGND sg13g2_nand2_1
X_3503_ _0314_ _0306_ _0308_ VPWR VGND sg13g2_nand2_1
Xhold504 DP_1.matrix\[78\] VPWR VGND net544 sg13g2_dlygate4sd3_1
X_4483_ _1256_ _1253_ _1257_ VPWR VGND sg13g2_xor2_1
X_3434_ _3010_ _3011_ _3012_ _3013_ VPWR VGND sg13g2_nor3_1
X_6222_ net1097 VGND VPWR net200 mac1.sum_lvl1_ff\[14\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_6153_ net1131 VGND VPWR _0102_ mac1.products_ff\[143\] clknet_leaf_53_clk sg13g2_dfrbpq_1
X_3365_ _2948_ _2947_ _2950_ VPWR VGND sg13g2_xor2_1
X_5104_ net824 net873 net828 _1850_ VPWR VGND net870 sg13g2_nand4_1
X_3296_ _2878_ VPWR _2883_ VGND _2880_ _2881_ sg13g2_o21ai_1
X_6084_ net1080 VGND VPWR net9 DP_3.Q_range.out_data\[2\] clknet_leaf_22_clk sg13g2_dfrbpq_2
X_5035_ net824 net877 net829 _1783_ VPWR VGND net875 sg13g2_nand4_1
Xheichips25_template_36 VPWR VGND uio_oe[3] sg13g2_tiehi
XFILLER_39_986 VPWR VGND sg13g2_decap_8
XFILLER_38_485 VPWR VGND sg13g2_fill_2
XFILLER_14_809 VPWR VGND sg13g2_fill_1
XFILLER_15_36 VPWR VGND sg13g2_fill_1
X_5937_ net282 net786 _2585_ VPWR VGND sg13g2_nor2_1
XFILLER_22_820 VPWR VGND sg13g2_fill_2
XFILLER_25_168 VPWR VGND sg13g2_fill_2
X_5868_ _2523_ net1050 net791 VPWR VGND sg13g2_nand2_1
X_5799_ VGND VPWR _2417_ _2453_ _2455_ _2454_ sg13g2_a21oi_1
X_4819_ _1579_ _1548_ _1577_ VPWR VGND sg13g2_xnor2_1
Xoutput24 net24 uio_out[7] VPWR VGND sg13g2_buf_1
XFILLER_45_901 VPWR VGND sg13g2_fill_1
XFILLER_16_102 VPWR VGND sg13g2_fill_1
XFILLER_17_658 VPWR VGND sg13g2_fill_2
XFILLER_9_813 VPWR VGND sg13g2_decap_8
XFILLER_12_363 VPWR VGND sg13g2_fill_1
XFILLER_9_868 VPWR VGND sg13g2_decap_8
X_3150_ _2740_ net926 net1003 net928 net1000 VPWR VGND sg13g2_a22oi_1
X_3081_ _2674_ _2662_ _2673_ VPWR VGND sg13g2_xnor2_1
XFILLER_48_772 VPWR VGND sg13g2_fill_2
XFILLER_36_934 VPWR VGND sg13g2_fill_1
XFILLER_47_293 VPWR VGND sg13g2_fill_1
XFILLER_22_116 VPWR VGND sg13g2_decap_8
X_3983_ _0736_ VPWR _0776_ VGND _0734_ _0737_ sg13g2_o21ai_1
XFILLER_22_127 VPWR VGND sg13g2_fill_2
X_5722_ net23 _2378_ _2381_ VPWR VGND sg13g2_xnor2_1
X_5653_ _0054_ _2326_ net438 VPWR VGND sg13g2_xnor2_1
X_5584_ mac2.sum_lvl3_ff\[21\] mac2.sum_lvl3_ff\[1\] _2273_ VPWR VGND sg13g2_nor2_1
X_4604_ net869 net863 net920 net918 _1370_ VPWR VGND sg13g2_and4_1
Xhold301 _2114_ VPWR VGND net341 sg13g2_dlygate4sd3_1
X_4535_ VGND VPWR _1307_ _1308_ _1306_ _1248_ sg13g2_a21oi_2
Xhold323 DP_2.matrix\[36\] VPWR VGND net363 sg13g2_dlygate4sd3_1
Xhold312 _0040_ VPWR VGND net352 sg13g2_dlygate4sd3_1
Xhold334 DP_4.matrix\[0\] VPWR VGND net374 sg13g2_dlygate4sd3_1
Xhold345 _0247_ VPWR VGND net385 sg13g2_dlygate4sd3_1
Xhold356 DP_1.matrix\[4\] VPWR VGND net396 sg13g2_dlygate4sd3_1
Xhold367 _0199_ VPWR VGND net407 sg13g2_dlygate4sd3_1
Xhold378 DP_1.matrix\[80\] VPWR VGND net418 sg13g2_dlygate4sd3_1
X_4466_ _1239_ _1215_ _1241_ VPWR VGND sg13g2_xor2_1
Xfanout825 net826 net825 VPWR VGND sg13g2_buf_8
Xfanout814 DP_4.matrix\[78\] net814 VPWR VGND sg13g2_buf_8
Xfanout803 net804 net803 VPWR VGND sg13g2_buf_8
X_3417_ _0099_ _2982_ _2998_ VPWR VGND sg13g2_xnor2_1
X_4397_ _1172_ _1127_ _0136_ VPWR VGND sg13g2_xor2_1
Xhold389 _2207_ VPWR VGND net429 sg13g2_dlygate4sd3_1
X_6205_ net1127 VGND VPWR _0220_ DP_3.matrix\[0\] clknet_leaf_34_clk sg13g2_dfrbpq_1
Xfanout858 DP_4.matrix\[4\] net858 VPWR VGND sg13g2_buf_1
X_6136_ net1091 VGND VPWR _0174_ DP_1.matrix\[2\] clknet_leaf_61_clk sg13g2_dfrbpq_2
X_3348_ _2933_ _2932_ _2930_ VPWR VGND sg13g2_nand2b_1
Xfanout847 net373 net847 VPWR VGND sg13g2_buf_8
Xfanout836 DP_4.matrix\[42\] net836 VPWR VGND sg13g2_buf_1
Xfanout869 net374 net869 VPWR VGND sg13g2_buf_8
X_6067_ net276 _0243_ VPWR VGND sg13g2_buf_1
X_3279_ _2841_ VPWR _2866_ VGND _2839_ _2842_ sg13g2_o21ai_1
X_5018_ _1767_ _1764_ _1766_ VPWR VGND sg13g2_nand2_1
XFILLER_39_783 VPWR VGND sg13g2_fill_1
XFILLER_26_455 VPWR VGND sg13g2_decap_8
XFILLER_26_477 VPWR VGND sg13g2_fill_2
XFILLER_10_812 VPWR VGND sg13g2_decap_8
XFILLER_22_683 VPWR VGND sg13g2_decap_8
XFILLER_10_889 VPWR VGND sg13g2_decap_8
XFILLER_27_1021 VPWR VGND sg13g2_decap_8
XFILLER_18_945 VPWR VGND sg13g2_decap_8
XFILLER_45_742 VPWR VGND sg13g2_fill_1
XFILLER_17_499 VPWR VGND sg13g2_decap_4
XFILLER_32_447 VPWR VGND sg13g2_decap_4
XFILLER_9_643 VPWR VGND sg13g2_fill_1
XFILLER_34_1025 VPWR VGND sg13g2_decap_4
XFILLER_8_131 VPWR VGND sg13g2_fill_2
X_4320_ _1098_ net899 net838 VPWR VGND sg13g2_nand2_1
X_4251_ _1031_ net906 net837 VPWR VGND sg13g2_nand2_1
X_3202_ _2791_ net932 net991 VPWR VGND sg13g2_nand2_2
X_4182_ _0968_ _0941_ _0969_ VPWR VGND sg13g2_xor2_1
XFILLER_41_1007 VPWR VGND sg13g2_decap_8
X_3133_ _2719_ VPWR _2724_ VGND _2720_ _2722_ sg13g2_o21ai_1
X_3064_ _0067_ _2644_ _2656_ VPWR VGND sg13g2_xnor2_1
XFILLER_24_926 VPWR VGND sg13g2_decap_8
X_3966_ _0759_ net1023 DP_2.matrix\[44\] VPWR VGND sg13g2_nand2_1
XFILLER_23_458 VPWR VGND sg13g2_fill_2
XFILLER_32_970 VPWR VGND sg13g2_decap_8
X_5705_ net20 _2366_ _2367_ VPWR VGND sg13g2_xnor2_1
X_3897_ _0692_ net1021 net951 VPWR VGND sg13g2_nand2_1
X_5636_ _2309_ VPWR _2314_ VGND _2305_ _2308_ sg13g2_o21ai_1
X_5567_ _0035_ _2257_ _2260_ VPWR VGND sg13g2_xnor2_1
XFILLER_2_318 VPWR VGND sg13g2_fill_2
Xhold153 mac1.sum_lvl2_ff\[43\] VPWR VGND net193 sg13g2_dlygate4sd3_1
Xhold142 mac1.sum_lvl1_ff\[9\] VPWR VGND net182 sg13g2_dlygate4sd3_1
X_5498_ VGND VPWR _2199_ _2204_ _2207_ net428 sg13g2_a21oi_1
X_4518_ _1288_ _1290_ _1291_ VPWR VGND sg13g2_nor2_1
Xhold120 mac2.products_ff\[7\] VPWR VGND net160 sg13g2_dlygate4sd3_1
Xhold131 mac2.sum_lvl1_ff\[76\] VPWR VGND net171 sg13g2_dlygate4sd3_1
Xhold175 mac1.sum_lvl1_ff\[73\] VPWR VGND net215 sg13g2_dlygate4sd3_1
Xhold186 mac1.sum_lvl1_ff\[11\] VPWR VGND net226 sg13g2_dlygate4sd3_1
Xhold164 mac1.sum_lvl1_ff\[12\] VPWR VGND net204 sg13g2_dlygate4sd3_1
X_4449_ _1224_ _1217_ _1223_ VPWR VGND sg13g2_xnor2_1
Xhold197 mac1.products_ff\[73\] VPWR VGND net237 sg13g2_dlygate4sd3_1
XFILLER_46_506 VPWR VGND sg13g2_fill_2
X_6119_ net1083 VGND VPWR _0122_ mac1.products_ff\[83\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_2_1001 VPWR VGND sg13g2_decap_8
XFILLER_37_67 VPWR VGND sg13g2_fill_1
XFILLER_15_904 VPWR VGND sg13g2_decap_8
XFILLER_27_786 VPWR VGND sg13g2_fill_2
XFILLER_41_211 VPWR VGND sg13g2_fill_2
XFILLER_41_233 VPWR VGND sg13g2_fill_2
XFILLER_22_491 VPWR VGND sg13g2_fill_1
XFILLER_6_624 VPWR VGND sg13g2_fill_1
XFILLER_49_333 VPWR VGND sg13g2_fill_2
XFILLER_2_896 VPWR VGND sg13g2_decap_8
XFILLER_49_344 VPWR VGND sg13g2_fill_2
XFILLER_18_753 VPWR VGND sg13g2_fill_1
XFILLER_18_775 VPWR VGND sg13g2_fill_2
XFILLER_32_211 VPWR VGND sg13g2_fill_1
X_3820_ net962 net1021 net958 net1018 _0619_ VPWR VGND sg13g2_and4_1
XFILLER_21_929 VPWR VGND sg13g2_decap_8
XFILLER_32_244 VPWR VGND sg13g2_fill_1
XFILLER_33_778 VPWR VGND sg13g2_fill_2
X_3751_ VGND VPWR _0516_ _0527_ _0556_ _0515_ sg13g2_a21oi_1
X_3682_ _0489_ net1026 net975 net1027 net973 VPWR VGND sg13g2_a22oi_1
X_6470_ net1086 VGND VPWR _0091_ mac2.products_ff\[138\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_5421_ VPWR VGND _2146_ _2145_ _2137_ mac1.sum_lvl2_ff\[30\] _2147_ mac1.sum_lvl2_ff\[11\]
+ sg13g2_a221oi_1
X_5352_ VGND VPWR _2091_ _2090_ _2077_ sg13g2_or2_1
X_4303_ VGND VPWR _1079_ _1080_ _1082_ _1062_ sg13g2_a21oi_1
X_5283_ _2024_ net1045 net819 net870 net816 VPWR VGND sg13g2_a22oi_1
X_4234_ _1015_ net902 net842 VPWR VGND sg13g2_nand2_1
X_4165_ _0953_ _0938_ _0952_ VPWR VGND sg13g2_nand2_1
X_3116_ _2684_ VPWR _2707_ VGND _2659_ _2682_ sg13g2_o21ai_1
XFILLER_28_528 VPWR VGND sg13g2_decap_4
X_4096_ _0885_ _0882_ _0886_ VPWR VGND sg13g2_xor2_1
X_3047_ _2638_ VPWR _2642_ VGND _2639_ _2640_ sg13g2_o21ai_1
X_4998_ _1748_ _1740_ _1747_ VPWR VGND sg13g2_nand2_1
X_3949_ _0732_ _0740_ _0742_ _0743_ VPWR VGND sg13g2_or3_1
X_5619_ _2296_ _2298_ _2300_ VPWR VGND sg13g2_nor2_1
XFILLER_24_1024 VPWR VGND sg13g2_decap_4
XFILLER_47_837 VPWR VGND sg13g2_fill_2
XFILLER_19_528 VPWR VGND sg13g2_fill_2
XFILLER_46_369 VPWR VGND sg13g2_fill_1
XFILLER_27_583 VPWR VGND sg13g2_fill_2
XFILLER_14_233 VPWR VGND sg13g2_fill_2
XFILLER_14_255 VPWR VGND sg13g2_fill_1
XFILLER_31_1006 VPWR VGND sg13g2_decap_8
XFILLER_10_450 VPWR VGND sg13g2_fill_2
XFILLER_7_933 VPWR VGND sg13g2_decap_8
XFILLER_11_973 VPWR VGND sg13g2_decap_8
XFILLER_2_671 VPWR VGND sg13g2_fill_1
XFILLER_49_163 VPWR VGND sg13g2_fill_1
XFILLER_49_185 VPWR VGND sg13g2_fill_1
X_5970_ _2606_ net923 net789 VPWR VGND sg13g2_nand2_1
X_4921_ VGND VPWR _1615_ _1646_ _1678_ _1647_ sg13g2_a21oi_1
X_4852_ _1611_ _1586_ _1610_ VPWR VGND sg13g2_nand2_1
XFILLER_21_726 VPWR VGND sg13g2_fill_2
X_3803_ _0604_ _0591_ _0606_ VPWR VGND sg13g2_xor2_1
XFILLER_21_748 VPWR VGND sg13g2_decap_4
X_4783_ _1496_ _1497_ _1541_ _1542_ _1544_ VPWR VGND sg13g2_and4_1
X_3734_ _0539_ net971 net1058 VPWR VGND sg13g2_nand2_1
X_6522_ net1141 VGND VPWR net82 mac2.sum_lvl2_ff\[6\] clknet_leaf_44_clk sg13g2_dfrbpq_1
X_3665_ _0461_ VPWR _0472_ VGND _0445_ _0462_ sg13g2_o21ai_1
X_6453_ net1105 VGND VPWR _0080_ mac2.products_ff\[69\] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_5404_ _2133_ _2132_ _2131_ VPWR VGND sg13g2_nand2b_1
X_3596_ _0405_ net977 net1028 VPWR VGND sg13g2_nand2_1
X_6384_ net1073 VGND VPWR net104 mac1.sum_lvl3_ff\[32\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_5335_ VPWR _2074_ _2073_ VGND sg13g2_inv_1
X_5266_ VGND VPWR _2008_ _2007_ _1962_ sg13g2_or2_1
X_4217_ net850 net847 net902 net900 _0999_ VPWR VGND sg13g2_and4_1
X_5197_ net826 net823 net870 net1045 _1941_ VPWR VGND sg13g2_and4_1
X_4148_ VGND VPWR _0877_ _0935_ _0937_ _0936_ sg13g2_a21oi_1
X_4079_ _0868_ _0844_ _0870_ VPWR VGND sg13g2_xor2_1
XFILLER_11_203 VPWR VGND sg13g2_decap_4
XFILLER_12_748 VPWR VGND sg13g2_fill_1
Xclkload1 clknet_4_2_0_clk clkload1/X VPWR VGND sg13g2_buf_8
XFILLER_4_936 VPWR VGND sg13g2_decap_8
XFILLER_46_122 VPWR VGND sg13g2_fill_2
XFILLER_35_807 VPWR VGND sg13g2_fill_1
XFILLER_11_792 VPWR VGND sg13g2_fill_2
X_3450_ _3027_ _3017_ _3028_ VPWR VGND sg13g2_xor2_1
X_3381_ _2965_ _2964_ _2961_ VPWR VGND sg13g2_nand2b_1
X_5120_ _1863_ _1862_ _1832_ _1866_ VPWR VGND sg13g2_a21o_1
X_5051_ _1796_ _1770_ _1799_ VPWR VGND sg13g2_xor2_1
X_4002_ VGND VPWR _0791_ _0792_ _0795_ _0757_ sg13g2_a21oi_1
XFILLER_18_380 VPWR VGND sg13g2_fill_1
XFILLER_19_881 VPWR VGND sg13g2_decap_8
X_5953_ net974 net783 _2595_ VPWR VGND sg13g2_nor2_1
X_4904_ VGND VPWR _1661_ _1659_ _1635_ sg13g2_or2_1
X_5884_ _2538_ net376 net798 VPWR VGND sg13g2_nand2_1
X_4835_ _1593_ _1589_ _1594_ VPWR VGND sg13g2_xor2_1
X_4766_ VGND VPWR _1523_ _1524_ _1527_ _1518_ sg13g2_a21oi_1
X_3717_ _0523_ _0476_ _0521_ VPWR VGND sg13g2_xnor2_1
X_6505_ net1118 VGND VPWR net184 mac2.sum_lvl1_ff\[41\] clknet_leaf_47_clk sg13g2_dfrbpq_1
X_4697_ _1459_ _1458_ _0145_ VPWR VGND sg13g2_xor2_1
X_3648_ _0456_ net1059 net980 net1025 net977 VPWR VGND sg13g2_a22oi_1
X_6436_ net1103 VGND VPWR _0084_ mac2.products_ff\[0\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_3579_ _0388_ net1037 net967 VPWR VGND sg13g2_nand2_1
X_6367_ net1077 VGND VPWR net108 mac2.sum_lvl1_ff\[83\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_5318_ _2057_ _2031_ _2058_ VPWR VGND sg13g2_xor2_1
XFILLER_1_928 VPWR VGND sg13g2_decap_8
X_6298_ net1092 VGND VPWR net52 mac1.sum_lvl2_ff\[25\] clknet_leaf_62_clk sg13g2_dfrbpq_1
Xhold13 mac2.sum_lvl1_ff\[43\] VPWR VGND net53 sg13g2_dlygate4sd3_1
Xhold46 mac1.products_ff\[5\] VPWR VGND net86 sg13g2_dlygate4sd3_1
Xhold24 mac2.sum_lvl1_ff\[80\] VPWR VGND net64 sg13g2_dlygate4sd3_1
XFILLER_29_601 VPWR VGND sg13g2_fill_1
Xhold35 mac2.sum_lvl1_ff\[51\] VPWR VGND net75 sg13g2_dlygate4sd3_1
X_5249_ _1989_ _1991_ _1992_ VPWR VGND sg13g2_nor2_1
Xhold79 mac1.sum_lvl2_ff\[39\] VPWR VGND net119 sg13g2_dlygate4sd3_1
XFILLER_21_1027 VPWR VGND sg13g2_fill_2
Xhold68 mac2.products_ff\[147\] VPWR VGND net108 sg13g2_dlygate4sd3_1
XFILLER_29_656 VPWR VGND sg13g2_fill_2
Xhold57 mac2.sum_lvl2_ff\[42\] VPWR VGND net97 sg13g2_dlygate4sd3_1
XFILLER_17_818 VPWR VGND sg13g2_decap_8
XFILLER_45_45 VPWR VGND sg13g2_fill_1
XFILLER_44_637 VPWR VGND sg13g2_fill_2
XFILLER_25_851 VPWR VGND sg13g2_fill_1
XFILLER_43_147 VPWR VGND sg13g2_fill_2
XFILLER_12_512 VPWR VGND sg13g2_decap_8
XFILLER_40_843 VPWR VGND sg13g2_fill_2
Xfanout1011 net1012 net1011 VPWR VGND sg13g2_buf_1
Xfanout1022 net448 net1022 VPWR VGND sg13g2_buf_8
Xfanout1000 net1001 net1000 VPWR VGND sg13g2_buf_8
Xfanout1044 net327 net1044 VPWR VGND sg13g2_buf_8
Xfanout1033 net396 net1033 VPWR VGND sg13g2_buf_8
Xfanout1055 DP_1.matrix\[80\] net1055 VPWR VGND sg13g2_buf_1
Xfanout1088 net1108 net1088 VPWR VGND sg13g2_buf_8
XFILLER_0_994 VPWR VGND sg13g2_decap_8
Xfanout1066 net1067 net1066 VPWR VGND sg13g2_buf_8
Xfanout1077 net1079 net1077 VPWR VGND sg13g2_buf_8
XFILLER_48_998 VPWR VGND sg13g2_decap_8
Xfanout1099 net1107 net1099 VPWR VGND sg13g2_buf_8
XFILLER_37_1023 VPWR VGND sg13g2_decap_4
XFILLER_15_383 VPWR VGND sg13g2_fill_1
XFILLER_30_342 VPWR VGND sg13g2_fill_2
X_4620_ _1371_ VPWR _1385_ VGND _1369_ _1372_ sg13g2_o21ai_1
X_4551_ _1323_ _1296_ _1321_ VPWR VGND sg13g2_xnor2_1
X_3502_ _0105_ _0286_ _0313_ VPWR VGND sg13g2_xnor2_1
Xhold505 mac2.sum_lvl3_ff\[7\] VPWR VGND net545 sg13g2_dlygate4sd3_1
X_4482_ _1256_ _1230_ _1254_ VPWR VGND sg13g2_xnor2_1
X_3433_ _3012_ net1036 net982 net978 net1038 VPWR VGND sg13g2_a22oi_1
X_6221_ net1129 VGND VPWR _0231_ DP_3.matrix\[39\] clknet_leaf_33_clk sg13g2_dfrbpq_1
X_6152_ net1090 VGND VPWR _0185_ DP_1.matrix\[41\] clknet_leaf_65_clk sg13g2_dfrbpq_1
X_5103_ net829 net824 net873 net870 _1849_ VPWR VGND sg13g2_and4_1
XFILLER_44_1027 VPWR VGND sg13g2_fill_2
X_3364_ _2948_ _2947_ _2949_ VPWR VGND sg13g2_nor2b_1
XFILLER_32_0 VPWR VGND sg13g2_fill_2
X_6083_ net813 _0267_ VPWR VGND sg13g2_buf_1
X_3295_ _2878_ _2880_ _2881_ _2882_ VPWR VGND sg13g2_nor3_1
X_5034_ net828 net824 net878 net875 _1782_ VPWR VGND sg13g2_and4_1
Xheichips25_template_37 VPWR VGND uio_oe[4] sg13g2_tiehi
XFILLER_26_626 VPWR VGND sg13g2_fill_1
X_5936_ VGND VPWR net786 _2584_ _0176_ _2583_ sg13g2_a21oi_1
X_5867_ VGND VPWR _2516_ _2521_ _2522_ net792 sg13g2_a21oi_1
X_5798_ net978 _2417_ _2454_ VPWR VGND sg13g2_nor2_1
X_4818_ _1578_ _1548_ _1577_ VPWR VGND sg13g2_nand2_1
X_4749_ _1510_ _1463_ _1509_ VPWR VGND sg13g2_xnor2_1
Xoutput25 net25 uo_out[0] VPWR VGND sg13g2_buf_1
X_6419_ net1103 VGND VPWR net167 mac2.sum_lvl3_ff\[35\] clknet_leaf_26_clk sg13g2_dfrbpq_1
XFILLER_0_279 VPWR VGND sg13g2_fill_1
XFILLER_5_1010 VPWR VGND sg13g2_decap_8
XFILLER_45_979 VPWR VGND sg13g2_decap_8
XFILLER_25_670 VPWR VGND sg13g2_fill_1
XFILLER_8_346 VPWR VGND sg13g2_fill_1
XFILLER_13_898 VPWR VGND sg13g2_decap_8
XFILLER_40_695 VPWR VGND sg13g2_fill_1
XFILLER_4_596 VPWR VGND sg13g2_fill_2
X_3080_ _2673_ _2670_ _2672_ VPWR VGND sg13g2_nand2_1
XFILLER_0_791 VPWR VGND sg13g2_decap_8
X_3982_ _0775_ _0770_ _0774_ VPWR VGND sg13g2_xnor2_1
X_5721_ mac2.total_sum\[14\] mac1.total_sum\[14\] _2381_ VPWR VGND sg13g2_xor2_1
X_5652_ _2327_ net437 mac2.sum_lvl3_ff\[15\] VPWR VGND sg13g2_xnor2_1
XFILLER_30_183 VPWR VGND sg13g2_fill_1
X_5583_ _2272_ mac2.sum_lvl3_ff\[21\] mac2.sum_lvl3_ff\[1\] VPWR VGND sg13g2_nand2_1
X_4603_ _1369_ net923 net861 VPWR VGND sg13g2_nand2_1
Xhold302 _0010_ VPWR VGND net342 sg13g2_dlygate4sd3_1
XFILLER_11_1015 VPWR VGND sg13g2_decap_8
X_4534_ VGND VPWR _1245_ _1274_ _1307_ _1276_ sg13g2_a21oi_1
Xhold313 DP_3.matrix\[76\] VPWR VGND net353 sg13g2_dlygate4sd3_1
Xhold335 _0244_ VPWR VGND net375 sg13g2_dlygate4sd3_1
Xhold324 DP_4.matrix\[41\] VPWR VGND net364 sg13g2_dlygate4sd3_1
Xhold357 _0176_ VPWR VGND net397 sg13g2_dlygate4sd3_1
Xhold346 DP_2.matrix\[80\] VPWR VGND net386 sg13g2_dlygate4sd3_1
Xhold368 DP_1.matrix\[6\] VPWR VGND net408 sg13g2_dlygate4sd3_1
X_4465_ _1240_ _1215_ _1239_ VPWR VGND sg13g2_nand2_1
Xfanout815 net419 net815 VPWR VGND sg13g2_buf_1
Xhold379 DP_4.matrix\[78\] VPWR VGND net419 sg13g2_dlygate4sd3_1
X_6204_ net1114 VGND VPWR net77 mac1.sum_lvl1_ff\[8\] clknet_leaf_59_clk sg13g2_dfrbpq_1
X_3416_ VPWR _2999_ _2998_ VGND sg13g2_inv_1
X_4396_ _1125_ _1126_ _1170_ _1171_ _1173_ VPWR VGND sg13g2_and4_1
Xfanout804 _2479_ net804 VPWR VGND sg13g2_buf_8
Xfanout826 net827 net826 VPWR VGND sg13g2_buf_8
X_6135_ net1062 VGND VPWR _0065_ mac1.products_ff\[137\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3347_ VGND VPWR _2932_ _2931_ _2879_ sg13g2_or2_1
Xfanout848 net849 net848 VPWR VGND sg13g2_buf_2
Xfanout837 net364 net837 VPWR VGND sg13g2_buf_8
X_6066_ net279 _0242_ VPWR VGND sg13g2_buf_1
Xfanout859 net384 net859 VPWR VGND sg13g2_buf_8
X_3278_ _2833_ VPWR _2865_ VGND _2780_ _2831_ sg13g2_o21ai_1
X_5017_ _1763_ _1762_ _1757_ _1766_ VPWR VGND sg13g2_a21o_1
XFILLER_38_250 VPWR VGND sg13g2_fill_1
XFILLER_26_423 VPWR VGND sg13g2_fill_1
XFILLER_27_979 VPWR VGND sg13g2_decap_8
X_5919_ VGND VPWR _2563_ _2568_ _2573_ net791 sg13g2_a21oi_1
XFILLER_10_868 VPWR VGND sg13g2_decap_8
XFILLER_6_839 VPWR VGND sg13g2_decap_8
XFILLER_1_522 VPWR VGND sg13g2_fill_1
XFILLER_27_1000 VPWR VGND sg13g2_decap_8
XFILLER_18_924 VPWR VGND sg13g2_decap_8
XFILLER_45_732 VPWR VGND sg13g2_fill_1
XFILLER_17_478 VPWR VGND sg13g2_fill_1
XFILLER_34_1004 VPWR VGND sg13g2_decap_8
XFILLER_41_993 VPWR VGND sg13g2_decap_8
XFILLER_8_198 VPWR VGND sg13g2_fill_2
XFILLER_4_393 VPWR VGND sg13g2_fill_1
X_4250_ _1021_ VPWR _1030_ VGND _1013_ _1022_ sg13g2_o21ai_1
X_4181_ _0968_ net949 net1056 VPWR VGND sg13g2_nand2_1
X_3201_ _2790_ net996 net930 VPWR VGND sg13g2_nand2_1
X_3132_ _2719_ _2720_ _2722_ _2723_ VPWR VGND sg13g2_or3_1
X_3063_ _2657_ _2656_ VPWR VGND _2644_ sg13g2_nand2b_2
XFILLER_36_765 VPWR VGND sg13g2_fill_2
X_3965_ _0729_ VPWR _0758_ VGND _0726_ _0730_ sg13g2_o21ai_1
X_3896_ _0674_ VPWR _0691_ VGND _0665_ _0675_ sg13g2_o21ai_1
X_5704_ _2367_ _2360_ _2364_ VPWR VGND sg13g2_nand2_1
XFILLER_12_27 VPWR VGND sg13g2_fill_2
X_5635_ net530 mac2.sum_lvl3_ff\[32\] _2313_ VPWR VGND sg13g2_xor2_1
Xhold110 mac1.sum_lvl1_ff\[74\] VPWR VGND net150 sg13g2_dlygate4sd3_1
X_5566_ VPWR VGND _2259_ _2258_ _2250_ mac2.sum_lvl2_ff\[30\] _2260_ mac2.sum_lvl2_ff\[11\]
+ sg13g2_a221oi_1
Xhold121 mac1.sum_lvl2_ff\[41\] VPWR VGND net161 sg13g2_dlygate4sd3_1
Xhold143 mac1.products_ff\[4\] VPWR VGND net183 sg13g2_dlygate4sd3_1
X_5497_ _2206_ mac1.sum_lvl3_ff\[33\] net427 VPWR VGND sg13g2_xnor2_1
X_4517_ _1290_ net834 net897 net836 net895 VPWR VGND sg13g2_a22oi_1
Xhold132 mac2.products_ff\[151\] VPWR VGND net172 sg13g2_dlygate4sd3_1
Xhold176 mac1.sum_lvl2_ff\[44\] VPWR VGND net216 sg13g2_dlygate4sd3_1
Xhold165 mac2.sum_lvl2_ff\[46\] VPWR VGND net205 sg13g2_dlygate4sd3_1
X_4448_ _1222_ _1218_ _1223_ VPWR VGND sg13g2_xor2_1
Xhold154 mac2.sum_lvl1_ff\[86\] VPWR VGND net194 sg13g2_dlygate4sd3_1
Xhold198 mac2.products_ff\[71\] VPWR VGND net238 sg13g2_dlygate4sd3_1
Xhold187 mac2.sum_lvl1_ff\[5\] VPWR VGND net227 sg13g2_dlygate4sd3_1
X_4379_ VGND VPWR _1152_ _1153_ _1156_ _1147_ sg13g2_a21oi_1
X_6118_ net1083 VGND VPWR _0121_ mac1.products_ff\[82\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_6049_ net931 _0217_ VPWR VGND sg13g2_buf_1
XFILLER_42_735 VPWR VGND sg13g2_fill_2
XFILLER_22_470 VPWR VGND sg13g2_fill_1
XFILLER_23_993 VPWR VGND sg13g2_decap_8
XFILLER_2_875 VPWR VGND sg13g2_decap_8
XFILLER_37_518 VPWR VGND sg13g2_fill_2
XFILLER_45_540 VPWR VGND sg13g2_fill_2
XFILLER_21_908 VPWR VGND sg13g2_decap_8
XFILLER_14_993 VPWR VGND sg13g2_decap_8
X_3750_ _0553_ _0541_ _0555_ VPWR VGND sg13g2_xor2_1
X_3681_ net975 net973 net1027 net1026 _0488_ VPWR VGND sg13g2_and4_1
X_5420_ _2136_ _2140_ _2146_ VPWR VGND sg13g2_nor2_1
X_5351_ _2088_ _2078_ _2090_ VPWR VGND sg13g2_xor2_1
X_5282_ _2010_ _2005_ _2012_ _2023_ VPWR VGND sg13g2_a21o_1
X_4302_ _1079_ _1080_ _1062_ _1081_ VPWR VGND sg13g2_nand3_1
X_4233_ _1000_ VPWR _1014_ VGND _0998_ _1001_ sg13g2_o21ai_1
X_4164_ _0952_ _0925_ _0950_ VPWR VGND sg13g2_xnor2_1
X_3115_ _2706_ _2698_ _2700_ VPWR VGND sg13g2_nand2_1
X_4095_ _0885_ _0859_ _0883_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_507 VPWR VGND sg13g2_decap_8
X_3046_ _2638_ _2639_ _2640_ _2641_ VPWR VGND sg13g2_nor3_1
XFILLER_24_779 VPWR VGND sg13g2_decap_8
X_4997_ _1745_ _1746_ _1747_ VPWR VGND sg13g2_nor2b_1
X_3948_ VGND VPWR _0738_ _0739_ _0742_ _0733_ sg13g2_a21oi_1
XFILLER_32_790 VPWR VGND sg13g2_fill_2
X_3879_ VGND VPWR _0671_ _0672_ _0675_ _0666_ sg13g2_a21oi_1
XFILLER_20_985 VPWR VGND sg13g2_decap_8
X_5618_ _2298_ net456 _0062_ VPWR VGND sg13g2_nor2b_1
X_5549_ _2246_ _2245_ _2244_ VPWR VGND sg13g2_nand2b_1
XFILLER_24_1003 VPWR VGND sg13g2_decap_8
XFILLER_11_952 VPWR VGND sg13g2_decap_8
XFILLER_7_912 VPWR VGND sg13g2_decap_8
XFILLER_7_989 VPWR VGND sg13g2_decap_8
XFILLER_6_488 VPWR VGND sg13g2_fill_1
XFILLER_9_1008 VPWR VGND sg13g2_decap_8
XFILLER_46_860 VPWR VGND sg13g2_decap_4
X_4920_ _1675_ _1674_ _1677_ VPWR VGND sg13g2_xor2_1
X_4851_ _1609_ _1597_ _1610_ VPWR VGND sg13g2_xor2_1
X_3802_ VGND VPWR _0605_ _0604_ _0591_ sg13g2_or2_1
X_4782_ _1543_ _1541_ _1542_ VPWR VGND sg13g2_nand2_1
X_3733_ _0538_ net1058 net973 net1026 net971 VPWR VGND sg13g2_a22oi_1
X_6521_ net1139 VGND VPWR net227 mac2.sum_lvl2_ff\[5\] clknet_leaf_33_clk sg13g2_dfrbpq_2
X_3664_ VGND VPWR _0436_ _0442_ _0471_ _0444_ sg13g2_a21oi_1
X_6452_ net1103 VGND VPWR _0079_ mac2.products_ff\[68\] clknet_leaf_29_clk sg13g2_dfrbpq_1
X_5403_ VGND VPWR _2132_ mac1.sum_lvl2_ff\[9\] mac1.sum_lvl2_ff\[28\] sg13g2_or2_1
X_3595_ _0364_ VPWR _0404_ VGND _0362_ _0365_ sg13g2_o21ai_1
X_6383_ net1137 VGND VPWR net125 mac1.sum_lvl3_ff\[31\] clknet_leaf_49_clk sg13g2_dfrbpq_2
X_5334_ _2073_ _2049_ _2071_ VPWR VGND sg13g2_nand2_1
X_5265_ _2007_ net876 net815 VPWR VGND sg13g2_nand2_1
X_5196_ _1940_ net823 net1045 VPWR VGND sg13g2_nand2_1
X_4216_ _0998_ net905 net842 VPWR VGND sg13g2_nand2_1
X_4147_ VGND VPWR _0874_ _0903_ _0936_ _0905_ sg13g2_a21oi_1
X_4078_ _0869_ _0844_ _0868_ VPWR VGND sg13g2_nand2_1
XFILLER_11_226 VPWR VGND sg13g2_fill_1
Xclkload2 clknet_4_3_0_clk clkload2/X VPWR VGND sg13g2_buf_8
XFILLER_4_915 VPWR VGND sg13g2_decap_8
X_3380_ _2963_ _2937_ _2964_ VPWR VGND sg13g2_xor2_1
X_5050_ VGND VPWR _1794_ _1795_ _1798_ _1770_ sg13g2_a21oi_1
X_4001_ _0791_ _0792_ _0757_ _0794_ VPWR VGND sg13g2_nand3_1
XFILLER_38_668 VPWR VGND sg13g2_fill_2
X_5952_ VGND VPWR net786 _2594_ _0198_ _2593_ sg13g2_a21oi_1
X_4903_ net914 net911 net854 net852 _1660_ VPWR VGND sg13g2_and4_1
X_5883_ VGND VPWR net270 net797 _2537_ _2536_ sg13g2_a21oi_1
X_4834_ _1593_ _1552_ _1591_ VPWR VGND sg13g2_xnor2_1
X_4765_ _1523_ _1524_ _1518_ _1526_ VPWR VGND sg13g2_nand3_1
X_3716_ VGND VPWR _0522_ _0521_ _0476_ sg13g2_or2_1
X_6504_ net1118 VGND VPWR net214 mac2.sum_lvl1_ff\[40\] clknet_leaf_46_clk sg13g2_dfrbpq_1
XFILLER_20_16 VPWR VGND sg13g2_fill_2
X_4696_ _1425_ VPWR _1459_ VGND _1400_ _1426_ sg13g2_o21ai_1
X_3647_ net981 net977 net1025 net1059 _0455_ VPWR VGND sg13g2_and4_1
X_6435_ net1074 VGND VPWR net291 mac1.total_sum\[15\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_1_907 VPWR VGND sg13g2_decap_8
X_3578_ _0387_ net1041 net1053 VPWR VGND sg13g2_nand2_1
X_6366_ net1077 VGND VPWR net236 mac2.sum_lvl1_ff\[82\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_5317_ _2057_ net815 net872 VPWR VGND sg13g2_nand2_1
Xhold14 mac1.products_ff\[70\] VPWR VGND net54 sg13g2_dlygate4sd3_1
X_6297_ net1109 VGND VPWR net211 mac1.sum_lvl2_ff\[24\] clknet_leaf_55_clk sg13g2_dfrbpq_1
X_5248_ VGND VPWR _1990_ _1991_ _1956_ _1916_ sg13g2_a21oi_2
Xhold47 mac1.sum_lvl2_ff\[52\] VPWR VGND net87 sg13g2_dlygate4sd3_1
XFILLER_29_69 VPWR VGND sg13g2_fill_2
Xhold36 mac2.sum_lvl2_ff\[41\] VPWR VGND net76 sg13g2_dlygate4sd3_1
Xhold25 mac2.sum_lvl1_ff\[1\] VPWR VGND net65 sg13g2_dlygate4sd3_1
X_5179_ _1923_ net887 net1042 VPWR VGND sg13g2_nand2_1
Xhold69 mac1.sum_lvl1_ff\[82\] VPWR VGND net109 sg13g2_dlygate4sd3_1
XFILLER_21_1006 VPWR VGND sg13g2_decap_8
Xhold58 mac1.products_ff\[83\] VPWR VGND net98 sg13g2_dlygate4sd3_1
XFILLER_45_13 VPWR VGND sg13g2_fill_2
XFILLER_40_811 VPWR VGND sg13g2_fill_1
XFILLER_4_723 VPWR VGND sg13g2_fill_2
XFILLER_4_745 VPWR VGND sg13g2_fill_2
XFILLER_3_266 VPWR VGND sg13g2_fill_2
Xfanout1001 net1002 net1001 VPWR VGND sg13g2_buf_1
Xfanout1012 net323 net1012 VPWR VGND sg13g2_buf_2
Xfanout1045 net1046 net1045 VPWR VGND sg13g2_buf_8
Xfanout1023 net328 net1023 VPWR VGND sg13g2_buf_8
XFILLER_0_973 VPWR VGND sg13g2_decap_8
Xfanout1056 net362 net1056 VPWR VGND sg13g2_buf_8
Xfanout1034 net453 net1034 VPWR VGND sg13g2_buf_8
Xfanout1089 net1108 net1089 VPWR VGND sg13g2_buf_8
Xfanout1067 net1068 net1067 VPWR VGND sg13g2_buf_8
Xfanout1078 net1079 net1078 VPWR VGND sg13g2_buf_2
XFILLER_48_977 VPWR VGND sg13g2_decap_8
XFILLER_19_134 VPWR VGND sg13g2_decap_8
XFILLER_19_167 VPWR VGND sg13g2_fill_1
XFILLER_37_1002 VPWR VGND sg13g2_decap_8
XFILLER_16_896 VPWR VGND sg13g2_decap_8
XFILLER_31_855 VPWR VGND sg13g2_fill_2
X_4550_ _1322_ _1321_ _1296_ VPWR VGND sg13g2_nand2b_1
X_3501_ _0310_ _0284_ _0313_ VPWR VGND sg13g2_xor2_1
Xhold506 mac1.sum_lvl3_ff\[5\] VPWR VGND net546 sg13g2_dlygate4sd3_1
X_4481_ VGND VPWR _1255_ _1254_ _1230_ sg13g2_or2_1
X_3432_ net982 net1038 net978 net1036 _3011_ VPWR VGND sg13g2_and4_1
X_6220_ net1126 VGND VPWR _0230_ DP_3.matrix\[38\] clknet_leaf_33_clk sg13g2_dfrbpq_2
X_6151_ net1090 VGND VPWR _0184_ DP_1.matrix\[40\] clknet_leaf_65_clk sg13g2_dfrbpq_1
X_3363_ VGND VPWR _2908_ _2919_ _2948_ _2907_ sg13g2_a21oi_1
X_5102_ _1848_ net822 net875 VPWR VGND sg13g2_nand2_1
XFILLER_44_1006 VPWR VGND sg13g2_decap_8
X_6082_ net815 _0266_ VPWR VGND sg13g2_buf_1
X_3294_ _2881_ net987 net935 net989 net932 VPWR VGND sg13g2_a22oi_1
X_5033_ _1781_ net822 net880 VPWR VGND sg13g2_nand2_1
XFILLER_39_922 VPWR VGND sg13g2_decap_4
Xheichips25_template_38 VPWR VGND uio_oe[5] sg13g2_tiehi
X_5935_ _2584_ _2425_ _2427_ VPWR VGND sg13g2_xnor2_1
XFILLER_34_660 VPWR VGND sg13g2_fill_1
X_5866_ VPWR _2521_ _2520_ VGND sg13g2_inv_1
XFILLER_21_343 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_60_clk clknet_4_9_0_clk clknet_leaf_60_clk VPWR VGND sg13g2_buf_8
X_4817_ _1576_ _1559_ _1577_ VPWR VGND sg13g2_xor2_1
X_5797_ _2453_ net799 net961 net808 net942 VPWR VGND sg13g2_a22oi_1
X_4748_ _1509_ _1500_ _1507_ VPWR VGND sg13g2_xnor2_1
X_4679_ net867 net865 net914 net913 _1442_ VPWR VGND sg13g2_and4_1
X_6418_ net1084 VGND VPWR net92 mac2.sum_lvl3_ff\[34\] clknet_leaf_20_clk sg13g2_dfrbpq_1
Xoutput26 net26 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_0_225 VPWR VGND sg13g2_fill_1
X_6349_ net1132 VGND VPWR net228 mac1.sum_lvl1_ff\[81\] clknet_leaf_51_clk sg13g2_dfrbpq_1
XFILLER_45_936 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_51_clk clknet_4_10_0_clk clknet_leaf_51_clk VPWR VGND sg13g2_buf_8
XFILLER_13_877 VPWR VGND sg13g2_decap_8
XFILLER_8_336 VPWR VGND sg13g2_fill_2
XFILLER_0_770 VPWR VGND sg13g2_decap_8
XFILLER_48_774 VPWR VGND sg13g2_fill_1
X_3981_ _0774_ _0727_ _0772_ VPWR VGND sg13g2_xnor2_1
X_5720_ mac1.total_sum\[14\] mac2.total_sum\[14\] _2380_ VPWR VGND sg13g2_nor2_1
XFILLER_15_192 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_42_clk clknet_4_14_0_clk clknet_leaf_42_clk VPWR VGND sg13g2_buf_8
XFILLER_31_685 VPWR VGND sg13g2_decap_4
X_5651_ _2323_ VPWR _2326_ VGND _2322_ _2324_ sg13g2_o21ai_1
X_4602_ VGND VPWR _1368_ _1363_ _1361_ sg13g2_or2_1
X_5582_ _2271_ net480 net325 VPWR VGND sg13g2_nand2_1
XFILLER_8_892 VPWR VGND sg13g2_decap_8
X_4533_ VGND VPWR _1244_ _1274_ _1306_ _1276_ sg13g2_a21oi_1
Xhold325 mac1.sum_lvl2_ff\[29\] VPWR VGND net365 sg13g2_dlygate4sd3_1
Xhold303 DP_4.matrix\[36\] VPWR VGND net343 sg13g2_dlygate4sd3_1
Xhold314 DP_3.matrix\[44\] VPWR VGND net354 sg13g2_dlygate4sd3_1
Xhold347 DP_3.matrix\[3\] VPWR VGND net387 sg13g2_dlygate4sd3_1
X_6203_ net1116 VGND VPWR _0219_ DP_2.matrix\[79\] clknet_leaf_58_clk sg13g2_dfrbpq_2
Xhold369 _0178_ VPWR VGND net409 sg13g2_dlygate4sd3_1
X_4464_ _1238_ _1226_ _1239_ VPWR VGND sg13g2_xor2_1
Xhold358 DP_4.matrix\[39\] VPWR VGND net398 sg13g2_dlygate4sd3_1
Xhold336 DP_4.matrix\[72\] VPWR VGND net376 sg13g2_dlygate4sd3_1
Xfanout816 net817 net816 VPWR VGND sg13g2_buf_8
X_3415_ _2996_ _2983_ _2998_ VPWR VGND sg13g2_xor2_1
X_4395_ _1172_ _1170_ _1171_ VPWR VGND sg13g2_nand2_1
Xfanout805 _2479_ net805 VPWR VGND sg13g2_buf_8
X_6134_ net1091 VGND VPWR _0173_ DP_1.matrix\[1\] clknet_leaf_62_clk sg13g2_dfrbpq_2
X_3346_ _2931_ net930 net1054 VPWR VGND sg13g2_nand2_1
Xfanout849 DP_4.matrix\[36\] net849 VPWR VGND sg13g2_buf_8
Xfanout838 net330 net838 VPWR VGND sg13g2_buf_8
Xfanout827 net473 net827 VPWR VGND sg13g2_buf_2
X_6065_ net277 _0241_ VPWR VGND sg13g2_buf_1
X_5016_ VGND VPWR _1762_ _1763_ _1765_ _1757_ sg13g2_a21oi_1
X_3277_ _2853_ VPWR _2864_ VGND _2837_ _2854_ sg13g2_o21ai_1
XFILLER_27_925 VPWR VGND sg13g2_fill_2
XFILLER_27_958 VPWR VGND sg13g2_decap_8
XFILLER_26_479 VPWR VGND sg13g2_fill_1
X_5918_ VGND VPWR net278 net798 _2572_ _2571_ sg13g2_a21oi_1
XFILLER_22_652 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_33_clk clknet_4_12_0_clk clknet_leaf_33_clk VPWR VGND sg13g2_buf_8
X_5849_ _2503_ _2499_ _2504_ VPWR VGND sg13g2_nor2b_1
XFILLER_10_847 VPWR VGND sg13g2_decap_8
XFILLER_21_184 VPWR VGND sg13g2_decap_8
XFILLER_21_195 VPWR VGND sg13g2_fill_2
XFILLER_18_903 VPWR VGND sg13g2_decap_8
XFILLER_45_755 VPWR VGND sg13g2_fill_2
XFILLER_29_284 VPWR VGND sg13g2_fill_1
XFILLER_32_427 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_24_clk clknet_4_7_0_clk clknet_leaf_24_clk VPWR VGND sg13g2_buf_8
XFILLER_41_972 VPWR VGND sg13g2_decap_8
XFILLER_12_184 VPWR VGND sg13g2_fill_1
XFILLER_9_689 VPWR VGND sg13g2_fill_2
XFILLER_5_884 VPWR VGND sg13g2_decap_8
X_3200_ _2761_ VPWR _2789_ VGND _2752_ _2762_ sg13g2_o21ai_1
X_4180_ _0967_ net947 net1056 VPWR VGND sg13g2_nand2_1
X_3131_ _2722_ net989 net943 net992 net939 VPWR VGND sg13g2_a22oi_1
X_3062_ _2655_ _2645_ _2656_ VPWR VGND sg13g2_xor2_1
XFILLER_23_427 VPWR VGND sg13g2_decap_8
X_3964_ _0746_ VPWR _0757_ VGND _0724_ _0747_ sg13g2_o21ai_1
XFILLER_16_490 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_15_clk clknet_4_4_0_clk clknet_leaf_15_clk VPWR VGND sg13g2_buf_8
X_3895_ _0688_ _0687_ _0690_ VPWR VGND sg13g2_xor2_1
X_5703_ _2366_ mac1.total_sum\[11\] mac2.total_sum\[11\] VPWR VGND sg13g2_xnor2_1
X_5634_ _2312_ mac2.sum_lvl3_ff\[32\] mac2.sum_lvl3_ff\[12\] VPWR VGND sg13g2_nand2_1
X_5565_ _2249_ _2253_ _2259_ VPWR VGND sg13g2_nor2_1
Xhold100 mac2.products_ff\[144\] VPWR VGND net140 sg13g2_dlygate4sd3_1
X_5496_ _2204_ _2205_ _0019_ VPWR VGND sg13g2_and2_1
Xhold144 mac2.products_ff\[73\] VPWR VGND net184 sg13g2_dlygate4sd3_1
Xhold133 mac2.sum_lvl1_ff\[40\] VPWR VGND net173 sg13g2_dlygate4sd3_1
Xhold111 mac1.products_ff\[13\] VPWR VGND net151 sg13g2_dlygate4sd3_1
X_4516_ VGND VPWR _1289_ _1287_ _1262_ sg13g2_or2_1
Xhold122 mac2.sum_lvl2_ff\[47\] VPWR VGND net162 sg13g2_dlygate4sd3_1
Xhold177 mac1.products_ff\[69\] VPWR VGND net217 sg13g2_dlygate4sd3_1
Xhold166 mac1.sum_lvl1_ff\[45\] VPWR VGND net206 sg13g2_dlygate4sd3_1
X_4447_ _1222_ _1181_ _1220_ VPWR VGND sg13g2_xnor2_1
Xhold155 mac2.sum_lvl2_ff\[40\] VPWR VGND net195 sg13g2_dlygate4sd3_1
Xhold199 mac1.products_ff\[68\] VPWR VGND net239 sg13g2_dlygate4sd3_1
Xhold188 mac1.products_ff\[145\] VPWR VGND net228 sg13g2_dlygate4sd3_1
X_6117_ net1096 VGND VPWR _0120_ mac1.products_ff\[81\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_4378_ _1152_ _1153_ _1147_ _1155_ VPWR VGND sg13g2_nand3_1
X_3329_ _2915_ _2868_ _2913_ VPWR VGND sg13g2_xnor2_1
XFILLER_46_508 VPWR VGND sg13g2_fill_1
X_6048_ net933 _0216_ VPWR VGND sg13g2_buf_1
XFILLER_27_744 VPWR VGND sg13g2_fill_2
XFILLER_27_755 VPWR VGND sg13g2_fill_1
XFILLER_27_777 VPWR VGND sg13g2_decap_4
XFILLER_15_939 VPWR VGND sg13g2_decap_8
XFILLER_41_235 VPWR VGND sg13g2_fill_1
XFILLER_42_769 VPWR VGND sg13g2_fill_1
XFILLER_23_972 VPWR VGND sg13g2_decap_8
XFILLER_5_103 VPWR VGND sg13g2_fill_2
XFILLER_2_854 VPWR VGND sg13g2_decap_8
XFILLER_18_777 VPWR VGND sg13g2_fill_1
XFILLER_33_747 VPWR VGND sg13g2_fill_2
XFILLER_14_972 VPWR VGND sg13g2_decap_8
XFILLER_13_493 VPWR VGND sg13g2_decap_4
X_3680_ _0487_ net973 net1026 VPWR VGND sg13g2_nand2_1
X_5350_ _2088_ _2078_ _2089_ VPWR VGND sg13g2_nor2b_1
X_4301_ _1078_ _1077_ _1068_ _1080_ VPWR VGND sg13g2_a21o_1
X_5281_ _0151_ _2021_ _2022_ VPWR VGND sg13g2_xnor2_1
X_4232_ VPWR _1013_ _1012_ VGND sg13g2_inv_1
Xclkbuf_leaf_4_clk clknet_4_1_0_clk clknet_leaf_4_clk VPWR VGND sg13g2_buf_8
X_4163_ _0951_ _0950_ _0925_ VPWR VGND sg13g2_nand2b_1
X_3114_ _0094_ _2678_ _2705_ VPWR VGND sg13g2_xnor2_1
X_4094_ VGND VPWR _0884_ _0883_ _0859_ sg13g2_or2_1
X_3045_ _2640_ net999 net946 net942 net1002 VPWR VGND sg13g2_a22oi_1
XFILLER_36_585 VPWR VGND sg13g2_fill_1
X_4996_ _1741_ VPWR _1746_ VGND _1742_ _1744_ sg13g2_o21ai_1
XFILLER_24_747 VPWR VGND sg13g2_decap_4
X_3947_ _0738_ _0739_ _0733_ _0741_ VPWR VGND sg13g2_nand3_1
X_3878_ _0671_ _0672_ _0666_ _0674_ VPWR VGND sg13g2_nand3_1
XFILLER_20_964 VPWR VGND sg13g2_decap_8
X_5617_ _2294_ _2297_ net455 _2299_ VPWR VGND sg13g2_nand3_1
X_5548_ VGND VPWR _2245_ mac2.sum_lvl2_ff\[9\] mac2.sum_lvl2_ff\[28\] sg13g2_or2_1
X_5479_ _2191_ _2188_ _2190_ VPWR VGND sg13g2_nand2_1
XFILLER_47_839 VPWR VGND sg13g2_fill_1
XFILLER_19_508 VPWR VGND sg13g2_fill_1
XFILLER_11_931 VPWR VGND sg13g2_decap_8
XFILLER_23_791 VPWR VGND sg13g2_fill_2
XFILLER_10_452 VPWR VGND sg13g2_fill_1
XFILLER_7_968 VPWR VGND sg13g2_decap_8
XFILLER_49_132 VPWR VGND sg13g2_fill_2
X_4850_ _1607_ _1598_ _1609_ VPWR VGND sg13g2_xor2_1
XFILLER_33_533 VPWR VGND sg13g2_fill_2
X_3801_ _0602_ _0592_ _0604_ VPWR VGND sg13g2_xor2_1
XFILLER_33_588 VPWR VGND sg13g2_fill_2
XFILLER_20_227 VPWR VGND sg13g2_decap_8
X_6520_ net1129 VGND VPWR net198 mac2.sum_lvl2_ff\[4\] clknet_leaf_33_clk sg13g2_dfrbpq_1
X_4781_ _1539_ _1538_ _1540_ _1542_ VPWR VGND sg13g2_a21o_1
X_3732_ _0524_ _0519_ _0526_ _0537_ VPWR VGND sg13g2_a21o_1
X_6451_ net1146 VGND VPWR _0144_ mac2.products_ff\[15\] clknet_leaf_38_clk sg13g2_dfrbpq_1
X_3663_ _0470_ _0431_ _0115_ VPWR VGND sg13g2_xor2_1
Xclkload20 clknet_leaf_44_clk clkload20/X VPWR VGND sg13g2_buf_8
X_5402_ mac1.sum_lvl2_ff\[28\] mac1.sum_lvl2_ff\[9\] _2131_ VPWR VGND sg13g2_and2_1
X_6382_ net1133 VGND VPWR net187 mac1.sum_lvl3_ff\[30\] clknet_leaf_49_clk sg13g2_dfrbpq_2
X_3594_ _0403_ _0398_ _0402_ VPWR VGND sg13g2_xnor2_1
X_5333_ _0153_ _2071_ _2072_ VPWR VGND sg13g2_xnor2_1
XFILLER_47_1015 VPWR VGND sg13g2_decap_8
X_5264_ _2006_ net882 net1042 VPWR VGND sg13g2_nand2_1
X_5195_ _1893_ VPWR _1939_ VGND _1891_ _1894_ sg13g2_o21ai_1
X_4215_ VGND VPWR _0997_ _0992_ _0990_ sg13g2_or2_1
X_4146_ VGND VPWR _0873_ _0903_ _0935_ _0905_ sg13g2_a21oi_1
XFILLER_28_338 VPWR VGND sg13g2_fill_1
X_4077_ _0867_ _0855_ _0868_ VPWR VGND sg13g2_xor2_1
XFILLER_37_850 VPWR VGND sg13g2_decap_4
XFILLER_24_555 VPWR VGND sg13g2_fill_2
X_4979_ _1731_ net827 net890 net888 net832 VPWR VGND sg13g2_a22oi_1
Xclkload3 clknet_4_5_0_clk clkload3/X VPWR VGND sg13g2_buf_8
XFILLER_27_371 VPWR VGND sg13g2_fill_1
XFILLER_6_220 VPWR VGND sg13g2_fill_1
XFILLER_3_993 VPWR VGND sg13g2_decap_8
X_4000_ _0793_ _0757_ _0791_ _0792_ VPWR VGND sg13g2_and3_1
X_5951_ _2458_ _2456_ _2594_ VPWR VGND sg13g2_xor2_1
X_4902_ _1659_ net912 net852 VPWR VGND sg13g2_nand2_1
XFILLER_34_831 VPWR VGND sg13g2_fill_1
X_5882_ net794 _2534_ _2535_ _2536_ VPWR VGND sg13g2_nor3_1
X_4833_ VGND VPWR _1592_ _1590_ _1553_ sg13g2_or2_1
XFILLER_14_1014 VPWR VGND sg13g2_decap_8
X_4764_ _1525_ _1518_ _1523_ _1524_ VPWR VGND sg13g2_and3_1
X_3715_ _0521_ net1031 net969 VPWR VGND sg13g2_nand2_1
X_6503_ net1120 VGND VPWR net238 mac2.sum_lvl1_ff\[39\] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_6434_ net1066 VGND VPWR net333 mac1.total_sum\[14\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_4695_ _1458_ _1428_ _1456_ VPWR VGND sg13g2_xnor2_1
X_3646_ _0454_ net977 net1059 VPWR VGND sg13g2_nand2_1
X_3577_ _0357_ VPWR _0386_ VGND _0354_ _0358_ sg13g2_o21ai_1
X_6365_ net1079 VGND VPWR net121 mac2.sum_lvl1_ff\[81\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_5316_ _2056_ net872 net811 VPWR VGND sg13g2_nand2_1
X_6296_ net1109 VGND VPWR net255 mac1.sum_lvl2_ff\[23\] clknet_leaf_55_clk sg13g2_dfrbpq_1
X_5247_ VGND VPWR _1913_ _1955_ _1990_ _1954_ sg13g2_a21oi_1
Xhold37 mac1.products_ff\[8\] VPWR VGND net77 sg13g2_dlygate4sd3_1
Xhold15 mac2.sum_lvl1_ff\[45\] VPWR VGND net55 sg13g2_dlygate4sd3_1
Xhold26 mac2.sum_lvl1_ff\[36\] VPWR VGND net66 sg13g2_dlygate4sd3_1
X_5178_ _1887_ VPWR _1922_ VGND _1884_ _1888_ sg13g2_o21ai_1
Xhold48 mac1.sum_lvl1_ff\[4\] VPWR VGND net88 sg13g2_dlygate4sd3_1
Xhold59 mac1.sum_lvl1_ff\[49\] VPWR VGND net99 sg13g2_dlygate4sd3_1
X_4129_ VGND VPWR _0918_ _0916_ _0891_ sg13g2_or2_1
XFILLER_43_149 VPWR VGND sg13g2_fill_1
XFILLER_8_518 VPWR VGND sg13g2_fill_2
XFILLER_3_212 VPWR VGND sg13g2_fill_2
Xfanout1013 net1015 net1013 VPWR VGND sg13g2_buf_8
Xfanout1002 net515 net1002 VPWR VGND sg13g2_buf_8
Xfanout1046 DP_3.matrix\[80\] net1046 VPWR VGND sg13g2_buf_1
XFILLER_48_912 VPWR VGND sg13g2_decap_8
Xfanout1035 DP_1.matrix\[3\] net1035 VPWR VGND sg13g2_buf_8
Xfanout1024 DP_1.matrix\[36\] net1024 VPWR VGND sg13g2_buf_1
XFILLER_0_952 VPWR VGND sg13g2_decap_8
Xfanout1057 DP_1.matrix\[44\] net1057 VPWR VGND sg13g2_buf_1
Xfanout1068 net1087 net1068 VPWR VGND sg13g2_buf_8
Xfanout1079 net1080 net1079 VPWR VGND sg13g2_buf_8
XFILLER_48_956 VPWR VGND sg13g2_decap_8
XFILLER_16_875 VPWR VGND sg13g2_decap_8
XFILLER_31_823 VPWR VGND sg13g2_fill_2
X_3500_ VGND VPWR _0308_ _0309_ _0312_ _0284_ sg13g2_a21oi_1
Xhold507 _2173_ VPWR VGND net547 sg13g2_dlygate4sd3_1
X_4480_ _1254_ net841 net1048 VPWR VGND sg13g2_nand2_1
X_3431_ _3010_ net1040 net976 VPWR VGND sg13g2_nand2_1
X_6150_ net1116 VGND VPWR _0101_ mac1.products_ff\[142\] clknet_leaf_52_clk sg13g2_dfrbpq_1
X_3362_ _2945_ _2933_ _2947_ VPWR VGND sg13g2_xor2_1
X_5101_ _1815_ VPWR _1847_ VGND _1813_ _1816_ sg13g2_o21ai_1
XFILLER_32_2 VPWR VGND sg13g2_fill_1
X_6081_ net817 _0265_ VPWR VGND sg13g2_buf_1
X_3293_ net935 net932 net989 net987 _2880_ VPWR VGND sg13g2_and4_1
X_5032_ _1760_ VPWR _1780_ VGND _1758_ _1761_ sg13g2_o21ai_1
Xheichips25_template_39 VPWR VGND uio_oe[6] sg13g2_tiehi
XFILLER_38_444 VPWR VGND sg13g2_fill_1
X_5934_ net1033 net786 _2583_ VPWR VGND sg13g2_nor2_1
X_5865_ VGND VPWR net276 net798 _2520_ _2519_ sg13g2_a21oi_1
X_4816_ _1576_ _1560_ _1574_ VPWR VGND sg13g2_xnor2_1
X_5796_ _2449_ VPWR _2452_ VGND _2450_ _2451_ sg13g2_o21ai_1
X_4747_ _1508_ _1500_ _1507_ VPWR VGND sg13g2_nand2_1
X_4678_ _1441_ net861 net917 VPWR VGND sg13g2_nand2_1
X_3629_ _0437_ net1039 net1053 VPWR VGND sg13g2_nand2_1
X_6417_ net1081 VGND VPWR net105 mac2.sum_lvl3_ff\[33\] clknet_leaf_20_clk sg13g2_dfrbpq_1
Xoutput27 net27 uo_out[2] VPWR VGND sg13g2_buf_1
X_6348_ net1111 VGND VPWR net176 mac1.sum_lvl1_ff\[80\] clknet_leaf_54_clk sg13g2_dfrbpq_1
X_6279_ net1088 VGND VPWR net62 mac1.sum_lvl2_ff\[3\] clknet_leaf_64_clk sg13g2_dfrbpq_1
XFILLER_44_414 VPWR VGND sg13g2_fill_2
XFILLER_29_488 VPWR VGND sg13g2_decap_4
XFILLER_44_458 VPWR VGND sg13g2_fill_1
XFILLER_25_661 VPWR VGND sg13g2_decap_8
XFILLER_12_300 VPWR VGND sg13g2_fill_2
XFILLER_9_827 VPWR VGND sg13g2_decap_8
XFILLER_13_856 VPWR VGND sg13g2_decap_8
XFILLER_4_554 VPWR VGND sg13g2_fill_1
XFILLER_48_742 VPWR VGND sg13g2_fill_2
X_3980_ VGND VPWR _0773_ _0771_ _0728_ sg13g2_or2_1
XFILLER_44_992 VPWR VGND sg13g2_decap_8
XFILLER_31_620 VPWR VGND sg13g2_fill_2
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
X_5650_ _0053_ _2322_ net298 VPWR VGND sg13g2_xnor2_1
X_4601_ _1367_ net924 net859 VPWR VGND sg13g2_nand2_1
X_5581_ net271 mac2.sum_lvl2_ff\[19\] _0032_ VPWR VGND sg13g2_xor2_1
XFILLER_8_871 VPWR VGND sg13g2_decap_8
X_4532_ _1303_ _1302_ _1305_ VPWR VGND sg13g2_xor2_1
Xhold315 DP_3.matrix\[0\] VPWR VGND net355 sg13g2_dlygate4sd3_1
Xhold326 _2134_ VPWR VGND net366 sg13g2_dlygate4sd3_1
X_4463_ _1236_ _1227_ _1238_ VPWR VGND sg13g2_xor2_1
Xhold304 DP_4.matrix\[44\] VPWR VGND net344 sg13g2_dlygate4sd3_1
Xhold348 _0223_ VPWR VGND net388 sg13g2_dlygate4sd3_1
X_6202_ net1116 VGND VPWR _0218_ DP_2.matrix\[78\] clknet_leaf_58_clk sg13g2_dfrbpq_2
Xhold359 DP_1.matrix\[43\] VPWR VGND net399 sg13g2_dlygate4sd3_1
Xhold337 DP_2.matrix\[7\] VPWR VGND net377 sg13g2_dlygate4sd3_1
X_3414_ VGND VPWR _2997_ _2996_ _2983_ sg13g2_or2_1
X_4394_ _1168_ _1167_ _1169_ _1171_ VPWR VGND sg13g2_a21o_1
Xfanout806 _2478_ net806 VPWR VGND sg13g2_buf_8
Xfanout817 net318 net817 VPWR VGND sg13g2_buf_2
X_6133_ net1093 VGND VPWR _0172_ DP_1.matrix\[0\] clknet_leaf_62_clk sg13g2_dfrbpq_1
X_3345_ _2930_ net1054 net932 net988 net930 VPWR VGND sg13g2_a22oi_1
Xfanout839 DP_4.matrix\[40\] net839 VPWR VGND sg13g2_buf_1
Xfanout828 net830 net828 VPWR VGND sg13g2_buf_8
X_6064_ net879 _0240_ VPWR VGND sg13g2_buf_1
X_3276_ VGND VPWR _2828_ _2834_ _2863_ _2836_ sg13g2_a21oi_1
X_5015_ _1762_ _1763_ _1757_ _1764_ VPWR VGND sg13g2_nand3_1
XFILLER_27_915 VPWR VGND sg13g2_fill_1
XFILLER_26_414 VPWR VGND sg13g2_decap_8
X_5917_ net796 _2569_ _2570_ _2571_ VPWR VGND sg13g2_nor3_1
XFILLER_35_992 VPWR VGND sg13g2_decap_8
XFILLER_41_439 VPWR VGND sg13g2_fill_1
XFILLER_10_826 VPWR VGND sg13g2_decap_8
XFILLER_21_141 VPWR VGND sg13g2_fill_1
XFILLER_21_152 VPWR VGND sg13g2_fill_1
XFILLER_22_675 VPWR VGND sg13g2_fill_2
X_5848_ VGND VPWR net885 net798 _2503_ _2502_ sg13g2_a21oi_1
X_5779_ net786 VPWR _2436_ VGND _2433_ _2435_ sg13g2_o21ai_1
XFILLER_17_414 VPWR VGND sg13g2_fill_2
XFILLER_18_959 VPWR VGND sg13g2_decap_8
XFILLER_26_992 VPWR VGND sg13g2_decap_8
XFILLER_8_101 VPWR VGND sg13g2_fill_2
XFILLER_12_152 VPWR VGND sg13g2_fill_2
XFILLER_5_863 VPWR VGND sg13g2_decap_8
XFILLER_4_340 VPWR VGND sg13g2_fill_2
XFILLER_4_362 VPWR VGND sg13g2_fill_1
X_3130_ net939 net992 net943 _2721_ VPWR VGND net989 sg13g2_nand4_1
X_3061_ _2655_ _2646_ _2653_ VPWR VGND sg13g2_xnor2_1
XFILLER_36_767 VPWR VGND sg13g2_fill_1
XFILLER_17_981 VPWR VGND sg13g2_decap_8
X_3963_ _0755_ _0754_ _0124_ VPWR VGND sg13g2_xor2_1
X_3894_ _0689_ _0687_ _0688_ VPWR VGND sg13g2_nand2b_1
X_5702_ mac1.total_sum\[11\] mac2.total_sum\[11\] _2365_ VPWR VGND sg13g2_nor2_1
XFILLER_31_450 VPWR VGND sg13g2_decap_8
XFILLER_31_461 VPWR VGND sg13g2_fill_1
XFILLER_32_984 VPWR VGND sg13g2_decap_8
X_5633_ _0050_ _2310_ net402 VPWR VGND sg13g2_xnor2_1
X_5564_ _2247_ _2252_ _2258_ VPWR VGND sg13g2_nor2_1
X_4515_ _1262_ _1287_ _1288_ VPWR VGND sg13g2_nor2_1
Xhold101 mac2.sum_lvl1_ff\[50\] VPWR VGND net141 sg13g2_dlygate4sd3_1
Xhold134 mac1.sum_lvl2_ff\[46\] VPWR VGND net174 sg13g2_dlygate4sd3_1
X_5495_ net541 _2201_ _2203_ _2205_ VPWR VGND sg13g2_or3_1
Xhold112 mac2.sum_lvl1_ff\[74\] VPWR VGND net152 sg13g2_dlygate4sd3_1
Xhold123 mac2.sum_lvl1_ff\[73\] VPWR VGND net163 sg13g2_dlygate4sd3_1
Xhold167 mac1.products_ff\[140\] VPWR VGND net207 sg13g2_dlygate4sd3_1
X_4446_ VGND VPWR _1221_ _1219_ _1182_ sg13g2_or2_1
Xhold156 mac2.products_ff\[143\] VPWR VGND net196 sg13g2_dlygate4sd3_1
Xhold145 mac2.products_ff\[0\] VPWR VGND net185 sg13g2_dlygate4sd3_1
Xhold189 mac1.sum_lvl1_ff\[86\] VPWR VGND net229 sg13g2_dlygate4sd3_1
X_4377_ _1154_ _1147_ _1152_ _1153_ VPWR VGND sg13g2_and3_1
Xhold178 mac2.products_ff\[69\] VPWR VGND net218 sg13g2_dlygate4sd3_1
X_3328_ VGND VPWR _2914_ _2913_ _2868_ sg13g2_or2_1
X_6116_ net1089 VGND VPWR _0119_ mac1.products_ff\[80\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_6047_ net934 _0215_ VPWR VGND sg13g2_buf_1
X_3259_ net938 net936 net986 net1055 _2847_ VPWR VGND sg13g2_and4_1
XFILLER_2_1015 VPWR VGND sg13g2_decap_8
XFILLER_15_918 VPWR VGND sg13g2_decap_8
XFILLER_26_266 VPWR VGND sg13g2_fill_1
XFILLER_42_737 VPWR VGND sg13g2_fill_1
XFILLER_23_951 VPWR VGND sg13g2_decap_8
XFILLER_42_759 VPWR VGND sg13g2_fill_2
XFILLER_10_612 VPWR VGND sg13g2_fill_1
XFILLER_22_483 VPWR VGND sg13g2_decap_4
XFILLER_2_833 VPWR VGND sg13g2_decap_8
XFILLER_18_734 VPWR VGND sg13g2_fill_1
XFILLER_45_542 VPWR VGND sg13g2_fill_1
XFILLER_17_233 VPWR VGND sg13g2_fill_2
XFILLER_14_951 VPWR VGND sg13g2_decap_8
XFILLER_9_421 VPWR VGND sg13g2_fill_2
XFILLER_9_487 VPWR VGND sg13g2_decap_8
X_4300_ _1077_ _1078_ _1068_ _1079_ VPWR VGND sg13g2_nand3_1
X_5280_ _1987_ _1992_ _2022_ VPWR VGND sg13g2_nor2_1
X_4231_ _1009_ _1011_ _1012_ VPWR VGND sg13g2_nor2_1
X_4162_ _0948_ _0910_ _0950_ VPWR VGND sg13g2_xor2_1
X_3113_ _2702_ _2676_ _2705_ VPWR VGND sg13g2_xor2_1
X_4093_ _0883_ net954 net1056 VPWR VGND sg13g2_nand2_1
X_3044_ net946 net1002 net942 net999 _2639_ VPWR VGND sg13g2_and4_1
X_4995_ _1741_ _1742_ _1744_ _1745_ VPWR VGND sg13g2_nor3_1
X_3946_ _0740_ _0733_ _0738_ _0739_ VPWR VGND sg13g2_and3_1
XFILLER_17_1023 VPWR VGND sg13g2_decap_4
XFILLER_20_943 VPWR VGND sg13g2_decap_8
XFILLER_32_792 VPWR VGND sg13g2_fill_1
X_3877_ _0673_ _0666_ _0671_ _0672_ VPWR VGND sg13g2_and3_1
X_5616_ VGND VPWR net455 _2294_ _2298_ _2297_ sg13g2_a21oi_1
XFILLER_3_608 VPWR VGND sg13g2_fill_2
X_5547_ mac2.sum_lvl2_ff\[28\] mac2.sum_lvl2_ff\[9\] _2244_ VPWR VGND sg13g2_and2_1
X_5478_ _0031_ _2187_ net510 VPWR VGND sg13g2_xnor2_1
X_4429_ _1205_ _1189_ _1203_ VPWR VGND sg13g2_xnor2_1
XFILLER_11_910 VPWR VGND sg13g2_decap_8
XFILLER_7_947 VPWR VGND sg13g2_decap_8
XFILLER_11_987 VPWR VGND sg13g2_decap_8
XFILLER_49_111 VPWR VGND sg13g2_fill_2
XFILLER_38_80 VPWR VGND sg13g2_fill_2
X_3800_ _0602_ _0592_ _0603_ VPWR VGND sg13g2_nor2b_1
X_4780_ _1539_ _1540_ _1538_ _1541_ VPWR VGND sg13g2_nand3_1
X_3731_ _0107_ _0535_ _0536_ VPWR VGND sg13g2_xnor2_1
XFILLER_9_251 VPWR VGND sg13g2_fill_2
X_6450_ net1145 VGND VPWR _0143_ mac2.products_ff\[14\] clknet_leaf_38_clk sg13g2_dfrbpq_1
X_3662_ _0468_ _0469_ _0470_ VPWR VGND sg13g2_nor2b_2
Xclkload10 clknet_4_14_0_clk clkload10/X VPWR VGND sg13g2_buf_8
X_5401_ net392 net458 net394 _2130_ VPWR VGND sg13g2_a21o_1
X_6381_ net1138 VGND VPWR net186 mac1.sum_lvl3_ff\[29\] clknet_leaf_51_clk sg13g2_dfrbpq_2
X_3593_ _0402_ _0355_ _0400_ VPWR VGND sg13g2_xnor2_1
Xclkload21 clkload21/Y clknet_leaf_45_clk VPWR VGND sg13g2_inv_2
X_5332_ VGND VPWR _2049_ _2052_ _2072_ _2048_ sg13g2_a21oi_1
X_5263_ VGND VPWR _2005_ _1976_ _1974_ sg13g2_or2_1
X_5194_ _1938_ _1933_ _1937_ VPWR VGND sg13g2_xnor2_1
X_4214_ _0996_ net906 net840 VPWR VGND sg13g2_nand2_1
X_4145_ _0932_ _0931_ _0934_ VPWR VGND sg13g2_xor2_1
X_4076_ _0865_ _0856_ _0867_ VPWR VGND sg13g2_xor2_1
XFILLER_24_501 VPWR VGND sg13g2_decap_4
XFILLER_12_718 VPWR VGND sg13g2_fill_1
X_4978_ _1730_ net888 net827 _0089_ VPWR VGND sg13g2_and3_2
X_3929_ _0723_ _0719_ _0722_ VPWR VGND sg13g2_nand2_1
Xclkload4 clknet_4_6_0_clk clkload4/X VPWR VGND sg13g2_buf_8
XFILLER_30_1020 VPWR VGND sg13g2_decap_8
X_6579_ net1065 VGND VPWR net403 mac2.total_sum\[11\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_46_103 VPWR VGND sg13g2_fill_2
XFILLER_43_821 VPWR VGND sg13g2_fill_2
XFILLER_15_512 VPWR VGND sg13g2_fill_2
XFILLER_15_523 VPWR VGND sg13g2_decap_4
XFILLER_11_740 VPWR VGND sg13g2_fill_2
XFILLER_11_773 VPWR VGND sg13g2_fill_2
XFILLER_6_276 VPWR VGND sg13g2_fill_2
XFILLER_40_81 VPWR VGND sg13g2_fill_1
XFILLER_3_972 VPWR VGND sg13g2_decap_8
X_5950_ net976 net786 _2593_ VPWR VGND sg13g2_nor2_1
X_4901_ _1658_ net917 net1044 VPWR VGND sg13g2_nand2_1
XFILLER_19_895 VPWR VGND sg13g2_decap_8
XFILLER_34_865 VPWR VGND sg13g2_decap_8
X_5881_ net840 net807 _2535_ VPWR VGND sg13g2_nor2_1
X_4832_ _1591_ net917 net854 VPWR VGND sg13g2_nand2_1
X_4763_ _1519_ VPWR _1524_ VGND _1520_ _1522_ sg13g2_o21ai_1
X_3714_ _0520_ net1035 net1053 VPWR VGND sg13g2_nand2_1
X_6502_ net1122 VGND VPWR net154 mac2.sum_lvl1_ff\[38\] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_4694_ _1456_ _1428_ _1457_ VPWR VGND sg13g2_nor2b_1
X_6433_ net1066 VGND VPWR net430 mac1.total_sum\[13\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_3645_ _0407_ VPWR _0453_ VGND _0405_ _0408_ sg13g2_o21ai_1
X_3576_ _0374_ VPWR _0385_ VGND _0352_ _0375_ sg13g2_o21ai_1
X_6364_ net1076 VGND VPWR net140 mac2.sum_lvl1_ff\[80\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_5315_ _2055_ net876 net1042 VPWR VGND sg13g2_nand2_1
X_6295_ net1088 VGND VPWR net147 mac1.sum_lvl2_ff\[22\] clknet_leaf_64_clk sg13g2_dfrbpq_1
X_5246_ _1989_ _1988_ _1987_ VPWR VGND sg13g2_nand2b_1
Xhold38 mac1.sum_lvl1_ff\[37\] VPWR VGND net78 sg13g2_dlygate4sd3_1
Xhold16 mac1.sum_lvl1_ff\[15\] VPWR VGND net56 sg13g2_dlygate4sd3_1
Xhold27 mac2.products_ff\[138\] VPWR VGND net67 sg13g2_dlygate4sd3_1
X_5177_ _1875_ _1878_ _1921_ VPWR VGND sg13g2_nor2_1
Xhold49 mac2.sum_lvl1_ff\[48\] VPWR VGND net89 sg13g2_dlygate4sd3_1
X_4128_ _0891_ _0916_ _0917_ VPWR VGND sg13g2_nor2_1
X_4059_ VGND VPWR _0850_ _0848_ _0811_ sg13g2_or2_1
XFILLER_37_670 VPWR VGND sg13g2_fill_2
XFILLER_43_139 VPWR VGND sg13g2_fill_2
XFILLER_24_397 VPWR VGND sg13g2_fill_1
XFILLER_25_898 VPWR VGND sg13g2_decap_4
XFILLER_40_868 VPWR VGND sg13g2_decap_8
Xfanout1003 net424 net1003 VPWR VGND sg13g2_buf_8
XFILLER_0_931 VPWR VGND sg13g2_decap_8
Xfanout1014 net1015 net1014 VPWR VGND sg13g2_buf_1
Xfanout1036 net425 net1036 VPWR VGND sg13g2_buf_8
Xfanout1025 DP_1.matrix\[7\] net1025 VPWR VGND sg13g2_buf_2
Xfanout1047 net354 net1047 VPWR VGND sg13g2_buf_8
XFILLER_48_935 VPWR VGND sg13g2_decap_8
XFILLER_47_423 VPWR VGND sg13g2_fill_2
Xfanout1069 net1072 net1069 VPWR VGND sg13g2_buf_8
Xfanout1058 DP_1.matrix\[8\] net1058 VPWR VGND sg13g2_buf_8
XFILLER_19_158 VPWR VGND sg13g2_decap_8
XFILLER_16_832 VPWR VGND sg13g2_decap_8
XFILLER_42_194 VPWR VGND sg13g2_fill_1
Xhold508 mac2.sum_lvl2_ff\[24\] VPWR VGND net548 sg13g2_dlygate4sd3_1
X_3430_ _3008_ _3009_ _0070_ VPWR VGND sg13g2_nor2_2
X_3361_ VGND VPWR _2946_ _2945_ _2933_ sg13g2_or2_1
X_5100_ _1846_ _1840_ _1845_ VPWR VGND sg13g2_xnor2_1
X_6080_ net269 _0264_ VPWR VGND sg13g2_buf_1
X_5031_ _1777_ _1774_ _1779_ VPWR VGND sg13g2_xor2_1
X_3292_ _2879_ net932 net988 VPWR VGND sg13g2_nand2_1
XFILLER_39_979 VPWR VGND sg13g2_decap_8
X_5933_ VGND VPWR net784 _2582_ _0175_ _2581_ sg13g2_a21oi_1
X_5864_ net796 _2517_ _2518_ _2519_ VPWR VGND sg13g2_nor3_1
XFILLER_33_150 VPWR VGND sg13g2_fill_2
X_4815_ _1575_ _1560_ _1574_ VPWR VGND sg13g2_nand2_1
X_5795_ net799 VPWR _2451_ VGND net965 net808 sg13g2_o21ai_1
X_4746_ _1505_ _1501_ _1507_ VPWR VGND sg13g2_xor2_1
X_4677_ _1411_ VPWR _1440_ VGND _1409_ _1412_ sg13g2_o21ai_1
X_3628_ _0401_ VPWR _0436_ VGND _0398_ _0402_ sg13g2_o21ai_1
X_6416_ net1077 VGND VPWR net50 mac2.sum_lvl3_ff\[32\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_6347_ net1132 VGND VPWR net90 mac1.sum_lvl1_ff\[79\] clknet_leaf_53_clk sg13g2_dfrbpq_1
Xoutput28 net28 uo_out[3] VPWR VGND sg13g2_buf_1
Xoutput17 net17 uio_out[0] VPWR VGND sg13g2_buf_1
XFILLER_0_205 VPWR VGND sg13g2_fill_1
X_3559_ _0366_ _0367_ _0361_ _0369_ VPWR VGND sg13g2_nand3_1
X_6278_ net1069 VGND VPWR net234 mac1.sum_lvl2_ff\[2\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_5229_ _1972_ net876 net816 VPWR VGND sg13g2_nand2_1
XFILLER_5_1024 VPWR VGND sg13g2_decap_4
XFILLER_8_338 VPWR VGND sg13g2_fill_1
XFILLER_47_275 VPWR VGND sg13g2_fill_2
XFILLER_16_640 VPWR VGND sg13g2_fill_1
XFILLER_44_971 VPWR VGND sg13g2_decap_8
XFILLER_22_109 VPWR VGND sg13g2_decap_8
XFILLER_43_492 VPWR VGND sg13g2_fill_1
X_4600_ _1365_ _1358_ _0086_ VPWR VGND sg13g2_xor2_1
X_5580_ _0038_ _2269_ net485 VPWR VGND sg13g2_xnor2_1
XFILLER_7_360 VPWR VGND sg13g2_fill_1
X_4531_ _1302_ _1303_ _1304_ VPWR VGND sg13g2_nor2_1
Xhold305 DP_3.matrix\[6\] VPWR VGND net345 sg13g2_dlygate4sd3_1
X_4462_ _1237_ _1227_ _1236_ VPWR VGND sg13g2_nand2b_1
Xhold316 DP_3.matrix\[41\] VPWR VGND net356 sg13g2_dlygate4sd3_1
Xhold349 mac1.sum_lvl2_ff\[2\] VPWR VGND net389 sg13g2_dlygate4sd3_1
X_6201_ net1115 VGND VPWR net81 mac1.sum_lvl1_ff\[7\] clknet_leaf_57_clk sg13g2_dfrbpq_1
Xhold338 _0203_ VPWR VGND net378 sg13g2_dlygate4sd3_1
X_3413_ _2994_ _2984_ _2996_ VPWR VGND sg13g2_xor2_1
Xhold327 _2141_ VPWR VGND net367 sg13g2_dlygate4sd3_1
X_4393_ _1168_ _1169_ _1167_ _1170_ VPWR VGND sg13g2_nand3_1
Xfanout807 _2478_ net807 VPWR VGND sg13g2_buf_1
Xfanout829 net830 net829 VPWR VGND sg13g2_buf_1
Xfanout818 net819 net818 VPWR VGND sg13g2_buf_8
X_6132_ net1062 VGND VPWR _0064_ mac1.products_ff\[136\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3344_ _2916_ _2911_ _2918_ _2929_ VPWR VGND sg13g2_a21o_1
X_6063_ net882 _0239_ VPWR VGND sg13g2_buf_1
X_3275_ _2862_ _2823_ _0104_ VPWR VGND sg13g2_xor2_1
X_5014_ _1758_ VPWR _1763_ VGND _1759_ _1761_ sg13g2_o21ai_1
XFILLER_27_927 VPWR VGND sg13g2_fill_1
X_5916_ net1043 net806 _2570_ VPWR VGND sg13g2_nor2_1
XFILLER_10_805 VPWR VGND sg13g2_decap_8
X_5847_ net795 _2500_ _2501_ _2502_ VPWR VGND sg13g2_nor3_1
X_5778_ _2435_ net800 _2434_ net802 DP_1.matrix\[79\] VPWR VGND sg13g2_a22oi_1
X_4729_ _1466_ VPWR _1491_ VGND _1487_ _1489_ sg13g2_o21ai_1
XFILLER_27_1014 VPWR VGND sg13g2_decap_8
XFILLER_17_404 VPWR VGND sg13g2_fill_2
XFILLER_18_938 VPWR VGND sg13g2_decap_8
XFILLER_44_234 VPWR VGND sg13g2_fill_1
XFILLER_26_971 VPWR VGND sg13g2_decap_8
XFILLER_32_429 VPWR VGND sg13g2_fill_1
XFILLER_34_1018 VPWR VGND sg13g2_decap_8
XFILLER_12_197 VPWR VGND sg13g2_fill_2
XFILLER_5_842 VPWR VGND sg13g2_decap_8
X_3060_ _2654_ _2646_ _2653_ VPWR VGND sg13g2_nand2_1
XFILLER_17_960 VPWR VGND sg13g2_decap_8
XFILLER_24_919 VPWR VGND sg13g2_decap_8
X_3962_ _0756_ _0754_ _0755_ VPWR VGND sg13g2_nand2_1
X_5701_ net19 _2362_ _2363_ VPWR VGND sg13g2_xnor2_1
X_3893_ _0688_ net1024 net950 VPWR VGND sg13g2_nand2_1
X_5632_ _2311_ _2305_ _2307_ VPWR VGND sg13g2_nand2_1
X_5563_ mac2.sum_lvl2_ff\[12\] mac2.sum_lvl2_ff\[31\] _2257_ VPWR VGND sg13g2_xor2_1
X_4514_ _1287_ net895 net834 VPWR VGND sg13g2_nand2_2
Xhold135 mac1.products_ff\[76\] VPWR VGND net175 sg13g2_dlygate4sd3_1
Xhold102 mac1.sum_lvl1_ff\[0\] VPWR VGND net142 sg13g2_dlygate4sd3_1
Xhold124 mac1.sum_lvl1_ff\[72\] VPWR VGND net164 sg13g2_dlygate4sd3_1
X_5494_ net541 VPWR _2204_ VGND _2201_ _2203_ sg13g2_o21ai_1
Xhold113 mac2.products_ff\[140\] VPWR VGND net153 sg13g2_dlygate4sd3_1
Xhold146 mac1.sum_lvl2_ff\[47\] VPWR VGND net186 sg13g2_dlygate4sd3_1
Xhold168 mac1.sum_lvl1_ff\[51\] VPWR VGND net208 sg13g2_dlygate4sd3_1
X_4445_ _1220_ net899 net836 VPWR VGND sg13g2_nand2_1
Xhold157 mac1.sum_lvl1_ff\[13\] VPWR VGND net197 sg13g2_dlygate4sd3_1
Xhold179 mac1.products_ff\[1\] VPWR VGND net219 sg13g2_dlygate4sd3_1
X_4376_ _1148_ VPWR _1153_ VGND _1149_ _1151_ sg13g2_o21ai_1
X_3327_ _2913_ net991 net928 VPWR VGND sg13g2_nand2_1
X_6115_ net1098 VGND VPWR _0118_ mac1.products_ff\[79\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_6046_ net936 _0214_ VPWR VGND sg13g2_buf_1
X_3258_ _2846_ net936 net1055 VPWR VGND sg13g2_nand2_1
XFILLER_39_540 VPWR VGND sg13g2_fill_2
X_3189_ _2749_ VPWR _2778_ VGND _2746_ _2750_ sg13g2_o21ai_1
XFILLER_27_746 VPWR VGND sg13g2_fill_1
XFILLER_23_930 VPWR VGND sg13g2_decap_8
XFILLER_5_105 VPWR VGND sg13g2_fill_1
XFILLER_2_812 VPWR VGND sg13g2_decap_8
XFILLER_2_889 VPWR VGND sg13g2_decap_8
XFILLER_40_1022 VPWR VGND sg13g2_decap_8
XFILLER_14_930 VPWR VGND sg13g2_decap_8
XFILLER_9_411 VPWR VGND sg13g2_fill_1
X_4230_ net906 net904 net840 net838 _1011_ VPWR VGND sg13g2_and4_1
X_4161_ _0910_ _0948_ _0949_ VPWR VGND sg13g2_nor2_1
X_3112_ VGND VPWR _2700_ _2701_ _2704_ _2676_ sg13g2_a21oi_1
X_4092_ _0882_ net951 net1008 VPWR VGND sg13g2_nand2_1
XFILLER_49_871 VPWR VGND sg13g2_decap_8
X_3043_ _2638_ net1003 net937 VPWR VGND sg13g2_nand2_1
X_4994_ _1744_ net880 net830 net883 net825 VPWR VGND sg13g2_a22oi_1
X_3945_ _0734_ VPWR _0739_ VGND _0735_ _0737_ sg13g2_o21ai_1
XFILLER_17_1002 VPWR VGND sg13g2_decap_8
XFILLER_20_922 VPWR VGND sg13g2_decap_8
X_3876_ _0667_ VPWR _0672_ VGND _0668_ _0670_ sg13g2_o21ai_1
X_5615_ _2297_ mac2.sum_lvl3_ff\[28\] mac2.sum_lvl3_ff\[8\] VPWR VGND sg13g2_xnor2_1
XFILLER_20_999 VPWR VGND sg13g2_decap_8
X_5546_ mac2.sum_lvl2_ff\[8\] mac2.sum_lvl2_ff\[27\] _2241_ _2243_ VPWR VGND sg13g2_a21o_1
X_5477_ _2189_ VPWR _2190_ VGND _2183_ _2185_ sg13g2_o21ai_1
X_4428_ _1204_ _1189_ _1203_ VPWR VGND sg13g2_nand2_1
XFILLER_24_1017 VPWR VGND sg13g2_decap_8
X_4359_ _1134_ _1130_ _1136_ VPWR VGND sg13g2_xor2_1
XFILLER_24_1028 VPWR VGND sg13g2_fill_1
X_6029_ net1001 _0189_ VPWR VGND sg13g2_buf_1
XFILLER_42_502 VPWR VGND sg13g2_fill_2
XFILLER_30_708 VPWR VGND sg13g2_fill_2
XFILLER_23_793 VPWR VGND sg13g2_fill_1
XFILLER_7_926 VPWR VGND sg13g2_decap_8
XFILLER_11_966 VPWR VGND sg13g2_decap_8
XFILLER_13_40 VPWR VGND sg13g2_fill_2
XFILLER_49_156 VPWR VGND sg13g2_fill_1
XFILLER_49_134 VPWR VGND sg13g2_fill_1
Xfanout990 net544 net990 VPWR VGND sg13g2_buf_8
XFILLER_46_841 VPWR VGND sg13g2_decap_4
XFILLER_18_565 VPWR VGND sg13g2_fill_2
XFILLER_33_513 VPWR VGND sg13g2_fill_2
XFILLER_33_535 VPWR VGND sg13g2_fill_1
X_3730_ _0501_ _0506_ _0536_ VPWR VGND sg13g2_nor2_1
X_3661_ _0469_ _0432_ _0467_ VPWR VGND sg13g2_nand2_1
X_5400_ net394 _2129_ _0014_ VPWR VGND sg13g2_nor2b_1
X_6380_ net1111 VGND VPWR net174 mac1.sum_lvl3_ff\[28\] clknet_leaf_54_clk sg13g2_dfrbpq_1
X_3592_ VGND VPWR _0401_ _0399_ _0356_ sg13g2_or2_1
Xclkload11 clknet_4_15_0_clk clkload11/X VPWR VGND sg13g2_buf_8
Xclkload22 clkload22/Y clknet_leaf_34_clk VPWR VGND sg13g2_inv_2
X_5331_ _2069_ _2070_ _2071_ VPWR VGND sg13g2_and2_1
X_5262_ _1964_ VPWR _2004_ VGND _1961_ _1965_ sg13g2_o21ai_1
X_5193_ _1937_ _1885_ _1934_ VPWR VGND sg13g2_xnor2_1
X_4213_ _0994_ _0987_ _0081_ VPWR VGND sg13g2_xor2_1
X_4144_ _0931_ _0932_ _0933_ VPWR VGND sg13g2_nor2_1
XFILLER_49_690 VPWR VGND sg13g2_fill_2
X_4075_ _0866_ _0856_ _0865_ VPWR VGND sg13g2_nand2b_1
X_4977_ net890 net832 _0089_ VPWR VGND sg13g2_and2_1
X_3928_ _0720_ _0721_ _0722_ VPWR VGND sg13g2_nor2b_1
Xclkload5 clknet_4_7_0_clk clkload5/X VPWR VGND sg13g2_buf_8
X_3859_ _0654_ _0655_ _0656_ VPWR VGND sg13g2_nor2b_2
X_6578_ net1065 VGND VPWR net348 mac2.total_sum\[10\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_4_929 VPWR VGND sg13g2_decap_8
X_5529_ net469 mac2.sum_lvl2_ff\[24\] _2230_ VPWR VGND sg13g2_xor2_1
XFILLER_8_1011 VPWR VGND sg13g2_decap_8
XFILLER_43_844 VPWR VGND sg13g2_fill_2
XFILLER_7_723 VPWR VGND sg13g2_fill_2
XFILLER_3_951 VPWR VGND sg13g2_decap_8
XFILLER_19_852 VPWR VGND sg13g2_fill_2
XFILLER_19_874 VPWR VGND sg13g2_decap_8
X_4900_ _1626_ VPWR _1657_ VGND _1624_ _1627_ sg13g2_o21ai_1
X_5880_ net859 net804 _2534_ VPWR VGND sg13g2_nor2_1
X_4831_ _1590_ net917 net852 VPWR VGND sg13g2_nand2_1
X_4762_ _1519_ _1520_ _1522_ _1523_ VPWR VGND sg13g2_or3_1
X_3713_ VGND VPWR _0519_ _0490_ _0488_ sg13g2_or2_1
X_6501_ net1105 VGND VPWR net218 mac2.sum_lvl1_ff\[37\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_4693_ _1456_ _1432_ _1455_ VPWR VGND sg13g2_xnor2_1
X_3644_ _0452_ _0447_ _0451_ VPWR VGND sg13g2_xnor2_1
X_6432_ net1065 VGND VPWR _0019_ mac1.total_sum\[12\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_3575_ _0383_ _0382_ _0113_ VPWR VGND sg13g2_xor2_1
X_6363_ net1079 VGND VPWR net196 mac2.sum_lvl1_ff\[79\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_5314_ _2033_ VPWR _2054_ VGND _2030_ _2034_ sg13g2_o21ai_1
X_6294_ net1069 VGND VPWR net68 mac1.sum_lvl2_ff\[21\] clknet_leaf_66_clk sg13g2_dfrbpq_1
X_5245_ _1952_ _1986_ _1950_ _1988_ VPWR VGND sg13g2_nand3_1
Xhold28 mac1.sum_lvl1_ff\[38\] VPWR VGND net68 sg13g2_dlygate4sd3_1
Xhold17 mac1.products_ff\[147\] VPWR VGND net57 sg13g2_dlygate4sd3_1
X_5176_ _1903_ VPWR _1920_ VGND _1882_ _1904_ sg13g2_o21ai_1
Xhold39 mac1.sum_lvl1_ff\[87\] VPWR VGND net79 sg13g2_dlygate4sd3_1
X_4127_ _0916_ net1008 net947 VPWR VGND sg13g2_nand2_2
X_4058_ _0849_ net1013 net949 VPWR VGND sg13g2_nand2_1
XFILLER_25_844 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_63_clk clknet_4_2_0_clk clknet_leaf_63_clk VPWR VGND sg13g2_buf_8
XFILLER_12_505 VPWR VGND sg13g2_decap_8
XFILLER_40_836 VPWR VGND sg13g2_decap_8
XFILLER_0_910 VPWR VGND sg13g2_decap_8
Xfanout1004 net424 net1004 VPWR VGND sg13g2_buf_1
Xfanout1037 DP_1.matrix\[2\] net1037 VPWR VGND sg13g2_buf_8
Xfanout1015 net313 net1015 VPWR VGND sg13g2_buf_2
Xfanout1026 DP_1.matrix\[7\] net1026 VPWR VGND sg13g2_buf_8
XFILLER_0_987 VPWR VGND sg13g2_decap_8
Xfanout1059 DP_1.matrix\[8\] net1059 VPWR VGND sg13g2_buf_1
Xfanout1048 DP_3.matrix\[44\] net1048 VPWR VGND sg13g2_buf_1
XFILLER_16_811 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_54_clk clknet_4_8_0_clk clknet_leaf_54_clk VPWR VGND sg13g2_buf_8
XFILLER_15_332 VPWR VGND sg13g2_fill_2
XFILLER_37_1016 VPWR VGND sg13g2_decap_8
XFILLER_31_825 VPWR VGND sg13g2_fill_1
XFILLER_37_1027 VPWR VGND sg13g2_fill_2
Xhold509 _2235_ VPWR VGND net549 sg13g2_dlygate4sd3_1
X_3360_ _2943_ _2934_ _2945_ VPWR VGND sg13g2_xor2_1
X_5030_ _1778_ _1777_ _1774_ VPWR VGND sg13g2_nand2b_1
X_3291_ _2878_ net991 net931 VPWR VGND sg13g2_nand2_1
XFILLER_19_660 VPWR VGND sg13g2_fill_2
XFILLER_20_1020 VPWR VGND sg13g2_decap_8
XFILLER_47_980 VPWR VGND sg13g2_decap_8
X_5932_ _2582_ _2412_ _2424_ VPWR VGND sg13g2_xnor2_1
XFILLER_18_181 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_45_clk clknet_4_14_0_clk clknet_leaf_45_clk VPWR VGND sg13g2_buf_8
X_5863_ net892 net807 _2518_ VPWR VGND sg13g2_nor2_1
X_4814_ _1573_ _1566_ _1574_ VPWR VGND sg13g2_xor2_1
X_5794_ net982 net809 _2450_ VPWR VGND sg13g2_nor2_1
X_4745_ _1501_ _1505_ _1506_ VPWR VGND sg13g2_nor2_1
XFILLER_21_379 VPWR VGND sg13g2_fill_1
XFILLER_30_880 VPWR VGND sg13g2_fill_1
X_4676_ _1439_ _1434_ _1437_ VPWR VGND sg13g2_xnor2_1
X_3627_ _0389_ _0392_ _0435_ VPWR VGND sg13g2_nor2_1
X_6415_ net1077 VGND VPWR net118 mac2.sum_lvl3_ff\[31\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_1_707 VPWR VGND sg13g2_fill_2
X_6346_ net1116 VGND VPWR net201 mac1.sum_lvl1_ff\[78\] clknet_leaf_52_clk sg13g2_dfrbpq_1
X_3558_ _0368_ _0361_ _0366_ _0367_ VPWR VGND sg13g2_and3_1
Xoutput29 net29 uo_out[4] VPWR VGND sg13g2_buf_1
Xoutput18 net18 uio_out[1] VPWR VGND sg13g2_buf_1
X_3489_ _0301_ _0294_ _0299_ _0300_ VPWR VGND sg13g2_and3_1
X_6277_ net1063 VGND VPWR net59 mac1.sum_lvl2_ff\[1\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_5228_ VGND VPWR net827 net871 _1971_ _1940_ sg13g2_a21oi_1
XFILLER_5_1003 VPWR VGND sg13g2_decap_8
X_5159_ VGND VPWR _1900_ _1901_ _1904_ _1883_ sg13g2_a21oi_1
XFILLER_44_416 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_36_clk clknet_4_13_0_clk clknet_leaf_36_clk VPWR VGND sg13g2_buf_8
XFILLER_12_302 VPWR VGND sg13g2_fill_1
XFILLER_24_173 VPWR VGND sg13g2_fill_1
XFILLER_0_784 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_27_clk clknet_4_7_0_clk clknet_leaf_27_clk VPWR VGND sg13g2_buf_8
XFILLER_11_1008 VPWR VGND sg13g2_decap_8
X_4530_ VGND VPWR _1251_ _1270_ _1303_ _1272_ sg13g2_a21oi_1
Xhold317 DP_4.matrix\[6\] VPWR VGND net357 sg13g2_dlygate4sd3_1
Xhold306 mac2.sum_lvl3_ff\[10\] VPWR VGND net346 sg13g2_dlygate4sd3_1
X_4461_ _1236_ _1228_ _1235_ VPWR VGND sg13g2_xnor2_1
Xhold339 DP_4.matrix\[2\] VPWR VGND net379 sg13g2_dlygate4sd3_1
X_6200_ net1114 VGND VPWR _0217_ DP_2.matrix\[77\] clknet_leaf_58_clk sg13g2_dfrbpq_1
X_3412_ _2994_ _2984_ _2995_ VPWR VGND sg13g2_nor2b_1
Xhold328 _0002_ VPWR VGND net368 sg13g2_dlygate4sd3_1
X_6131_ net1124 VGND VPWR _0171_ DP_4.matrix\[80\] clknet_leaf_36_clk sg13g2_dfrbpq_2
X_4392_ _1121_ VPWR _1169_ VGND _1060_ _1122_ sg13g2_o21ai_1
Xfanout819 DP_4.matrix\[76\] net819 VPWR VGND sg13g2_buf_1
Xfanout808 _2397_ net808 VPWR VGND sg13g2_buf_8
X_3343_ _0096_ _2927_ _2928_ VPWR VGND sg13g2_xnor2_1
X_6062_ net885 _0238_ VPWR VGND sg13g2_buf_1
X_3274_ _2860_ _2861_ _2862_ VPWR VGND sg13g2_nor2b_1
X_5013_ _1758_ _1759_ _1761_ _1762_ VPWR VGND sg13g2_or3_1
XFILLER_26_438 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_18_clk clknet_4_5_0_clk clknet_leaf_18_clk VPWR VGND sg13g2_buf_8
X_5915_ net1044 net803 _2569_ VPWR VGND sg13g2_nor2_1
X_5846_ net902 net806 _2501_ VPWR VGND sg13g2_nor2_1
XFILLER_22_677 VPWR VGND sg13g2_fill_1
X_5777_ net1026 DP_1.matrix\[43\] net810 _2434_ VPWR VGND sg13g2_mux2_1
X_4728_ _1466_ _1487_ _1489_ _1490_ VPWR VGND sg13g2_or3_1
X_4659_ _1421_ _1420_ _1382_ _1423_ VPWR VGND sg13g2_a21o_1
X_6329_ net1082 VGND VPWR net112 mac2.sum_lvl2_ff\[43\] clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_18_917 VPWR VGND sg13g2_decap_8
XFILLER_26_950 VPWR VGND sg13g2_decap_8
XFILLER_41_986 VPWR VGND sg13g2_decap_8
XFILLER_5_821 VPWR VGND sg13g2_decap_8
XFILLER_5_898 VPWR VGND sg13g2_decap_8
XFILLER_35_202 VPWR VGND sg13g2_fill_1
X_3961_ _0717_ _0716_ _0715_ _0755_ VPWR VGND sg13g2_a21o_2
X_5700_ _2364_ _2361_ _2363_ VPWR VGND sg13g2_nand2_1
X_3892_ _0664_ VPWR _0687_ VGND _0639_ _0662_ sg13g2_o21ai_1
X_5631_ _2310_ _2309_ _2308_ VPWR VGND sg13g2_nand2b_1
X_5562_ mac2.sum_lvl2_ff\[31\] mac2.sum_lvl2_ff\[12\] _2256_ VPWR VGND sg13g2_nor2_1
X_4513_ _1286_ net899 net1043 VPWR VGND sg13g2_nand2_1
Xhold103 mac1.sum_lvl2_ff\[53\] VPWR VGND net143 sg13g2_dlygate4sd3_1
X_5493_ VGND VPWR _2202_ _2203_ _2190_ _2188_ sg13g2_a21oi_2
Xhold114 mac2.products_ff\[70\] VPWR VGND net154 sg13g2_dlygate4sd3_1
Xhold125 mac2.sum_lvl1_ff\[75\] VPWR VGND net165 sg13g2_dlygate4sd3_1
Xhold136 mac1.products_ff\[144\] VPWR VGND net176 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_4_3_0_clk clknet_leaf_7_clk VPWR VGND sg13g2_buf_8
Xhold147 mac1.sum_lvl2_ff\[48\] VPWR VGND net187 sg13g2_dlygate4sd3_1
X_4444_ _1219_ net899 net834 VPWR VGND sg13g2_nand2_1
Xhold158 mac2.sum_lvl1_ff\[4\] VPWR VGND net198 sg13g2_dlygate4sd3_1
Xhold169 mac1.sum_lvl2_ff\[45\] VPWR VGND net209 sg13g2_dlygate4sd3_1
X_4375_ _1148_ _1149_ _1151_ _1152_ VPWR VGND sg13g2_or3_1
X_3326_ _2912_ net996 net1051 VPWR VGND sg13g2_nand2_1
X_6114_ net1089 VGND VPWR _0117_ mac1.products_ff\[78\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_6045_ net940 _0213_ VPWR VGND sg13g2_buf_1
X_3257_ _2799_ VPWR _2845_ VGND _2797_ _2800_ sg13g2_o21ai_1
X_3188_ _2766_ VPWR _2777_ VGND _2744_ _2767_ sg13g2_o21ai_1
XFILLER_42_717 VPWR VGND sg13g2_fill_1
X_5829_ net794 _2482_ _2483_ _2484_ VPWR VGND sg13g2_nor3_1
XFILLER_23_986 VPWR VGND sg13g2_decap_8
XFILLER_2_868 VPWR VGND sg13g2_decap_8
XFILLER_40_1001 VPWR VGND sg13g2_decap_8
XFILLER_45_500 VPWR VGND sg13g2_fill_1
XFILLER_17_213 VPWR VGND sg13g2_fill_1
XFILLER_45_566 VPWR VGND sg13g2_fill_2
XFILLER_13_474 VPWR VGND sg13g2_decap_8
XFILLER_14_986 VPWR VGND sg13g2_decap_8
XFILLER_9_467 VPWR VGND sg13g2_fill_2
X_4160_ _0948_ _0939_ _0947_ VPWR VGND sg13g2_xnor2_1
X_3111_ _2700_ _2701_ _2676_ _2703_ VPWR VGND sg13g2_nand3_1
XFILLER_49_850 VPWR VGND sg13g2_fill_1
X_4091_ _0864_ _0857_ _0827_ _0881_ VPWR VGND sg13g2_a21o_1
X_3042_ _2636_ net516 _0065_ VPWR VGND sg13g2_nor2_2
XFILLER_24_706 VPWR VGND sg13g2_fill_2
X_4993_ net825 net883 net830 _1743_ VPWR VGND net880 sg13g2_nand4_1
X_3944_ _0734_ _0735_ _0737_ _0738_ VPWR VGND sg13g2_or3_1
XFILLER_20_901 VPWR VGND sg13g2_decap_8
X_3875_ _0667_ _0668_ _0670_ _0671_ VPWR VGND sg13g2_or3_1
X_5614_ mac2.sum_lvl3_ff\[28\] mac2.sum_lvl3_ff\[8\] _2296_ VPWR VGND sg13g2_and2_1
XFILLER_20_978 VPWR VGND sg13g2_decap_8
X_5545_ net519 _2242_ _0046_ VPWR VGND sg13g2_nor2b_2
X_5476_ net509 mac1.sum_lvl3_ff\[29\] _2189_ VPWR VGND sg13g2_xor2_1
X_4427_ _1202_ _1195_ _1203_ VPWR VGND sg13g2_xor2_1
X_4358_ _1130_ _1134_ _1135_ VPWR VGND sg13g2_nor2_1
X_3309_ VGND VPWR _2819_ _2861_ _2896_ _2860_ sg13g2_a21oi_1
X_4289_ _1068_ _1063_ _1066_ VPWR VGND sg13g2_xnor2_1
X_6028_ net1004 _0188_ VPWR VGND sg13g2_buf_1
XFILLER_14_216 VPWR VGND sg13g2_fill_1
XFILLER_23_750 VPWR VGND sg13g2_fill_2
XFILLER_10_444 VPWR VGND sg13g2_fill_1
XFILLER_10_433 VPWR VGND sg13g2_fill_1
XFILLER_7_905 VPWR VGND sg13g2_decap_8
XFILLER_11_945 VPWR VGND sg13g2_decap_8
Xfanout991 net993 net991 VPWR VGND sg13g2_buf_8
Xfanout980 net981 net980 VPWR VGND sg13g2_buf_1
XFILLER_46_853 VPWR VGND sg13g2_decap_8
XFILLER_46_897 VPWR VGND sg13g2_decap_8
XFILLER_33_569 VPWR VGND sg13g2_fill_2
XFILLER_9_231 VPWR VGND sg13g2_fill_2
X_3660_ _0432_ _0467_ _0468_ VPWR VGND sg13g2_nor2_1
Xclkload12 clknet_leaf_67_clk clkload12/Y VPWR VGND sg13g2_inv_4
X_3591_ _0400_ net975 net1031 VPWR VGND sg13g2_nand2_1
X_5330_ _2043_ _2045_ _2068_ _2070_ VPWR VGND sg13g2_or3_1
X_5261_ _2003_ _1995_ _2000_ VPWR VGND sg13g2_xnor2_1
XFILLER_6_993 VPWR VGND sg13g2_decap_8
X_4212_ _0995_ _0987_ _0994_ VPWR VGND sg13g2_nand2_1
X_5192_ _1885_ _1934_ _1936_ VPWR VGND sg13g2_and2_1
X_4143_ VGND VPWR _0880_ _0899_ _0932_ _0901_ sg13g2_a21oi_1
X_4074_ _0865_ _0857_ _0864_ VPWR VGND sg13g2_xnor2_1
XFILLER_12_709 VPWR VGND sg13g2_fill_1
XFILLER_34_29 VPWR VGND sg13g2_fill_1
X_4976_ _0144_ _1722_ _1729_ VPWR VGND sg13g2_xnor2_1
X_3927_ net1022 net950 net1024 _0721_ VPWR VGND net948 sg13g2_nand4_1
X_3858_ _0634_ VPWR _0655_ VGND _0625_ _0635_ sg13g2_o21ai_1
Xclkload6 clknet_4_9_0_clk clkload6/X VPWR VGND sg13g2_buf_8
XFILLER_4_908 VPWR VGND sg13g2_decap_8
X_3789_ _0576_ _0568_ _0575_ _0592_ VPWR VGND sg13g2_a21o_1
X_6577_ net1066 VGND VPWR net317 mac2.total_sum\[9\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_5528_ net548 net469 _2229_ VPWR VGND sg13g2_nor2_1
X_5459_ _2175_ mac1.sum_lvl3_ff\[26\] net532 VPWR VGND sg13g2_xnor2_1
XFILLER_28_842 VPWR VGND sg13g2_fill_2
XFILLER_43_823 VPWR VGND sg13g2_fill_1
XFILLER_42_311 VPWR VGND sg13g2_fill_1
XFILLER_43_889 VPWR VGND sg13g2_decap_4
XFILLER_11_742 VPWR VGND sg13g2_fill_1
XFILLER_10_263 VPWR VGND sg13g2_fill_2
XFILLER_10_296 VPWR VGND sg13g2_fill_2
XFILLER_6_256 VPWR VGND sg13g2_fill_2
XFILLER_3_930 VPWR VGND sg13g2_decap_8
X_4830_ _1589_ net921 net1044 VPWR VGND sg13g2_nand2_1
X_4761_ _1522_ net1049 net867 net909 net864 VPWR VGND sg13g2_a22oi_1
XFILLER_14_1028 VPWR VGND sg13g2_fill_1
X_3712_ _0478_ VPWR _0518_ VGND _0475_ _0479_ sg13g2_o21ai_1
X_6500_ net1103 VGND VPWR net49 mac2.sum_lvl1_ff\[36\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_4692_ _1455_ _1452_ _1454_ VPWR VGND sg13g2_nand2_1
X_3643_ _0451_ _0399_ _0448_ VPWR VGND sg13g2_xnor2_1
X_6431_ net1065 VGND VPWR net526 mac1.total_sum\[11\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_6362_ net1079 VGND VPWR net60 mac2.sum_lvl1_ff\[78\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_5313_ _2036_ _2029_ _2038_ _2053_ VPWR VGND sg13g2_a21o_1
X_3574_ _0384_ _0382_ _0383_ VPWR VGND sg13g2_nand2_1
X_6293_ net1063 VGND VPWR net78 mac1.sum_lvl2_ff\[20\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_5244_ VGND VPWR _1950_ _1952_ _1987_ _1986_ sg13g2_a21oi_1
X_5175_ _1880_ VPWR _1919_ VGND _1835_ _1881_ sg13g2_o21ai_1
Xhold29 mac2.sum_lvl1_ff\[83\] VPWR VGND net69 sg13g2_dlygate4sd3_1
Xhold18 mac1.sum_lvl1_ff\[14\] VPWR VGND net58 sg13g2_dlygate4sd3_1
X_4126_ _0915_ net1013 net1052 VPWR VGND sg13g2_nand2_1
XFILLER_44_609 VPWR VGND sg13g2_fill_1
X_4057_ _0848_ net1013 net947 VPWR VGND sg13g2_nand2_1
XFILLER_24_300 VPWR VGND sg13g2_fill_2
XFILLER_25_823 VPWR VGND sg13g2_fill_2
XFILLER_37_672 VPWR VGND sg13g2_fill_1
XFILLER_24_388 VPWR VGND sg13g2_fill_1
X_4959_ _1714_ _1707_ _1713_ VPWR VGND sg13g2_nand2_1
XFILLER_3_204 VPWR VGND sg13g2_fill_2
Xfanout1038 net1039 net1038 VPWR VGND sg13g2_buf_8
Xfanout1016 net1017 net1016 VPWR VGND sg13g2_buf_8
XFILLER_0_966 VPWR VGND sg13g2_decap_8
Xfanout1005 net1006 net1005 VPWR VGND sg13g2_buf_2
Xfanout1027 net1029 net1027 VPWR VGND sg13g2_buf_8
Xfanout1049 net1050 net1049 VPWR VGND sg13g2_buf_8
XFILLER_47_425 VPWR VGND sg13g2_fill_1
XFILLER_16_889 VPWR VGND sg13g2_decap_8
XFILLER_30_303 VPWR VGND sg13g2_fill_2
XFILLER_11_561 VPWR VGND sg13g2_fill_1
X_3290_ VGND VPWR net938 net986 _2877_ _2846_ sg13g2_a21oi_1
XFILLER_2_270 VPWR VGND sg13g2_fill_2
XFILLER_38_403 VPWR VGND sg13g2_fill_1
XFILLER_39_926 VPWR VGND sg13g2_fill_2
X_5931_ net1034 net784 _2581_ VPWR VGND sg13g2_nor2_1
XFILLER_19_694 VPWR VGND sg13g2_decap_8
XFILLER_34_642 VPWR VGND sg13g2_fill_2
X_5862_ net910 net803 _2517_ VPWR VGND sg13g2_nor2_1
XFILLER_33_152 VPWR VGND sg13g2_fill_1
X_4813_ _1573_ _1567_ _1571_ VPWR VGND sg13g2_xnor2_1
X_5793_ _2449_ net946 net801 VPWR VGND sg13g2_nand2_1
X_4744_ VGND VPWR _1505_ _1504_ _1503_ sg13g2_or2_1
X_4675_ _1438_ _1437_ _1434_ VPWR VGND sg13g2_nand2b_1
X_3626_ _0417_ VPWR _0434_ VGND _0396_ _0418_ sg13g2_o21ai_1
X_6414_ net1067 VGND VPWR net101 mac2.sum_lvl3_ff\[30\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_6345_ net1131 VGND VPWR net135 mac1.sum_lvl1_ff\[77\] clknet_leaf_52_clk sg13g2_dfrbpq_1
X_3557_ _0362_ VPWR _0367_ VGND _0363_ _0365_ sg13g2_o21ai_1
Xoutput19 net19 uio_out[2] VPWR VGND sg13g2_buf_1
X_6276_ net1064 VGND VPWR net142 mac1.sum_lvl2_ff\[0\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_5227_ _1944_ VPWR _1970_ VGND _1938_ _1945_ sg13g2_o21ai_1
X_3488_ _0295_ VPWR _0300_ VGND _0296_ _0298_ sg13g2_o21ai_1
X_5158_ _1900_ _1901_ _1883_ _1903_ VPWR VGND sg13g2_nand3_1
XFILLER_45_929 VPWR VGND sg13g2_decap_8
X_5089_ net886 net814 net889 _1835_ VPWR VGND net811 sg13g2_nand4_1
X_4109_ _0897_ _0887_ _0899_ VPWR VGND sg13g2_xor2_1
XFILLER_38_981 VPWR VGND sg13g2_decap_8
XFILLER_21_30 VPWR VGND sg13g2_fill_1
XFILLER_43_1021 VPWR VGND sg13g2_decap_8
XFILLER_0_763 VPWR VGND sg13g2_decap_8
XFILLER_47_277 VPWR VGND sg13g2_fill_1
XFILLER_16_686 VPWR VGND sg13g2_fill_2
XFILLER_15_196 VPWR VGND sg13g2_fill_1
XFILLER_30_100 VPWR VGND sg13g2_fill_1
XFILLER_31_678 VPWR VGND sg13g2_fill_2
XFILLER_12_892 VPWR VGND sg13g2_decap_8
XFILLER_31_689 VPWR VGND sg13g2_fill_2
XFILLER_8_885 VPWR VGND sg13g2_decap_8
Xhold307 _2306_ VPWR VGND net347 sg13g2_dlygate4sd3_1
X_4460_ _1233_ _1234_ _1235_ VPWR VGND sg13g2_nor2b_1
Xhold318 _0250_ VPWR VGND net358 sg13g2_dlygate4sd3_1
Xhold329 DP_1.matrix\[42\] VPWR VGND net369 sg13g2_dlygate4sd3_1
X_3411_ _2994_ _2970_ _2993_ VPWR VGND sg13g2_xnor2_1
X_4391_ _1094_ VPWR _1168_ VGND _1164_ _1166_ sg13g2_o21ai_1
X_3342_ _2893_ _2898_ _2928_ VPWR VGND sg13g2_nor2_1
X_6130_ net1129 VGND VPWR _0170_ DP_4.matrix\[44\] clknet_leaf_45_clk sg13g2_dfrbpq_2
Xfanout809 net810 net809 VPWR VGND sg13g2_buf_8
X_6061_ net888 _0237_ VPWR VGND sg13g2_buf_1
X_3273_ _2861_ _2824_ _2859_ VPWR VGND sg13g2_nand2_1
X_5012_ _1761_ net877 net828 net881 net825 VPWR VGND sg13g2_a22oi_1
XFILLER_38_211 VPWR VGND sg13g2_fill_1
X_5914_ VPWR _2568_ _2567_ VGND sg13g2_inv_1
X_5845_ net920 net805 _2500_ VPWR VGND sg13g2_nor2_1
XFILLER_22_645 VPWR VGND sg13g2_decap_8
X_5776_ VPWR _2433_ _2432_ VGND sg13g2_inv_1
XFILLER_21_177 VPWR VGND sg13g2_decap_8
X_4727_ VGND VPWR _1485_ _1486_ _1489_ _1467_ sg13g2_a21oi_1
X_4658_ _1420_ _1421_ _1382_ _1422_ VPWR VGND sg13g2_nand3_1
X_3609_ VGND VPWR _0414_ _0415_ _0418_ _0397_ sg13g2_a21oi_1
X_4589_ net924 net869 _0084_ VPWR VGND sg13g2_and2_1
X_6328_ net1084 VGND VPWR net171 mac2.sum_lvl2_ff\[42\] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_6259_ net1125 VGND VPWR _0267_ DP_4.matrix\[79\] clknet_leaf_35_clk sg13g2_dfrbpq_1
XFILLER_29_200 VPWR VGND sg13g2_fill_1
XFILLER_45_737 VPWR VGND sg13g2_fill_1
XFILLER_17_439 VPWR VGND sg13g2_fill_2
XFILLER_44_269 VPWR VGND sg13g2_fill_1
XFILLER_40_442 VPWR VGND sg13g2_fill_2
XFILLER_8_115 VPWR VGND sg13g2_fill_2
XFILLER_12_166 VPWR VGND sg13g2_decap_8
XFILLER_5_877 VPWR VGND sg13g2_decap_8
XFILLER_36_715 VPWR VGND sg13g2_fill_1
X_3960_ _0753_ _0689_ _0754_ VPWR VGND sg13g2_xor2_1
XFILLER_17_995 VPWR VGND sg13g2_decap_8
X_3891_ _0686_ _0678_ _0680_ VPWR VGND sg13g2_nand2_1
X_5630_ _2309_ mac2.sum_lvl3_ff\[31\] mac2.sum_lvl3_ff\[11\] VPWR VGND sg13g2_nand2_1
XFILLER_32_998 VPWR VGND sg13g2_decap_8
X_5561_ _2255_ mac2.sum_lvl2_ff\[31\] mac2.sum_lvl2_ff\[12\] VPWR VGND sg13g2_nand2_1
XFILLER_8_660 VPWR VGND sg13g2_fill_2
X_5492_ _2196_ _2193_ _2202_ VPWR VGND _2195_ sg13g2_nand3b_1
X_4512_ _1255_ VPWR _1285_ VGND _1253_ _1256_ sg13g2_o21ai_1
Xhold115 mac1.products_ff\[146\] VPWR VGND net155 sg13g2_dlygate4sd3_1
Xhold126 mac1.sum_lvl1_ff\[85\] VPWR VGND net166 sg13g2_dlygate4sd3_1
Xhold104 mac2.products_ff\[139\] VPWR VGND net144 sg13g2_dlygate4sd3_1
Xhold159 mac2.products_ff\[76\] VPWR VGND net199 sg13g2_dlygate4sd3_1
Xhold137 mac1.products_ff\[82\] VPWR VGND net177 sg13g2_dlygate4sd3_1
Xhold148 mac1.sum_lvl1_ff\[50\] VPWR VGND net188 sg13g2_dlygate4sd3_1
X_4443_ _1218_ net903 net1043 VPWR VGND sg13g2_nand2_1
X_4374_ _1151_ net1047 net848 net891 net845 VPWR VGND sg13g2_a22oi_1
X_6113_ net1092 VGND VPWR _0126_ mac1.products_ff\[77\] clknet_leaf_56_clk sg13g2_dfrbpq_1
X_3325_ VGND VPWR _2911_ _2882_ _2880_ sg13g2_or2_1
X_6044_ net943 _0212_ VPWR VGND sg13g2_buf_1
X_3256_ _2844_ _2839_ _2843_ VPWR VGND sg13g2_xnor2_1
XFILLER_39_520 VPWR VGND sg13g2_fill_1
XFILLER_39_542 VPWR VGND sg13g2_fill_1
X_3187_ _2775_ _2774_ _0102_ VPWR VGND sg13g2_xor2_1
XFILLER_27_726 VPWR VGND sg13g2_decap_4
XFILLER_39_575 VPWR VGND sg13g2_fill_1
XFILLER_35_781 VPWR VGND sg13g2_fill_2
XFILLER_23_965 VPWR VGND sg13g2_decap_8
X_5828_ net915 net804 _2483_ VPWR VGND sg13g2_nor2_1
X_5759_ _2413_ VPWR _2416_ VGND _2414_ _2415_ sg13g2_o21ai_1
XFILLER_2_847 VPWR VGND sg13g2_decap_8
XFILLER_17_269 VPWR VGND sg13g2_fill_2
XFILLER_14_965 VPWR VGND sg13g2_decap_8
XFILLER_43_50 VPWR VGND sg13g2_fill_1
XFILLER_13_464 VPWR VGND sg13g2_decap_4
XFILLER_4_173 VPWR VGND sg13g2_fill_1
XFILLER_4_195 VPWR VGND sg13g2_fill_2
X_3110_ _2700_ _2701_ _2702_ VPWR VGND sg13g2_and2_1
X_4090_ _0866_ VPWR _0880_ VGND _0855_ _0867_ sg13g2_o21ai_1
X_3041_ _2637_ net942 net1003 net1002 net946 VPWR VGND sg13g2_a22oi_1
X_4992_ net828 net825 net883 net880 _1742_ VPWR VGND sg13g2_and4_1
X_3943_ _0737_ net1005 net963 net1009 net960 VPWR VGND sg13g2_a22oi_1
XFILLER_23_239 VPWR VGND sg13g2_fill_2
XFILLER_32_740 VPWR VGND sg13g2_fill_2
X_3874_ _0670_ net1011 net962 net1014 net958 VPWR VGND sg13g2_a22oi_1
XFILLER_20_957 VPWR VGND sg13g2_decap_8
X_5613_ _2294_ _2295_ _0061_ VPWR VGND sg13g2_and2_1
XFILLER_9_980 VPWR VGND sg13g2_decap_8
X_5544_ _2238_ _2240_ _2236_ _2242_ VPWR VGND sg13g2_nand3_1
X_5475_ _2188_ mac1.sum_lvl3_ff\[29\] net509 VPWR VGND sg13g2_nand2_1
X_4426_ _1202_ _1196_ _1200_ VPWR VGND sg13g2_xnor2_1
X_4357_ VGND VPWR _1134_ _1133_ _1132_ sg13g2_or2_1
X_3308_ _2895_ _2894_ _2893_ VPWR VGND sg13g2_nand2b_1
X_4288_ _1067_ _1066_ _1063_ VPWR VGND sg13g2_nand2b_1
X_6027_ net1007 _0187_ VPWR VGND sg13g2_buf_1
X_3239_ _2781_ _2784_ _2827_ VPWR VGND sg13g2_nor2_2
XFILLER_27_556 VPWR VGND sg13g2_fill_1
XFILLER_11_924 VPWR VGND sg13g2_decap_8
XFILLER_23_784 VPWR VGND sg13g2_decap_8
XFILLER_10_423 VPWR VGND sg13g2_fill_1
XFILLER_13_42 VPWR VGND sg13g2_fill_1
Xhold490 mac2.sum_lvl3_ff\[12\] VPWR VGND net530 sg13g2_dlygate4sd3_1
Xfanout970 DP_2.matrix\[6\] net970 VPWR VGND sg13g2_buf_1
Xfanout981 DP_2.matrix\[1\] net981 VPWR VGND sg13g2_buf_1
Xfanout992 net993 net992 VPWR VGND sg13g2_buf_1
XFILLER_33_515 VPWR VGND sg13g2_fill_1
XFILLER_14_751 VPWR VGND sg13g2_fill_1
XFILLER_14_784 VPWR VGND sg13g2_fill_1
Xclkload13 clknet_leaf_65_clk clkload13/X VPWR VGND sg13g2_buf_8
X_3590_ _0399_ net973 net1030 VPWR VGND sg13g2_nand2_2
XFILLER_6_972 VPWR VGND sg13g2_decap_8
XFILLER_47_1008 VPWR VGND sg13g2_decap_8
X_5260_ VGND VPWR _2002_ _2000_ _1995_ sg13g2_or2_1
XFILLER_5_493 VPWR VGND sg13g2_fill_2
X_4211_ _0992_ _0993_ _0994_ VPWR VGND sg13g2_nor2b_1
X_5191_ VGND VPWR _1935_ _1934_ _1885_ sg13g2_or2_1
X_4142_ _0929_ _0908_ _0931_ VPWR VGND sg13g2_xor2_1
X_4073_ _0862_ _0863_ _0864_ VPWR VGND sg13g2_nor2b_1
XFILLER_49_692 VPWR VGND sg13g2_fill_1
XFILLER_37_854 VPWR VGND sg13g2_fill_2
XFILLER_24_537 VPWR VGND sg13g2_fill_1
X_4975_ _1729_ _1723_ _1728_ VPWR VGND sg13g2_xnor2_1
X_3926_ _0720_ net948 net1024 net950 net1022 VPWR VGND sg13g2_a22oi_1
XFILLER_32_581 VPWR VGND sg13g2_fill_1
X_3857_ _0654_ _0642_ _0653_ VPWR VGND sg13g2_xnor2_1
Xclkload7 clknet_4_10_0_clk clkload7/X VPWR VGND sg13g2_buf_8
X_6576_ net1065 VGND VPWR net457 mac2.total_sum\[8\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_3788_ VGND VPWR _0567_ _0581_ _0591_ _0580_ sg13g2_a21oi_1
X_5527_ VGND VPWR _2225_ _2227_ _2228_ _2226_ sg13g2_a21oi_1
X_5458_ mac1.sum_lvl3_ff\[26\] mac1.sum_lvl3_ff\[6\] _2174_ VPWR VGND sg13g2_and2_1
X_5389_ _2116_ net462 _2120_ _2121_ VPWR VGND sg13g2_nor3_1
X_4409_ _1185_ _1180_ _1183_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_810 VPWR VGND sg13g2_decap_4
XFILLER_28_821 VPWR VGND sg13g2_decap_4
XFILLER_43_846 VPWR VGND sg13g2_fill_1
XFILLER_27_397 VPWR VGND sg13g2_fill_2
XFILLER_7_725 VPWR VGND sg13g2_fill_1
XFILLER_6_213 VPWR VGND sg13g2_decap_8
XFILLER_11_798 VPWR VGND sg13g2_fill_1
XFILLER_3_986 VPWR VGND sg13g2_decap_8
XFILLER_18_331 VPWR VGND sg13g2_fill_1
X_4760_ net864 net909 net867 _1521_ VPWR VGND net1049 sg13g2_nand4_1
XFILLER_14_1007 VPWR VGND sg13g2_decap_8
X_3711_ _0517_ _0509_ _0514_ VPWR VGND sg13g2_xnor2_1
X_4691_ _1451_ _1450_ _1433_ _1454_ VPWR VGND sg13g2_a21o_1
X_3642_ _0399_ _0448_ _0450_ VPWR VGND sg13g2_and2_1
X_6430_ net1065 VGND VPWR _0017_ mac1.total_sum\[10\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_6361_ net1081 VGND VPWR net128 mac2.sum_lvl1_ff\[77\] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_3573_ _0345_ _0344_ _0343_ _0383_ VPWR VGND sg13g2_a21o_2
X_5312_ _2052_ _2049_ _0152_ VPWR VGND sg13g2_xor2_1
X_6292_ net1064 VGND VPWR net212 mac1.sum_lvl2_ff\[19\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_5243_ _1984_ _1957_ _1986_ VPWR VGND sg13g2_xor2_1
X_5174_ _1908_ VPWR _1918_ VGND _1837_ _1909_ sg13g2_o21ai_1
Xhold19 mac1.sum_lvl1_ff\[1\] VPWR VGND net59 sg13g2_dlygate4sd3_1
X_4125_ _0884_ VPWR _0914_ VGND _0882_ _0885_ sg13g2_o21ai_1
X_4056_ _0847_ net1018 net1052 VPWR VGND sg13g2_nand2_1
XFILLER_24_367 VPWR VGND sg13g2_fill_2
X_4958_ _1713_ _1708_ _1711_ VPWR VGND sg13g2_xnor2_1
X_4889_ VGND VPWR _1611_ _1613_ _1647_ _1645_ sg13g2_a21oi_1
X_3909_ _0699_ VPWR _0704_ VGND _0700_ _0702_ sg13g2_o21ai_1
X_6559_ net1082 VGND VPWR _0045_ mac2.sum_lvl3_ff\[7\] clknet_leaf_19_clk sg13g2_dfrbpq_1
Xfanout1017 net312 net1017 VPWR VGND sg13g2_buf_8
XFILLER_0_945 VPWR VGND sg13g2_decap_8
Xfanout1006 net1007 net1006 VPWR VGND sg13g2_buf_1
Xfanout1028 net1029 net1028 VPWR VGND sg13g2_buf_1
XFILLER_48_905 VPWR VGND sg13g2_decap_8
Xfanout1039 net504 net1039 VPWR VGND sg13g2_buf_8
XFILLER_48_949 VPWR VGND sg13g2_decap_8
XFILLER_19_106 VPWR VGND sg13g2_decap_8
XFILLER_28_651 VPWR VGND sg13g2_decap_8
XFILLER_28_662 VPWR VGND sg13g2_fill_2
XFILLER_15_334 VPWR VGND sg13g2_fill_1
XFILLER_16_846 VPWR VGND sg13g2_decap_4
XFILLER_16_868 VPWR VGND sg13g2_decap_8
XFILLER_28_695 VPWR VGND sg13g2_decap_4
XFILLER_7_555 VPWR VGND sg13g2_fill_1
XFILLER_18_4 VPWR VGND sg13g2_fill_2
X_5930_ VGND VPWR net785 _2580_ _0174_ _2579_ sg13g2_a21oi_1
XFILLER_19_662 VPWR VGND sg13g2_fill_1
XFILLER_18_194 VPWR VGND sg13g2_decap_4
X_5861_ _2511_ _2515_ _2516_ VPWR VGND sg13g2_nor2b_1
X_4812_ _1572_ _1567_ _1571_ VPWR VGND sg13g2_nand2_1
X_5792_ _2447_ VPWR _2448_ VGND _2402_ _2446_ sg13g2_o21ai_1
XFILLER_15_890 VPWR VGND sg13g2_decap_8
XFILLER_33_197 VPWR VGND sg13g2_fill_2
X_4743_ _1504_ net851 net922 net854 net921 VPWR VGND sg13g2_a22oi_1
X_6413_ net1078 VGND VPWR net162 mac2.sum_lvl3_ff\[29\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_4674_ _1436_ _1403_ _1437_ VPWR VGND sg13g2_xor2_1
X_3625_ _0394_ VPWR _0433_ VGND _0349_ _0395_ sg13g2_o21ai_1
X_6344_ net1116 VGND VPWR net207 mac1.sum_lvl1_ff\[76\] clknet_leaf_53_clk sg13g2_dfrbpq_1
X_3556_ _0362_ _0363_ _0365_ _0366_ VPWR VGND sg13g2_or3_1
X_6275_ net1096 VGND VPWR net98 mac1.sum_lvl1_ff\[51\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_5226_ _1967_ _1959_ _1969_ VPWR VGND sg13g2_xor2_1
X_3487_ _0295_ _0296_ _0298_ _0299_ VPWR VGND sg13g2_or3_1
X_5157_ _1902_ _1883_ _1900_ _1901_ VPWR VGND sg13g2_and3_1
X_5088_ _1834_ net811 net889 net814 net886 VPWR VGND sg13g2_a22oi_1
X_4108_ _0887_ _0897_ _0898_ VPWR VGND sg13g2_nor2_1
X_4039_ _0831_ _0825_ _0829_ VPWR VGND sg13g2_xnor2_1
XFILLER_25_654 VPWR VGND sg13g2_decap_8
XFILLER_13_827 VPWR VGND sg13g2_fill_2
XFILLER_25_698 VPWR VGND sg13g2_fill_1
XFILLER_21_871 VPWR VGND sg13g2_fill_2
XFILLER_43_1000 VPWR VGND sg13g2_decap_8
XFILLER_29_982 VPWR VGND sg13g2_decap_8
XFILLER_28_470 VPWR VGND sg13g2_fill_1
XFILLER_44_985 VPWR VGND sg13g2_decap_8
XFILLER_31_657 VPWR VGND sg13g2_fill_2
XFILLER_12_871 VPWR VGND sg13g2_decap_8
XFILLER_8_864 VPWR VGND sg13g2_decap_8
Xhold308 _0049_ VPWR VGND net348 sg13g2_dlygate4sd3_1
X_3410_ _2991_ _2985_ _2993_ VPWR VGND sg13g2_xor2_1
X_4390_ _1094_ _1164_ _1166_ _1167_ VPWR VGND sg13g2_or3_1
Xhold319 mac2.sum_lvl3_ff\[5\] VPWR VGND net359 sg13g2_dlygate4sd3_1
X_3341_ _2925_ _2926_ _2927_ VPWR VGND sg13g2_nor2_1
X_6060_ net275 _0236_ VPWR VGND sg13g2_buf_1
X_3272_ _2824_ _2859_ _2860_ VPWR VGND sg13g2_nor2_1
X_5011_ net825 net880 net828 _1760_ VPWR VGND net877 sg13g2_nand4_1
XFILLER_39_724 VPWR VGND sg13g2_fill_2
X_5913_ VGND VPWR net813 net798 _2567_ _2566_ sg13g2_a21oi_1
XFILLER_34_440 VPWR VGND sg13g2_fill_2
XFILLER_35_985 VPWR VGND sg13g2_decap_8
X_5844_ _2493_ _2498_ _2499_ VPWR VGND sg13g2_and2_1
XFILLER_21_134 VPWR VGND sg13g2_decap_8
XFILLER_10_819 VPWR VGND sg13g2_decap_8
X_5775_ _2429_ _2431_ _2432_ VPWR VGND sg13g2_nor2_1
X_4726_ _1485_ _1486_ _1467_ _1488_ VPWR VGND sg13g2_nand3_1
X_4657_ _1419_ _1418_ _1401_ _1421_ VPWR VGND sg13g2_a21o_1
X_3608_ _0414_ _0415_ _0397_ _0417_ VPWR VGND sg13g2_nand3_1
X_4588_ _0133_ _1350_ _1357_ VPWR VGND sg13g2_xnor2_1
X_6327_ net1100 VGND VPWR net165 mac2.sum_lvl2_ff\[41\] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_3539_ DP_1.matrix\[1\] net970 net1041 _0349_ VPWR VGND net966 sg13g2_nand4_1
XFILLER_27_1028 VPWR VGND sg13g2_fill_1
X_6258_ net1100 VGND VPWR _0266_ DP_4.matrix\[78\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_5209_ _1953_ _1919_ _1951_ VPWR VGND sg13g2_xnor2_1
X_6189_ net1088 VGND VPWR net96 mac1.sum_lvl1_ff\[3\] clknet_leaf_64_clk sg13g2_dfrbpq_1
XFILLER_45_749 VPWR VGND sg13g2_fill_1
XFILLER_26_985 VPWR VGND sg13g2_decap_8
XFILLER_12_101 VPWR VGND sg13g2_fill_1
XFILLER_16_64 VPWR VGND sg13g2_fill_1
XFILLER_40_487 VPWR VGND sg13g2_fill_1
XFILLER_5_801 VPWR VGND sg13g2_decap_4
XFILLER_5_856 VPWR VGND sg13g2_decap_8
XFILLER_16_451 VPWR VGND sg13g2_fill_1
XFILLER_17_974 VPWR VGND sg13g2_decap_8
XFILLER_16_473 VPWR VGND sg13g2_fill_2
X_3890_ _0116_ _0658_ _0685_ VPWR VGND sg13g2_xnor2_1
XFILLER_32_977 VPWR VGND sg13g2_decap_8
X_5560_ _0034_ _2253_ _2254_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_498 VPWR VGND sg13g2_fill_1
X_5491_ _2196_ VPWR _2201_ VGND _2192_ _2195_ sg13g2_o21ai_1
X_4511_ _1263_ VPWR _1284_ VGND _1261_ _1264_ sg13g2_o21ai_1
Xhold116 mac1.sum_lvl1_ff\[8\] VPWR VGND net156 sg13g2_dlygate4sd3_1
X_4442_ _1192_ VPWR _1217_ VGND _1190_ _1193_ sg13g2_o21ai_1
Xhold105 mac2.products_ff\[136\] VPWR VGND net145 sg13g2_dlygate4sd3_1
Xhold149 mac1.products_ff\[74\] VPWR VGND net189 sg13g2_dlygate4sd3_1
Xhold138 mac2.products_ff\[81\] VPWR VGND net178 sg13g2_dlygate4sd3_1
Xhold127 mac2.sum_lvl2_ff\[53\] VPWR VGND net167 sg13g2_dlygate4sd3_1
X_4373_ net845 net891 net848 _1150_ VPWR VGND net1047 sg13g2_nand4_1
X_6112_ net1092 VGND VPWR _0125_ mac1.products_ff\[76\] clknet_leaf_56_clk sg13g2_dfrbpq_1
X_3324_ _2870_ VPWR _2910_ VGND _2867_ _2871_ sg13g2_o21ai_1
X_6043_ net948 _0211_ VPWR VGND sg13g2_buf_1
X_3255_ _2843_ _2791_ _2840_ VPWR VGND sg13g2_xnor2_1
X_3186_ _2776_ _2774_ _2775_ VPWR VGND sg13g2_nand2_1
XFILLER_2_1008 VPWR VGND sg13g2_decap_8
XFILLER_42_708 VPWR VGND sg13g2_fill_1
XFILLER_23_944 VPWR VGND sg13g2_decap_8
XFILLER_22_476 VPWR VGND sg13g2_decap_8
X_5827_ net896 net807 _2482_ VPWR VGND sg13g2_nor2_1
X_5758_ net799 VPWR _2415_ VGND net1023 net808 sg13g2_o21ai_1
X_4709_ VGND VPWR _1471_ _1469_ _1436_ sg13g2_or2_1
X_5689_ _2351_ _2353_ _2349_ _2355_ VPWR VGND sg13g2_nand3_1
XFILLER_2_826 VPWR VGND sg13g2_decap_8
XFILLER_26_771 VPWR VGND sg13g2_decap_8
XFILLER_26_782 VPWR VGND sg13g2_fill_1
XFILLER_14_944 VPWR VGND sg13g2_decap_8
XFILLER_41_730 VPWR VGND sg13g2_decap_4
XFILLER_9_469 VPWR VGND sg13g2_fill_1
XFILLER_4_78 VPWR VGND sg13g2_fill_1
X_3040_ _2636_ net1002 net942 _0064_ VPWR VGND sg13g2_and3_2
XFILLER_49_896 VPWR VGND sg13g2_decap_8
X_4991_ _1741_ net887 net822 VPWR VGND sg13g2_nand2_1
X_3942_ net959 net1009 net963 _0736_ VPWR VGND net1005 sg13g2_nand4_1
X_3873_ net958 net1014 net965 _0669_ VPWR VGND net1011 sg13g2_nand4_1
XFILLER_17_1016 VPWR VGND sg13g2_decap_8
XFILLER_17_1027 VPWR VGND sg13g2_fill_2
XFILLER_20_936 VPWR VGND sg13g2_decap_8
X_5612_ _2287_ _2290_ _2293_ _2295_ VPWR VGND sg13g2_or3_1
X_5543_ VGND VPWR _2236_ _2238_ _2241_ net518 sg13g2_a21oi_1
X_5474_ _2183_ _2185_ _2187_ VPWR VGND sg13g2_nor2_1
X_4425_ _1201_ _1196_ _1200_ VPWR VGND sg13g2_nand2_1
X_4356_ _1133_ net833 net904 net835 net903 VPWR VGND sg13g2_a22oi_1
X_3307_ _2858_ _2892_ _2856_ _2894_ VPWR VGND sg13g2_nand3_1
X_4287_ _1065_ _1032_ _1066_ VPWR VGND sg13g2_xor2_1
X_6026_ net1008 _0186_ VPWR VGND sg13g2_buf_1
X_3238_ _2809_ VPWR _2826_ VGND _2788_ _2810_ sg13g2_o21ai_1
X_3169_ _2754_ VPWR _2759_ VGND _2755_ _2757_ sg13g2_o21ai_1
XFILLER_11_903 VPWR VGND sg13g2_decap_8
XFILLER_13_10 VPWR VGND sg13g2_fill_2
Xhold480 _0046_ VPWR VGND net520 sg13g2_dlygate4sd3_1
Xhold491 _2313_ VPWR VGND net531 sg13g2_dlygate4sd3_1
Xfanout960 net961 net960 VPWR VGND sg13g2_buf_2
XFILLER_46_800 VPWR VGND sg13g2_fill_1
Xfanout982 net322 net982 VPWR VGND sg13g2_buf_8
Xfanout971 net460 net971 VPWR VGND sg13g2_buf_8
Xfanout993 net542 net993 VPWR VGND sg13g2_buf_2
XFILLER_46_833 VPWR VGND sg13g2_fill_2
XFILLER_9_233 VPWR VGND sg13g2_fill_1
XFILLER_9_211 VPWR VGND sg13g2_decap_8
XFILLER_9_277 VPWR VGND sg13g2_fill_2
Xclkload14 clknet_leaf_24_clk clkload14/X VPWR VGND sg13g2_buf_8
XFILLER_10_980 VPWR VGND sg13g2_decap_8
XFILLER_6_951 VPWR VGND sg13g2_decap_8
XFILLER_5_472 VPWR VGND sg13g2_fill_2
X_4210_ _0989_ VPWR _0993_ VGND _0990_ _0991_ sg13g2_o21ai_1
X_5190_ _1934_ net820 net873 VPWR VGND sg13g2_nand2_1
X_4141_ _0929_ _0908_ _0930_ VPWR VGND sg13g2_nor2b_1
X_4072_ _0858_ VPWR _0863_ VGND _0860_ _0861_ sg13g2_o21ai_1
XFILLER_48_192 VPWR VGND sg13g2_fill_1
XFILLER_36_332 VPWR VGND sg13g2_fill_2
XFILLER_24_505 VPWR VGND sg13g2_fill_1
X_4974_ _1728_ _1714_ _1727_ VPWR VGND sg13g2_xnor2_1
X_3925_ _0696_ VPWR _0719_ VGND _0661_ _0694_ sg13g2_o21ai_1
XFILLER_20_722 VPWR VGND sg13g2_decap_8
XFILLER_20_733 VPWR VGND sg13g2_fill_2
X_3856_ _0653_ _0650_ _0652_ VPWR VGND sg13g2_nand2_1
Xclkload8 clknet_4_11_0_clk clkload8/X VPWR VGND sg13g2_buf_8
X_6575_ net1065 VGND VPWR _0061_ mac2.total_sum\[7\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_3787_ _0590_ _0589_ _0584_ _0588_ _0566_ VPWR VGND sg13g2_a22oi_1
XFILLER_30_1013 VPWR VGND sg13g2_decap_8
X_5526_ net513 _2225_ _0042_ VPWR VGND sg13g2_xor2_1
X_5457_ _0027_ _2171_ net547 VPWR VGND sg13g2_xnor2_1
X_4408_ _1184_ _1183_ _1180_ VPWR VGND sg13g2_nand2b_1
X_5388_ VPWR VGND _2114_ _2113_ _2112_ mac1.sum_lvl2_ff\[24\] _2120_ net294 sg13g2_a221oi_1
XFILLER_8_1025 VPWR VGND sg13g2_decap_4
X_4339_ _1114_ _1115_ _1096_ _1117_ VPWR VGND sg13g2_nand3_1
X_6009_ _2631_ _2567_ _2563_ VPWR VGND sg13g2_nand2b_1
Xclkbuf_leaf_66_clk clknet_4_0_0_clk clknet_leaf_66_clk VPWR VGND sg13g2_buf_8
XFILLER_15_527 VPWR VGND sg13g2_fill_2
XFILLER_24_75 VPWR VGND sg13g2_fill_1
XFILLER_11_755 VPWR VGND sg13g2_fill_2
XFILLER_10_265 VPWR VGND sg13g2_fill_1
XFILLER_6_258 VPWR VGND sg13g2_fill_1
XFILLER_3_965 VPWR VGND sg13g2_decap_8
XFILLER_49_50 VPWR VGND sg13g2_fill_2
Xfanout790 _2475_ net790 VPWR VGND sg13g2_buf_1
Xclkbuf_leaf_57_clk clknet_4_8_0_clk clknet_leaf_57_clk VPWR VGND sg13g2_buf_8
XFILLER_19_888 VPWR VGND sg13g2_decap_8
X_3710_ VGND VPWR _0516_ _0514_ _0509_ sg13g2_or2_1
X_4690_ VGND VPWR _1450_ _1451_ _1453_ _1433_ sg13g2_a21oi_1
X_3641_ VGND VPWR _0449_ _0448_ _0399_ sg13g2_or2_1
X_3572_ _0381_ _0317_ _0382_ VPWR VGND sg13g2_xor2_1
X_6360_ net1081 VGND VPWR net153 mac2.sum_lvl1_ff\[76\] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_5311_ VGND VPWR _2051_ _2052_ _2050_ _1991_ sg13g2_a21oi_2
X_6291_ net1097 VGND VPWR net56 mac1.sum_lvl2_ff\[15\] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_5242_ _1985_ _1984_ _1957_ VPWR VGND sg13g2_nand2b_1
X_5173_ _1913_ VPWR _1917_ VGND _1870_ _1915_ sg13g2_o21ai_1
XFILLER_39_0 VPWR VGND sg13g2_fill_2
X_4124_ _0892_ VPWR _0913_ VGND _0890_ _0893_ sg13g2_o21ai_1
XFILLER_28_129 VPWR VGND sg13g2_fill_2
Xinput1 ui_in[0] net1 VPWR VGND sg13g2_buf_1
X_4055_ _0821_ VPWR _0846_ VGND _0819_ _0822_ sg13g2_o21ai_1
Xclkbuf_leaf_48_clk clknet_4_11_0_clk clknet_leaf_48_clk VPWR VGND sg13g2_buf_8
XFILLER_25_825 VPWR VGND sg13g2_fill_1
XFILLER_12_519 VPWR VGND sg13g2_decap_4
X_4957_ _1712_ _1711_ _1708_ VPWR VGND sg13g2_nand2b_1
X_4888_ _1613_ _1645_ _1611_ _1646_ VPWR VGND sg13g2_nand3_1
X_3908_ _0699_ _0700_ _0702_ _0703_ VPWR VGND sg13g2_or3_1
X_3839_ _0637_ _0636_ _0624_ VPWR VGND sg13g2_nand2b_1
X_6558_ net1083 VGND VPWR _0044_ mac2.sum_lvl3_ff\[6\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_3_206 VPWR VGND sg13g2_fill_1
X_5509_ net265 mac1.sum_lvl3_ff\[20\] _0016_ VPWR VGND sg13g2_xor2_1
X_6489_ net1139 VGND VPWR net249 mac2.sum_lvl1_ff\[5\] clknet_leaf_33_clk sg13g2_dfrbpq_1
Xfanout1018 net1020 net1018 VPWR VGND sg13g2_buf_8
XFILLER_0_924 VPWR VGND sg13g2_decap_8
Xfanout1007 net399 net1007 VPWR VGND sg13g2_buf_2
Xfanout1029 net408 net1029 VPWR VGND sg13g2_buf_8
XFILLER_48_928 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_39_clk clknet_4_15_0_clk clknet_leaf_39_clk VPWR VGND sg13g2_buf_8
XFILLER_16_825 VPWR VGND sg13g2_decap_8
XFILLER_30_305 VPWR VGND sg13g2_fill_1
XFILLER_3_773 VPWR VGND sg13g2_fill_2
XFILLER_47_994 VPWR VGND sg13g2_decap_8
XFILLER_19_652 VPWR VGND sg13g2_decap_4
X_5860_ _2512_ VPWR _2515_ VGND net794 _2514_ sg13g2_o21ai_1
XFILLER_34_644 VPWR VGND sg13g2_fill_1
X_4811_ _1569_ _1570_ _1571_ VPWR VGND sg13g2_nor2_1
X_5791_ net808 _2402_ DP_2.matrix\[75\] _2447_ VPWR VGND sg13g2_nand3_1
X_4742_ net922 net921 net854 net851 _1503_ VPWR VGND sg13g2_and4_1
X_4673_ _1436_ net919 net859 VPWR VGND sg13g2_nand2_1
X_3624_ _0422_ VPWR _0432_ VGND _0351_ _0423_ sg13g2_o21ai_1
X_6412_ net1078 VGND VPWR net205 mac2.sum_lvl3_ff\[28\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_6343_ net1071 VGND VPWR net126 mac1.sum_lvl1_ff\[75\] clknet_leaf_66_clk sg13g2_dfrbpq_1
X_3555_ _0365_ net1025 net983 net1028 net980 VPWR VGND sg13g2_a22oi_1
X_3486_ _0298_ net1030 net983 net1032 net979 VPWR VGND sg13g2_a22oi_1
X_6274_ net1096 VGND VPWR net177 mac1.sum_lvl1_ff\[50\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_5225_ _1967_ _1959_ _1968_ VPWR VGND sg13g2_nor2b_1
X_5156_ _1889_ VPWR _1901_ VGND _1897_ _1899_ sg13g2_o21ai_1
XFILLER_5_1028 VPWR VGND sg13g2_fill_1
XFILLER_5_1017 VPWR VGND sg13g2_decap_8
XFILLER_29_416 VPWR VGND sg13g2_fill_1
X_5087_ _1810_ VPWR _1833_ VGND _1775_ _1808_ sg13g2_o21ai_1
X_4107_ _0895_ _0888_ _0897_ VPWR VGND sg13g2_xor2_1
X_4038_ _0830_ _0825_ _0829_ VPWR VGND sg13g2_nand2_1
X_5989_ VPWR _0227_ _2618_ VGND sg13g2_inv_1
XFILLER_24_187 VPWR VGND sg13g2_fill_2
XFILLER_4_526 VPWR VGND sg13g2_fill_2
XFILLER_21_98 VPWR VGND sg13g2_decap_8
XFILLER_0_798 VPWR VGND sg13g2_decap_8
XFILLER_29_961 VPWR VGND sg13g2_decap_8
XFILLER_44_964 VPWR VGND sg13g2_decap_8
XFILLER_16_688 VPWR VGND sg13g2_fill_1
XFILLER_16_699 VPWR VGND sg13g2_fill_2
XFILLER_12_850 VPWR VGND sg13g2_decap_8
XFILLER_7_320 VPWR VGND sg13g2_fill_2
Xhold309 DP_3.matrix\[36\] VPWR VGND net349 sg13g2_dlygate4sd3_1
X_3340_ VGND VPWR _2889_ _2891_ _2926_ _2923_ sg13g2_a21oi_1
X_5010_ net828 net825 net881 net877 _1759_ VPWR VGND sg13g2_and4_1
X_3271_ _2859_ _2825_ _2857_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_4 VPWR VGND sg13g2_fill_1
X_5912_ net796 _2564_ _2565_ _2566_ VPWR VGND sg13g2_nor3_1
X_5843_ VGND VPWR _2494_ _2496_ _2498_ _2497_ sg13g2_a21oi_1
X_5774_ _2431_ net800 _2430_ net802 DP_1.matrix\[78\] VPWR VGND sg13g2_a22oi_1
X_4725_ _1487_ _1467_ _1485_ _1486_ VPWR VGND sg13g2_and3_1
X_4656_ _1418_ _1419_ _1401_ _1420_ VPWR VGND sg13g2_nand3_1
X_3607_ _0416_ _0397_ _0414_ _0415_ VPWR VGND sg13g2_and3_1
X_4587_ _1357_ _1351_ _1356_ VPWR VGND sg13g2_xnor2_1
X_3538_ _0348_ net966 net1041 net970 net1039 VPWR VGND sg13g2_a22oi_1
X_6326_ net1100 VGND VPWR net152 mac2.sum_lvl2_ff\[40\] clknet_leaf_28_clk sg13g2_dfrbpq_1
XFILLER_27_1007 VPWR VGND sg13g2_decap_8
X_6257_ net1123 VGND VPWR _0265_ DP_4.matrix\[77\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_3469_ _0282_ _0270_ _0281_ VPWR VGND sg13g2_xnor2_1
X_5208_ _1952_ _1919_ _1951_ VPWR VGND sg13g2_nand2b_1
X_6188_ net1070 VGND VPWR _0209_ DP_2.matrix\[41\] clknet_leaf_2_clk sg13g2_dfrbpq_2
X_5139_ _1884_ net880 net816 VPWR VGND sg13g2_nand2_1
XFILLER_38_791 VPWR VGND sg13g2_fill_2
XFILLER_26_964 VPWR VGND sg13g2_decap_8
XFILLER_41_912 VPWR VGND sg13g2_fill_2
XFILLER_40_444 VPWR VGND sg13g2_fill_1
XFILLER_8_117 VPWR VGND sg13g2_fill_1
XFILLER_5_835 VPWR VGND sg13g2_decap_8
XFILLER_10_1022 VPWR VGND sg13g2_decap_8
XFILLER_29_780 VPWR VGND sg13g2_fill_1
XFILLER_17_953 VPWR VGND sg13g2_decap_8
XFILLER_31_411 VPWR VGND sg13g2_decap_8
XFILLER_8_662 VPWR VGND sg13g2_fill_1
X_5490_ net540 mac1.sum_lvl3_ff\[32\] _2200_ VPWR VGND sg13g2_xor2_1
X_4510_ _1283_ _1282_ _1280_ VPWR VGND sg13g2_nand2b_1
Xhold106 mac1.products_ff\[75\] VPWR VGND net146 sg13g2_dlygate4sd3_1
Xhold117 mac1.sum_lvl1_ff\[75\] VPWR VGND net157 sg13g2_dlygate4sd3_1
X_4441_ _1184_ VPWR _1216_ VGND _1131_ _1182_ sg13g2_o21ai_1
Xhold128 mac1.sum_lvl1_ff\[7\] VPWR VGND net168 sg13g2_dlygate4sd3_1
Xhold139 mac2.products_ff\[3\] VPWR VGND net179 sg13g2_dlygate4sd3_1
X_6111_ net1090 VGND VPWR _0124_ mac1.products_ff\[75\] clknet_leaf_63_clk sg13g2_dfrbpq_1
X_4372_ net849 net844 net891 net1047 _1149_ VPWR VGND sg13g2_and4_1
X_3323_ _2909_ _2901_ _2906_ VPWR VGND sg13g2_xnor2_1
X_6042_ net950 _0210_ VPWR VGND sg13g2_buf_1
X_3254_ _2791_ _2840_ _2842_ VPWR VGND sg13g2_and2_1
XFILLER_21_0 VPWR VGND sg13g2_fill_1
X_3185_ _2737_ _2736_ _2735_ _2775_ VPWR VGND sg13g2_a21o_2
XFILLER_23_923 VPWR VGND sg13g2_decap_8
XFILLER_35_783 VPWR VGND sg13g2_fill_1
X_5826_ _2481_ _2476_ _2477_ VPWR VGND sg13g2_xnor2_1
X_5757_ net1040 net809 _2414_ VPWR VGND sg13g2_nor2_1
X_4708_ _1470_ net859 net917 VPWR VGND sg13g2_nand2_1
X_5688_ VGND VPWR _2349_ _2351_ _2354_ _2353_ sg13g2_a21oi_1
X_4639_ _1403_ net921 net858 VPWR VGND sg13g2_nand2_1
XFILLER_2_805 VPWR VGND sg13g2_decap_8
X_6309_ net1062 VGND VPWR net215 mac1.sum_lvl2_ff\[39\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_40_1015 VPWR VGND sg13g2_decap_8
XFILLER_14_923 VPWR VGND sg13g2_decap_8
XFILLER_43_63 VPWR VGND sg13g2_fill_2
XFILLER_4_197 VPWR VGND sg13g2_fill_1
XFILLER_49_820 VPWR VGND sg13g2_fill_2
XFILLER_1_893 VPWR VGND sg13g2_decap_8
XFILLER_49_864 VPWR VGND sg13g2_fill_2
X_4990_ VGND VPWR _1740_ _1735_ _1733_ sg13g2_or2_1
X_3941_ net962 net959 net1009 net1005 _0735_ VPWR VGND sg13g2_and4_1
X_3872_ net962 net958 net1013 net1010 _0668_ VPWR VGND sg13g2_and4_1
XFILLER_20_915 VPWR VGND sg13g2_decap_8
XFILLER_31_263 VPWR VGND sg13g2_fill_2
X_6591_ net1086 VGND VPWR DP_3.I_range.data_plus_4\[6\] DP_3.I_range.out_data\[5\]
+ clknet_leaf_21_clk sg13g2_dfrbpq_1
X_5611_ _2293_ VPWR _2294_ VGND _2287_ _2290_ sg13g2_o21ai_1
X_5542_ _2240_ mac2.sum_lvl2_ff\[27\] net517 VPWR VGND sg13g2_xnor2_1
X_5473_ net496 _2186_ _0030_ VPWR VGND sg13g2_nor2b_2
X_4424_ _1198_ _1199_ _1200_ VPWR VGND sg13g2_nor2_1
X_4355_ net904 net903 net835 net833 _1132_ VPWR VGND sg13g2_and4_1
X_3306_ VGND VPWR _2856_ _2858_ _2893_ _2892_ sg13g2_a21oi_1
X_4286_ _1065_ net901 net840 VPWR VGND sg13g2_nand2_2
X_6025_ net1012 _0185_ VPWR VGND sg13g2_buf_1
X_3237_ _2786_ VPWR _2825_ VGND _2741_ _2787_ sg13g2_o21ai_1
X_3168_ _2754_ _2755_ _2757_ _2758_ VPWR VGND sg13g2_or3_1
X_3099_ _2687_ _2688_ _2690_ _2691_ VPWR VGND sg13g2_or3_1
XFILLER_11_959 VPWR VGND sg13g2_decap_8
X_5809_ net969 net950 _2396_ _2465_ VPWR VGND sg13g2_mux2_1
XFILLER_7_919 VPWR VGND sg13g2_decap_8
Xhold470 _2189_ VPWR VGND net510 sg13g2_dlygate4sd3_1
Xhold481 mac1.sum_lvl3_ff\[10\] VPWR VGND net521 sg13g2_dlygate4sd3_1
Xhold492 mac1.sum_lvl3_ff\[6\] VPWR VGND net532 sg13g2_dlygate4sd3_1
Xfanout950 net415 net950 VPWR VGND sg13g2_buf_1
Xfanout961 net524 net961 VPWR VGND sg13g2_buf_8
Xfanout994 net995 net994 VPWR VGND sg13g2_buf_8
Xfanout983 net984 net983 VPWR VGND sg13g2_buf_2
Xfanout972 net414 net972 VPWR VGND sg13g2_buf_8
XFILLER_45_333 VPWR VGND sg13g2_fill_1
XFILLER_26_580 VPWR VGND sg13g2_fill_1
XFILLER_6_930 VPWR VGND sg13g2_decap_8
Xclkload15 clkload15/Y clknet_leaf_47_clk VPWR VGND sg13g2_inv_2
XFILLER_5_495 VPWR VGND sg13g2_fill_1
X_4140_ _0927_ _0926_ _0929_ VPWR VGND sg13g2_xor2_1
X_4071_ _0858_ _0860_ _0861_ _0862_ VPWR VGND sg13g2_nor3_1
XFILLER_23_1021 VPWR VGND sg13g2_decap_8
X_4973_ _1727_ _1724_ _1726_ VPWR VGND sg13g2_xnor2_1
X_3924_ _0710_ VPWR _0718_ VGND _0690_ _0711_ sg13g2_o21ai_1
X_3855_ _0649_ _0648_ _0643_ _0652_ VPWR VGND sg13g2_a21o_1
Xclkload9 clknet_4_13_0_clk clkload9/X VPWR VGND sg13g2_buf_8
X_6574_ net1061 VGND VPWR net490 mac2.total_sum\[6\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_3786_ _0583_ VPWR _0589_ VGND _0560_ _0561_ sg13g2_o21ai_1
X_5525_ net512 mac2.sum_lvl2_ff\[23\] _2227_ VPWR VGND sg13g2_xor2_1
X_5456_ net546 mac1.sum_lvl3_ff\[25\] _2173_ VPWR VGND sg13g2_xor2_1
X_4407_ _1182_ _1131_ _1183_ VPWR VGND sg13g2_xor2_1
XFILLER_8_1004 VPWR VGND sg13g2_decap_8
X_5387_ _2119_ mac1.sum_lvl2_ff\[25\] net461 VPWR VGND sg13g2_xnor2_1
X_4338_ _1116_ _1096_ _1114_ _1115_ VPWR VGND sg13g2_and3_1
X_4269_ _1047_ _1048_ _1030_ _1049_ VPWR VGND sg13g2_nand3_1
X_6008_ _2629_ VPWR _0250_ VGND net791 _2630_ sg13g2_o21ai_1
XFILLER_43_837 VPWR VGND sg13g2_fill_2
XFILLER_11_734 VPWR VGND sg13g2_fill_1
XFILLER_23_583 VPWR VGND sg13g2_fill_1
XFILLER_11_767 VPWR VGND sg13g2_fill_1
XFILLER_3_944 VPWR VGND sg13g2_decap_8
Xfanout791 net792 net791 VPWR VGND sg13g2_buf_8
XFILLER_46_642 VPWR VGND sg13g2_fill_1
XFILLER_19_867 VPWR VGND sg13g2_decap_8
X_3640_ _0448_ net975 net1027 VPWR VGND sg13g2_nand2_1
X_3571_ _0381_ _0378_ _0380_ VPWR VGND sg13g2_nand2_1
X_5310_ VGND VPWR _1988_ _2018_ _2051_ _2020_ sg13g2_a21oi_1
X_6290_ net1097 VGND VPWR net58 mac1.sum_lvl2_ff\[14\] clknet_leaf_29_clk sg13g2_dfrbpq_1
X_5241_ _1982_ _1958_ _1984_ VPWR VGND sg13g2_xor2_1
X_5172_ _1915_ _1870_ _0158_ VPWR VGND sg13g2_xor2_1
X_4123_ _0912_ _0911_ _0909_ VPWR VGND sg13g2_nand2b_1
X_4054_ _0813_ VPWR _0845_ VGND _0760_ _0811_ sg13g2_o21ai_1
Xinput2 ui_in[1] net2 VPWR VGND sg13g2_buf_1
XFILLER_24_369 VPWR VGND sg13g2_fill_1
X_4956_ _1710_ _1684_ _1711_ VPWR VGND sg13g2_xor2_1
X_4887_ _1643_ _1621_ _1645_ VPWR VGND sg13g2_xor2_1
X_3907_ _0702_ net1009 DP_2.matrix\[36\] net1011 net958 VPWR VGND sg13g2_a22oi_1
X_3838_ _0635_ _0625_ _0636_ VPWR VGND sg13g2_xor2_1
X_6557_ net1083 VGND VPWR net471 mac2.sum_lvl3_ff\[5\] clknet_leaf_12_clk sg13g2_dfrbpq_2
X_3769_ _0573_ _0572_ _0569_ VPWR VGND sg13g2_nand2b_1
X_5508_ _0022_ _2213_ net290 VPWR VGND sg13g2_xnor2_1
X_6488_ net1127 VGND VPWR net133 mac2.sum_lvl1_ff\[4\] clknet_leaf_33_clk sg13g2_dfrbpq_1
XFILLER_0_903 VPWR VGND sg13g2_decap_8
X_5439_ mac1.sum_lvl3_ff\[21\] mac1.sum_lvl3_ff\[1\] _2160_ VPWR VGND sg13g2_nor2_1
Xfanout1019 net1020 net1019 VPWR VGND sg13g2_buf_1
Xfanout1008 net369 net1008 VPWR VGND sg13g2_buf_8
XFILLER_19_32 VPWR VGND sg13g2_fill_1
XFILLER_28_631 VPWR VGND sg13g2_decap_4
XFILLER_16_804 VPWR VGND sg13g2_decap_8
XFILLER_37_1009 VPWR VGND sg13g2_decap_8
XFILLER_20_1013 VPWR VGND sg13g2_decap_8
XFILLER_47_973 VPWR VGND sg13g2_decap_8
XFILLER_18_163 VPWR VGND sg13g2_fill_2
X_4810_ _1570_ net1049 net866 net908 net862 VPWR VGND sg13g2_a22oi_1
X_5790_ VGND VPWR net955 net809 _2446_ _2445_ sg13g2_a21oi_1
X_4741_ _1502_ net921 net851 VPWR VGND sg13g2_nand2_1
X_4672_ _1435_ net919 net857 VPWR VGND sg13g2_nand2_1
X_3623_ _0427_ VPWR _0431_ VGND _0384_ _0429_ sg13g2_o21ai_1
X_6411_ net1082 VGND VPWR net85 mac2.sum_lvl3_ff\[27\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_6342_ net1069 VGND VPWR net43 mac1.sum_lvl1_ff\[74\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3554_ net980 net1028 net983 _0364_ VPWR VGND net1025 sg13g2_nand4_1
X_3485_ net979 net1033 net983 _0297_ VPWR VGND net1030 sg13g2_nand4_1
X_6273_ net1097 VGND VPWR net253 mac1.sum_lvl1_ff\[49\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_5224_ _1967_ _1960_ _1966_ VPWR VGND sg13g2_xnor2_1
X_5155_ _1889_ _1897_ _1899_ _1900_ VPWR VGND sg13g2_or3_1
X_5086_ _1824_ VPWR _1832_ VGND _1804_ _1825_ sg13g2_o21ai_1
X_4106_ _0895_ _0888_ _0896_ VPWR VGND sg13g2_nor2b_1
X_4037_ _0827_ _0828_ _0829_ VPWR VGND sg13g2_nor2_1
XFILLER_38_995 VPWR VGND sg13g2_decap_8
X_5988_ _2618_ _2522_ _2617_ net792 net910 VPWR VGND sg13g2_a22oi_1
X_4939_ _1693_ _1668_ _1695_ VPWR VGND sg13g2_xor2_1
XFILLER_24_199 VPWR VGND sg13g2_fill_1
XFILLER_0_722 VPWR VGND sg13g2_decap_8
XFILLER_0_777 VPWR VGND sg13g2_decap_8
XFILLER_47_225 VPWR VGND sg13g2_fill_2
XFILLER_16_667 VPWR VGND sg13g2_fill_2
XFILLER_11_350 VPWR VGND sg13g2_fill_2
XFILLER_8_899 VPWR VGND sg13g2_decap_8
X_3270_ _2858_ _2825_ _2857_ VPWR VGND sg13g2_nand2b_1
X_5911_ net833 net807 _2565_ VPWR VGND sg13g2_nor2_1
XFILLER_34_442 VPWR VGND sg13g2_fill_1
X_5842_ net923 _2495_ _2497_ VPWR VGND sg13g2_nor2_1
X_5773_ net1029 DP_1.matrix\[42\] net810 _2430_ VPWR VGND sg13g2_mux2_1
XFILLER_22_659 VPWR VGND sg13g2_decap_8
X_4724_ _1474_ VPWR _1486_ VGND _1482_ _1484_ sg13g2_o21ai_1
X_4655_ _1407_ VPWR _1419_ VGND _1415_ _1417_ sg13g2_o21ai_1
X_3606_ _0403_ VPWR _0415_ VGND _0411_ _0413_ sg13g2_o21ai_1
X_4586_ _1356_ _1343_ _1355_ VPWR VGND sg13g2_xnor2_1
X_3537_ _0324_ VPWR _0347_ VGND _0289_ _0322_ sg13g2_o21ai_1
X_6325_ net1101 VGND VPWR net163 mac2.sum_lvl2_ff\[39\] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_6256_ net1123 VGND VPWR _0264_ DP_4.matrix\[76\] clknet_leaf_25_clk sg13g2_dfrbpq_2
X_3468_ _0281_ _0278_ _0280_ VPWR VGND sg13g2_nand2_1
X_5207_ _1951_ _1920_ _1949_ VPWR VGND sg13g2_xnor2_1
X_6187_ net1088 VGND VPWR _0208_ DP_2.matrix\[40\] clknet_leaf_65_clk sg13g2_dfrbpq_1
X_3399_ _2982_ _2981_ _2976_ _2980_ _2958_ VPWR VGND sg13g2_a22oi_1
X_5138_ _1855_ VPWR _1883_ VGND _1846_ _1856_ sg13g2_o21ai_1
X_5069_ _1816_ net873 net829 net875 net824 VPWR VGND sg13g2_a22oi_1
XFILLER_26_943 VPWR VGND sg13g2_decap_8
XFILLER_41_979 VPWR VGND sg13g2_decap_8
XFILLER_32_43 VPWR VGND sg13g2_fill_1
XFILLER_5_814 VPWR VGND sg13g2_decap_8
XFILLER_10_1001 VPWR VGND sg13g2_decap_8
XFILLER_17_932 VPWR VGND sg13g2_decap_8
XFILLER_16_464 VPWR VGND sg13g2_decap_4
XFILLER_32_924 VPWR VGND sg13g2_fill_2
XFILLER_7_140 VPWR VGND sg13g2_fill_1
Xhold107 mac1.sum_lvl1_ff\[39\] VPWR VGND net147 sg13g2_dlygate4sd3_1
X_4440_ _1204_ VPWR _1215_ VGND _1188_ _1205_ sg13g2_o21ai_1
Xhold118 mac2.sum_lvl1_ff\[2\] VPWR VGND net158 sg13g2_dlygate4sd3_1
Xhold129 mac2.products_ff\[2\] VPWR VGND net169 sg13g2_dlygate4sd3_1
XFILLER_4_880 VPWR VGND sg13g2_decap_8
X_6110_ net1090 VGND VPWR _0123_ mac1.products_ff\[74\] clknet_leaf_63_clk sg13g2_dfrbpq_1
X_4371_ _1148_ net842 net894 VPWR VGND sg13g2_nand2_1
X_3322_ VGND VPWR _2908_ _2906_ _2901_ sg13g2_or2_1
X_6041_ net951 _0209_ VPWR VGND sg13g2_buf_1
X_3253_ VGND VPWR _2841_ _2840_ _2791_ sg13g2_or2_1
X_3184_ _2773_ _2709_ _2774_ VPWR VGND sg13g2_xor2_1
XFILLER_35_762 VPWR VGND sg13g2_fill_1
XFILLER_22_434 VPWR VGND sg13g2_fill_2
X_5825_ _2476_ net805 _2480_ VPWR VGND sg13g2_nor2_1
XFILLER_23_979 VPWR VGND sg13g2_decap_8
X_5756_ _2413_ net1003 net801 VPWR VGND sg13g2_nand2_1
XFILLER_33_1023 VPWR VGND sg13g2_decap_4
X_4707_ _1469_ net917 net857 VPWR VGND sg13g2_nand2_1
X_5687_ _2353_ mac1.total_sum\[8\] mac2.total_sum\[8\] VPWR VGND sg13g2_xnor2_1
X_4638_ _1402_ net925 net856 VPWR VGND sg13g2_nand2_1
X_4569_ _1339_ _1312_ _1340_ VPWR VGND sg13g2_xor2_1
X_6308_ net1064 VGND VPWR net164 mac1.sum_lvl2_ff\[38\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_6239_ net1124 VGND VPWR net385 DP_4.matrix\[3\] clknet_leaf_35_clk sg13g2_dfrbpq_2
XFILLER_13_401 VPWR VGND sg13g2_fill_1
XFILLER_14_902 VPWR VGND sg13g2_decap_8
XFILLER_14_979 VPWR VGND sg13g2_decap_8
XFILLER_1_872 VPWR VGND sg13g2_decap_8
XFILLER_49_843 VPWR VGND sg13g2_decap_8
XFILLER_48_386 VPWR VGND sg13g2_fill_1
XFILLER_36_548 VPWR VGND sg13g2_fill_1
X_3940_ _0734_ net956 net1010 VPWR VGND sg13g2_nand2_1
XFILLER_17_784 VPWR VGND sg13g2_fill_1
X_3871_ _0667_ net956 net1016 VPWR VGND sg13g2_nand2_1
X_6590_ net1086 VGND VPWR net15 DP_3.I_range.out_data\[4\] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_5610_ net545 net454 _2293_ VPWR VGND sg13g2_xor2_1
X_5541_ _2238_ _2239_ _0045_ VPWR VGND sg13g2_and2_1
XFILLER_9_994 VPWR VGND sg13g2_decap_8
X_5472_ _2181_ _2184_ _2179_ _2186_ VPWR VGND sg13g2_nand3_1
X_4423_ _1199_ net1047 net845 net891 net843 VPWR VGND sg13g2_a22oi_1
X_4354_ _1131_ net903 net833 VPWR VGND sg13g2_nand2_1
X_3305_ _2890_ _2863_ _2892_ VPWR VGND sg13g2_xor2_1
X_6024_ net1015 _0184_ VPWR VGND sg13g2_buf_1
X_4285_ _1064_ net901 net839 VPWR VGND sg13g2_nand2_1
X_3236_ _2814_ VPWR _2824_ VGND _2743_ _2815_ sg13g2_o21ai_1
X_3167_ _2757_ net986 net943 net990 net938 VPWR VGND sg13g2_a22oi_1
X_3098_ _2690_ net991 net944 net994 net940 VPWR VGND sg13g2_a22oi_1
XFILLER_23_710 VPWR VGND sg13g2_fill_1
XFILLER_22_220 VPWR VGND sg13g2_decap_4
X_5808_ VGND VPWR _2464_ _2463_ _2444_ sg13g2_or2_1
XFILLER_11_938 VPWR VGND sg13g2_decap_8
XFILLER_13_12 VPWR VGND sg13g2_fill_1
XFILLER_23_798 VPWR VGND sg13g2_fill_1
X_5739_ DP_1.Q_range.out_data\[2\] DP_1.I_range.out_data\[2\] _2396_ VPWR VGND sg13g2_xor2_1
Xhold471 _0031_ VPWR VGND net511 sg13g2_dlygate4sd3_1
Xhold460 _0056_ VPWR VGND net500 sg13g2_dlygate4sd3_1
Xhold493 _2175_ VPWR VGND net533 sg13g2_dlygate4sd3_1
Xhold482 _2193_ VPWR VGND net522 sg13g2_dlygate4sd3_1
Xfanout940 net941 net940 VPWR VGND sg13g2_buf_1
Xfanout951 net400 net951 VPWR VGND sg13g2_buf_8
XFILLER_1_179 VPWR VGND sg13g2_fill_1
Xfanout995 net528 net995 VPWR VGND sg13g2_buf_8
Xfanout984 net985 net984 VPWR VGND sg13g2_buf_1
Xfanout962 net964 net962 VPWR VGND sg13g2_buf_2
Xfanout973 DP_2.matrix\[4\] net973 VPWR VGND sg13g2_buf_1
XFILLER_46_835 VPWR VGND sg13g2_fill_1
XFILLER_45_301 VPWR VGND sg13g2_fill_1
XFILLER_45_367 VPWR VGND sg13g2_fill_2
XFILLER_13_275 VPWR VGND sg13g2_fill_2
XFILLER_14_798 VPWR VGND sg13g2_decap_8
XFILLER_9_268 VPWR VGND sg13g2_fill_1
Xclkload16 clknet_leaf_60_clk clkload16/Y VPWR VGND sg13g2_inv_4
XFILLER_6_986 VPWR VGND sg13g2_decap_8
XFILLER_5_474 VPWR VGND sg13g2_fill_1
X_4070_ _0861_ net1006 net954 net1008 net952 VPWR VGND sg13g2_a22oi_1
XFILLER_23_1000 VPWR VGND sg13g2_decap_8
XFILLER_37_835 VPWR VGND sg13g2_fill_2
X_4972_ _1725_ _1709_ _1726_ VPWR VGND sg13g2_xor2_1
X_3923_ _0717_ _0716_ _0123_ VPWR VGND sg13g2_xor2_1
X_3854_ VGND VPWR _0648_ _0649_ _0651_ _0643_ sg13g2_a21oi_1
X_6573_ net1060 VGND VPWR net361 mac2.total_sum\[5\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_3785_ VPWR _0588_ _0587_ VGND sg13g2_inv_1
X_5524_ mac2.sum_lvl2_ff\[23\] mac2.sum_lvl2_ff\[4\] _2226_ VPWR VGND sg13g2_and2_1
X_5455_ mac1.sum_lvl3_ff\[25\] mac1.sum_lvl3_ff\[5\] _2172_ VPWR VGND sg13g2_nor2_1
X_4406_ _1182_ net901 net836 VPWR VGND sg13g2_nand2_1
X_5386_ mac1.sum_lvl2_ff\[25\] net461 _2118_ VPWR VGND sg13g2_and2_1
X_4337_ _1103_ VPWR _1115_ VGND _1111_ _1113_ sg13g2_o21ai_1
X_4268_ _1036_ VPWR _1048_ VGND _1044_ _1046_ sg13g2_o21ai_1
X_6007_ _2562_ _2558_ _2630_ VPWR VGND sg13g2_xor2_1
X_3219_ _2808_ _2789_ _2806_ _2807_ VPWR VGND sg13g2_and3_1
X_4199_ _0985_ _0972_ _0984_ VPWR VGND sg13g2_xnor2_1
XFILLER_42_326 VPWR VGND sg13g2_fill_1
XFILLER_23_540 VPWR VGND sg13g2_fill_1
XFILLER_10_223 VPWR VGND sg13g2_fill_1
XFILLER_40_43 VPWR VGND sg13g2_fill_2
XFILLER_3_923 VPWR VGND sg13g2_decap_8
XFILLER_46_1022 VPWR VGND sg13g2_decap_8
Xhold290 DP_4.matrix\[40\] VPWR VGND net330 sg13g2_dlygate4sd3_1
Xfanout792 net793 net792 VPWR VGND sg13g2_buf_8
XFILLER_19_824 VPWR VGND sg13g2_fill_1
X_3570_ _0377_ _0376_ _0346_ _0380_ VPWR VGND sg13g2_a21o_1
X_5240_ _1983_ _1958_ _1982_ VPWR VGND sg13g2_nand2_1
XFILLER_5_293 VPWR VGND sg13g2_fill_1
X_5171_ _1868_ _1869_ _1913_ _1914_ _1916_ VPWR VGND sg13g2_and4_1
X_4122_ VGND VPWR _0911_ _0910_ _0859_ sg13g2_or2_1
X_4053_ _0833_ VPWR _0844_ VGND _0817_ _0834_ sg13g2_o21ai_1
Xinput3 ui_in[2] net3 VPWR VGND sg13g2_buf_1
XFILLER_37_632 VPWR VGND sg13g2_fill_2
XFILLER_25_816 VPWR VGND sg13g2_decap_8
X_4955_ _1710_ net855 net1050 VPWR VGND sg13g2_nand2_1
XFILLER_24_337 VPWR VGND sg13g2_fill_1
XFILLER_40_819 VPWR VGND sg13g2_fill_1
X_3906_ net958 net1011 net965 _0701_ VPWR VGND net1009 sg13g2_nand4_1
XFILLER_33_860 VPWR VGND sg13g2_fill_2
X_4886_ _1643_ _1621_ _1644_ VPWR VGND sg13g2_nor2b_1
X_3837_ _0635_ _0626_ _0633_ VPWR VGND sg13g2_xnor2_1
X_3768_ _0571_ _0545_ _0572_ VPWR VGND sg13g2_xor2_1
X_6556_ net1083 VGND VPWR net514 mac2.sum_lvl3_ff\[4\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_5507_ _2214_ mac1.sum_lvl3_ff\[35\] net289 VPWR VGND sg13g2_xnor2_1
XFILLER_3_219 VPWR VGND sg13g2_decap_8
X_3699_ _0503_ _0505_ _0506_ VPWR VGND sg13g2_nor2_1
X_6487_ net1124 VGND VPWR net179 mac2.sum_lvl1_ff\[3\] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_5438_ _2159_ mac1.sum_lvl3_ff\[21\] mac1.sum_lvl3_ff\[1\] VPWR VGND sg13g2_nand2_1
Xfanout1009 DP_1.matrix\[42\] net1009 VPWR VGND sg13g2_buf_1
X_5369_ _0007_ _2102_ _2105_ VPWR VGND sg13g2_xnor2_1
XFILLER_0_959 VPWR VGND sg13g2_decap_8
XFILLER_28_621 VPWR VGND sg13g2_fill_2
XFILLER_31_808 VPWR VGND sg13g2_fill_2
XFILLER_7_514 VPWR VGND sg13g2_fill_2
XFILLER_13_1010 VPWR VGND sg13g2_decap_8
XFILLER_3_775 VPWR VGND sg13g2_fill_1
XFILLER_25_8 VPWR VGND sg13g2_fill_1
XFILLER_47_952 VPWR VGND sg13g2_decap_8
XFILLER_33_123 VPWR VGND sg13g2_fill_2
X_4740_ _1501_ net925 net1044 VPWR VGND sg13g2_nand2_1
X_4671_ _1434_ net922 DP_4.matrix\[5\] VPWR VGND sg13g2_nand2_1
X_3622_ _0429_ _0384_ _0114_ VPWR VGND sg13g2_xor2_1
X_6410_ net1082 VGND VPWR net113 mac2.sum_lvl3_ff\[26\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_6341_ net1062 VGND VPWR net95 mac1.sum_lvl1_ff\[73\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_3553_ net984 net980 net1028 net1025 _0363_ VPWR VGND sg13g2_and4_1
X_3484_ net984 net979 net1032 net1030 _0296_ VPWR VGND sg13g2_and4_1
X_6272_ net1096 VGND VPWR net230 mac1.sum_lvl1_ff\[48\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_5223_ _1965_ _1961_ _1966_ VPWR VGND sg13g2_xor2_1
X_5154_ VGND VPWR _1895_ _1896_ _1899_ _1890_ sg13g2_a21oi_1
X_4105_ _0895_ _0889_ _0894_ VPWR VGND sg13g2_xnor2_1
X_5085_ _1831_ _1830_ _0156_ VPWR VGND sg13g2_xor2_1
X_4036_ _0828_ net1057 net960 net1005 net956 VPWR VGND sg13g2_a22oi_1
XFILLER_25_668 VPWR VGND sg13g2_fill_2
X_5987_ _2617_ _2520_ _2516_ VPWR VGND sg13g2_nand2b_1
X_4938_ _1668_ _1693_ _1694_ VPWR VGND sg13g2_nor2_1
XFILLER_24_189 VPWR VGND sg13g2_fill_1
X_4869_ _1627_ _1601_ _1625_ VPWR VGND sg13g2_xnor2_1
X_6539_ net1137 VGND VPWR net53 mac2.sum_lvl2_ff\[26\] clknet_leaf_43_clk sg13g2_dfrbpq_1
XFILLER_43_1014 VPWR VGND sg13g2_decap_8
XFILLER_0_756 VPWR VGND sg13g2_decap_8
XFILLER_29_930 VPWR VGND sg13g2_fill_1
XFILLER_29_996 VPWR VGND sg13g2_decap_8
XFILLER_44_999 VPWR VGND sg13g2_decap_8
XFILLER_7_322 VPWR VGND sg13g2_fill_1
XFILLER_12_885 VPWR VGND sg13g2_decap_8
XFILLER_8_878 VPWR VGND sg13g2_decap_8
XFILLER_39_738 VPWR VGND sg13g2_fill_1
XFILLER_47_760 VPWR VGND sg13g2_fill_2
XFILLER_19_451 VPWR VGND sg13g2_fill_1
XFILLER_38_248 VPWR VGND sg13g2_fill_2
XFILLER_47_771 VPWR VGND sg13g2_fill_2
X_5910_ net853 net803 _2564_ VPWR VGND sg13g2_nor2_1
XFILLER_35_911 VPWR VGND sg13g2_fill_2
XFILLER_19_495 VPWR VGND sg13g2_decap_8
X_5841_ net806 VPWR _2496_ VGND net888 _2476_ sg13g2_o21ai_1
XFILLER_35_999 VPWR VGND sg13g2_decap_8
X_5772_ VGND VPWR _2429_ _2428_ _2408_ sg13g2_or2_1
XFILLER_22_638 VPWR VGND sg13g2_decap_8
X_4723_ _1474_ _1482_ _1484_ _1485_ VPWR VGND sg13g2_or3_1
X_4654_ _1407_ _1415_ _1417_ _1418_ VPWR VGND sg13g2_or3_1
X_3605_ _0403_ _0411_ _0413_ _0414_ VPWR VGND sg13g2_or3_1
X_4585_ _1355_ _1352_ _1354_ VPWR VGND sg13g2_xnor2_1
X_3536_ _0338_ VPWR _0346_ VGND _0318_ _0339_ sg13g2_o21ai_1
X_6324_ net1102 VGND VPWR net190 mac2.sum_lvl2_ff\[38\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_6255_ net1104 VGND VPWR _0263_ DP_4.matrix\[75\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_5206_ _1950_ _1920_ _1949_ VPWR VGND sg13g2_nand2_1
X_3467_ _0277_ _0276_ _0271_ _0280_ VPWR VGND sg13g2_a21o_1
X_6186_ net1070 VGND VPWR net103 mac1.sum_lvl1_ff\[2\] clknet_leaf_66_clk sg13g2_dfrbpq_1
X_3398_ _2975_ VPWR _2981_ VGND _2952_ _2953_ sg13g2_o21ai_1
X_5137_ _1882_ _1835_ _1881_ VPWR VGND sg13g2_xnor2_1
X_5068_ net824 net875 net828 _1815_ VPWR VGND net873 sg13g2_nand4_1
X_4019_ _0811_ net1016 net949 VPWR VGND sg13g2_nand2_1
XFILLER_25_432 VPWR VGND sg13g2_decap_4
XFILLER_16_78 VPWR VGND sg13g2_fill_1
XFILLER_26_999 VPWR VGND sg13g2_decap_8
XFILLER_21_693 VPWR VGND sg13g2_fill_2
XFILLER_17_911 VPWR VGND sg13g2_decap_8
XFILLER_17_988 VPWR VGND sg13g2_decap_8
XFILLER_43_262 VPWR VGND sg13g2_fill_2
XFILLER_40_980 VPWR VGND sg13g2_decap_8
XFILLER_7_130 VPWR VGND sg13g2_fill_1
Xhold108 mac1.sum_lvl1_ff\[48\] VPWR VGND net148 sg13g2_dlygate4sd3_1
Xhold119 mac1.sum_lvl1_ff\[78\] VPWR VGND net159 sg13g2_dlygate4sd3_1
X_4370_ _1107_ VPWR _1147_ VGND _1105_ _1108_ sg13g2_o21ai_1
X_3321_ _2901_ _2906_ _2907_ VPWR VGND sg13g2_and2_1
X_6040_ net953 _0208_ VPWR VGND sg13g2_buf_1
X_3252_ _2840_ net934 net989 VPWR VGND sg13g2_nand2_1
XFILLER_26_1020 VPWR VGND sg13g2_decap_8
X_3183_ _2773_ _2770_ _2772_ VPWR VGND sg13g2_nand2_1
XFILLER_26_207 VPWR VGND sg13g2_fill_1
XFILLER_23_958 VPWR VGND sg13g2_decap_8
X_5824_ DP_3.Q_range.out_data\[2\] DP_3.I_range.out_data\[2\] _2479_ VPWR VGND sg13g2_xor2_1
XFILLER_22_446 VPWR VGND sg13g2_fill_2
XFILLER_33_1002 VPWR VGND sg13g2_decap_8
X_5755_ _2411_ VPWR _2412_ VGND _2402_ _2410_ sg13g2_o21ai_1
X_4706_ _1468_ net921 DP_4.matrix\[5\] VPWR VGND sg13g2_nand2_1
X_5686_ _2351_ _2352_ net32 VPWR VGND sg13g2_and2_1
X_4637_ _1392_ VPWR _1401_ VGND _1384_ _1393_ sg13g2_o21ai_1
X_4568_ _1339_ net835 net1048 VPWR VGND sg13g2_nand2_1
X_3519_ _0330_ net1029 net983 net1030 net979 VPWR VGND sg13g2_a22oi_1
X_6307_ net1096 VGND VPWR net208 mac1.sum_lvl2_ff\[34\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_4499_ _1271_ _1250_ _1273_ VPWR VGND sg13g2_xor2_1
X_6238_ net1122 VGND VPWR net380 DP_4.matrix\[2\] clknet_leaf_35_clk sg13g2_dfrbpq_1
X_6169_ net1091 VGND VPWR _0196_ DP_2.matrix\[0\] clknet_leaf_62_clk sg13g2_dfrbpq_2
XFILLER_14_958 VPWR VGND sg13g2_decap_8
XFILLER_40_210 VPWR VGND sg13g2_fill_1
XFILLER_43_32 VPWR VGND sg13g2_fill_2
XFILLER_13_468 VPWR VGND sg13g2_fill_1
XFILLER_41_744 VPWR VGND sg13g2_fill_2
XFILLER_41_777 VPWR VGND sg13g2_fill_2
XFILLER_22_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_20_clk clknet_4_5_0_clk clknet_leaf_20_clk VPWR VGND sg13g2_buf_8
XFILLER_1_851 VPWR VGND sg13g2_decap_8
X_3870_ _0646_ VPWR _0666_ VGND _0644_ _0647_ sg13g2_o21ai_1
Xclkbuf_leaf_11_clk clknet_4_6_0_clk clknet_leaf_11_clk VPWR VGND sg13g2_buf_8
X_5540_ _2231_ _2234_ _2237_ _2239_ VPWR VGND sg13g2_or3_1
XFILLER_9_973 VPWR VGND sg13g2_decap_8
X_5471_ VGND VPWR net495 _2185_ _2181_ _2179_ sg13g2_a21oi_2
X_4422_ net844 net842 net892 net1047 _1198_ VPWR VGND sg13g2_and4_1
X_4353_ _1130_ net907 net1043 VPWR VGND sg13g2_nand2_1
X_3304_ _2891_ _2890_ _2863_ VPWR VGND sg13g2_nand2b_1
X_4284_ _1063_ net904 net837 VPWR VGND sg13g2_nand2_1
X_3235_ _2819_ VPWR _2823_ VGND _2776_ _2821_ sg13g2_o21ai_1
X_6023_ net1017 _0183_ VPWR VGND sg13g2_buf_1
X_3166_ net938 net990 net943 _2756_ VPWR VGND net986 sg13g2_nand4_1
X_3097_ net940 net994 net944 _2689_ VPWR VGND net991 sg13g2_nand4_1
XFILLER_23_722 VPWR VGND sg13g2_fill_2
X_3999_ _0768_ VPWR _0792_ VGND _0788_ _0790_ sg13g2_o21ai_1
XFILLER_11_917 VPWR VGND sg13g2_decap_8
X_5807_ VGND VPWR _2463_ _2462_ _2460_ sg13g2_or2_1
X_5738_ DP_1.Q_range.out_data\[3\] DP_1.I_range.out_data\[3\] _2395_ VPWR VGND sg13g2_xor2_1
X_5669_ mac1.total_sum\[4\] mac2.total_sum\[4\] _2339_ VPWR VGND sg13g2_and2_1
XFILLER_2_637 VPWR VGND sg13g2_fill_1
Xhold450 _0060_ VPWR VGND net490 sg13g2_dlygate4sd3_1
Xhold472 mac2.sum_lvl2_ff\[4\] VPWR VGND net512 sg13g2_dlygate4sd3_1
Xhold461 mac2.sum_lvl3_ff\[3\] VPWR VGND net501 sg13g2_dlygate4sd3_1
Xhold494 _2178_ VPWR VGND net534 sg13g2_dlygate4sd3_1
Xhold483 DP_2.matrix\[79\] VPWR VGND net523 sg13g2_dlygate4sd3_1
Xfanout952 DP_2.matrix\[40\] net952 VPWR VGND sg13g2_buf_8
Xfanout941 net543 net941 VPWR VGND sg13g2_buf_1
Xfanout930 net931 net930 VPWR VGND sg13g2_buf_8
Xfanout985 DP_2.matrix\[0\] net985 VPWR VGND sg13g2_buf_1
Xfanout963 net964 net963 VPWR VGND sg13g2_buf_1
Xfanout974 net406 net974 VPWR VGND sg13g2_buf_8
Xfanout996 net997 net996 VPWR VGND sg13g2_buf_8
XFILLER_18_527 VPWR VGND sg13g2_decap_4
XFILLER_13_232 VPWR VGND sg13g2_fill_1
Xclkload17 VPWR clkload17/Y clknet_leaf_51_clk VGND sg13g2_inv_1
XFILLER_10_994 VPWR VGND sg13g2_decap_8
XFILLER_6_965 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_0_clk clknet_4_0_0_clk clknet_leaf_0_clk VPWR VGND sg13g2_buf_8
XFILLER_0_191 VPWR VGND sg13g2_fill_1
X_4971_ _1725_ net908 DP_4.matrix\[8\] VPWR VGND sg13g2_nand2_1
X_3922_ _0683_ VPWR _0717_ VGND _0658_ _0684_ sg13g2_o21ai_1
X_3853_ _0648_ _0649_ _0643_ _0650_ VPWR VGND sg13g2_nand3_1
X_6572_ net1060 VGND VPWR net446 mac2.total_sum\[4\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_3784_ _0587_ _0563_ _0585_ VPWR VGND sg13g2_nand2_1
XFILLER_30_1027 VPWR VGND sg13g2_fill_2
X_5523_ _2223_ VPWR _2225_ VGND _2222_ _2224_ sg13g2_o21ai_1
X_5454_ VGND VPWR _2168_ _2170_ _2171_ _2169_ sg13g2_a21oi_1
X_5385_ _0011_ _2115_ net295 VPWR VGND sg13g2_xnor2_1
X_4405_ _1181_ net901 net834 VPWR VGND sg13g2_nand2_1
X_4336_ _1103_ _1111_ _1113_ _1114_ VPWR VGND sg13g2_or3_1
X_4267_ _1036_ _1044_ _1046_ _1047_ VPWR VGND sg13g2_or3_1
X_6006_ _2629_ net855 net791 VPWR VGND sg13g2_nand2_1
X_3218_ _2795_ VPWR _2807_ VGND _2803_ _2805_ sg13g2_o21ai_1
X_4198_ _0984_ _0981_ _0983_ VPWR VGND sg13g2_xnor2_1
XFILLER_27_302 VPWR VGND sg13g2_fill_2
XFILLER_28_814 VPWR VGND sg13g2_fill_2
X_3149_ _2716_ VPWR _2739_ VGND _2681_ _2714_ sg13g2_o21ai_1
XFILLER_3_902 VPWR VGND sg13g2_decap_8
XFILLER_46_1001 VPWR VGND sg13g2_decap_8
XFILLER_3_979 VPWR VGND sg13g2_decap_8
Xhold280 _2144_ VPWR VGND net320 sg13g2_dlygate4sd3_1
XFILLER_49_31 VPWR VGND sg13g2_fill_2
Xhold291 mac1.sum_lvl3_ff\[14\] VPWR VGND net331 sg13g2_dlygate4sd3_1
XFILLER_1_27 VPWR VGND sg13g2_fill_2
Xfanout793 _2475_ net793 VPWR VGND sg13g2_buf_8
XFILLER_33_349 VPWR VGND sg13g2_fill_1
X_5170_ _1915_ _1913_ _1914_ VPWR VGND sg13g2_nand2_1
X_4121_ _0910_ net951 net1056 VPWR VGND sg13g2_nand2_1
X_4052_ VGND VPWR _0808_ _0814_ _0843_ _0816_ sg13g2_a21oi_1
Xinput4 ui_in[3] net4 VPWR VGND sg13g2_buf_1
X_4954_ _1709_ net851 net1050 VPWR VGND sg13g2_nand2_1
XFILLER_40_809 VPWR VGND sg13g2_fill_2
X_3905_ net962 net959 net1011 net1009 _0700_ VPWR VGND sg13g2_and4_1
X_4885_ _1643_ _1622_ _1642_ VPWR VGND sg13g2_xnor2_1
X_3836_ _0634_ _0626_ _0633_ VPWR VGND sg13g2_nand2_1
X_3767_ _0571_ net969 net1026 VPWR VGND sg13g2_nand2_1
X_6555_ net1096 VGND VPWR net434 mac2.sum_lvl3_ff\[3\] clknet_leaf_29_clk sg13g2_dfrbpq_1
X_5506_ _2210_ VPWR _2213_ VGND _2209_ _2211_ sg13g2_o21ai_1
X_3698_ VGND VPWR _0504_ _0505_ _0470_ _0430_ sg13g2_a21oi_2
X_6486_ net1122 VGND VPWR net169 mac2.sum_lvl1_ff\[2\] clknet_leaf_26_clk sg13g2_dfrbpq_1
X_5437_ _2158_ net292 net265 VPWR VGND sg13g2_nand2_1
X_5368_ mac1.sum_lvl2_ff\[1\] mac1.sum_lvl2_ff\[20\] _2105_ VPWR VGND sg13g2_xor2_1
XFILLER_0_938 VPWR VGND sg13g2_decap_8
X_4319_ _1097_ net903 net837 VPWR VGND sg13g2_nand2_1
X_5299_ VGND VPWR _2040_ _2039_ _2027_ sg13g2_or2_1
XFILLER_19_45 VPWR VGND sg13g2_fill_1
XFILLER_15_316 VPWR VGND sg13g2_fill_1
XFILLER_16_839 VPWR VGND sg13g2_decap_8
XFILLER_11_544 VPWR VGND sg13g2_fill_1
XFILLER_4_0 VPWR VGND sg13g2_fill_2
XFILLER_18_165 VPWR VGND sg13g2_fill_1
XFILLER_18_198 VPWR VGND sg13g2_fill_1
XFILLER_33_135 VPWR VGND sg13g2_fill_2
XFILLER_34_658 VPWR VGND sg13g2_fill_2
XFILLER_15_883 VPWR VGND sg13g2_decap_8
X_4670_ _1416_ VPWR _1433_ VGND _1407_ _1417_ sg13g2_o21ai_1
X_3621_ _0382_ _0383_ _0427_ _0428_ _0430_ VPWR VGND sg13g2_and4_1
X_3552_ _0362_ net976 net1030 VPWR VGND sg13g2_nand2_1
X_6340_ net1062 VGND VPWR net91 mac1.sum_lvl1_ff\[72\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_3483_ _0295_ net976 net1035 VPWR VGND sg13g2_nand2_1
X_6271_ net1098 VGND VPWR net63 mac1.sum_lvl1_ff\[47\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_5222_ _1965_ _1924_ _1963_ VPWR VGND sg13g2_xnor2_1
X_5153_ _1895_ _1896_ _1890_ _1898_ VPWR VGND sg13g2_nand3_1
X_4104_ _0893_ _0890_ _0894_ VPWR VGND sg13g2_xor2_1
X_5084_ _1797_ VPWR _1831_ VGND _1772_ _1798_ sg13g2_o21ai_1
X_4035_ net960 net956 net1005 net1057 _0827_ VPWR VGND sg13g2_and4_1
XFILLER_25_603 VPWR VGND sg13g2_decap_4
X_5986_ _2615_ VPWR _0226_ VGND net792 _2616_ sg13g2_o21ai_1
X_4937_ _1693_ _1653_ _1691_ VPWR VGND sg13g2_xnor2_1
XFILLER_36_1022 VPWR VGND sg13g2_decap_8
X_4868_ VGND VPWR _1626_ _1625_ _1601_ sg13g2_or2_1
X_3819_ _0618_ net1023 net956 VPWR VGND sg13g2_nand2_1
X_4799_ _1559_ _1549_ _1557_ VPWR VGND sg13g2_xnor2_1
X_6538_ net1136 VGND VPWR net180 mac2.sum_lvl2_ff\[25\] clknet_leaf_43_clk sg13g2_dfrbpq_1
X_6469_ net1100 VGND VPWR _0090_ mac2.products_ff\[137\] clknet_leaf_23_clk sg13g2_dfrbpq_1
XFILLER_29_975 VPWR VGND sg13g2_decap_8
XFILLER_28_463 VPWR VGND sg13g2_decap_8
XFILLER_46_87 VPWR VGND sg13g2_fill_1
XFILLER_44_978 VPWR VGND sg13g2_decap_8
XFILLER_43_455 VPWR VGND sg13g2_fill_1
XFILLER_12_820 VPWR VGND sg13g2_decap_8
XFILLER_12_864 VPWR VGND sg13g2_decap_8
XFILLER_8_857 VPWR VGND sg13g2_decap_8
XFILLER_7_367 VPWR VGND sg13g2_fill_2
XFILLER_39_717 VPWR VGND sg13g2_decap_8
XFILLER_4_1020 VPWR VGND sg13g2_decap_8
X_5840_ _2495_ _2476_ net806 VPWR VGND sg13g2_nand2_1
X_5771_ VGND VPWR _2428_ _2427_ _2425_ sg13g2_or2_1
XFILLER_21_105 VPWR VGND sg13g2_decap_4
XFILLER_21_127 VPWR VGND sg13g2_decap_8
X_4722_ VGND VPWR _1480_ _1481_ _1484_ _1475_ sg13g2_a21oi_1
XFILLER_30_694 VPWR VGND sg13g2_fill_2
X_4653_ VGND VPWR _1413_ _1414_ _1417_ _1408_ sg13g2_a21oi_1
X_3604_ VGND VPWR _0409_ _0410_ _0413_ _0404_ sg13g2_a21oi_1
X_4584_ _1354_ _1338_ _1353_ VPWR VGND sg13g2_xnor2_1
X_3535_ _0345_ _0344_ _0112_ VPWR VGND sg13g2_xor2_1
X_6323_ net1089 VGND VPWR net79 mac1.sum_lvl2_ff\[53\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_3466_ VGND VPWR _0276_ _0277_ _0279_ _0271_ sg13g2_a21oi_1
X_6254_ net1101 VGND VPWR _0262_ DP_4.matrix\[74\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_5205_ _1948_ _1931_ _1949_ VPWR VGND sg13g2_xor2_1
X_6185_ net1090 VGND VPWR _0207_ DP_2.matrix\[39\] clknet_leaf_64_clk sg13g2_dfrbpq_1
X_3397_ VPWR _2980_ _2979_ VGND sg13g2_inv_1
X_5136_ _1881_ _1872_ _1879_ VPWR VGND sg13g2_xnor2_1
X_5067_ net829 net824 net875 net873 _1814_ VPWR VGND sg13g2_and4_1
X_4018_ _0810_ net1016 net947 VPWR VGND sg13g2_nand2_1
XFILLER_26_978 VPWR VGND sg13g2_decap_8
X_5969_ _2605_ _2493_ _2498_ VPWR VGND sg13g2_xnor2_1
XFILLER_32_89 VPWR VGND sg13g2_fill_1
XFILLER_5_849 VPWR VGND sg13g2_decap_8
XFILLER_48_503 VPWR VGND sg13g2_fill_1
XFILLER_17_967 VPWR VGND sg13g2_decap_8
XFILLER_16_488 VPWR VGND sg13g2_fill_2
XFILLER_16_499 VPWR VGND sg13g2_decap_8
XFILLER_31_425 VPWR VGND sg13g2_decap_4
XFILLER_32_926 VPWR VGND sg13g2_fill_1
Xhold109 mac1.products_ff\[6\] VPWR VGND net149 sg13g2_dlygate4sd3_1
X_3320_ _2905_ _2902_ _2906_ VPWR VGND sg13g2_xor2_1
X_3251_ _2839_ net994 net930 VPWR VGND sg13g2_nand2_1
X_3182_ _2769_ _2768_ _2738_ _2772_ VPWR VGND sg13g2_a21o_1
XFILLER_23_937 VPWR VGND sg13g2_decap_8
XFILLER_34_274 VPWR VGND sg13g2_fill_2
X_5823_ _2478_ DP_3.I_range.out_data\[2\] DP_3.Q_range.out_data\[2\] VPWR VGND sg13g2_xnor2_1
X_5754_ net808 _2402_ net997 _2411_ VPWR VGND sg13g2_nand3_1
X_5685_ _2344_ _2347_ _2350_ _2352_ VPWR VGND sg13g2_or3_1
XFILLER_31_992 VPWR VGND sg13g2_decap_8
X_4705_ _1449_ _1439_ _1447_ _1467_ VPWR VGND sg13g2_a21o_1
X_4636_ _1399_ _1379_ _0088_ VPWR VGND sg13g2_xor2_1
XFILLER_2_819 VPWR VGND sg13g2_decap_8
X_6306_ net1096 VGND VPWR net188 mac1.sum_lvl2_ff\[33\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_4567_ _1338_ net833 net1048 VPWR VGND sg13g2_nand2_1
X_3518_ net979 net1030 net983 _0329_ VPWR VGND net1029 sg13g2_nand4_1
X_4498_ _1271_ _1250_ _1272_ VPWR VGND sg13g2_nor2b_1
X_6237_ net1105 VGND VPWR net508 DP_4.matrix\[1\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_3449_ _3027_ _3018_ _3025_ VPWR VGND sg13g2_xnor2_1
X_6168_ net1119 VGND VPWR _0097_ mac1.products_ff\[148\] clknet_leaf_47_clk sg13g2_dfrbpq_2
X_5119_ VGND VPWR _1862_ _1863_ _1865_ _1832_ sg13g2_a21oi_1
X_6099_ net1121 VGND VPWR _0107_ mac1.products_ff\[11\] clknet_leaf_31_clk sg13g2_dfrbpq_1
XFILLER_14_937 VPWR VGND sg13g2_decap_8
XFILLER_43_11 VPWR VGND sg13g2_fill_1
XFILLER_13_458 VPWR VGND sg13g2_fill_1
XFILLER_5_624 VPWR VGND sg13g2_fill_1
XFILLER_49_801 VPWR VGND sg13g2_fill_1
XFILLER_1_830 VPWR VGND sg13g2_decap_8
XFILLER_49_856 VPWR VGND sg13g2_decap_4
XFILLER_49_889 VPWR VGND sg13g2_decap_8
XFILLER_49_878 VPWR VGND sg13g2_fill_2
XFILLER_1_1012 VPWR VGND sg13g2_decap_8
XFILLER_17_797 VPWR VGND sg13g2_decap_8
XFILLER_17_1009 VPWR VGND sg13g2_decap_8
XFILLER_20_929 VPWR VGND sg13g2_decap_8
XFILLER_9_952 VPWR VGND sg13g2_decap_8
X_5470_ _2184_ mac1.sum_lvl3_ff\[28\] net494 VPWR VGND sg13g2_xnor2_1
XFILLER_8_484 VPWR VGND sg13g2_fill_2
X_4421_ _1197_ net843 net1047 VPWR VGND sg13g2_nand2_1
X_4352_ _1100_ VPWR _1129_ VGND _1097_ _1101_ sg13g2_o21ai_1
X_3303_ _2888_ _2864_ _2890_ VPWR VGND sg13g2_xor2_1
X_4283_ _1045_ VPWR _1062_ VGND _1036_ _1046_ sg13g2_o21ai_1
X_3234_ _2821_ _2776_ _0103_ VPWR VGND sg13g2_xor2_1
X_6022_ net1018 _0182_ VPWR VGND sg13g2_buf_1
X_3165_ net943 net938 DP_1.matrix\[78\] net986 _2755_ VPWR VGND sg13g2_and4_1
XFILLER_27_517 VPWR VGND sg13g2_decap_4
X_3096_ net945 net940 net994 net993 _2688_ VPWR VGND sg13g2_and4_1
X_3998_ _0768_ _0788_ _0790_ _0791_ VPWR VGND sg13g2_or3_1
X_5806_ _2462_ net799 _2461_ net801 net404 VPWR VGND sg13g2_a22oi_1
X_5737_ net1059 net786 _2394_ VPWR VGND sg13g2_nor2_1
X_5668_ _2336_ VPWR _2338_ VGND _2335_ _2337_ sg13g2_o21ai_1
X_4619_ VPWR _1384_ _1383_ VGND sg13g2_inv_1
X_5599_ VGND VPWR _2281_ _2283_ _2284_ _2282_ sg13g2_a21oi_1
Xhold440 mac2.sum_lvl3_ff\[20\] VPWR VGND net480 sg13g2_dlygate4sd3_1
Xhold451 DP_2.matrix\[72\] VPWR VGND net491 sg13g2_dlygate4sd3_1
Xhold462 _2280_ VPWR VGND net502 sg13g2_dlygate4sd3_1
Xhold495 mac1.sum_lvl2_ff\[7\] VPWR VGND net535 sg13g2_dlygate4sd3_1
Xhold484 DP_2.matrix\[37\] VPWR VGND net524 sg13g2_dlygate4sd3_1
Xhold473 _2227_ VPWR VGND net513 sg13g2_dlygate4sd3_1
Xfanout942 DP_2.matrix\[73\] net942 VPWR VGND sg13g2_buf_8
Xfanout931 net311 net931 VPWR VGND sg13g2_buf_8
Xfanout920 net435 net920 VPWR VGND sg13g2_buf_8
Xfanout953 net452 net953 VPWR VGND sg13g2_buf_1
Xfanout964 net965 net964 VPWR VGND sg13g2_buf_1
Xfanout975 DP_2.matrix\[3\] net975 VPWR VGND sg13g2_buf_1
Xfanout986 net987 net986 VPWR VGND sg13g2_buf_2
Xfanout997 net314 net997 VPWR VGND sg13g2_buf_8
XFILLER_9_204 VPWR VGND sg13g2_decap_8
XFILLER_10_973 VPWR VGND sg13g2_decap_8
XFILLER_6_944 VPWR VGND sg13g2_decap_8
Xclkload18 clknet_leaf_50_clk clkload18/Y VPWR VGND sg13g2_inv_4
XFILLER_48_8 VPWR VGND sg13g2_fill_2
XFILLER_48_174 VPWR VGND sg13g2_fill_1
XFILLER_37_837 VPWR VGND sg13g2_fill_1
X_4970_ _1712_ VPWR _1724_ VGND _1684_ _1710_ sg13g2_o21ai_1
XFILLER_17_583 VPWR VGND sg13g2_fill_2
X_3921_ _0716_ _0686_ _0714_ VPWR VGND sg13g2_xnor2_1
X_3852_ _0644_ VPWR _0649_ VGND _0645_ _0647_ sg13g2_o21ai_1
X_6571_ net1060 VGND VPWR net503 mac2.total_sum\[3\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_30_1006 VPWR VGND sg13g2_decap_8
X_3783_ _0109_ _0585_ _0586_ VPWR VGND sg13g2_xnor2_1
X_5522_ net433 _2222_ _0041_ VPWR VGND sg13g2_xor2_1
X_5453_ _2170_ _2168_ _0026_ VPWR VGND sg13g2_xor2_1
X_5384_ net294 mac1.sum_lvl2_ff\[24\] _2117_ VPWR VGND sg13g2_xor2_1
X_4404_ _1180_ net904 net1043 VPWR VGND sg13g2_nand2_1
X_4335_ VGND VPWR _1109_ _1110_ _1113_ _1104_ sg13g2_a21oi_1
XFILLER_8_1018 VPWR VGND sg13g2_decap_8
X_4266_ VGND VPWR _1042_ _1043_ _1046_ _1037_ sg13g2_a21oi_1
X_6005_ _2627_ VPWR _0249_ VGND net792 _2628_ sg13g2_o21ai_1
X_3217_ _2795_ _2803_ _2805_ _2806_ VPWR VGND sg13g2_or3_1
X_4197_ _0983_ _0967_ _0982_ VPWR VGND sg13g2_xnor2_1
X_3148_ _2730_ VPWR _2738_ VGND _2710_ _2731_ sg13g2_o21ai_1
XFILLER_27_369 VPWR VGND sg13g2_fill_2
X_3079_ _2669_ _2668_ _2663_ _2672_ VPWR VGND sg13g2_a21o_1
XFILLER_3_958 VPWR VGND sg13g2_decap_8
Xhold270 DP_3.matrix\[73\] VPWR VGND net310 sg13g2_dlygate4sd3_1
Xhold281 _0003_ VPWR VGND net321 sg13g2_dlygate4sd3_1
Xhold292 _2212_ VPWR VGND net332 sg13g2_dlygate4sd3_1
XFILLER_49_87 VPWR VGND sg13g2_fill_2
XFILLER_49_76 VPWR VGND sg13g2_fill_1
Xfanout794 net796 net794 VPWR VGND sg13g2_buf_8
Xfanout783 net788 net783 VPWR VGND sg13g2_buf_2
XFILLER_45_166 VPWR VGND sg13g2_fill_2
XFILLER_2_980 VPWR VGND sg13g2_decap_8
X_4120_ _0909_ net1056 net952 net1007 net951 VPWR VGND sg13g2_a22oi_1
X_4051_ _0842_ _0803_ _0126_ VPWR VGND sg13g2_xor2_1
Xinput5 ui_in[4] net5 VPWR VGND sg13g2_buf_1
XFILLER_37_634 VPWR VGND sg13g2_fill_1
XFILLER_36_122 VPWR VGND sg13g2_fill_2
X_4953_ _1708_ net912 DP_4.matrix\[8\] VPWR VGND sg13g2_nand2_1
X_3904_ _0699_ net956 net1013 VPWR VGND sg13g2_nand2_1
X_4884_ _1642_ _1631_ _1641_ VPWR VGND sg13g2_xnor2_1
X_3835_ _0631_ _0632_ _0633_ VPWR VGND sg13g2_nor2b_1
X_3766_ _0570_ net1026 net966 VPWR VGND sg13g2_nand2_1
X_6554_ net1101 VGND VPWR net352 mac2.sum_lvl3_ff\[2\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_5505_ _0021_ _2209_ net332 VPWR VGND sg13g2_xnor2_1
X_6485_ net1105 VGND VPWR net220 mac2.sum_lvl1_ff\[1\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_5436_ net267 mac1.sum_lvl2_ff\[19\] _0000_ VPWR VGND sg13g2_xor2_1
X_3697_ VGND VPWR _0427_ _0469_ _0504_ _0468_ sg13g2_a21oi_1
X_5367_ mac1.sum_lvl2_ff\[20\] mac1.sum_lvl2_ff\[1\] _2104_ VPWR VGND sg13g2_nor2_1
XFILLER_0_917 VPWR VGND sg13g2_decap_8
X_5298_ _2037_ _2028_ _2039_ VPWR VGND sg13g2_xor2_1
X_4318_ _1078_ _1068_ _1076_ _1096_ VPWR VGND sg13g2_a21o_1
X_4249_ _1028_ _1008_ _0083_ VPWR VGND sg13g2_xor2_1
XFILLER_16_818 VPWR VGND sg13g2_decap_8
XFILLER_42_136 VPWR VGND sg13g2_fill_1
XFILLER_11_512 VPWR VGND sg13g2_decap_4
XFILLER_18_133 VPWR VGND sg13g2_fill_1
XFILLER_19_634 VPWR VGND sg13g2_fill_1
XFILLER_20_1027 VPWR VGND sg13g2_fill_2
XFILLER_47_987 VPWR VGND sg13g2_decap_8
XFILLER_33_125 VPWR VGND sg13g2_fill_1
X_3620_ _0429_ _0427_ _0428_ VPWR VGND sg13g2_nand2_1
X_3551_ _0329_ VPWR _0361_ VGND _0327_ _0330_ sg13g2_o21ai_1
X_3482_ _0274_ VPWR _0294_ VGND _0272_ _0275_ sg13g2_o21ai_1
X_6270_ net1089 VGND VPWR net124 mac1.sum_lvl1_ff\[46\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_5221_ VGND VPWR _1964_ _1962_ _1925_ sg13g2_or2_1
X_5152_ _1897_ _1890_ _1895_ _1896_ VPWR VGND sg13g2_and3_1
X_4103_ _0893_ _0848_ _0891_ VPWR VGND sg13g2_xnor2_1
X_5083_ _1830_ _1800_ _1828_ VPWR VGND sg13g2_xnor2_1
X_4034_ _0826_ net956 net1056 VPWR VGND sg13g2_nand2_1
X_5985_ _2515_ _2511_ _2616_ VPWR VGND sg13g2_xor2_1
XFILLER_36_1001 VPWR VGND sg13g2_decap_8
X_4936_ _1653_ _1691_ _1692_ VPWR VGND sg13g2_nor2_1
XFILLER_40_629 VPWR VGND sg13g2_fill_1
X_4867_ _1625_ net860 net1049 VPWR VGND sg13g2_nand2_1
X_3818_ _0616_ net449 _0075_ VPWR VGND sg13g2_nor2_1
X_6537_ net1135 VGND VPWR net231 mac2.sum_lvl2_ff\[24\] clknet_leaf_47_clk sg13g2_dfrbpq_2
X_4798_ _1549_ _1557_ _1558_ VPWR VGND sg13g2_nor2_1
X_3749_ VGND VPWR _0554_ _0553_ _0541_ sg13g2_or2_1
X_6468_ net1100 VGND VPWR _0089_ mac2.products_ff\[136\] clknet_leaf_24_clk sg13g2_dfrbpq_1
XFILLER_0_714 VPWR VGND sg13g2_fill_2
X_6399_ net1118 VGND VPWR net368 mac1.sum_lvl3_ff\[11\] clknet_leaf_47_clk sg13g2_dfrbpq_1
X_5419_ _2134_ _2139_ _2145_ VPWR VGND sg13g2_nor2_1
XFILLER_28_442 VPWR VGND sg13g2_decap_8
XFILLER_29_954 VPWR VGND sg13g2_decap_8
XFILLER_15_169 VPWR VGND sg13g2_fill_2
XFILLER_8_814 VPWR VGND sg13g2_decap_4
XFILLER_12_843 VPWR VGND sg13g2_decap_8
XFILLER_11_386 VPWR VGND sg13g2_fill_1
XFILLER_7_379 VPWR VGND sg13g2_fill_2
XFILLER_3_596 VPWR VGND sg13g2_fill_2
Xclkbuf_4_9_0_clk clknet_0_clk clknet_4_9_0_clk VPWR VGND sg13g2_buf_8
XFILLER_47_762 VPWR VGND sg13g2_fill_1
X_5770_ _2427_ net800 _2426_ net802 DP_1.matrix\[76\] VPWR VGND sg13g2_a22oi_1
XFILLER_15_681 VPWR VGND sg13g2_fill_2
X_4721_ _1480_ _1481_ _1475_ _1483_ VPWR VGND sg13g2_nand3_1
X_4652_ _1413_ _1414_ _1408_ _1416_ VPWR VGND sg13g2_nand3_1
X_3603_ _0409_ _0410_ _0404_ _0412_ VPWR VGND sg13g2_nand3_1
X_4583_ _1353_ net893 net1043 VPWR VGND sg13g2_nand2_1
XFILLER_7_891 VPWR VGND sg13g2_decap_8
X_3534_ _0311_ VPWR _0345_ VGND _0286_ _0312_ sg13g2_o21ai_1
X_6322_ net1073 VGND VPWR net229 mac1.sum_lvl2_ff\[52\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_3465_ _0276_ _0277_ _0271_ _0278_ VPWR VGND sg13g2_nand3_1
X_6253_ net1085 VGND VPWR _0261_ DP_4.matrix\[73\] clknet_leaf_24_clk sg13g2_dfrbpq_1
X_5204_ _1948_ _1932_ _1946_ VPWR VGND sg13g2_xnor2_1
X_6184_ net1090 VGND VPWR _0206_ DP_2.matrix\[38\] clknet_leaf_63_clk sg13g2_dfrbpq_1
X_3396_ _2979_ _2955_ _2977_ VPWR VGND sg13g2_nand2_1
X_5135_ _1880_ _1872_ _1879_ VPWR VGND sg13g2_nand2_1
X_5066_ _1813_ net822 net877 VPWR VGND sg13g2_nand2_1
X_4017_ _0809_ net1021 net1052 VPWR VGND sg13g2_nand2_1
XFILLER_26_957 VPWR VGND sg13g2_decap_8
X_5968_ _0220_ net924 net792 VPWR VGND sg13g2_xnor2_1
XFILLER_34_990 VPWR VGND sg13g2_decap_8
X_4919_ _1674_ _1675_ _1676_ VPWR VGND sg13g2_nor2_1
X_5899_ _2553_ net269 net797 VPWR VGND sg13g2_nand2_1
XFILLER_20_172 VPWR VGND sg13g2_decap_4
XFILLER_21_695 VPWR VGND sg13g2_fill_1
XFILLER_5_828 VPWR VGND sg13g2_decap_8
XFILLER_10_1015 VPWR VGND sg13g2_decap_8
XFILLER_48_537 VPWR VGND sg13g2_fill_1
XFILLER_29_762 VPWR VGND sg13g2_fill_1
XFILLER_17_946 VPWR VGND sg13g2_decap_8
XFILLER_8_699 VPWR VGND sg13g2_fill_2
XFILLER_4_894 VPWR VGND sg13g2_decap_8
X_3250_ _2804_ VPWR _2838_ VGND _2795_ _2805_ sg13g2_o21ai_1
X_3181_ VGND VPWR _2768_ _2769_ _2771_ _2738_ sg13g2_a21oi_1
XFILLER_23_916 VPWR VGND sg13g2_decap_8
X_5822_ DP_3.Q_range.out_data\[2\] DP_3.I_range.out_data\[2\] _2477_ VPWR VGND sg13g2_nor2b_1
X_5753_ VGND VPWR net1017 net809 _2410_ _2409_ sg13g2_a21oi_1
XFILLER_31_971 VPWR VGND sg13g2_decap_8
X_4704_ _1466_ _1461_ _1464_ VPWR VGND sg13g2_xnor2_1
X_5684_ _2350_ VPWR _2351_ VGND _2344_ _2347_ sg13g2_o21ai_1
X_4635_ VGND VPWR _1400_ _1399_ _1379_ sg13g2_or2_1
X_4566_ _1337_ net895 DP_4.matrix\[44\] VPWR VGND sg13g2_nand2_1
X_3517_ net983 net979 net1030 net1029 _0328_ VPWR VGND sg13g2_and4_1
X_6305_ net1097 VGND VPWR net99 mac1.sum_lvl2_ff\[32\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_4497_ _1271_ _1251_ _1270_ VPWR VGND sg13g2_xnor2_1
X_3448_ _3026_ _3018_ _3025_ VPWR VGND sg13g2_nand2_1
X_6236_ net1127 VGND VPWR net375 DP_4.matrix\[0\] clknet_leaf_37_clk sg13g2_dfrbpq_2
X_3379_ _2963_ net928 net988 VPWR VGND sg13g2_nand2_1
X_6167_ net1135 VGND VPWR _0195_ DP_1.matrix\[79\] clknet_leaf_48_clk sg13g2_dfrbpq_2
X_5118_ _1862_ _1863_ _1832_ _1864_ VPWR VGND sg13g2_nand3_1
XFILLER_40_1008 VPWR VGND sg13g2_decap_8
X_6098_ net1121 VGND VPWR _0106_ mac1.products_ff\[10\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_5049_ _1794_ _1795_ _1770_ _1797_ VPWR VGND sg13g2_nand3_1
XFILLER_14_916 VPWR VGND sg13g2_decap_8
XFILLER_41_746 VPWR VGND sg13g2_fill_1
XFILLER_43_34 VPWR VGND sg13g2_fill_1
XFILLER_41_779 VPWR VGND sg13g2_fill_1
XFILLER_49_1022 VPWR VGND sg13g2_decap_8
XFILLER_1_886 VPWR VGND sg13g2_decap_8
XFILLER_44_562 VPWR VGND sg13g2_fill_2
XFILLER_20_908 VPWR VGND sg13g2_decap_8
XFILLER_9_931 VPWR VGND sg13g2_decap_8
XFILLER_8_430 VPWR VGND sg13g2_fill_2
XFILLER_13_982 VPWR VGND sg13g2_decap_8
X_4420_ _1150_ VPWR _1196_ VGND _1148_ _1151_ sg13g2_o21ai_1
X_4351_ _1117_ VPWR _1128_ VGND _1095_ _1118_ sg13g2_o21ai_1
X_3302_ _2889_ _2864_ _2888_ VPWR VGND sg13g2_nand2_1
X_4282_ _1059_ _1058_ _1061_ VPWR VGND sg13g2_xor2_1
X_3233_ _2774_ _2775_ _2819_ _2820_ _2822_ VPWR VGND sg13g2_and4_1
X_6021_ net1021 _0181_ VPWR VGND sg13g2_buf_1
X_3164_ _2754_ net936 net991 VPWR VGND sg13g2_nand2_1
X_3095_ _2687_ net936 net997 VPWR VGND sg13g2_nand2_1
XFILLER_23_702 VPWR VGND sg13g2_fill_1
X_5805_ net972 net953 net810 _2461_ VPWR VGND sg13g2_mux2_1
X_3997_ VGND VPWR _0786_ _0787_ _0790_ _0769_ sg13g2_a21oi_1
X_5736_ DP_1.I_range.out_data\[2\] DP_1.Q_range.out_data\[2\] _2385_ _2393_ VGND VPWR
+ _2392_ sg13g2_nor4_2
X_5667_ _2337_ _2335_ net28 VPWR VGND sg13g2_xor2_1
X_4618_ _1380_ _1382_ _1383_ VPWR VGND sg13g2_nor2_1
X_5598_ net445 _2281_ _0058_ VPWR VGND sg13g2_xor2_1
Xhold452 DP_1.matrix\[74\] VPWR VGND net492 sg13g2_dlygate4sd3_1
Xhold441 _0055_ VPWR VGND net481 sg13g2_dlygate4sd3_1
Xhold463 _0057_ VPWR VGND net503 sg13g2_dlygate4sd3_1
Xhold430 _2230_ VPWR VGND net470 sg13g2_dlygate4sd3_1
X_4549_ _1319_ _1281_ _1321_ VPWR VGND sg13g2_xor2_1
Xhold496 _2124_ VPWR VGND net536 sg13g2_dlygate4sd3_1
Xhold485 mac1.sum_lvl3_ff\[30\] VPWR VGND net525 sg13g2_dlygate4sd3_1
Xhold474 _0042_ VPWR VGND net514 sg13g2_dlygate4sd3_1
Xfanout910 net451 net910 VPWR VGND sg13g2_buf_2
Xfanout943 net944 net943 VPWR VGND sg13g2_buf_8
Xfanout932 net933 net932 VPWR VGND sg13g2_buf_8
X_6219_ net1098 VGND VPWR net151 mac1.sum_lvl1_ff\[13\] clknet_leaf_29_clk sg13g2_dfrbpq_1
Xfanout921 DP_3.matrix\[2\] net921 VPWR VGND sg13g2_buf_8
Xfanout965 net363 net965 VPWR VGND sg13g2_buf_8
Xfanout954 DP_2.matrix\[39\] net954 VPWR VGND sg13g2_buf_8
Xfanout976 net440 net976 VPWR VGND sg13g2_buf_8
Xfanout998 net999 net998 VPWR VGND sg13g2_buf_8
Xfanout987 net988 net987 VPWR VGND sg13g2_buf_1
XFILLER_45_315 VPWR VGND sg13g2_fill_2
XFILLER_10_952 VPWR VGND sg13g2_decap_8
Xclkload19 clknet_leaf_37_clk clkload19/Y VPWR VGND sg13g2_inv_4
XFILLER_6_923 VPWR VGND sg13g2_decap_8
XFILLER_23_1014 VPWR VGND sg13g2_decap_8
XFILLER_49_665 VPWR VGND sg13g2_fill_2
XFILLER_37_805 VPWR VGND sg13g2_fill_2
XFILLER_37_816 VPWR VGND sg13g2_fill_1
XFILLER_48_164 VPWR VGND sg13g2_fill_2
X_3920_ _0714_ _0686_ _0715_ VPWR VGND sg13g2_nor2b_1
X_3851_ _0644_ _0645_ _0647_ _0648_ VPWR VGND sg13g2_or3_1
XFILLER_32_565 VPWR VGND sg13g2_fill_2
X_6570_ net1061 VGND VPWR net500 mac2.total_sum\[2\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_3782_ VGND VPWR _0563_ _0566_ _0586_ _0562_ sg13g2_a21oi_1
XFILLER_9_772 VPWR VGND sg13g2_fill_2
X_5521_ _2224_ mac2.sum_lvl2_ff\[22\] net432 VPWR VGND sg13g2_xnor2_1
X_5452_ net551 mac1.sum_lvl3_ff\[24\] _2170_ VPWR VGND sg13g2_xor2_1
X_5383_ mac1.sum_lvl2_ff\[24\] net294 _2116_ VPWR VGND sg13g2_nor2_1
X_4403_ _1144_ VPWR _1179_ VGND _1141_ _1145_ sg13g2_o21ai_1
X_4334_ _1109_ _1110_ _1104_ _1112_ VPWR VGND sg13g2_nand3_1
X_6004_ _2557_ _2533_ _2628_ VPWR VGND sg13g2_xor2_1
X_4265_ _1042_ _1043_ _1037_ _1045_ VPWR VGND sg13g2_nand3_1
X_4196_ _0982_ net1007 net1052 VPWR VGND sg13g2_nand2_1
X_3216_ VGND VPWR _2801_ _2802_ _2805_ _2796_ sg13g2_a21oi_1
X_3147_ _2737_ _2736_ _0101_ VPWR VGND sg13g2_xor2_1
XFILLER_28_838 VPWR VGND sg13g2_decap_4
X_3078_ VGND VPWR _2668_ _2669_ _2671_ _2663_ sg13g2_a21oi_1
XFILLER_39_1021 VPWR VGND sg13g2_decap_8
XFILLER_10_204 VPWR VGND sg13g2_fill_2
XFILLER_10_237 VPWR VGND sg13g2_fill_1
X_5719_ _2379_ mac1.total_sum\[14\] mac2.total_sum\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_3_937 VPWR VGND sg13g2_decap_8
Xhold260 DP_2.matrix\[43\] VPWR VGND net300 sg13g2_dlygate4sd3_1
Xhold271 DP_2.matrix\[77\] VPWR VGND net311 sg13g2_dlygate4sd3_1
XFILLER_49_44 VPWR VGND sg13g2_fill_1
XFILLER_49_33 VPWR VGND sg13g2_fill_1
Xhold282 DP_2.matrix\[0\] VPWR VGND net322 sg13g2_dlygate4sd3_1
Xhold293 _0021_ VPWR VGND net333 sg13g2_dlygate4sd3_1
Xfanout784 net785 net784 VPWR VGND sg13g2_buf_1
XFILLER_1_29 VPWR VGND sg13g2_fill_1
Xfanout795 _2481_ net795 VPWR VGND sg13g2_buf_8
XFILLER_30_90 VPWR VGND sg13g2_fill_1
X_4050_ _0840_ _0841_ _0842_ VPWR VGND sg13g2_nor2b_2
XFILLER_49_484 VPWR VGND sg13g2_fill_1
Xinput6 ui_in[5] net6 VPWR VGND sg13g2_buf_1
X_4952_ _1687_ VPWR _1707_ VGND _1659_ _1685_ sg13g2_o21ai_1
XFILLER_18_882 VPWR VGND sg13g2_decap_8
XFILLER_33_830 VPWR VGND sg13g2_decap_4
X_4883_ _1641_ _1632_ _1639_ VPWR VGND sg13g2_xnor2_1
X_3903_ _0669_ VPWR _0698_ VGND _0667_ _0670_ sg13g2_o21ai_1
X_3834_ _0627_ VPWR _0632_ VGND _0628_ _0630_ sg13g2_o21ai_1
XFILLER_20_557 VPWR VGND sg13g2_fill_2
X_3765_ _0569_ net1031 DP_2.matrix\[8\] VPWR VGND sg13g2_nand2_1
X_6553_ net1101 VGND VPWR net309 mac2.sum_lvl3_ff\[1\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_3696_ _0503_ _0502_ _0501_ VPWR VGND sg13g2_nand2b_1
X_5504_ net331 mac1.sum_lvl3_ff\[34\] _2212_ VPWR VGND sg13g2_xor2_1
X_6484_ net1103 VGND VPWR net185 mac2.sum_lvl1_ff\[0\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_5435_ _0006_ _2156_ net285 VPWR VGND sg13g2_xnor2_1
X_5366_ _2103_ mac1.sum_lvl2_ff\[20\] mac1.sum_lvl2_ff\[1\] VPWR VGND sg13g2_nand2_1
X_5297_ _2037_ _2028_ _2038_ VPWR VGND sg13g2_nor2b_1
X_4317_ _1095_ _1090_ _1093_ VPWR VGND sg13g2_xnor2_1
X_4248_ VGND VPWR _1029_ _1028_ _1008_ sg13g2_or2_1
X_4179_ _0966_ net1008 net1052 VPWR VGND sg13g2_nand2_1
XFILLER_28_635 VPWR VGND sg13g2_fill_2
XFILLER_43_605 VPWR VGND sg13g2_fill_2
XFILLER_43_627 VPWR VGND sg13g2_fill_1
XFILLER_24_830 VPWR VGND sg13g2_fill_1
XFILLER_13_1024 VPWR VGND sg13g2_decap_4
XFILLER_4_2 VPWR VGND sg13g2_fill_1
XFILLER_2_299 VPWR VGND sg13g2_fill_2
XFILLER_47_922 VPWR VGND sg13g2_fill_2
XFILLER_47_966 VPWR VGND sg13g2_decap_8
XFILLER_20_1006 VPWR VGND sg13g2_decap_8
XFILLER_27_690 VPWR VGND sg13g2_fill_2
XFILLER_30_899 VPWR VGND sg13g2_fill_2
X_3550_ _0360_ _0354_ _0359_ VPWR VGND sg13g2_xnor2_1
X_5220_ _1963_ net878 net814 VPWR VGND sg13g2_nand2_1
X_3481_ _0291_ _0288_ _0293_ VPWR VGND sg13g2_xor2_1
X_5151_ _1891_ VPWR _1896_ VGND _1892_ _1894_ sg13g2_o21ai_1
X_4102_ VGND VPWR _0892_ _0891_ _0848_ sg13g2_or2_1
X_5082_ _1828_ _1800_ _1829_ VPWR VGND sg13g2_nor2b_1
X_4033_ _0779_ VPWR _0825_ VGND _0777_ _0780_ sg13g2_o21ai_1
XFILLER_38_988 VPWR VGND sg13g2_decap_8
X_5984_ _2615_ net913 net792 VPWR VGND sg13g2_nand2_1
XFILLER_24_148 VPWR VGND sg13g2_decap_4
X_4935_ _1691_ _1682_ _1690_ VPWR VGND sg13g2_xnor2_1
X_4866_ _1624_ net856 net912 VPWR VGND sg13g2_nand2_1
XFILLER_32_170 VPWR VGND sg13g2_fill_1
X_4797_ _1557_ _1550_ _1556_ VPWR VGND sg13g2_xnor2_1
X_3817_ _0617_ net960 net1023 net1021 net964 VPWR VGND sg13g2_a22oi_1
X_6536_ net1118 VGND VPWR net173 mac2.sum_lvl2_ff\[23\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_3748_ _0551_ _0542_ _0553_ VPWR VGND sg13g2_xor2_1
X_3679_ _0486_ net1031 net971 VPWR VGND sg13g2_nand2_1
X_6467_ net1140 VGND VPWR _0133_ mac2.products_ff\[83\] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_6398_ net1118 VGND VPWR net479 mac1.sum_lvl3_ff\[10\] clknet_leaf_47_clk sg13g2_dfrbpq_1
X_5418_ net319 mac1.sum_lvl2_ff\[31\] _2144_ VPWR VGND sg13g2_xor2_1
X_5349_ _2088_ _2064_ _2087_ VPWR VGND sg13g2_xnor2_1
XFILLER_43_1028 VPWR VGND sg13g2_fill_1
XFILLER_15_137 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_50_clk clknet_4_11_0_clk clknet_leaf_50_clk VPWR VGND sg13g2_buf_8
XFILLER_12_899 VPWR VGND sg13g2_decap_8
XFILLER_7_369 VPWR VGND sg13g2_fill_1
XFILLER_14_192 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_41_clk clknet_4_14_0_clk clknet_leaf_41_clk VPWR VGND sg13g2_buf_8
X_4720_ _1482_ _1475_ _1480_ _1481_ VPWR VGND sg13g2_and3_1
X_4651_ _1415_ _1408_ _1413_ _1414_ VPWR VGND sg13g2_and3_1
X_3602_ _0411_ _0404_ _0409_ _0410_ VPWR VGND sg13g2_and3_1
XFILLER_7_870 VPWR VGND sg13g2_decap_8
X_4582_ _1341_ VPWR _1352_ VGND _1312_ _1339_ sg13g2_o21ai_1
X_3533_ _0344_ _0314_ _0342_ VPWR VGND sg13g2_xnor2_1
X_6321_ net1074 VGND VPWR net166 mac1.sum_lvl2_ff\[51\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_3464_ _0272_ VPWR _0277_ VGND _0273_ _0275_ sg13g2_o21ai_1
X_6252_ net1085 VGND VPWR _0260_ DP_4.matrix\[72\] clknet_leaf_23_clk sg13g2_dfrbpq_1
XFILLER_42_0 VPWR VGND sg13g2_fill_2
X_5203_ _1947_ _1932_ _1946_ VPWR VGND sg13g2_nand2_1
X_6183_ net1063 VGND VPWR net219 mac1.sum_lvl1_ff\[1\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_5134_ _1877_ _1873_ _1879_ VPWR VGND sg13g2_xor2_1
X_3395_ _0098_ _2977_ _2978_ VPWR VGND sg13g2_xnor2_1
X_5065_ _1783_ VPWR _1812_ VGND _1781_ _1784_ sg13g2_o21ai_1
X_4016_ _0773_ VPWR _0808_ VGND _0770_ _0774_ sg13g2_o21ai_1
XFILLER_37_240 VPWR VGND sg13g2_fill_1
XFILLER_26_936 VPWR VGND sg13g2_decap_8
X_5967_ _2603_ VPWR _0203_ VGND _2471_ _2604_ sg13g2_o21ai_1
X_4918_ VGND VPWR _1622_ _1642_ _1675_ _1644_ sg13g2_a21oi_1
Xclkbuf_leaf_32_clk clknet_4_12_0_clk clknet_leaf_32_clk VPWR VGND sg13g2_buf_8
X_5898_ _2552_ _2551_ _2537_ VPWR VGND sg13g2_nand2b_1
X_4849_ _1608_ _1598_ _1607_ VPWR VGND sg13g2_nand2b_1
X_6519_ net1126 VGND VPWR net222 mac2.sum_lvl2_ff\[3\] clknet_leaf_33_clk sg13g2_dfrbpq_1
XFILLER_17_925 VPWR VGND sg13g2_decap_8
XFILLER_28_284 VPWR VGND sg13g2_fill_1
XFILLER_29_796 VPWR VGND sg13g2_decap_8
XFILLER_16_457 VPWR VGND sg13g2_decap_8
XFILLER_44_799 VPWR VGND sg13g2_fill_2
XFILLER_16_468 VPWR VGND sg13g2_fill_1
XFILLER_43_254 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_23_clk clknet_4_7_0_clk clknet_leaf_23_clk VPWR VGND sg13g2_buf_8
XFILLER_40_994 VPWR VGND sg13g2_decap_8
XFILLER_4_873 VPWR VGND sg13g2_decap_8
X_3180_ _2768_ _2769_ _2738_ _2770_ VPWR VGND sg13g2_nand3_1
Xfanout1140 net1144 net1140 VPWR VGND sg13g2_buf_8
XFILLER_39_516 VPWR VGND sg13g2_decap_4
XFILLER_16_980 VPWR VGND sg13g2_decap_8
X_5821_ DP_3.Q_range.out_data\[3\] DP_3.I_range.out_data\[3\] _2476_ VPWR VGND sg13g2_xor2_1
X_5752_ net1034 _2397_ _2409_ VPWR VGND sg13g2_and2_1
Xclkbuf_leaf_14_clk clknet_4_4_0_clk clknet_leaf_14_clk VPWR VGND sg13g2_buf_8
XFILLER_33_1016 VPWR VGND sg13g2_decap_8
X_4703_ _1465_ _1461_ _1464_ VPWR VGND sg13g2_nand2_1
X_5683_ mac2.total_sum\[7\] mac1.total_sum\[7\] _2350_ VPWR VGND sg13g2_xor2_1
XFILLER_33_1027 VPWR VGND sg13g2_fill_2
XFILLER_8_71 VPWR VGND sg13g2_fill_2
X_4634_ _1397_ _1396_ _1399_ VPWR VGND sg13g2_xor2_1
X_4565_ _1315_ VPWR _1336_ VGND _1287_ _1313_ sg13g2_o21ai_1
X_3516_ _0327_ net976 net1033 VPWR VGND sg13g2_nand2_1
X_6304_ net1098 VGND VPWR net148 mac1.sum_lvl2_ff\[31\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_4496_ _1268_ _1258_ _1270_ VPWR VGND sg13g2_xor2_1
X_6235_ net1123 VGND VPWR _0243_ DP_3.matrix\[79\] clknet_leaf_25_clk sg13g2_dfrbpq_2
X_3447_ _3023_ _3024_ _3025_ VPWR VGND sg13g2_nor2b_1
X_6166_ net1132 VGND VPWR _0194_ DP_1.matrix\[78\] clknet_leaf_51_clk sg13g2_dfrbpq_2
X_3378_ _2962_ net988 net927 VPWR VGND sg13g2_nand2_1
X_5117_ _1838_ VPWR _1863_ VGND _1859_ _1861_ sg13g2_o21ai_1
X_6097_ net1115 VGND VPWR _0115_ mac1.products_ff\[9\] clknet_leaf_59_clk sg13g2_dfrbpq_1
X_5048_ _1794_ _1795_ _1796_ VPWR VGND sg13g2_and2_1
XFILLER_26_700 VPWR VGND sg13g2_decap_4
XFILLER_26_711 VPWR VGND sg13g2_fill_2
XFILLER_26_799 VPWR VGND sg13g2_fill_1
XFILLER_41_703 VPWR VGND sg13g2_fill_1
Xclkbuf_4_8_0_clk clknet_0_clk clknet_4_8_0_clk VPWR VGND sg13g2_buf_8
XFILLER_43_79 VPWR VGND sg13g2_fill_2
XFILLER_22_994 VPWR VGND sg13g2_decap_8
XFILLER_49_1001 VPWR VGND sg13g2_decap_8
XFILLER_1_865 VPWR VGND sg13g2_decap_8
XFILLER_48_346 VPWR VGND sg13g2_fill_2
XFILLER_16_221 VPWR VGND sg13g2_fill_1
XFILLER_44_585 VPWR VGND sg13g2_fill_1
XFILLER_16_287 VPWR VGND sg13g2_fill_2
XFILLER_31_213 VPWR VGND sg13g2_fill_1
XFILLER_9_910 VPWR VGND sg13g2_decap_8
XFILLER_13_961 VPWR VGND sg13g2_decap_8
XFILLER_9_987 VPWR VGND sg13g2_decap_8
XFILLER_8_486 VPWR VGND sg13g2_fill_1
X_4350_ _1126_ _1125_ _0135_ VPWR VGND sg13g2_xor2_1
X_3301_ _2887_ _2875_ _2888_ VPWR VGND sg13g2_xor2_1
X_4281_ _1060_ _1058_ _1059_ VPWR VGND sg13g2_nand2b_1
X_6020_ net1023 _0180_ VPWR VGND sg13g2_buf_1
X_3232_ _2821_ _2819_ _2820_ VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_3_clk clknet_4_1_0_clk clknet_leaf_3_clk VPWR VGND sg13g2_buf_8
X_3163_ _2721_ VPWR _2753_ VGND _2719_ _2722_ sg13g2_o21ai_1
X_3094_ _2666_ VPWR _2686_ VGND _2664_ _2667_ sg13g2_o21ai_1
X_5804_ _2460_ _2448_ _2459_ VPWR VGND sg13g2_nand2_1
XFILLER_22_213 VPWR VGND sg13g2_decap_8
XFILLER_22_224 VPWR VGND sg13g2_fill_2
X_3996_ _0786_ _0787_ _0769_ _0789_ VPWR VGND sg13g2_nand3_1
X_5735_ _2392_ _2389_ _2391_ VPWR VGND sg13g2_nand2_1
X_5666_ _2337_ mac1.total_sum\[3\] mac2.total_sum\[3\] VPWR VGND sg13g2_xnor2_1
X_4617_ net924 net922 net859 net857 _1382_ VPWR VGND sg13g2_and4_1
Xhold420 DP_2.matrix\[5\] VPWR VGND net460 sg13g2_dlygate4sd3_1
X_5597_ net444 mac2.sum_lvl3_ff\[24\] _2283_ VPWR VGND sg13g2_xor2_1
Xhold442 DP_2.matrix\[74\] VPWR VGND net482 sg13g2_dlygate4sd3_1
Xhold453 DP_1.matrix\[38\] VPWR VGND net493 sg13g2_dlygate4sd3_1
X_4548_ _1281_ _1319_ _1320_ VPWR VGND sg13g2_nor2_1
Xhold431 _0043_ VPWR VGND net471 sg13g2_dlygate4sd3_1
Xhold464 DP_1.matrix\[1\] VPWR VGND net504 sg13g2_dlygate4sd3_1
Xhold475 DP_1.matrix\[73\] VPWR VGND net515 sg13g2_dlygate4sd3_1
Xhold486 _0018_ VPWR VGND net526 sg13g2_dlygate4sd3_1
Xfanout900 net901 net900 VPWR VGND sg13g2_buf_8
X_4479_ _1253_ net837 DP_3.matrix\[42\] VPWR VGND sg13g2_nand2_2
Xfanout911 net913 net911 VPWR VGND sg13g2_buf_8
Xhold497 _2125_ VPWR VGND net537 sg13g2_dlygate4sd3_1
Xfanout933 net404 net933 VPWR VGND sg13g2_buf_2
X_6218_ net1122 VGND VPWR _0229_ DP_3.matrix\[37\] clknet_leaf_32_clk sg13g2_dfrbpq_2
Xfanout922 net923 net922 VPWR VGND sg13g2_buf_8
Xfanout944 net945 net944 VPWR VGND sg13g2_buf_1
Xfanout955 net431 net955 VPWR VGND sg13g2_buf_1
Xfanout977 DP_2.matrix\[2\] net977 VPWR VGND sg13g2_buf_1
Xfanout966 net968 net966 VPWR VGND sg13g2_buf_8
XFILLER_46_806 VPWR VGND sg13g2_fill_2
Xfanout999 net492 net999 VPWR VGND sg13g2_buf_8
X_6149_ net1088 VGND VPWR _0183_ DP_1.matrix\[39\] clknet_leaf_63_clk sg13g2_dfrbpq_1
Xfanout988 DP_1.matrix\[79\] net988 VPWR VGND sg13g2_buf_1
XFILLER_26_552 VPWR VGND sg13g2_fill_1
XFILLER_13_246 VPWR VGND sg13g2_fill_2
XFILLER_9_239 VPWR VGND sg13g2_fill_2
XFILLER_16_1022 VPWR VGND sg13g2_decap_8
XFILLER_10_931 VPWR VGND sg13g2_decap_8
XFILLER_6_902 VPWR VGND sg13g2_decap_8
XFILLER_6_979 VPWR VGND sg13g2_decap_8
XFILLER_49_622 VPWR VGND sg13g2_fill_2
XFILLER_45_894 VPWR VGND sg13g2_decap_8
XFILLER_17_585 VPWR VGND sg13g2_fill_1
X_3850_ _0647_ net1014 net965 net1017 net961 VPWR VGND sg13g2_a22oi_1
XFILLER_13_780 VPWR VGND sg13g2_fill_2
X_3781_ _0583_ _0584_ _0585_ VPWR VGND sg13g2_and2_1
X_5520_ _2223_ mac2.sum_lvl2_ff\[22\] net432 VPWR VGND sg13g2_nand2_1
X_5451_ mac1.sum_lvl3_ff\[24\] mac1.sum_lvl3_ff\[4\] _2169_ VPWR VGND sg13g2_and2_1
X_5382_ VGND VPWR _2112_ _2114_ _2115_ _2113_ sg13g2_a21oi_1
X_4402_ _1132_ _1135_ _1178_ VPWR VGND sg13g2_nor2_1
X_4333_ _1111_ _1104_ _1109_ _1110_ VPWR VGND sg13g2_and3_1
X_4264_ _1044_ _1037_ _1042_ _1043_ VPWR VGND sg13g2_and3_1
X_6003_ _2627_ net856 net792 VPWR VGND sg13g2_nand2_1
X_3215_ _2801_ _2802_ _2796_ _2804_ VPWR VGND sg13g2_nand3_1
X_4195_ _0970_ VPWR _0981_ VGND _0941_ _0968_ sg13g2_o21ai_1
X_3146_ _2703_ VPWR _2737_ VGND _2678_ _2704_ sg13g2_o21ai_1
X_3077_ _2668_ _2669_ _2663_ _2670_ VPWR VGND sg13g2_nand3_1
XFILLER_39_187 VPWR VGND sg13g2_fill_2
XFILLER_39_1000 VPWR VGND sg13g2_decap_8
X_3979_ _0772_ net954 net1010 VPWR VGND sg13g2_nand2_1
X_5718_ VGND VPWR _2374_ _2376_ _2378_ _2375_ sg13g2_a21oi_1
X_5649_ net297 mac2.sum_lvl3_ff\[34\] _2325_ VPWR VGND sg13g2_xor2_1
XFILLER_3_916 VPWR VGND sg13g2_decap_8
XFILLER_46_1015 VPWR VGND sg13g2_decap_8
Xhold261 DP_3.matrix\[75\] VPWR VGND net301 sg13g2_dlygate4sd3_1
Xhold250 _2214_ VPWR VGND net290 sg13g2_dlygate4sd3_1
XFILLER_49_23 VPWR VGND sg13g2_fill_2
Xhold283 DP_1.matrix\[41\] VPWR VGND net323 sg13g2_dlygate4sd3_1
Xhold272 DP_1.matrix\[39\] VPWR VGND net312 sg13g2_dlygate4sd3_1
Xhold294 DP_4.matrix\[43\] VPWR VGND net334 sg13g2_dlygate4sd3_1
XFILLER_49_89 VPWR VGND sg13g2_fill_1
Xfanout785 net788 net785 VPWR VGND sg13g2_buf_8
Xfanout796 _2481_ net796 VPWR VGND sg13g2_buf_1
XFILLER_34_809 VPWR VGND sg13g2_fill_1
XFILLER_45_168 VPWR VGND sg13g2_fill_1
XFILLER_14_555 VPWR VGND sg13g2_fill_1
XFILLER_5_220 VPWR VGND sg13g2_fill_2
XFILLER_6_776 VPWR VGND sg13g2_fill_2
XFILLER_5_253 VPWR VGND sg13g2_fill_1
Xinput7 ui_in[6] net7 VPWR VGND sg13g2_buf_1
XFILLER_36_124 VPWR VGND sg13g2_fill_1
XFILLER_18_861 VPWR VGND sg13g2_decap_8
X_4951_ _1690_ _1682_ _1689_ _1706_ VPWR VGND sg13g2_a21o_1
XFILLER_36_179 VPWR VGND sg13g2_fill_1
X_4882_ _1639_ _1632_ _1640_ VPWR VGND sg13g2_nor2b_1
X_3902_ _0697_ _0692_ _0695_ VPWR VGND sg13g2_xnor2_1
X_3833_ _0627_ _0628_ _0630_ _0631_ VPWR VGND sg13g2_nor3_1
XFILLER_20_503 VPWR VGND sg13g2_fill_1
X_3764_ _0547_ VPWR _0568_ VGND _0544_ _0548_ sg13g2_o21ai_1
X_6552_ net1102 VGND VPWR net272 mac2.sum_lvl3_ff\[0\] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_3695_ _0466_ _0500_ _0464_ _0502_ VPWR VGND sg13g2_nand3_1
X_5503_ mac1.sum_lvl3_ff\[34\] mac1.sum_lvl3_ff\[14\] _2211_ VPWR VGND sg13g2_nor2_1
X_6483_ net1101 VGND VPWR _0155_ mac2.products_ff\[151\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_5434_ _2157_ mac1.sum_lvl2_ff\[34\] net284 VPWR VGND sg13g2_xnor2_1
X_5365_ _2102_ net287 net267 VPWR VGND sg13g2_nand2_1
X_5296_ _2037_ _2029_ _2036_ VPWR VGND sg13g2_xnor2_1
X_4316_ _1094_ _1090_ _1093_ VPWR VGND sg13g2_nand2_1
X_4247_ _1026_ _1025_ _1028_ VPWR VGND sg13g2_xor2_1
X_4178_ _0944_ VPWR _0965_ VGND _0916_ _0942_ sg13g2_o21ai_1
XFILLER_28_658 VPWR VGND sg13g2_decap_4
X_3129_ net944 net939 net992 net989 _2720_ VPWR VGND sg13g2_and4_1
XFILLER_13_1003 VPWR VGND sg13g2_decap_8
XFILLER_47_945 VPWR VGND sg13g2_decap_8
XFILLER_15_831 VPWR VGND sg13g2_decap_8
XFILLER_18_179 VPWR VGND sg13g2_fill_2
XFILLER_15_897 VPWR VGND sg13g2_decap_8
XFILLER_30_834 VPWR VGND sg13g2_decap_4
XFILLER_30_878 VPWR VGND sg13g2_fill_2
X_3480_ _0292_ _0291_ _0288_ VPWR VGND sg13g2_nand2b_1
XFILLER_29_1010 VPWR VGND sg13g2_decap_8
X_5150_ _1891_ _1892_ _1894_ _1895_ VPWR VGND sg13g2_or3_1
X_5081_ _1828_ _1804_ _1827_ VPWR VGND sg13g2_xnor2_1
X_4101_ _0891_ net1010 net949 VPWR VGND sg13g2_nand2_2
X_4032_ _0824_ _0819_ _0823_ VPWR VGND sg13g2_xnor2_1
X_5983_ net793 net915 _2614_ _0225_ VPWR VGND sg13g2_a21o_1
XFILLER_24_105 VPWR VGND sg13g2_fill_2
X_4934_ _1690_ _1654_ _1688_ VPWR VGND sg13g2_xnor2_1
XFILLER_17_190 VPWR VGND sg13g2_fill_2
X_4865_ _1606_ _1599_ _1569_ _1623_ VPWR VGND sg13g2_a21o_2
X_4796_ _1556_ _1551_ _1554_ VPWR VGND sg13g2_xnor2_1
X_3816_ _0616_ net1021 net960 _0074_ VPWR VGND sg13g2_and3_2
X_3747_ _0551_ _0542_ _0552_ VPWR VGND sg13g2_nor2b_1
X_6535_ net1120 VGND VPWR net203 mac2.sum_lvl2_ff\[22\] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_3678_ VGND VPWR net981 net1025 _0485_ _0454_ sg13g2_a21oi_1
X_6466_ net1140 VGND VPWR _0132_ mac2.products_ff\[82\] clknet_leaf_41_clk sg13g2_dfrbpq_1
X_6397_ net1114 VGND VPWR net459 mac1.sum_lvl3_ff\[9\] clknet_leaf_60_clk sg13g2_dfrbpq_1
X_5417_ mac1.sum_lvl2_ff\[31\] net319 _2143_ VPWR VGND sg13g2_nor2_1
X_5348_ _2085_ _2079_ _2087_ VPWR VGND sg13g2_xor2_1
XFILLER_0_716 VPWR VGND sg13g2_fill_1
XFILLER_43_1007 VPWR VGND sg13g2_decap_8
X_5279_ _2019_ _2020_ _2021_ VPWR VGND sg13g2_nor2_1
XFILLER_29_989 VPWR VGND sg13g2_decap_8
XFILLER_43_447 VPWR VGND sg13g2_fill_2
XFILLER_43_469 VPWR VGND sg13g2_fill_2
XFILLER_7_304 VPWR VGND sg13g2_fill_2
XFILLER_12_878 VPWR VGND sg13g2_decap_8
XFILLER_2_0 VPWR VGND sg13g2_fill_1
XFILLER_3_598 VPWR VGND sg13g2_fill_1
XFILLER_47_731 VPWR VGND sg13g2_fill_2
XFILLER_47_753 VPWR VGND sg13g2_fill_2
XFILLER_15_683 VPWR VGND sg13g2_fill_1
X_4650_ _1409_ VPWR _1414_ VGND _1410_ _1412_ sg13g2_o21ai_1
X_3601_ _0405_ VPWR _0410_ VGND _0406_ _0408_ sg13g2_o21ai_1
Xinput10 uio_in[1] net10 VPWR VGND sg13g2_buf_1
X_6320_ net1073 VGND VPWR net248 mac1.sum_lvl2_ff\[50\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_4581_ VGND VPWR _1320_ _1344_ _1351_ _1346_ sg13g2_a21oi_1
X_3532_ _0342_ _0314_ _0343_ VPWR VGND sg13g2_nor2b_1
X_3463_ _0272_ _0273_ _0275_ _0276_ VPWR VGND sg13g2_or3_1
X_6251_ net1139 VGND VPWR _0259_ DP_4.matrix\[43\] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_5202_ _1945_ _1938_ _1946_ VPWR VGND sg13g2_xor2_1
X_6182_ net1072 VGND VPWR _0205_ DP_2.matrix\[37\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_5133_ _1873_ _1877_ _1878_ VPWR VGND sg13g2_nor2_1
X_3394_ VGND VPWR _2955_ _2958_ _2978_ _2954_ sg13g2_a21oi_1
XFILLER_35_0 VPWR VGND sg13g2_fill_2
X_5064_ _1811_ _1806_ _1809_ VPWR VGND sg13g2_xnor2_1
XFILLER_29_219 VPWR VGND sg13g2_fill_2
XFILLER_38_720 VPWR VGND sg13g2_fill_1
X_4015_ _0761_ _0764_ _0807_ VPWR VGND sg13g2_nor2_1
XFILLER_25_403 VPWR VGND sg13g2_fill_2
XFILLER_25_414 VPWR VGND sg13g2_fill_1
XFILLER_25_425 VPWR VGND sg13g2_decap_8
XFILLER_16_27 VPWR VGND sg13g2_fill_2
XFILLER_25_436 VPWR VGND sg13g2_fill_2
XFILLER_25_458 VPWR VGND sg13g2_fill_2
X_5966_ _2467_ _2470_ _2604_ VPWR VGND sg13g2_nor2b_1
X_4917_ _1672_ _1651_ _1674_ VPWR VGND sg13g2_xor2_1
X_5897_ _2550_ _2546_ _2551_ VPWR VGND sg13g2_nor2b_1
X_4848_ _1607_ _1599_ _1606_ VPWR VGND sg13g2_xnor2_1
X_4779_ _1492_ VPWR _1540_ VGND _1431_ _1493_ sg13g2_o21ai_1
X_6518_ net1124 VGND VPWR net158 mac2.sum_lvl2_ff\[2\] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_6449_ net1145 VGND VPWR _0142_ mac2.products_ff\[13\] clknet_leaf_38_clk sg13g2_dfrbpq_1
XFILLER_17_904 VPWR VGND sg13g2_decap_8
XFILLER_40_973 VPWR VGND sg13g2_decap_8
XFILLER_4_852 VPWR VGND sg13g2_decap_8
XFILLER_26_1013 VPWR VGND sg13g2_decap_8
Xfanout1130 net1148 net1130 VPWR VGND sg13g2_buf_8
Xfanout1141 net1144 net1141 VPWR VGND sg13g2_buf_8
XFILLER_34_244 VPWR VGND sg13g2_fill_2
X_5820_ _2475_ net506 _2474_ VPWR VGND sg13g2_nand2_2
X_5751_ _2408_ net800 _2407_ net802 DP_1.matrix\[77\] VPWR VGND sg13g2_a22oi_1
X_4702_ _1462_ _1463_ _1464_ VPWR VGND sg13g2_nor2b_1
X_5682_ _2349_ mac1.total_sum\[7\] mac2.total_sum\[7\] VPWR VGND sg13g2_nand2_1
X_4633_ _1396_ _1397_ _1398_ VPWR VGND sg13g2_nor2b_2
X_4564_ _1318_ _1310_ _1317_ _1335_ VPWR VGND sg13g2_a21o_1
X_3515_ _0297_ VPWR _0326_ VGND _0295_ _0298_ sg13g2_o21ai_1
X_6303_ net1107 VGND VPWR net42 mac1.sum_lvl2_ff\[30\] clknet_leaf_10_clk sg13g2_dfrbpq_2
X_6234_ net1104 VGND VPWR _0242_ DP_3.matrix\[78\] clknet_leaf_25_clk sg13g2_dfrbpq_2
X_4495_ _1258_ _1268_ _1269_ VPWR VGND sg13g2_nor2_1
X_3446_ _3019_ VPWR _3024_ VGND _3020_ _3022_ sg13g2_o21ai_1
X_3377_ _2961_ net993 DP_2.matrix\[80\] VPWR VGND sg13g2_nand2_1
X_6165_ net1133 VGND VPWR _0096_ mac1.products_ff\[147\] clknet_leaf_48_clk sg13g2_dfrbpq_1
X_5116_ _1838_ _1859_ _1861_ _1862_ VPWR VGND sg13g2_or3_1
X_6096_ net1114 VGND VPWR _0114_ mac1.products_ff\[8\] clknet_leaf_59_clk sg13g2_dfrbpq_1
X_5047_ _1793_ _1792_ _1754_ _1795_ VPWR VGND sg13g2_a21o_1
XFILLER_26_778 VPWR VGND sg13g2_decap_4
X_5949_ VGND VPWR net785 _2592_ _0197_ _2591_ sg13g2_a21oi_1
XFILLER_13_428 VPWR VGND sg13g2_fill_1
XFILLER_22_973 VPWR VGND sg13g2_decap_8
XFILLER_4_115 VPWR VGND sg13g2_fill_2
XFILLER_1_844 VPWR VGND sg13g2_decap_8
XFILLER_0_343 VPWR VGND sg13g2_fill_1
XFILLER_1_1026 VPWR VGND sg13g2_fill_2
XFILLER_17_92 VPWR VGND sg13g2_fill_2
XFILLER_17_767 VPWR VGND sg13g2_fill_2
XFILLER_13_940 VPWR VGND sg13g2_decap_8
XFILLER_12_461 VPWR VGND sg13g2_fill_1
XFILLER_9_966 VPWR VGND sg13g2_decap_8
X_3300_ _2885_ _2876_ _2887_ VPWR VGND sg13g2_xor2_1
X_4280_ _1059_ net907 net835 VPWR VGND sg13g2_nand2_1
X_3231_ _2817_ _2816_ _2818_ _2820_ VPWR VGND sg13g2_a21o_1
X_3162_ _2752_ _2746_ _2751_ VPWR VGND sg13g2_xnor2_1
X_3093_ _2683_ _2680_ _2685_ VPWR VGND sg13g2_xor2_1
XFILLER_39_369 VPWR VGND sg13g2_fill_2
X_5803_ _2458_ _2456_ _2459_ VPWR VGND sg13g2_nor2b_1
X_3995_ _0788_ _0769_ _0786_ _0787_ VPWR VGND sg13g2_and3_1
X_5734_ VGND VPWR _2386_ _2387_ _2391_ _2390_ sg13g2_a21oi_1
X_5665_ _2336_ mac1.total_sum\[3\] mac2.total_sum\[3\] VPWR VGND sg13g2_nand2_1
X_4616_ _1381_ net922 net857 VPWR VGND sg13g2_nand2_1
Xhold410 DP_4.matrix\[5\] VPWR VGND net450 sg13g2_dlygate4sd3_1
X_5596_ mac2.sum_lvl3_ff\[24\] net444 _2282_ VPWR VGND sg13g2_and2_1
Xhold454 mac1.sum_lvl3_ff\[8\] VPWR VGND net494 sg13g2_dlygate4sd3_1
Xhold432 DP_2.matrix\[1\] VPWR VGND net472 sg13g2_dlygate4sd3_1
Xhold421 mac1.sum_lvl2_ff\[6\] VPWR VGND net461 sg13g2_dlygate4sd3_1
Xhold443 DP_3.matrix\[39\] VPWR VGND net483 sg13g2_dlygate4sd3_1
X_4547_ _1319_ _1310_ _1318_ VPWR VGND sg13g2_xnor2_1
Xhold476 _2637_ VPWR VGND net516 sg13g2_dlygate4sd3_1
Xhold487 DP_2.matrix\[8\] VPWR VGND net527 sg13g2_dlygate4sd3_1
X_4478_ _1235_ _1228_ _1198_ _1252_ VPWR VGND sg13g2_a21o_1
Xhold465 DP_3.Q_range.out_data\[4\] VPWR VGND net505 sg13g2_dlygate4sd3_1
Xfanout912 net913 net912 VPWR VGND sg13g2_buf_1
X_3429_ _3009_ net978 net1040 net1038 net982 VPWR VGND sg13g2_a22oi_1
Xhold498 _0013_ VPWR VGND net538 sg13g2_dlygate4sd3_1
Xfanout934 net935 net934 VPWR VGND sg13g2_buf_8
X_6217_ net1121 VGND VPWR _0228_ DP_3.matrix\[36\] clknet_leaf_46_clk sg13g2_dfrbpq_1
Xfanout901 net483 net901 VPWR VGND sg13g2_buf_8
Xfanout923 net422 net923 VPWR VGND sg13g2_buf_8
Xfanout956 net957 net956 VPWR VGND sg13g2_buf_8
X_6148_ net1088 VGND VPWR _0182_ DP_1.matrix\[38\] clknet_leaf_64_clk sg13g2_dfrbpq_1
Xfanout945 DP_2.matrix\[72\] net945 VPWR VGND sg13g2_buf_1
Xfanout967 net968 net967 VPWR VGND sg13g2_buf_1
Xfanout978 net472 net978 VPWR VGND sg13g2_buf_2
Xfanout989 net990 net989 VPWR VGND sg13g2_buf_8
X_6079_ net270 _0263_ VPWR VGND sg13g2_buf_1
XFILLER_16_1001 VPWR VGND sg13g2_decap_8
XFILLER_41_556 VPWR VGND sg13g2_fill_1
XFILLER_10_910 VPWR VGND sg13g2_decap_8
XFILLER_9_218 VPWR VGND sg13g2_fill_1
XFILLER_10_987 VPWR VGND sg13g2_decap_8
XFILLER_6_958 VPWR VGND sg13g2_decap_8
XFILLER_5_446 VPWR VGND sg13g2_fill_2
XFILLER_49_667 VPWR VGND sg13g2_fill_1
XFILLER_48_111 VPWR VGND sg13g2_fill_2
XFILLER_0_173 VPWR VGND sg13g2_fill_1
XFILLER_29_391 VPWR VGND sg13g2_fill_1
XFILLER_45_884 VPWR VGND sg13g2_fill_2
XFILLER_32_523 VPWR VGND sg13g2_fill_2
XFILLER_32_567 VPWR VGND sg13g2_fill_1
XFILLER_20_729 VPWR VGND sg13g2_decap_4
X_3780_ _0557_ _0559_ _0582_ _0584_ VPWR VGND sg13g2_or3_1
XFILLER_9_774 VPWR VGND sg13g2_fill_1
X_5450_ _2166_ VPWR _2168_ VGND _2165_ _2167_ sg13g2_o21ai_1
X_4401_ _1160_ VPWR _1177_ VGND _1139_ _1161_ sg13g2_o21ai_1
X_5381_ net341 _2112_ _0010_ VPWR VGND sg13g2_xor2_1
X_4332_ _1105_ VPWR _1110_ VGND _1106_ _1108_ sg13g2_o21ai_1
X_4263_ _1038_ VPWR _1043_ VGND _1039_ _1041_ sg13g2_o21ai_1
X_6002_ _2625_ VPWR _0248_ VGND net793 _2626_ sg13g2_o21ai_1
X_3214_ _2803_ _2796_ _2801_ _2802_ VPWR VGND sg13g2_and3_1
Xclkbuf_4_7_0_clk clknet_0_clk clknet_4_7_0_clk VPWR VGND sg13g2_buf_8
X_4194_ VGND VPWR _0949_ _0973_ _0980_ _0975_ sg13g2_a21oi_1
X_3145_ _2736_ _2706_ _2734_ VPWR VGND sg13g2_xnor2_1
X_3076_ _2664_ VPWR _2669_ VGND _2665_ _2667_ sg13g2_o21ai_1
XFILLER_36_840 VPWR VGND sg13g2_fill_1
X_3978_ _0771_ net952 net1010 VPWR VGND sg13g2_nand2_2
XFILLER_23_567 VPWR VGND sg13g2_fill_2
X_5717_ net22 _2374_ _2377_ VPWR VGND sg13g2_xnor2_1
X_5648_ mac2.sum_lvl3_ff\[34\] net297 _2324_ VPWR VGND sg13g2_nor2_1
X_5579_ _2270_ mac2.sum_lvl2_ff\[34\] net484 VPWR VGND sg13g2_xnor2_1
Xhold262 DP_3.matrix\[8\] VPWR VGND net302 sg13g2_dlygate4sd3_1
Xhold240 DP_1.matrix\[7\] VPWR VGND net280 sg13g2_dlygate4sd3_1
Xhold251 _0022_ VPWR VGND net291 sg13g2_dlygate4sd3_1
Xhold284 DP_4.matrix\[79\] VPWR VGND net324 sg13g2_dlygate4sd3_1
Xhold273 DP_1.matrix\[40\] VPWR VGND net313 sg13g2_dlygate4sd3_1
Xhold295 DP_4.matrix\[42\] VPWR VGND net335 sg13g2_dlygate4sd3_1
XFILLER_49_57 VPWR VGND sg13g2_fill_1
Xfanout797 net798 net797 VPWR VGND sg13g2_buf_8
Xfanout786 net788 net786 VPWR VGND sg13g2_buf_8
XFILLER_26_383 VPWR VGND sg13g2_fill_2
XFILLER_26_394 VPWR VGND sg13g2_fill_2
XFILLER_7_1010 VPWR VGND sg13g2_decap_8
XFILLER_2_994 VPWR VGND sg13g2_decap_8
Xinput8 ui_in[7] net8 VPWR VGND sg13g2_buf_1
X_4950_ VGND VPWR _1681_ _1695_ _1705_ _1694_ sg13g2_a21oi_1
X_4881_ _1639_ _1633_ _1638_ VPWR VGND sg13g2_xnor2_1
XFILLER_45_692 VPWR VGND sg13g2_fill_2
X_3901_ _0696_ _0695_ _0692_ VPWR VGND sg13g2_nand2b_1
X_3832_ _0630_ net1016 net962 net1018 net959 VPWR VGND sg13g2_a22oi_1
X_6551_ net1075 VGND VPWR DP_1.I_range.data_plus_4\[6\] DP_1.I_range.out_data\[5\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_32_397 VPWR VGND sg13g2_fill_2
XFILLER_20_559 VPWR VGND sg13g2_fill_1
X_3763_ _0550_ _0543_ _0552_ _0567_ VPWR VGND sg13g2_a21o_1
X_5502_ _2210_ mac1.sum_lvl3_ff\[34\] mac1.sum_lvl3_ff\[14\] VPWR VGND sg13g2_nand2_1
X_3694_ VGND VPWR _0464_ _0466_ _0501_ _0500_ sg13g2_a21oi_1
X_6482_ net1085 VGND VPWR _0154_ mac2.products_ff\[150\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_5433_ _2153_ VPWR _2156_ VGND _2152_ _2154_ sg13g2_o21ai_1
X_5364_ _0155_ _2094_ _2101_ VPWR VGND sg13g2_xnor2_1
X_4315_ _1091_ _1092_ _1093_ VPWR VGND sg13g2_nor2b_1
X_5295_ _2036_ _2030_ _2035_ VPWR VGND sg13g2_xnor2_1
X_4246_ _1025_ _1026_ _1027_ VPWR VGND sg13g2_nor2b_2
X_4177_ _0947_ _0939_ _0946_ _0964_ VPWR VGND sg13g2_a21o_1
X_3128_ _2719_ net937 net995 VPWR VGND sg13g2_nand2_1
XFILLER_43_607 VPWR VGND sg13g2_fill_1
XFILLER_27_158 VPWR VGND sg13g2_fill_2
X_3059_ _2651_ _2652_ _2653_ VPWR VGND sg13g2_nor2b_2
XFILLER_11_559 VPWR VGND sg13g2_fill_2
XFILLER_3_714 VPWR VGND sg13g2_fill_1
XFILLER_47_924 VPWR VGND sg13g2_fill_1
XFILLER_18_125 VPWR VGND sg13g2_fill_2
XFILLER_15_810 VPWR VGND sg13g2_fill_1
XFILLER_27_692 VPWR VGND sg13g2_fill_1
XFILLER_15_876 VPWR VGND sg13g2_decap_8
XFILLER_30_857 VPWR VGND sg13g2_fill_1
XFILLER_6_552 VPWR VGND sg13g2_fill_1
XFILLER_2_780 VPWR VGND sg13g2_decap_8
X_4100_ _0890_ net1016 net1052 VPWR VGND sg13g2_nand2_1
X_5080_ _1827_ _1824_ _1826_ VPWR VGND sg13g2_nand2_1
X_4031_ _0823_ _0771_ _0820_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_913 VPWR VGND sg13g2_fill_2
XFILLER_37_401 VPWR VGND sg13g2_fill_2
X_5982_ VGND VPWR _2485_ _2510_ _2614_ _2613_ sg13g2_a21oi_1
X_4933_ _1654_ _1688_ _1689_ VPWR VGND sg13g2_nor2b_1
XFILLER_24_139 VPWR VGND sg13g2_fill_1
XFILLER_36_1015 VPWR VGND sg13g2_decap_8
X_4864_ _1608_ VPWR _1622_ VGND _1597_ _1609_ sg13g2_o21ai_1
X_4795_ _1555_ _1554_ _1551_ VPWR VGND sg13g2_nand2b_1
X_3815_ net1023 net964 _0074_ VPWR VGND sg13g2_and2_1
XFILLER_21_28 VPWR VGND sg13g2_fill_2
X_3746_ _0551_ _0543_ _0550_ VPWR VGND sg13g2_xnor2_1
X_6534_ net1124 VGND VPWR net210 mac2.sum_lvl2_ff\[21\] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_6465_ net1141 VGND VPWR _0131_ mac2.products_ff\[81\] clknet_leaf_41_clk sg13g2_dfrbpq_1
X_3677_ _0458_ VPWR _0484_ VGND _0452_ _0459_ sg13g2_o21ai_1
X_5416_ _2142_ mac1.sum_lvl2_ff\[31\] net319 VPWR VGND sg13g2_nand2_1
X_6396_ net1112 VGND VPWR net395 mac1.sum_lvl3_ff\[8\] clknet_leaf_57_clk sg13g2_dfrbpq_1
X_5347_ _2086_ _2079_ _2085_ VPWR VGND sg13g2_nand2_1
X_5278_ VGND VPWR _1983_ _1985_ _2020_ _2017_ sg13g2_a21oi_1
X_4229_ _1010_ net904 net838 VPWR VGND sg13g2_nand2_1
XFILLER_28_456 VPWR VGND sg13g2_decap_8
XFILLER_29_968 VPWR VGND sg13g2_decap_8
XFILLER_12_813 VPWR VGND sg13g2_decap_8
XFILLER_24_662 VPWR VGND sg13g2_fill_1
XFILLER_12_857 VPWR VGND sg13g2_decap_8
XFILLER_11_50 VPWR VGND sg13g2_fill_2
XFILLER_11_61 VPWR VGND sg13g2_fill_2
XFILLER_38_209 VPWR VGND sg13g2_fill_2
XFILLER_4_1013 VPWR VGND sg13g2_decap_8
XFILLER_21_109 VPWR VGND sg13g2_fill_1
XFILLER_43_993 VPWR VGND sg13g2_decap_8
Xinput11 uio_in[2] net11 VPWR VGND sg13g2_buf_1
X_3600_ _0405_ _0406_ _0408_ _0409_ VPWR VGND sg13g2_or3_1
X_4580_ VGND VPWR _1333_ _1349_ _1350_ _1348_ sg13g2_a21oi_1
X_3531_ _0342_ _0318_ _0341_ VPWR VGND sg13g2_xnor2_1
X_3462_ _0275_ net1033 net985 net1034 net981 VPWR VGND sg13g2_a22oi_1
X_6250_ net1139 VGND VPWR _0258_ DP_4.matrix\[42\] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_5201_ _1945_ _1939_ _1943_ VPWR VGND sg13g2_xnor2_1
X_6181_ net1071 VGND VPWR _0204_ DP_2.matrix\[36\] clknet_leaf_66_clk sg13g2_dfrbpq_1
X_3393_ _2975_ _2976_ _2977_ VPWR VGND sg13g2_and2_1
X_5132_ VGND VPWR _1877_ _1876_ _1875_ sg13g2_or2_1
X_5063_ _1810_ _1809_ _1806_ VPWR VGND sg13g2_nand2b_1
X_4014_ _0789_ VPWR _0806_ VGND _0768_ _0790_ sg13g2_o21ai_1
X_5965_ _2603_ net968 net784 VPWR VGND sg13g2_nand2b_1
X_4916_ _1672_ _1651_ _1673_ VPWR VGND sg13g2_nor2b_1
X_5896_ VGND VPWR net370 net798 _2550_ _2549_ sg13g2_a21oi_1
X_4847_ _1604_ _1605_ _1606_ VPWR VGND sg13g2_nor2b_1
X_4778_ _1465_ VPWR _1539_ VGND _1535_ _1537_ sg13g2_o21ai_1
X_3729_ _0533_ _0534_ _0535_ VPWR VGND sg13g2_nor2_1
X_6517_ net1105 VGND VPWR net65 mac2.sum_lvl2_ff\[1\] clknet_leaf_30_clk sg13g2_dfrbpq_1
X_6448_ net1145 VGND VPWR _0141_ mac2.products_ff\[12\] clknet_leaf_38_clk sg13g2_dfrbpq_1
X_6379_ net1138 VGND VPWR net209 mac1.sum_lvl3_ff\[27\] clknet_leaf_51_clk sg13g2_dfrbpq_2
XFILLER_0_569 VPWR VGND sg13g2_fill_2
XFILLER_16_404 VPWR VGND sg13g2_fill_2
XFILLER_43_212 VPWR VGND sg13g2_fill_1
XFILLER_19_1021 VPWR VGND sg13g2_decap_8
XFILLER_25_982 VPWR VGND sg13g2_decap_8
XFILLER_31_418 VPWR VGND sg13g2_decap_8
XFILLER_31_429 VPWR VGND sg13g2_fill_1
XFILLER_11_153 VPWR VGND sg13g2_fill_2
XFILLER_11_175 VPWR VGND sg13g2_fill_2
XFILLER_11_197 VPWR VGND sg13g2_fill_2
XFILLER_4_831 VPWR VGND sg13g2_decap_8
Xfanout1131 net1132 net1131 VPWR VGND sg13g2_buf_8
Xfanout1120 net1121 net1120 VPWR VGND sg13g2_buf_8
Xfanout1142 net1143 net1142 VPWR VGND sg13g2_buf_8
X_5750_ DP_1.matrix\[5\] net1012 net810 _2407_ VPWR VGND sg13g2_mux2_1
XFILLER_31_930 VPWR VGND sg13g2_decap_8
XFILLER_15_492 VPWR VGND sg13g2_fill_1
X_5681_ _2347_ _2348_ net31 VPWR VGND sg13g2_nor2b_2
X_4701_ DP_3.matrix\[1\] net854 net925 _1463_ VPWR VGND net851 sg13g2_nand4_1
XFILLER_31_985 VPWR VGND sg13g2_decap_8
X_4632_ _1376_ VPWR _1397_ VGND _1367_ _1377_ sg13g2_o21ai_1
XFILLER_8_73 VPWR VGND sg13g2_fill_1
X_4563_ _1322_ _1324_ _1334_ VPWR VGND sg13g2_and2_1
XFILLER_7_691 VPWR VGND sg13g2_fill_2
X_3514_ _0325_ _0320_ _0323_ VPWR VGND sg13g2_xnor2_1
X_6302_ net1120 VGND VPWR net262 mac1.sum_lvl2_ff\[29\] clknet_leaf_60_clk sg13g2_dfrbpq_1
X_4494_ _1266_ _1259_ _1268_ VPWR VGND sg13g2_xor2_1
X_6233_ net1124 VGND VPWR _0241_ DP_3.matrix\[77\] clknet_leaf_35_clk sg13g2_dfrbpq_2
X_3445_ _3019_ _3020_ _3022_ _3023_ VPWR VGND sg13g2_nor3_1
X_6164_ net1117 VGND VPWR _0193_ DP_1.matrix\[77\] clknet_leaf_58_clk sg13g2_dfrbpq_2
X_3376_ _2939_ VPWR _2960_ VGND _2936_ _2940_ sg13g2_o21ai_1
X_5115_ VGND VPWR _1857_ _1858_ _1861_ _1839_ sg13g2_a21oi_1
X_6095_ net1115 VGND VPWR _0113_ mac1.products_ff\[7\] clknet_leaf_57_clk sg13g2_dfrbpq_1
X_5046_ _1792_ _1793_ _1754_ _1794_ VPWR VGND sg13g2_nand3_1
XFILLER_26_735 VPWR VGND sg13g2_fill_2
XFILLER_41_716 VPWR VGND sg13g2_fill_2
X_5948_ _2592_ _2452_ _2455_ VPWR VGND sg13g2_xnor2_1
XFILLER_22_952 VPWR VGND sg13g2_decap_8
XFILLER_43_48 VPWR VGND sg13g2_fill_2
X_5879_ _2530_ VPWR _2533_ VGND net794 _2532_ sg13g2_o21ai_1
XFILLER_21_484 VPWR VGND sg13g2_fill_2
XFILLER_1_823 VPWR VGND sg13g2_decap_8
XFILLER_48_348 VPWR VGND sg13g2_fill_1
XFILLER_1_1005 VPWR VGND sg13g2_decap_8
XFILLER_16_245 VPWR VGND sg13g2_fill_1
XFILLER_9_945 VPWR VGND sg13g2_decap_8
XFILLER_13_996 VPWR VGND sg13g2_decap_8
X_3230_ _2817_ _2818_ _2816_ _2819_ VPWR VGND sg13g2_nand3_1
X_3161_ _2751_ _2713_ _2748_ VPWR VGND sg13g2_xnor2_1
X_3092_ _2684_ _2683_ _2680_ VPWR VGND sg13g2_nand2b_1
X_5802_ _2458_ net800 _2457_ net801 net937 VPWR VGND sg13g2_a22oi_1
X_3994_ _0775_ VPWR _0787_ VGND _0783_ _0785_ sg13g2_o21ai_1
X_5733_ DP_1.I_range.out_data\[4\] _2386_ _2388_ _2390_ VPWR VGND sg13g2_nor3_1
X_5664_ VGND VPWR _2332_ _2334_ _2335_ _2333_ sg13g2_a21oi_1
XFILLER_31_793 VPWR VGND sg13g2_fill_2
X_5595_ _2279_ VPWR _2281_ VGND _2278_ _2280_ sg13g2_o21ai_1
X_4615_ _1380_ net857 net924 net859 net922 VPWR VGND sg13g2_a22oi_1
Xhold411 DP_3.matrix\[7\] VPWR VGND net451 sg13g2_dlygate4sd3_1
Xhold400 DP_2.matrix\[2\] VPWR VGND net440 sg13g2_dlygate4sd3_1
X_4546_ _1318_ _1282_ _1316_ VPWR VGND sg13g2_xnor2_1
Xhold444 mac2.sum_lvl2_ff\[15\] VPWR VGND net484 sg13g2_dlygate4sd3_1
Xhold422 _2119_ VPWR VGND net462 sg13g2_dlygate4sd3_1
XFILLER_2_609 VPWR VGND sg13g2_fill_1
Xhold433 DP_4.matrix\[73\] VPWR VGND net473 sg13g2_dlygate4sd3_1
Xhold455 _2184_ VPWR VGND net495 sg13g2_dlygate4sd3_1
Xhold477 mac2.sum_lvl2_ff\[8\] VPWR VGND net517 sg13g2_dlygate4sd3_1
X_4477_ _1237_ VPWR _1251_ VGND _1226_ _1238_ sg13g2_o21ai_1
Xhold466 _2473_ VPWR VGND net506 sg13g2_dlygate4sd3_1
Xfanout913 net345 net913 VPWR VGND sg13g2_buf_8
Xhold488 DP_1.matrix\[76\] VPWR VGND net528 sg13g2_dlygate4sd3_1
X_3428_ _3008_ net1038 net978 _0069_ VPWR VGND sg13g2_and3_2
X_6216_ net1098 VGND VPWR net71 mac1.sum_lvl1_ff\[12\] clknet_leaf_10_clk sg13g2_dfrbpq_1
Xhold499 DP_3.matrix\[42\] VPWR VGND net539 sg13g2_dlygate4sd3_1
Xfanout902 net339 net902 VPWR VGND sg13g2_buf_8
Xfanout924 net355 net924 VPWR VGND sg13g2_buf_8
Xfanout935 net550 net935 VPWR VGND sg13g2_buf_1
Xfanout946 net491 net946 VPWR VGND sg13g2_buf_8
Xfanout957 net306 net957 VPWR VGND sg13g2_buf_8
X_6147_ net1116 VGND VPWR _0094_ mac1.products_ff\[141\] clknet_leaf_52_clk sg13g2_dfrbpq_1
Xfanout968 net377 net968 VPWR VGND sg13g2_buf_2
X_3359_ _2943_ _2934_ _2944_ VPWR VGND sg13g2_nor2b_1
Xfanout979 net981 net979 VPWR VGND sg13g2_buf_2
X_6078_ net823 _0262_ VPWR VGND sg13g2_buf_1
X_5029_ _1776_ _1753_ _1777_ VPWR VGND sg13g2_xor2_1
XFILLER_26_510 VPWR VGND sg13g2_decap_4
XFILLER_14_749 VPWR VGND sg13g2_fill_2
XFILLER_22_760 VPWR VGND sg13g2_fill_1
XFILLER_10_966 VPWR VGND sg13g2_decap_8
XFILLER_6_937 VPWR VGND sg13g2_decap_8
XFILLER_0_163 VPWR VGND sg13g2_fill_1
XFILLER_23_1028 VPWR VGND sg13g2_fill_1
XFILLER_44_395 VPWR VGND sg13g2_fill_2
XFILLER_13_771 VPWR VGND sg13g2_fill_2
XFILLER_9_742 VPWR VGND sg13g2_fill_1
XFILLER_40_590 VPWR VGND sg13g2_fill_1
X_4400_ _1137_ VPWR _1176_ VGND _1092_ _1138_ sg13g2_o21ai_1
X_5380_ net340 mac1.sum_lvl2_ff\[23\] _2114_ VPWR VGND sg13g2_xor2_1
X_4331_ _1105_ _1106_ _1108_ _1109_ VPWR VGND sg13g2_or3_1
X_4262_ _1038_ _1039_ _1041_ _1042_ VPWR VGND sg13g2_or3_1
X_6001_ _2556_ _2552_ _2626_ VPWR VGND sg13g2_xor2_1
X_3213_ _2797_ VPWR _2802_ VGND _2798_ _2800_ sg13g2_o21ai_1
X_4193_ VGND VPWR _0962_ _0978_ _0979_ _0977_ sg13g2_a21oi_1
X_3144_ _2734_ _2706_ _2735_ VPWR VGND sg13g2_nor2b_1
X_3075_ _2664_ _2665_ _2667_ _2668_ VPWR VGND sg13g2_or3_1
X_3977_ _0770_ net1017 DP_2.matrix\[41\] VPWR VGND sg13g2_nand2_1
XFILLER_11_719 VPWR VGND sg13g2_fill_2
X_5716_ _2377_ _2376_ _2375_ VPWR VGND sg13g2_nand2b_1
X_5647_ _2323_ mac2.sum_lvl3_ff\[34\] net297 VPWR VGND sg13g2_nand2_1
X_5578_ _2266_ VPWR _2269_ VGND _2265_ _2267_ sg13g2_o21ai_1
Xhold230 DP_4.matrix\[75\] VPWR VGND net270 sg13g2_dlygate4sd3_1
Xhold252 mac1.sum_lvl3_ff\[20\] VPWR VGND net292 sg13g2_dlygate4sd3_1
Xhold241 _0179_ VPWR VGND net281 sg13g2_dlygate4sd3_1
X_4529_ _1300_ _1279_ _1302_ VPWR VGND sg13g2_xor2_1
XFILLER_49_25 VPWR VGND sg13g2_fill_1
Xhold296 DP_1.matrix\[0\] VPWR VGND net336 sg13g2_dlygate4sd3_1
Xhold274 DP_1.matrix\[75\] VPWR VGND net314 sg13g2_dlygate4sd3_1
Xhold263 mac1.sum_lvl2_ff\[14\] VPWR VGND net303 sg13g2_dlygate4sd3_1
Xhold285 mac2.sum_lvl3_ff\[0\] VPWR VGND net325 sg13g2_dlygate4sd3_1
Xfanout787 net788 net787 VPWR VGND sg13g2_buf_1
Xfanout798 _2480_ net798 VPWR VGND sg13g2_buf_8
XFILLER_18_329 VPWR VGND sg13g2_fill_2
XFILLER_27_885 VPWR VGND sg13g2_fill_2
XFILLER_14_524 VPWR VGND sg13g2_decap_4
XFILLER_42_888 VPWR VGND sg13g2_fill_1
XFILLER_5_211 VPWR VGND sg13g2_decap_4
XFILLER_6_756 VPWR VGND sg13g2_fill_2
XFILLER_2_973 VPWR VGND sg13g2_decap_8
Xinput9 uio_in[0] net9 VPWR VGND sg13g2_buf_1
XFILLER_18_841 VPWR VGND sg13g2_decap_8
XFILLER_18_896 VPWR VGND sg13g2_decap_8
X_4880_ _1637_ _1634_ _1638_ VPWR VGND sg13g2_xor2_1
X_3900_ _0694_ _0661_ _0695_ VPWR VGND sg13g2_xor2_1
X_3831_ net961 net1018 net965 _0629_ VPWR VGND net1016 sg13g2_nand4_1
X_6550_ net1076 VGND VPWR net3 DP_1.I_range.out_data\[4\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_3762_ _0566_ _0563_ _0108_ VPWR VGND sg13g2_xor2_1
X_5501_ VGND VPWR mac1.sum_lvl3_ff\[33\] mac1.sum_lvl3_ff\[13\] _2209_ _2207_ sg13g2_a21oi_1
X_3693_ _0498_ _0471_ _0500_ VPWR VGND sg13g2_xor2_1
X_6481_ net1085 VGND VPWR _0153_ mac2.products_ff\[149\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_5432_ _0005_ _2152_ net304 VPWR VGND sg13g2_xnor2_1
X_5363_ _2101_ _2095_ _2100_ VPWR VGND sg13g2_xnor2_1
X_4314_ DP_3.matrix\[37\] net835 net907 _1092_ VPWR VGND net833 sg13g2_nand4_1
X_5294_ _2032_ _2034_ _2035_ VPWR VGND sg13g2_nor2_1
X_4245_ _1005_ VPWR _1026_ VGND _0996_ _1006_ sg13g2_o21ai_1
X_4176_ _0951_ _0953_ _0963_ VPWR VGND sg13g2_and2_1
X_3127_ _2689_ VPWR _2718_ VGND _2687_ _2690_ sg13g2_o21ai_1
X_3058_ _2647_ VPWR _2652_ VGND _2648_ _2650_ sg13g2_o21ai_1
Xclkbuf_leaf_62_clk clknet_4_2_0_clk clknet_leaf_62_clk VPWR VGND sg13g2_buf_8
XFILLER_35_181 VPWR VGND sg13g2_fill_2
XFILLER_11_516 VPWR VGND sg13g2_fill_2
XFILLER_11_527 VPWR VGND sg13g2_decap_4
XFILLER_3_704 VPWR VGND sg13g2_fill_2
XFILLER_2_214 VPWR VGND sg13g2_fill_2
XFILLER_46_457 VPWR VGND sg13g2_fill_2
XFILLER_33_107 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_53_clk clknet_4_10_0_clk clknet_leaf_53_clk VPWR VGND sg13g2_buf_8
Xclkbuf_4_6_0_clk clknet_0_clk clknet_4_6_0_clk VPWR VGND sg13g2_buf_8
X_4030_ _0771_ _0820_ _0822_ VPWR VGND sg13g2_and2_1
X_5981_ _2613_ _2511_ net793 VPWR VGND sg13g2_nand2b_1
XFILLER_46_980 VPWR VGND sg13g2_decap_8
X_4932_ _1688_ _1683_ _1686_ VPWR VGND sg13g2_xnor2_1
Xclkbuf_leaf_44_clk clknet_4_14_0_clk clknet_leaf_44_clk VPWR VGND sg13g2_buf_8
XFILLER_17_192 VPWR VGND sg13g2_fill_1
X_4863_ _1594_ _1588_ _1596_ _1621_ VPWR VGND sg13g2_a21o_1
XFILLER_33_696 VPWR VGND sg13g2_fill_2
X_4794_ _1553_ _1502_ _1554_ VPWR VGND sg13g2_xor2_1
X_3814_ _0111_ _0608_ _0615_ VPWR VGND sg13g2_xnor2_1
X_3745_ _0550_ _0544_ _0549_ VPWR VGND sg13g2_xnor2_1
X_6533_ net1105 VGND VPWR net122 mac2.sum_lvl2_ff\[20\] clknet_leaf_31_clk sg13g2_dfrbpq_1
X_6464_ net1141 VGND VPWR _0130_ mac2.products_ff\[80\] clknet_leaf_42_clk sg13g2_dfrbpq_1
X_3676_ _0481_ _0473_ _0483_ VPWR VGND sg13g2_xor2_1
X_5415_ _0002_ _2140_ net367 VPWR VGND sg13g2_xnor2_1
X_6395_ net1112 VGND VPWR net538 mac1.sum_lvl3_ff\[7\] clknet_leaf_57_clk sg13g2_dfrbpq_1
X_5346_ _2085_ _2080_ _2083_ VPWR VGND sg13g2_xnor2_1
XFILLER_0_707 VPWR VGND sg13g2_decap_8
X_5277_ VPWR _2019_ _2018_ VGND sg13g2_inv_1
X_4228_ _1009_ net838 net906 net840 net904 VPWR VGND sg13g2_a22oi_1
XFILLER_29_947 VPWR VGND sg13g2_decap_8
X_4159_ _0947_ _0911_ _0945_ VPWR VGND sg13g2_xnor2_1
XFILLER_43_449 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_35_clk clknet_4_12_0_clk clknet_leaf_35_clk VPWR VGND sg13g2_buf_8
XFILLER_8_818 VPWR VGND sg13g2_fill_2
XFILLER_8_807 VPWR VGND sg13g2_decap_8
XFILLER_7_306 VPWR VGND sg13g2_fill_1
XFILLER_46_221 VPWR VGND sg13g2_fill_1
XFILLER_19_435 VPWR VGND sg13g2_fill_2
XFILLER_36_81 VPWR VGND sg13g2_fill_1
XFILLER_43_972 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_26_clk clknet_4_13_0_clk clknet_leaf_26_clk VPWR VGND sg13g2_buf_8
XFILLER_30_622 VPWR VGND sg13g2_fill_2
Xinput12 uio_in[3] net12 VPWR VGND sg13g2_buf_1
XFILLER_30_688 VPWR VGND sg13g2_fill_2
X_3530_ _0341_ _0338_ _0340_ VPWR VGND sg13g2_nand2_1
XFILLER_7_884 VPWR VGND sg13g2_decap_8
X_3461_ net979 net1034 net985 _0274_ VPWR VGND net1033 sg13g2_nand4_1
X_5200_ _1944_ _1939_ _1943_ VPWR VGND sg13g2_nand2_1
X_6180_ net1063 VGND VPWR net107 mac1.sum_lvl1_ff\[0\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3392_ _2949_ _2951_ _2974_ _2976_ VPWR VGND sg13g2_or3_1
X_5131_ _1876_ net811 net886 net814 net884 VPWR VGND sg13g2_a22oi_1
X_5062_ _1808_ _1775_ _1809_ VPWR VGND sg13g2_xor2_1
X_4013_ _0766_ VPWR _0805_ VGND _0721_ _0767_ sg13g2_o21ai_1
XFILLER_25_405 VPWR VGND sg13g2_fill_1
X_5964_ VGND VPWR net783 _2602_ _0202_ _2601_ sg13g2_a21oi_1
Xclkbuf_leaf_17_clk clknet_4_4_0_clk clknet_leaf_17_clk VPWR VGND sg13g2_buf_8
X_4915_ _1670_ _1669_ _1672_ VPWR VGND sg13g2_xor2_1
XFILLER_34_983 VPWR VGND sg13g2_decap_8
X_5895_ net795 _2547_ _2548_ _2549_ VPWR VGND sg13g2_nor3_1
X_4846_ _1600_ VPWR _1605_ VGND _1602_ _1603_ sg13g2_o21ai_1
XFILLER_20_165 VPWR VGND sg13g2_decap_8
XFILLER_20_176 VPWR VGND sg13g2_fill_1
X_6516_ net1103 VGND VPWR net100 mac2.sum_lvl2_ff\[0\] clknet_leaf_26_clk sg13g2_dfrbpq_1
X_4777_ _1465_ _1535_ _1537_ _1538_ VPWR VGND sg13g2_or3_1
XFILLER_10_1008 VPWR VGND sg13g2_decap_8
X_3728_ VGND VPWR _0497_ _0499_ _0534_ _0531_ sg13g2_a21oi_1
X_3659_ _0467_ _0433_ _0465_ VPWR VGND sg13g2_xnor2_1
X_6447_ net1140 VGND VPWR _0140_ mac2.products_ff\[11\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_6378_ net1131 VGND VPWR net216 mac1.sum_lvl3_ff\[26\] clknet_leaf_52_clk sg13g2_dfrbpq_2
X_5329_ _2068_ VPWR _2069_ VGND _2043_ _2045_ sg13g2_o21ai_1
XFILLER_29_755 VPWR VGND sg13g2_fill_2
XFILLER_17_939 VPWR VGND sg13g2_decap_8
XFILLER_28_265 VPWR VGND sg13g2_fill_2
XFILLER_16_449 VPWR VGND sg13g2_fill_2
XFILLER_19_1000 VPWR VGND sg13g2_decap_8
XFILLER_25_961 VPWR VGND sg13g2_decap_8
XFILLER_24_460 VPWR VGND sg13g2_decap_4
XFILLER_12_644 VPWR VGND sg13g2_fill_1
XFILLER_11_165 VPWR VGND sg13g2_decap_4
XFILLER_4_887 VPWR VGND sg13g2_decap_8
XFILLER_3_397 VPWR VGND sg13g2_fill_1
Xfanout1110 net1113 net1110 VPWR VGND sg13g2_buf_1
Xfanout1132 net1147 net1132 VPWR VGND sg13g2_buf_8
Xfanout1121 net1130 net1121 VPWR VGND sg13g2_buf_8
Xfanout1143 net1144 net1143 VPWR VGND sg13g2_buf_8
XFILLER_23_909 VPWR VGND sg13g2_decap_8
XFILLER_34_246 VPWR VGND sg13g2_fill_1
XFILLER_16_994 VPWR VGND sg13g2_decap_8
X_4700_ _1462_ net851 net925 net854 net922 VPWR VGND sg13g2_a22oi_1
X_5680_ _2345_ VPWR _2348_ VGND _2342_ _2346_ sg13g2_o21ai_1
XFILLER_31_964 VPWR VGND sg13g2_decap_8
X_4631_ _1396_ _1384_ _1395_ VPWR VGND sg13g2_xnor2_1
X_4562_ _1330_ _1308_ _1332_ _1333_ VPWR VGND sg13g2_a21o_1
X_3513_ _0324_ _0323_ _0320_ VPWR VGND sg13g2_nand2b_1
X_6301_ net1115 VGND VPWR net206 mac1.sum_lvl2_ff\[28\] clknet_leaf_59_clk sg13g2_dfrbpq_1
X_4493_ _1266_ _1259_ _1267_ VPWR VGND sg13g2_nor2b_1
X_6232_ net1123 VGND VPWR _0240_ DP_3.matrix\[76\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_3444_ _3022_ net1034 DP_2.matrix\[0\] net1036 DP_2.matrix\[1\] VPWR VGND sg13g2_a22oi_1
Xclkbuf_leaf_6_clk clknet_4_1_0_clk clknet_leaf_6_clk VPWR VGND sg13g2_buf_8
XFILLER_40_0 VPWR VGND sg13g2_fill_2
X_6163_ net1117 VGND VPWR _0192_ DP_1.matrix\[76\] clknet_leaf_58_clk sg13g2_dfrbpq_2
X_3375_ _2942_ _2935_ _2944_ _2959_ VPWR VGND sg13g2_a21o_1
X_5114_ _1857_ _1858_ _1839_ _1860_ VPWR VGND sg13g2_nand3_1
X_6094_ net1109 VGND VPWR _0112_ mac1.products_ff\[6\] clknet_leaf_56_clk sg13g2_dfrbpq_1
X_5045_ _1791_ _1790_ _1773_ _1793_ VPWR VGND sg13g2_a21o_1
XFILLER_14_909 VPWR VGND sg13g2_decap_8
X_5947_ net978 net785 _2591_ VPWR VGND sg13g2_nor2_1
XFILLER_22_931 VPWR VGND sg13g2_decap_8
X_5878_ _2531_ VPWR _2532_ VGND net856 net803 sg13g2_o21ai_1
X_4829_ _1563_ VPWR _1588_ VGND _1561_ _1564_ sg13g2_o21ai_1
XFILLER_49_1015 VPWR VGND sg13g2_decap_8
XFILLER_1_802 VPWR VGND sg13g2_decap_8
XFILLER_1_879 VPWR VGND sg13g2_decap_8
XFILLER_48_327 VPWR VGND sg13g2_fill_1
XFILLER_1_1028 VPWR VGND sg13g2_fill_1
XFILLER_9_924 VPWR VGND sg13g2_decap_8
XFILLER_13_975 VPWR VGND sg13g2_decap_8
XFILLER_40_783 VPWR VGND sg13g2_fill_2
X_3160_ _2713_ _2748_ _2750_ VPWR VGND sg13g2_and2_1
X_3091_ _2682_ _2659_ _2683_ VPWR VGND sg13g2_xor2_1
Xhold1 mac2.sum_lvl1_ff\[46\] VPWR VGND net41 sg13g2_dlygate4sd3_1
XFILLER_35_522 VPWR VGND sg13g2_fill_1
X_5801_ net976 net957 net810 _2457_ VPWR VGND sg13g2_mux2_1
X_3993_ _0775_ _0783_ _0785_ _0786_ VPWR VGND sg13g2_or3_1
X_5732_ DP_1.I_range.out_data\[4\] VPWR _2389_ VGND _2386_ _2388_ sg13g2_o21ai_1
X_5663_ _2334_ _2332_ net27 VPWR VGND sg13g2_xor2_1
X_4614_ _0087_ _1366_ _1378_ VPWR VGND sg13g2_xnor2_1
X_5594_ net502 _2278_ _0057_ VPWR VGND sg13g2_xor2_1
XFILLER_8_990 VPWR VGND sg13g2_decap_8
Xhold401 mac1.sum_lvl3_ff\[3\] VPWR VGND net441 sg13g2_dlygate4sd3_1
X_4545_ _1282_ _1316_ _1317_ VPWR VGND sg13g2_nor2b_1
Xhold434 DP_4.matrix\[1\] VPWR VGND net474 sg13g2_dlygate4sd3_1
Xhold412 DP_2.matrix\[40\] VPWR VGND net452 sg13g2_dlygate4sd3_1
Xhold423 _2122_ VPWR VGND net463 sg13g2_dlygate4sd3_1
Xhold445 _2270_ VPWR VGND net485 sg13g2_dlygate4sd3_1
Xhold456 _2185_ VPWR VGND net496 sg13g2_dlygate4sd3_1
X_4476_ _1223_ _1217_ _1225_ _1250_ VPWR VGND sg13g2_a21o_1
Xhold478 _2240_ VPWR VGND net518 sg13g2_dlygate4sd3_1
Xhold467 _2475_ VPWR VGND net507 sg13g2_dlygate4sd3_1
X_6215_ net1126 VGND VPWR _0227_ DP_3.matrix\[7\] clknet_leaf_36_clk sg13g2_dfrbpq_1
Xfanout914 net915 net914 VPWR VGND sg13g2_buf_8
X_3427_ net1040 net982 _0069_ VPWR VGND sg13g2_and2_1
Xfanout903 DP_3.matrix\[38\] net903 VPWR VGND sg13g2_buf_8
Xfanout925 DP_3.matrix\[0\] net925 VPWR VGND sg13g2_buf_1
Xhold489 DP_3.matrix\[43\] VPWR VGND net529 sg13g2_dlygate4sd3_1
Xfanout936 net937 net936 VPWR VGND sg13g2_buf_8
X_6146_ net1071 VGND VPWR _0181_ DP_1.matrix\[37\] clknet_leaf_65_clk sg13g2_dfrbpq_1
Xfanout958 net959 net958 VPWR VGND sg13g2_buf_2
Xfanout947 net948 net947 VPWR VGND sg13g2_buf_8
X_3358_ _2943_ _2935_ _2942_ VPWR VGND sg13g2_xnor2_1
Xfanout969 net416 net969 VPWR VGND sg13g2_buf_8
X_6077_ net826 _0261_ VPWR VGND sg13g2_buf_1
X_3289_ _2850_ VPWR _2876_ VGND _2844_ _2851_ sg13g2_o21ai_1
X_5028_ _1776_ net883 net820 VPWR VGND sg13g2_nand2_1
XFILLER_10_945 VPWR VGND sg13g2_decap_8
XFILLER_6_916 VPWR VGND sg13g2_decap_8
XFILLER_5_448 VPWR VGND sg13g2_fill_1
XFILLER_0_197 VPWR VGND sg13g2_fill_2
XFILLER_23_1007 VPWR VGND sg13g2_decap_8
XFILLER_17_522 VPWR VGND sg13g2_fill_2
XFILLER_5_982 VPWR VGND sg13g2_decap_8
XFILLER_4_470 VPWR VGND sg13g2_fill_2
X_4330_ _1108_ net891 net848 net894 net845 VPWR VGND sg13g2_a22oi_1
XFILLER_5_75 VPWR VGND sg13g2_fill_1
X_4261_ _1041_ net896 net849 net898 net846 VPWR VGND sg13g2_a22oi_1
X_3212_ _2797_ _2798_ _2800_ _2801_ VPWR VGND sg13g2_or3_1
X_6000_ _2625_ net857 net793 VPWR VGND sg13g2_nand2_1
X_4192_ _0978_ _0962_ _0121_ VPWR VGND sg13g2_xor2_1
X_3143_ _2734_ _2710_ _2733_ VPWR VGND sg13g2_xnor2_1
X_3074_ _2667_ net995 net945 net996 net941 VPWR VGND sg13g2_a22oi_1
XFILLER_39_1014 VPWR VGND sg13g2_decap_8
X_3976_ _0741_ VPWR _0769_ VGND _0732_ _0742_ sg13g2_o21ai_1
X_5715_ VGND VPWR _2376_ mac2.total_sum\[13\] mac1.total_sum\[13\] sg13g2_or2_1
X_5646_ VGND VPWR mac2.sum_lvl3_ff\[33\] net410 _2322_ _2320_ sg13g2_a21oi_1
Xhold220 mac1.sum_lvl1_ff\[43\] VPWR VGND net260 sg13g2_dlygate4sd3_1
X_5577_ _0037_ _2265_ _2268_ VPWR VGND sg13g2_xnor2_1
Xhold253 _0023_ VPWR VGND net293 sg13g2_dlygate4sd3_1
Xhold242 DP_1.matrix\[5\] VPWR VGND net282 sg13g2_dlygate4sd3_1
X_4528_ _1300_ _1279_ _1301_ VPWR VGND sg13g2_nor2b_1
Xhold231 mac2.sum_lvl2_ff\[0\] VPWR VGND net271 sg13g2_dlygate4sd3_1
Xhold286 _0048_ VPWR VGND net326 sg13g2_dlygate4sd3_1
Xhold264 _2155_ VPWR VGND net304 sg13g2_dlygate4sd3_1
Xhold275 mac2.sum_lvl3_ff\[9\] VPWR VGND net315 sg13g2_dlygate4sd3_1
X_4459_ _1229_ VPWR _1234_ VGND _1231_ _1232_ sg13g2_o21ai_1
Xhold297 DP_3.matrix\[40\] VPWR VGND net337 sg13g2_dlygate4sd3_1
X_6129_ net1127 VGND VPWR _0169_ DP_4.matrix\[8\] clknet_leaf_36_clk sg13g2_dfrbpq_2
Xfanout799 _2401_ net799 VPWR VGND sg13g2_buf_8
Xfanout788 _2393_ net788 VPWR VGND sg13g2_buf_2
XFILLER_26_330 VPWR VGND sg13g2_fill_1
XFILLER_26_396 VPWR VGND sg13g2_fill_1
XFILLER_42_856 VPWR VGND sg13g2_fill_1
XFILLER_10_775 VPWR VGND sg13g2_decap_4
XFILLER_2_952 VPWR VGND sg13g2_decap_8
XFILLER_49_455 VPWR VGND sg13g2_fill_1
XFILLER_18_875 VPWR VGND sg13g2_decap_8
XFILLER_45_694 VPWR VGND sg13g2_fill_1
XFILLER_33_834 VPWR VGND sg13g2_fill_2
X_3830_ net962 net958 net1018 net1016 _0628_ VPWR VGND sg13g2_and4_1
XFILLER_33_889 VPWR VGND sg13g2_fill_2
X_3761_ VGND VPWR _0565_ _0566_ _0564_ _0505_ sg13g2_a21oi_2
XFILLER_32_399 VPWR VGND sg13g2_fill_1
X_5500_ net429 _2208_ _0020_ VPWR VGND sg13g2_nor2b_1
X_3692_ _0499_ _0498_ _0471_ VPWR VGND sg13g2_nand2b_1
X_6480_ net1075 VGND VPWR _0152_ mac2.products_ff\[148\] clknet_leaf_22_clk sg13g2_dfrbpq_1
X_5431_ net303 mac1.sum_lvl2_ff\[33\] _2155_ VPWR VGND sg13g2_xor2_1
X_5362_ _2100_ _2086_ _2099_ VPWR VGND sg13g2_xnor2_1
X_4313_ _1091_ net833 net907 net835 net904 VPWR VGND sg13g2_a22oi_1
X_5293_ _2034_ net812 net876 net814 net874 VPWR VGND sg13g2_a22oi_1
X_4244_ _1025_ _1013_ _1024_ VPWR VGND sg13g2_xnor2_1
X_4175_ _0959_ _0937_ _0961_ _0962_ VPWR VGND sg13g2_a21o_1
X_3126_ _2717_ _2712_ _2715_ VPWR VGND sg13g2_xnor2_1
X_3057_ _2647_ _2648_ _2650_ _2651_ VPWR VGND sg13g2_nor3_1
XFILLER_23_300 VPWR VGND sg13g2_fill_1
XFILLER_23_344 VPWR VGND sg13g2_fill_2
XFILLER_23_377 VPWR VGND sg13g2_fill_2
X_3959_ _0753_ _0750_ _0752_ VPWR VGND sg13g2_nand2_1
XFILLER_13_1017 VPWR VGND sg13g2_decap_8
XFILLER_13_1028 VPWR VGND sg13g2_fill_1
X_5629_ mac2.sum_lvl3_ff\[31\] mac2.sum_lvl3_ff\[11\] _2308_ VPWR VGND sg13g2_nor2_1
XFILLER_47_959 VPWR VGND sg13g2_decap_8
XFILLER_18_127 VPWR VGND sg13g2_fill_1
XFILLER_27_650 VPWR VGND sg13g2_decap_8
XFILLER_15_845 VPWR VGND sg13g2_fill_2
XFILLER_42_686 VPWR VGND sg13g2_fill_2
XFILLER_29_1024 VPWR VGND sg13g2_decap_4
XFILLER_1_270 VPWR VGND sg13g2_fill_1
XFILLER_37_403 VPWR VGND sg13g2_fill_1
X_5980_ _2611_ VPWR _0224_ VGND net793 _2612_ sg13g2_o21ai_1
X_4931_ _1687_ _1686_ _1683_ VPWR VGND sg13g2_nand2b_1
X_4862_ _1619_ _1617_ _0139_ VPWR VGND sg13g2_xor2_1
X_3813_ _0615_ _0609_ _0614_ VPWR VGND sg13g2_xnor2_1
X_4793_ _1553_ net919 net854 VPWR VGND sg13g2_nand2_1
X_3744_ _0546_ _0548_ _0549_ VPWR VGND sg13g2_nor2_1
X_6532_ net1103 VGND VPWR net66 mac2.sum_lvl2_ff\[19\] clknet_leaf_30_clk sg13g2_dfrbpq_1
XFILLER_9_381 VPWR VGND sg13g2_fill_2
X_3675_ _0481_ _0473_ _0482_ VPWR VGND sg13g2_nor2b_1
X_6463_ net1134 VGND VPWR _0129_ mac2.products_ff\[79\] clknet_leaf_44_clk sg13g2_dfrbpq_1
X_5414_ _2141_ net366 _2138_ VPWR VGND sg13g2_nand2_1
X_6394_ net1111 VGND VPWR net464 mac1.sum_lvl3_ff\[6\] clknet_leaf_54_clk sg13g2_dfrbpq_1
X_5345_ _2084_ _2083_ _2080_ VPWR VGND sg13g2_nand2b_1
X_5276_ _1985_ _2017_ _1983_ _2018_ VPWR VGND sg13g2_nand3_1
X_4227_ _0082_ _0995_ _1007_ VPWR VGND sg13g2_xnor2_1
X_4158_ _0911_ _0945_ _0946_ VPWR VGND sg13g2_nor2b_1
X_3109_ _2699_ _2698_ _2660_ _2701_ VPWR VGND sg13g2_a21o_1
X_4089_ _0852_ _0846_ _0854_ _0879_ VPWR VGND sg13g2_a21o_1
XFILLER_37_981 VPWR VGND sg13g2_decap_8
XFILLER_46_288 VPWR VGND sg13g2_fill_1
XFILLER_28_981 VPWR VGND sg13g2_decap_8
XFILLER_14_152 VPWR VGND sg13g2_fill_2
Xinput13 uio_in[4] net13 VPWR VGND sg13g2_buf_1
XFILLER_7_863 VPWR VGND sg13g2_decap_8
X_3460_ net985 net981 net1034 net1033 _0273_ VPWR VGND sg13g2_and4_1
X_3391_ _2974_ VPWR _2975_ VGND _2949_ _2951_ sg13g2_o21ai_1
X_5130_ net886 net883 net814 net811 _1875_ VPWR VGND sg13g2_and4_1
X_5061_ _1808_ net880 net820 VPWR VGND sg13g2_nand2_1
X_4012_ _0794_ VPWR _0804_ VGND _0723_ _0795_ sg13g2_o21ai_1
XFILLER_38_756 VPWR VGND sg13g2_fill_1
XFILLER_26_929 VPWR VGND sg13g2_decap_8
X_5963_ _2602_ _2464_ _2466_ VPWR VGND sg13g2_xnor2_1
X_4914_ _1670_ _1669_ _1671_ VPWR VGND sg13g2_nor2b_1
X_5894_ net842 net806 _2548_ VPWR VGND sg13g2_nor2_1
X_4845_ _1600_ _1602_ _1603_ _1604_ VPWR VGND sg13g2_nor3_1
XFILLER_21_656 VPWR VGND sg13g2_fill_2
XFILLER_21_667 VPWR VGND sg13g2_fill_2
X_4776_ VGND VPWR _1533_ _1534_ _1537_ _1499_ sg13g2_a21oi_1
X_3727_ VPWR _0533_ _0532_ VGND sg13g2_inv_1
X_6515_ net1142 VGND VPWR net240 mac2.sum_lvl1_ff\[51\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_3658_ _0466_ _0433_ _0465_ VPWR VGND sg13g2_nand2b_1
X_6446_ net1140 VGND VPWR _0139_ mac2.products_ff\[10\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_6377_ net1132 VGND VPWR net193 mac1.sum_lvl3_ff\[25\] clknet_leaf_52_clk sg13g2_dfrbpq_2
X_3589_ _0398_ net1035 net971 VPWR VGND sg13g2_nand2_1
X_5328_ _2067_ _2053_ _2068_ VPWR VGND sg13g2_xor2_1
X_5259_ _1995_ _2000_ _2001_ VPWR VGND sg13g2_and2_1
Xclkbuf_4_5_0_clk clknet_0_clk clknet_4_5_0_clk VPWR VGND sg13g2_buf_8
XFILLER_17_918 VPWR VGND sg13g2_decap_8
XFILLER_25_940 VPWR VGND sg13g2_decap_8
XFILLER_24_494 VPWR VGND sg13g2_decap_8
XFILLER_11_155 VPWR VGND sg13g2_fill_1
XFILLER_40_987 VPWR VGND sg13g2_decap_8
XFILLER_11_177 VPWR VGND sg13g2_fill_1
XFILLER_4_866 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_fill_2
Xfanout1122 net1125 net1122 VPWR VGND sg13g2_buf_8
Xfanout1111 net1113 net1111 VPWR VGND sg13g2_buf_8
XFILLER_26_1027 VPWR VGND sg13g2_fill_2
Xfanout1100 net1102 net1100 VPWR VGND sg13g2_buf_8
Xfanout1133 net1135 net1133 VPWR VGND sg13g2_buf_8
Xfanout1144 net1146 net1144 VPWR VGND sg13g2_buf_8
XFILLER_39_509 VPWR VGND sg13g2_fill_2
XFILLER_34_203 VPWR VGND sg13g2_fill_1
XFILLER_16_973 VPWR VGND sg13g2_decap_8
X_4630_ _1395_ _1392_ _1394_ VPWR VGND sg13g2_nand2_1
XFILLER_33_1009 VPWR VGND sg13g2_decap_8
X_6300_ net1110 VGND VPWR net139 mac1.sum_lvl2_ff\[27\] clknet_leaf_56_clk sg13g2_dfrbpq_1
X_4561_ _1332_ _1326_ _1331_ VPWR VGND sg13g2_nand2_1
XFILLER_7_693 VPWR VGND sg13g2_fill_1
X_3512_ _0322_ _0289_ _0323_ VPWR VGND sg13g2_xor2_1
X_4492_ _1266_ _1260_ _1265_ VPWR VGND sg13g2_xnor2_1
X_6231_ net1104 VGND VPWR _0239_ DP_3.matrix\[75\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_3443_ net978 net1036 net982 _3021_ VPWR VGND net1034 sg13g2_nand4_1
X_6162_ net1133 VGND VPWR _0095_ mac1.products_ff\[146\] clknet_leaf_48_clk sg13g2_dfrbpq_1
X_5113_ _1859_ _1839_ _1857_ _1858_ VPWR VGND sg13g2_and3_1
X_3374_ _2958_ _2955_ _0097_ VPWR VGND sg13g2_xor2_1
XFILLER_33_0 VPWR VGND sg13g2_fill_1
X_6093_ net1109 VGND VPWR _0105_ mac1.products_ff\[5\] clknet_leaf_56_clk sg13g2_dfrbpq_1
X_5044_ _1790_ _1791_ _1773_ _1792_ VPWR VGND sg13g2_nand3_1
XFILLER_26_704 VPWR VGND sg13g2_fill_2
X_5946_ net785 net982 _0196_ VPWR VGND sg13g2_xor2_1
XFILLER_22_910 VPWR VGND sg13g2_decap_8
X_5877_ _2531_ net804 net837 VPWR VGND sg13g2_nand2b_1
X_4828_ _1555_ VPWR _1587_ VGND _1502_ _1553_ sg13g2_o21ai_1
XFILLER_22_987 VPWR VGND sg13g2_decap_8
XFILLER_21_475 VPWR VGND sg13g2_fill_1
XFILLER_21_486 VPWR VGND sg13g2_fill_1
X_4759_ net867 net866 net909 net1049 _1520_ VPWR VGND sg13g2_and4_1
X_6429_ net1065 VGND VPWR net511 mac1.total_sum\[9\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_49_807 VPWR VGND sg13g2_fill_2
XFILLER_1_858 VPWR VGND sg13g2_decap_8
XFILLER_17_715 VPWR VGND sg13g2_fill_2
XFILLER_32_729 VPWR VGND sg13g2_fill_2
XFILLER_9_903 VPWR VGND sg13g2_decap_8
XFILLER_13_954 VPWR VGND sg13g2_decap_8
XFILLER_40_795 VPWR VGND sg13g2_fill_2
XFILLER_3_173 VPWR VGND sg13g2_fill_2
XFILLER_39_317 VPWR VGND sg13g2_fill_2
X_3090_ _2682_ net999 net934 VPWR VGND sg13g2_nand2_1
Xhold2 mac1.sum_lvl1_ff\[47\] VPWR VGND net42 sg13g2_dlygate4sd3_1
XFILLER_48_840 VPWR VGND sg13g2_fill_2
X_3992_ VGND VPWR _0781_ _0782_ _0785_ _0776_ sg13g2_a21oi_1
X_5800_ _2452_ _2455_ _2456_ VPWR VGND sg13g2_and2_1
XFILLER_22_206 VPWR VGND sg13g2_decap_8
XFILLER_23_718 VPWR VGND sg13g2_decap_4
XFILLER_23_729 VPWR VGND sg13g2_fill_2
X_5731_ DP_1.Q_range.out_data\[3\] DP_1.I_range.out_data\[3\] _2388_ VPWR VGND sg13g2_nor2b_1
X_5662_ mac2.total_sum\[2\] mac1.total_sum\[2\] _2334_ VPWR VGND sg13g2_xor2_1
XFILLER_31_784 VPWR VGND sg13g2_fill_1
XFILLER_31_795 VPWR VGND sg13g2_fill_1
X_5593_ _2280_ mac2.sum_lvl3_ff\[23\] net501 VPWR VGND sg13g2_xnor2_1
X_4613_ _1379_ _1378_ _1366_ VPWR VGND sg13g2_nand2b_1
Xhold402 _2167_ VPWR VGND net442 sg13g2_dlygate4sd3_1
X_4544_ _1316_ _1311_ _1314_ VPWR VGND sg13g2_xnor2_1
Xhold424 _0012_ VPWR VGND net464 sg13g2_dlygate4sd3_1
Xhold435 mac1.sum_lvl2_ff\[3\] VPWR VGND net475 sg13g2_dlygate4sd3_1
Xhold413 DP_1.matrix\[3\] VPWR VGND net453 sg13g2_dlygate4sd3_1
X_6214_ net1126 VGND VPWR _0226_ DP_3.matrix\[6\] clknet_leaf_36_clk sg13g2_dfrbpq_1
Xhold468 _0245_ VPWR VGND net508 sg13g2_dlygate4sd3_1
Xhold457 _0030_ VPWR VGND net497 sg13g2_dlygate4sd3_1
X_4475_ _1248_ _1246_ _0128_ VPWR VGND sg13g2_xor2_1
Xhold446 _0038_ VPWR VGND net486 sg13g2_dlygate4sd3_1
Xfanout915 net447 net915 VPWR VGND sg13g2_buf_8
X_3426_ _0100_ _3000_ _3007_ VPWR VGND sg13g2_xnor2_1
Xfanout904 net905 net904 VPWR VGND sg13g2_buf_8
Xhold479 _2241_ VPWR VGND net519 sg13g2_dlygate4sd3_1
X_6145_ net1072 VGND VPWR _0180_ DP_1.matrix\[36\] clknet_leaf_2_clk sg13g2_dfrbpq_1
Xfanout937 net482 net937 VPWR VGND sg13g2_buf_8
Xfanout926 net927 net926 VPWR VGND sg13g2_buf_8
Xfanout948 net300 net948 VPWR VGND sg13g2_buf_8
X_3357_ _2942_ _2936_ _2941_ VPWR VGND sg13g2_xnor2_1
X_6076_ net832 _0260_ VPWR VGND sg13g2_buf_1
Xfanout959 net960 net959 VPWR VGND sg13g2_buf_2
X_5027_ _1775_ net883 net818 VPWR VGND sg13g2_nand2_1
X_3288_ _2873_ _2865_ _2875_ VPWR VGND sg13g2_xor2_1
XFILLER_26_523 VPWR VGND sg13g2_fill_2
X_5929_ _2423_ _2421_ _2580_ VPWR VGND sg13g2_xor2_1
XFILLER_16_1015 VPWR VGND sg13g2_decap_8
XFILLER_22_751 VPWR VGND sg13g2_fill_2
XFILLER_10_924 VPWR VGND sg13g2_decap_8
XFILLER_45_810 VPWR VGND sg13g2_fill_2
XFILLER_45_865 VPWR VGND sg13g2_decap_8
XFILLER_45_843 VPWR VGND sg13g2_fill_1
XFILLER_5_961 VPWR VGND sg13g2_decap_8
X_4260_ net846 net898 net848 _1040_ VPWR VGND net896 sg13g2_nand4_1
X_3211_ _2800_ net1055 net943 net986 net938 VPWR VGND sg13g2_a22oi_1
X_4191_ _0976_ _0963_ _0978_ VPWR VGND sg13g2_xor2_1
X_3142_ _2733_ _2730_ _2732_ VPWR VGND sg13g2_nand2_1
X_3073_ net941 net996 net945 _2666_ VPWR VGND net995 sg13g2_nand4_1
XFILLER_36_810 VPWR VGND sg13g2_fill_2
XFILLER_36_821 VPWR VGND sg13g2_fill_1
XFILLER_36_876 VPWR VGND sg13g2_fill_1
X_3975_ _0768_ _0721_ _0767_ VPWR VGND sg13g2_xnor2_1
X_5714_ mac1.total_sum\[13\] mac2.total_sum\[13\] _2375_ VPWR VGND sg13g2_and2_1
X_5645_ net412 _2321_ _0052_ VPWR VGND sg13g2_nor2b_1
XFILLER_3_909 VPWR VGND sg13g2_decap_8
X_5576_ net552 mac2.sum_lvl2_ff\[33\] _2268_ VPWR VGND sg13g2_xor2_1
Xhold210 mac2.sum_lvl1_ff\[13\] VPWR VGND net250 sg13g2_dlygate4sd3_1
Xhold243 _0177_ VPWR VGND net283 sg13g2_dlygate4sd3_1
X_4527_ _1298_ _1297_ _1300_ VPWR VGND sg13g2_xor2_1
Xhold221 mac2.products_ff\[6\] VPWR VGND net261 sg13g2_dlygate4sd3_1
Xhold232 _0032_ VPWR VGND net272 sg13g2_dlygate4sd3_1
Xhold287 DP_4.matrix\[8\] VPWR VGND net327 sg13g2_dlygate4sd3_1
XFILLER_46_1008 VPWR VGND sg13g2_decap_8
Xhold254 mac1.sum_lvl2_ff\[5\] VPWR VGND net294 sg13g2_dlygate4sd3_1
Xhold276 _2302_ VPWR VGND net316 sg13g2_dlygate4sd3_1
Xhold265 _0005_ VPWR VGND net305 sg13g2_dlygate4sd3_1
X_4458_ _1229_ _1231_ _1232_ _1233_ VPWR VGND sg13g2_nor3_1
X_3409_ _2992_ _2985_ _2991_ VPWR VGND sg13g2_nand2_1
Xhold298 DP_3.matrix\[37\] VPWR VGND net338 sg13g2_dlygate4sd3_1
X_6128_ net1106 VGND VPWR _0168_ DP_3.matrix\[80\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_4389_ VGND VPWR _1162_ _1163_ _1166_ _1128_ sg13g2_a21oi_1
XFILLER_46_607 VPWR VGND sg13g2_fill_1
Xfanout789 net507 net789 VPWR VGND sg13g2_buf_8
X_6059_ net892 _0235_ VPWR VGND sg13g2_buf_1
XFILLER_27_876 VPWR VGND sg13g2_decap_4
XFILLER_27_887 VPWR VGND sg13g2_fill_1
XFILLER_42_824 VPWR VGND sg13g2_decap_4
XFILLER_10_743 VPWR VGND sg13g2_fill_1
XFILLER_10_765 VPWR VGND sg13g2_decap_4
XFILLER_2_931 VPWR VGND sg13g2_decap_8
XFILLER_7_1024 VPWR VGND sg13g2_decap_4
XFILLER_18_821 VPWR VGND sg13g2_decap_4
X_3760_ VGND VPWR _0502_ _0532_ _0565_ _0534_ sg13g2_a21oi_1
XFILLER_9_596 VPWR VGND sg13g2_fill_2
XFILLER_9_585 VPWR VGND sg13g2_fill_2
X_3691_ _0496_ _0472_ _0498_ VPWR VGND sg13g2_xor2_1
X_5430_ mac1.sum_lvl2_ff\[33\] mac1.sum_lvl2_ff\[14\] _2154_ VPWR VGND sg13g2_nor2_1
X_5361_ _2099_ _2096_ _2098_ VPWR VGND sg13g2_xnor2_1
X_5292_ VGND VPWR _2033_ _2031_ _2007_ sg13g2_or2_1
XFILLER_5_780 VPWR VGND sg13g2_decap_8
X_4312_ _1067_ VPWR _1090_ VGND _1032_ _1065_ sg13g2_o21ai_1
X_4243_ _1024_ _1021_ _1023_ VPWR VGND sg13g2_nand2_1
X_4174_ _0961_ _0955_ _0960_ VPWR VGND sg13g2_nand2_1
X_3125_ _2716_ _2715_ _2712_ VPWR VGND sg13g2_nand2b_1
X_3056_ _2650_ net997 net946 net999 net942 VPWR VGND sg13g2_a22oi_1
XFILLER_35_183 VPWR VGND sg13g2_fill_1
XFILLER_23_389 VPWR VGND sg13g2_fill_2
X_3958_ _0749_ _0748_ _0718_ _0752_ VPWR VGND sg13g2_a21o_1
X_3889_ _0682_ _0656_ _0685_ VPWR VGND sg13g2_xor2_1
X_5628_ net347 _2304_ _0049_ VPWR VGND sg13g2_xor2_1
X_5559_ _2254_ _2247_ _2251_ VPWR VGND sg13g2_nand2_1
XFILLER_2_216 VPWR VGND sg13g2_fill_1
XFILLER_47_938 VPWR VGND sg13g2_decap_8
XFILLER_46_459 VPWR VGND sg13g2_fill_1
XFILLER_18_139 VPWR VGND sg13g2_fill_1
XFILLER_27_640 VPWR VGND sg13g2_fill_2
XFILLER_15_824 VPWR VGND sg13g2_decap_8
XFILLER_42_621 VPWR VGND sg13g2_fill_2
XFILLER_25_73 VPWR VGND sg13g2_fill_2
XFILLER_30_816 VPWR VGND sg13g2_fill_1
XFILLER_30_838 VPWR VGND sg13g2_fill_2
XFILLER_29_1003 VPWR VGND sg13g2_decap_8
XFILLER_37_426 VPWR VGND sg13g2_fill_1
X_4930_ _1685_ _1659_ _1686_ VPWR VGND sg13g2_xor2_1
XFILLER_33_632 VPWR VGND sg13g2_fill_2
X_4861_ _1617_ _1619_ _1620_ VPWR VGND sg13g2_nor2_1
XFILLER_20_315 VPWR VGND sg13g2_fill_2
X_3812_ _0614_ _0600_ _0613_ VPWR VGND sg13g2_xnor2_1
X_4792_ _1552_ net919 net851 VPWR VGND sg13g2_nand2_1
X_6531_ net1145 VGND VPWR net137 mac2.sum_lvl2_ff\[15\] clknet_leaf_38_clk sg13g2_dfrbpq_1
X_3743_ _0548_ net966 net1031 net969 net1027 VPWR VGND sg13g2_a22oi_1
X_3674_ _0481_ _0474_ _0480_ VPWR VGND sg13g2_xnor2_1
X_6462_ net1133 VGND VPWR _0128_ mac2.products_ff\[78\] clknet_leaf_49_clk sg13g2_dfrbpq_1
X_6393_ net1111 VGND VPWR net296 mac1.sum_lvl3_ff\[5\] clknet_leaf_55_clk sg13g2_dfrbpq_1
X_5413_ _2140_ mac1.sum_lvl2_ff\[30\] mac1.sum_lvl2_ff\[11\] VPWR VGND sg13g2_xnor2_1
X_5344_ _2082_ _2056_ _2083_ VPWR VGND sg13g2_xor2_1
X_5275_ _2015_ _1993_ _2017_ VPWR VGND sg13g2_xor2_1
X_4226_ _1008_ _1007_ _0995_ VPWR VGND sg13g2_nand2b_1
X_4157_ _0945_ _0940_ _0943_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_415 VPWR VGND sg13g2_decap_4
X_3108_ _2698_ _2699_ _2660_ _2700_ VPWR VGND sg13g2_nand3_1
X_4088_ _0877_ _0875_ _0117_ VPWR VGND sg13g2_xor2_1
X_3039_ net1003 net946 _0064_ VPWR VGND sg13g2_and2_1
XFILLER_23_120 VPWR VGND sg13g2_fill_2
XFILLER_24_643 VPWR VGND sg13g2_fill_2
XFILLER_3_536 VPWR VGND sg13g2_fill_2
XFILLER_19_404 VPWR VGND sg13g2_fill_2
XFILLER_4_1027 VPWR VGND sg13g2_fill_2
XFILLER_28_960 VPWR VGND sg13g2_decap_8
XFILLER_43_930 VPWR VGND sg13g2_decap_4
XFILLER_30_624 VPWR VGND sg13g2_fill_1
XFILLER_7_842 VPWR VGND sg13g2_decap_8
XFILLER_11_882 VPWR VGND sg13g2_decap_8
Xinput14 uio_in[5] net14 VPWR VGND sg13g2_buf_1
XFILLER_6_363 VPWR VGND sg13g2_fill_2
X_3390_ _2973_ _2959_ _2974_ VPWR VGND sg13g2_xor2_1
X_5060_ _1807_ net880 net818 VPWR VGND sg13g2_nand2_1
X_4011_ _0799_ VPWR _0803_ VGND _0756_ _0801_ sg13g2_o21ai_1
XFILLER_42_1011 VPWR VGND sg13g2_decap_8
X_5962_ net969 net783 _2601_ VPWR VGND sg13g2_nor2_1
XFILLER_19_993 VPWR VGND sg13g2_decap_8
X_4913_ VGND VPWR _1630_ _1641_ _1670_ _1629_ sg13g2_a21oi_1
X_5893_ net861 net805 _2547_ VPWR VGND sg13g2_nor2_1
X_4844_ _1603_ net910 net860 net911 net858 VPWR VGND sg13g2_a22oi_1
X_4775_ _1533_ _1534_ _1499_ _1536_ VPWR VGND sg13g2_nand3_1
XFILLER_20_189 VPWR VGND sg13g2_fill_1
X_3726_ _0499_ _0531_ _0497_ _0532_ VPWR VGND sg13g2_nand3_1
X_6514_ net1142 VGND VPWR net45 mac2.sum_lvl1_ff\[50\] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_3657_ _0465_ _0434_ _0463_ VPWR VGND sg13g2_xnor2_1
X_6445_ net1140 VGND VPWR _0148_ mac2.products_ff\[9\] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_6376_ net1117 VGND VPWR net136 mac1.sum_lvl3_ff\[24\] clknet_leaf_54_clk sg13g2_dfrbpq_1
X_3588_ _0369_ VPWR _0397_ VGND _0360_ _0370_ sg13g2_o21ai_1
X_5327_ _2065_ _2040_ _2067_ VPWR VGND sg13g2_xor2_1
X_5258_ _1999_ _1996_ _2000_ VPWR VGND sg13g2_xor2_1
X_5189_ _1933_ net878 net816 VPWR VGND sg13g2_nand2_1
X_4209_ _0989_ _0990_ _0991_ _0992_ VPWR VGND sg13g2_nor3_1
XFILLER_29_757 VPWR VGND sg13g2_fill_1
XFILLER_24_451 VPWR VGND sg13g2_fill_1
XFILLER_25_996 VPWR VGND sg13g2_decap_8
XFILLER_40_911 VPWR VGND sg13g2_fill_1
XFILLER_8_617 VPWR VGND sg13g2_fill_1
XFILLER_40_966 VPWR VGND sg13g2_decap_8
XFILLER_20_690 VPWR VGND sg13g2_decap_8
XFILLER_4_845 VPWR VGND sg13g2_decap_8
Xfanout1112 net1113 net1112 VPWR VGND sg13g2_buf_8
XFILLER_26_1006 VPWR VGND sg13g2_decap_8
Xfanout1101 net1102 net1101 VPWR VGND sg13g2_buf_8
Xfanout1134 net1135 net1134 VPWR VGND sg13g2_buf_1
Xfanout1123 net1125 net1123 VPWR VGND sg13g2_buf_1
Xfanout1145 net1146 net1145 VPWR VGND sg13g2_buf_8
XFILLER_47_598 VPWR VGND sg13g2_fill_2
XFILLER_35_738 VPWR VGND sg13g2_fill_2
XFILLER_16_952 VPWR VGND sg13g2_decap_8
XFILLER_8_43 VPWR VGND sg13g2_fill_2
XFILLER_31_999 VPWR VGND sg13g2_decap_8
X_4560_ _1331_ _1304_ _1327_ VPWR VGND sg13g2_nand2_1
X_3511_ _0322_ net1035 net974 VPWR VGND sg13g2_nand2_2
X_4491_ _1264_ _1261_ _1265_ VPWR VGND sg13g2_xor2_1
X_6230_ net1104 VGND VPWR _0238_ DP_3.matrix\[74\] clknet_leaf_26_clk sg13g2_dfrbpq_1
X_3442_ net982 net978 net1036 net1034 _3020_ VPWR VGND sg13g2_and4_1
X_6161_ net1112 VGND VPWR _0191_ DP_1.matrix\[75\] clknet_leaf_57_clk sg13g2_dfrbpq_1
X_3373_ VGND VPWR _2957_ _2958_ _2956_ _2897_ sg13g2_a21oi_2
X_5112_ _1846_ VPWR _1858_ VGND _1854_ _1856_ sg13g2_o21ai_1
X_6092_ net1092 VGND VPWR _0073_ mac1.products_ff\[4\] clknet_leaf_62_clk sg13g2_dfrbpq_1
X_5043_ _1779_ VPWR _1791_ VGND _1787_ _1789_ sg13g2_o21ai_1
XFILLER_38_543 VPWR VGND sg13g2_fill_2
XFILLER_38_576 VPWR VGND sg13g2_fill_1
XFILLER_25_226 VPWR VGND sg13g2_fill_2
X_5945_ _2589_ VPWR _0179_ VGND _2436_ _2590_ sg13g2_o21ai_1
X_5876_ _2530_ net817 net797 VPWR VGND sg13g2_nand2_1
X_4827_ _1575_ VPWR _1586_ VGND _1559_ _1576_ sg13g2_o21ai_1
XFILLER_22_966 VPWR VGND sg13g2_decap_8
X_4758_ _1519_ net861 net911 VPWR VGND sg13g2_nand2_1
X_3709_ _0509_ _0514_ _0515_ VPWR VGND sg13g2_and2_1
X_4689_ _1450_ _1451_ _1433_ _1452_ VPWR VGND sg13g2_nand3_1
X_6428_ net1060 VGND VPWR net497 mac1.total_sum\[8\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_1_837 VPWR VGND sg13g2_decap_8
X_6359_ net1086 VGND VPWR net144 mac2.sum_lvl1_ff\[75\] clknet_leaf_23_clk sg13g2_dfrbpq_1
XFILLER_0_369 VPWR VGND sg13g2_decap_8
XFILLER_1_1019 VPWR VGND sg13g2_decap_8
XFILLER_13_933 VPWR VGND sg13g2_decap_8
XFILLER_9_959 VPWR VGND sg13g2_decap_8
XFILLER_12_487 VPWR VGND sg13g2_fill_1
XFILLER_40_785 VPWR VGND sg13g2_fill_1
XFILLER_8_447 VPWR VGND sg13g2_fill_2
Xhold3 mac1.products_ff\[138\] VPWR VGND net43 sg13g2_dlygate4sd3_1
X_3991_ _0781_ _0782_ _0776_ _0784_ VPWR VGND sg13g2_nand3_1
XFILLER_23_708 VPWR VGND sg13g2_fill_2
X_5730_ DP_1.Q_range.out_data\[3\] DP_1.Q_range.out_data\[5\] _2387_ VPWR VGND DP_1.I_range.out_data\[3\]
+ sg13g2_nand3b_1
XFILLER_31_730 VPWR VGND sg13g2_fill_2
X_5661_ mac1.total_sum\[2\] mac2.total_sum\[2\] _2333_ VPWR VGND sg13g2_and2_1
X_5592_ _2279_ mac2.sum_lvl3_ff\[23\] mac2.sum_lvl3_ff\[3\] VPWR VGND sg13g2_nand2_1
Xclkbuf_4_4_0_clk clknet_0_clk clknet_4_4_0_clk VPWR VGND sg13g2_buf_8
X_4612_ _1377_ _1367_ _1378_ VPWR VGND sg13g2_xor2_1
X_4543_ _1315_ _1314_ _1311_ VPWR VGND sg13g2_nand2b_1
Xhold436 _2111_ VPWR VGND net476 sg13g2_dlygate4sd3_1
Xhold403 _0025_ VPWR VGND net443 sg13g2_dlygate4sd3_1
Xhold414 mac2.sum_lvl3_ff\[27\] VPWR VGND net454 sg13g2_dlygate4sd3_1
Xhold425 mac1.sum_lvl2_ff\[13\] VPWR VGND net465 sg13g2_dlygate4sd3_1
Xhold469 mac1.sum_lvl3_ff\[9\] VPWR VGND net509 sg13g2_dlygate4sd3_1
X_4474_ _1246_ _1248_ _1249_ VPWR VGND sg13g2_nor2_1
X_6213_ net1121 VGND VPWR net134 mac1.sum_lvl1_ff\[11\] clknet_leaf_31_clk sg13g2_dfrbpq_1
Xhold447 mac2.sum_lvl3_ff\[26\] VPWR VGND net487 sg13g2_dlygate4sd3_1
Xhold458 mac2.sum_lvl3_ff\[2\] VPWR VGND net498 sg13g2_dlygate4sd3_1
Xfanout916 net420 net916 VPWR VGND sg13g2_buf_8
X_3425_ _3007_ _3001_ _3006_ VPWR VGND sg13g2_xnor2_1
Xfanout905 net338 net905 VPWR VGND sg13g2_buf_8
X_6144_ net1116 VGND VPWR _0068_ mac1.products_ff\[140\] clknet_leaf_53_clk sg13g2_dfrbpq_1
Xfanout938 net939 net938 VPWR VGND sg13g2_buf_2
Xfanout927 net523 net927 VPWR VGND sg13g2_buf_8
Xfanout949 DP_2.matrix\[42\] net949 VPWR VGND sg13g2_buf_8
X_3356_ _2938_ _2940_ _2941_ VPWR VGND sg13g2_nor2_1
X_3287_ _2873_ _2865_ _2874_ VPWR VGND sg13g2_nor2b_1
X_6075_ net833 _0259_ VPWR VGND sg13g2_buf_1
X_5026_ _1774_ net889 net816 VPWR VGND sg13g2_nand2_1
X_5928_ net1036 net785 _2579_ VPWR VGND sg13g2_nor2_1
XFILLER_41_538 VPWR VGND sg13g2_fill_1
XFILLER_10_903 VPWR VGND sg13g2_decap_8
X_5859_ _2513_ VPWR _2514_ VGND net913 net803 sg13g2_o21ai_1
XFILLER_1_678 VPWR VGND sg13g2_fill_2
XFILLER_0_155 VPWR VGND sg13g2_fill_2
XFILLER_0_199 VPWR VGND sg13g2_fill_1
XFILLER_45_800 VPWR VGND sg13g2_fill_2
XFILLER_45_833 VPWR VGND sg13g2_fill_2
XFILLER_5_940 VPWR VGND sg13g2_decap_8
X_3210_ net938 net986 net943 _2799_ VPWR VGND net1054 sg13g2_nand4_1
X_4190_ _0963_ _0976_ _0977_ VPWR VGND sg13g2_nor2_1
X_3141_ _2729_ _2728_ _2711_ _2732_ VPWR VGND sg13g2_a21o_1
XFILLER_39_159 VPWR VGND sg13g2_fill_2
X_3072_ net945 net941 net996 net995 _2665_ VPWR VGND sg13g2_and4_1
X_3974_ _0767_ _0758_ _0765_ VPWR VGND sg13g2_xnor2_1
X_5713_ _2368_ VPWR _2374_ VGND _2369_ _2373_ sg13g2_o21ai_1
X_5644_ _2317_ net411 _2312_ _2321_ VPWR VGND sg13g2_nand3_1
X_5575_ mac2.sum_lvl2_ff\[33\] mac2.sum_lvl2_ff\[14\] _2267_ VPWR VGND sg13g2_nor2_1
Xhold211 mac2.sum_lvl1_ff\[12\] VPWR VGND net251 sg13g2_dlygate4sd3_1
Xhold200 mac2.products_ff\[83\] VPWR VGND net240 sg13g2_dlygate4sd3_1
Xhold233 DP_3.matrix\[80\] VPWR VGND net273 sg13g2_dlygate4sd3_1
Xhold222 mac1.sum_lvl1_ff\[46\] VPWR VGND net262 sg13g2_dlygate4sd3_1
X_4526_ _1298_ _1297_ _1299_ VPWR VGND sg13g2_nor2b_1
Xhold244 mac1.sum_lvl2_ff\[15\] VPWR VGND net284 sg13g2_dlygate4sd3_1
Xhold266 DP_2.matrix\[38\] VPWR VGND net306 sg13g2_dlygate4sd3_1
Xhold255 _2117_ VPWR VGND net295 sg13g2_dlygate4sd3_1
Xhold277 _0063_ VPWR VGND net317 sg13g2_dlygate4sd3_1
X_4457_ _1232_ net893 net841 net895 net838 VPWR VGND sg13g2_a22oi_1
Xhold288 DP_1.matrix\[36\] VPWR VGND net328 sg13g2_dlygate4sd3_1
X_3408_ _2991_ _2986_ _2989_ VPWR VGND sg13g2_xnor2_1
Xhold299 DP_3.matrix\[38\] VPWR VGND net339 sg13g2_dlygate4sd3_1
X_4388_ _1162_ _1163_ _1128_ _1165_ VPWR VGND sg13g2_nand3_1
X_6127_ net1127 VGND VPWR _0167_ DP_3.matrix\[44\] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_3339_ VPWR _2925_ _2924_ VGND sg13g2_inv_1
XFILLER_27_811 VPWR VGND sg13g2_decap_8
X_6058_ net894 _0234_ VPWR VGND sg13g2_buf_1
XFILLER_39_671 VPWR VGND sg13g2_fill_1
X_5009_ _1758_ net883 net822 VPWR VGND sg13g2_nand2_1
XFILLER_45_129 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_65_clk clknet_4_2_0_clk clknet_leaf_65_clk VPWR VGND sg13g2_buf_8
XFILLER_42_814 VPWR VGND sg13g2_fill_1
XFILLER_26_376 VPWR VGND sg13g2_fill_2
XFILLER_6_726 VPWR VGND sg13g2_fill_2
XFILLER_2_910 VPWR VGND sg13g2_decap_8
XFILLER_49_413 VPWR VGND sg13g2_fill_1
XFILLER_7_1003 VPWR VGND sg13g2_decap_8
XFILLER_2_987 VPWR VGND sg13g2_decap_8
XFILLER_18_800 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_56_clk clknet_4_8_0_clk clknet_leaf_56_clk VPWR VGND sg13g2_buf_8
XFILLER_17_354 VPWR VGND sg13g2_fill_2
XFILLER_44_151 VPWR VGND sg13g2_fill_1
X_3690_ _0497_ _0472_ _0496_ VPWR VGND sg13g2_nand2_1
X_5360_ _2097_ _2081_ _2098_ VPWR VGND sg13g2_xor2_1
X_5291_ net876 net874 net815 net812 _2032_ VPWR VGND sg13g2_and4_1
X_4311_ _1081_ VPWR _1089_ VGND _1061_ _1082_ sg13g2_o21ai_1
X_4242_ _1020_ _1019_ _1014_ _1023_ VPWR VGND sg13g2_a21o_1
X_4173_ _0960_ _0933_ _0956_ VPWR VGND sg13g2_nand2_1
XFILLER_49_980 VPWR VGND sg13g2_decap_8
X_3124_ _2714_ _2681_ _2715_ VPWR VGND sg13g2_xor2_1
X_3055_ net942 net999 net946 _2649_ VPWR VGND net996 sg13g2_nand4_1
Xclkbuf_leaf_47_clk clknet_4_9_0_clk clknet_leaf_47_clk VPWR VGND sg13g2_buf_8
XFILLER_35_162 VPWR VGND sg13g2_fill_1
X_3957_ VGND VPWR _0748_ _0749_ _0751_ _0718_ sg13g2_a21oi_1
XFILLER_23_379 VPWR VGND sg13g2_fill_1
X_3888_ VGND VPWR _0680_ _0681_ _0684_ _0656_ sg13g2_a21oi_1
X_5627_ _2307_ _2304_ net347 VPWR VGND sg13g2_nand2_1
X_5558_ _2253_ mac2.sum_lvl2_ff\[30\] mac2.sum_lvl2_ff\[11\] VPWR VGND sg13g2_xnor2_1
X_4509_ VGND VPWR _1282_ _1281_ _1230_ sg13g2_or2_1
X_5489_ _2199_ mac1.sum_lvl3_ff\[32\] mac1.sum_lvl3_ff\[12\] VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_38_clk clknet_4_15_0_clk clknet_leaf_38_clk VPWR VGND sg13g2_buf_8
XFILLER_15_803 VPWR VGND sg13g2_decap_8
XFILLER_25_30 VPWR VGND sg13g2_fill_2
XFILLER_15_847 VPWR VGND sg13g2_fill_1
XFILLER_1_250 VPWR VGND sg13g2_decap_4
XFILLER_49_221 VPWR VGND sg13g2_fill_2
XFILLER_49_298 VPWR VGND sg13g2_fill_1
XFILLER_49_276 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_29_clk clknet_4_6_0_clk clknet_leaf_29_clk VPWR VGND sg13g2_buf_8
XFILLER_46_994 VPWR VGND sg13g2_decap_8
XFILLER_18_696 VPWR VGND sg13g2_fill_1
XFILLER_36_1008 VPWR VGND sg13g2_decap_8
X_4860_ VGND VPWR _1618_ _1619_ _1584_ _1544_ sg13g2_a21oi_2
X_3811_ _0613_ _0610_ _0612_ VPWR VGND sg13g2_xnor2_1
X_6530_ net1145 VGND VPWR net117 mac2.sum_lvl2_ff\[14\] clknet_leaf_38_clk sg13g2_dfrbpq_2
X_4791_ _1551_ net922 net1044 VPWR VGND sg13g2_nand2_1
X_3742_ VGND VPWR _0547_ _0545_ _0521_ sg13g2_or2_1
X_3673_ _0479_ _0475_ _0480_ VPWR VGND sg13g2_xor2_1
X_6461_ net1133 VGND VPWR _0137_ mac2.products_ff\[77\] clknet_leaf_48_clk sg13g2_dfrbpq_1
X_6392_ net1111 VGND VPWR net342 mac1.sum_lvl3_ff\[4\] clknet_leaf_55_clk sg13g2_dfrbpq_1
X_5412_ mac1.sum_lvl2_ff\[30\] mac1.sum_lvl2_ff\[11\] _2139_ VPWR VGND sg13g2_nor2_1
X_5343_ _2082_ net815 net1046 VPWR VGND sg13g2_nand2_1
X_5274_ _2015_ _1993_ _2016_ VPWR VGND sg13g2_nor2b_1
X_4225_ _1006_ _0996_ _1007_ VPWR VGND sg13g2_xor2_1
X_4156_ _0944_ _0943_ _0940_ VPWR VGND sg13g2_nand2b_1
X_3107_ _2697_ _2696_ _2679_ _2699_ VPWR VGND sg13g2_a21o_1
XFILLER_28_449 VPWR VGND sg13g2_decap_8
X_4087_ _0875_ _0877_ _0878_ VPWR VGND sg13g2_nor2_1
X_3038_ VPWR _2635_ net850 VGND sg13g2_inv_1
XFILLER_23_110 VPWR VGND sg13g2_fill_2
XFILLER_12_806 VPWR VGND sg13g2_decap_8
X_4989_ _1739_ net889 net820 VPWR VGND sg13g2_nand2_1
XFILLER_24_699 VPWR VGND sg13g2_decap_8
XFILLER_20_850 VPWR VGND sg13g2_fill_1
XFILLER_20_894 VPWR VGND sg13g2_decap_8
XFILLER_11_76 VPWR VGND sg13g2_fill_1
XFILLER_4_1006 VPWR VGND sg13g2_decap_8
XFILLER_47_747 VPWR VGND sg13g2_fill_1
XFILLER_19_449 VPWR VGND sg13g2_fill_2
XFILLER_43_986 VPWR VGND sg13g2_decap_8
XFILLER_30_636 VPWR VGND sg13g2_fill_2
XFILLER_11_861 VPWR VGND sg13g2_decap_8
Xinput15 uio_in[6] net15 VPWR VGND sg13g2_buf_1
XFILLER_7_898 VPWR VGND sg13g2_decap_8
X_4010_ _0801_ _0756_ _0125_ VPWR VGND sg13g2_xor2_1
XFILLER_28_4 VPWR VGND sg13g2_fill_1
X_5961_ VGND VPWR net783 _2600_ _0201_ _2599_ sg13g2_a21oi_1
XFILLER_19_972 VPWR VGND sg13g2_decap_8
X_4912_ _1667_ _1655_ _1669_ VPWR VGND sg13g2_xor2_1
X_5892_ _2541_ _2545_ _2546_ VPWR VGND sg13g2_and2_1
XFILLER_34_997 VPWR VGND sg13g2_decap_8
X_4843_ net860 net858 net911 net908 _1602_ VPWR VGND sg13g2_and4_1
XFILLER_20_102 VPWR VGND sg13g2_fill_2
XFILLER_21_658 VPWR VGND sg13g2_fill_1
X_4774_ _1535_ _1499_ _1533_ _1534_ VPWR VGND sg13g2_and3_1
X_3725_ _0529_ _0507_ _0531_ VPWR VGND sg13g2_xor2_1
X_6513_ net1141 VGND VPWR net178 mac2.sum_lvl1_ff\[49\] clknet_leaf_41_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_9_clk clknet_4_3_0_clk clknet_leaf_9_clk VPWR VGND sg13g2_buf_8
X_6444_ net1140 VGND VPWR _0147_ mac2.products_ff\[8\] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_3656_ _0464_ _0434_ _0463_ VPWR VGND sg13g2_nand2_1
X_6375_ net1071 VGND VPWR net161 mac1.sum_lvl3_ff\[23\] clknet_leaf_66_clk sg13g2_dfrbpq_1
X_3587_ _0396_ _0349_ _0395_ VPWR VGND sg13g2_xnor2_1
X_5326_ _2040_ _2065_ _2066_ VPWR VGND sg13g2_nor2_1
X_5257_ _1999_ _1973_ _1997_ VPWR VGND sg13g2_xnor2_1
X_4208_ _0991_ net902 net850 net847 net905 VPWR VGND sg13g2_a22oi_1
X_5188_ _1898_ VPWR _1932_ VGND _1889_ _1899_ sg13g2_o21ai_1
X_4139_ _0927_ _0926_ _0928_ VPWR VGND sg13g2_nor2b_1
XFILLER_16_419 VPWR VGND sg13g2_fill_1
XFILLER_19_1014 VPWR VGND sg13g2_decap_8
XFILLER_25_975 VPWR VGND sg13g2_decap_8
XFILLER_4_824 VPWR VGND sg13g2_decap_8
XFILLER_0_2 VPWR VGND sg13g2_fill_1
Xfanout1113 net1130 net1113 VPWR VGND sg13g2_buf_8
Xfanout1102 net1107 net1102 VPWR VGND sg13g2_buf_8
Xfanout1124 net1125 net1124 VPWR VGND sg13g2_buf_8
Xfanout1135 net1147 net1135 VPWR VGND sg13g2_buf_8
Xfanout1146 net1147 net1146 VPWR VGND sg13g2_buf_8
XFILLER_47_83 VPWR VGND sg13g2_fill_2
XFILLER_19_257 VPWR VGND sg13g2_fill_2
XFILLER_16_931 VPWR VGND sg13g2_decap_8
XFILLER_42_282 VPWR VGND sg13g2_fill_2
XFILLER_31_978 VPWR VGND sg13g2_decap_8
XFILLER_8_55 VPWR VGND sg13g2_fill_2
XFILLER_7_640 VPWR VGND sg13g2_fill_1
X_3510_ _0321_ net1035 net972 VPWR VGND sg13g2_nand2_1
X_4490_ _1264_ _1219_ _1262_ VPWR VGND sg13g2_xnor2_1
X_3441_ _3019_ net1038 net976 VPWR VGND sg13g2_nand2_1
X_6160_ net1112 VGND VPWR _0190_ DP_1.matrix\[74\] clknet_leaf_58_clk sg13g2_dfrbpq_1
X_3372_ VGND VPWR _2894_ _2924_ _2957_ _2926_ sg13g2_a21oi_1
X_5111_ _1846_ _1854_ _1856_ _1857_ VPWR VGND sg13g2_or3_1
X_6091_ net1071 VGND VPWR _0072_ mac1.products_ff\[3\] clknet_leaf_64_clk sg13g2_dfrbpq_1
X_5042_ _1779_ _1787_ _1789_ _1790_ VPWR VGND sg13g2_or3_1
XFILLER_38_566 VPWR VGND sg13g2_fill_2
XFILLER_38_588 VPWR VGND sg13g2_fill_1
X_5944_ _2432_ _2435_ _2590_ VPWR VGND sg13g2_nor2b_1
X_5875_ VGND VPWR _2522_ _2527_ _0166_ _2529_ sg13g2_a21oi_1
XFILLER_22_945 VPWR VGND sg13g2_decap_8
X_4826_ VGND VPWR _1550_ _1556_ _1585_ _1558_ sg13g2_a21oi_1
X_4757_ _1478_ VPWR _1518_ VGND _1476_ _1479_ sg13g2_o21ai_1
X_3708_ _0513_ _0510_ _0514_ VPWR VGND sg13g2_xor2_1
X_4688_ _1449_ _1448_ _1439_ _1451_ VPWR VGND sg13g2_a21o_1
X_3639_ _0447_ net1032 net971 VPWR VGND sg13g2_nand2_1
X_6427_ net1060 VGND VPWR _0029_ mac1.total_sum\[7\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_1_816 VPWR VGND sg13g2_decap_8
X_6358_ net1100 VGND VPWR net67 mac2.sum_lvl1_ff\[74\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_5309_ VGND VPWR _1987_ _2018_ _2050_ _2020_ sg13g2_a21oi_1
X_6289_ net1099 VGND VPWR net197 mac1.sum_lvl2_ff\[13\] clknet_leaf_29_clk sg13g2_dfrbpq_1
XFILLER_17_717 VPWR VGND sg13g2_fill_1
XFILLER_16_238 VPWR VGND sg13g2_fill_2
XFILLER_29_599 VPWR VGND sg13g2_fill_2
XFILLER_13_912 VPWR VGND sg13g2_decap_8
XFILLER_9_938 VPWR VGND sg13g2_decap_8
XFILLER_13_989 VPWR VGND sg13g2_decap_8
XFILLER_3_120 VPWR VGND sg13g2_fill_2
XFILLER_3_131 VPWR VGND sg13g2_fill_1
XFILLER_3_175 VPWR VGND sg13g2_fill_1
Xhold4 mac2.sum_lvl1_ff\[87\] VPWR VGND net44 sg13g2_dlygate4sd3_1
XFILLER_0_882 VPWR VGND sg13g2_decap_8
XFILLER_39_319 VPWR VGND sg13g2_fill_1
XFILLER_35_503 VPWR VGND sg13g2_fill_2
X_3990_ _0783_ _0776_ _0781_ _0782_ VPWR VGND sg13g2_and3_1
X_5660_ _2329_ VPWR _2332_ VGND _2328_ _2330_ sg13g2_o21ai_1
X_4611_ _1377_ _1368_ _1375_ VPWR VGND sg13g2_xnor2_1
X_5591_ VGND VPWR _2275_ _2277_ _2278_ _2276_ sg13g2_a21oi_1
X_4542_ _1313_ _1287_ _1314_ VPWR VGND sg13g2_xor2_1
X_4473_ VGND VPWR _1247_ _1248_ _1213_ _1173_ sg13g2_a21oi_2
Xhold426 _2150_ VPWR VGND net466 sg13g2_dlygate4sd3_1
Xhold415 _2292_ VPWR VGND net455 sg13g2_dlygate4sd3_1
Xhold404 mac2.sum_lvl3_ff\[4\] VPWR VGND net444 sg13g2_dlygate4sd3_1
X_6212_ net1128 VGND VPWR _0225_ DP_3.matrix\[5\] clknet_leaf_36_clk sg13g2_dfrbpq_2
Xhold437 _0009_ VPWR VGND net477 sg13g2_dlygate4sd3_1
X_3424_ _3006_ _2992_ _3005_ VPWR VGND sg13g2_xnor2_1
Xhold448 _2288_ VPWR VGND net488 sg13g2_dlygate4sd3_1
Xhold459 _2277_ VPWR VGND net499 sg13g2_dlygate4sd3_1
Xfanout906 net349 net906 VPWR VGND sg13g2_buf_8
Xfanout917 DP_3.matrix\[4\] net917 VPWR VGND sg13g2_buf_8
Xfanout939 net940 net939 VPWR VGND sg13g2_buf_1
Xfanout928 net929 net928 VPWR VGND sg13g2_buf_8
X_3355_ _2940_ net926 net991 net928 net990 VPWR VGND sg13g2_a22oi_1
X_6143_ net1095 VGND VPWR net281 DP_1.matrix\[7\] clknet_leaf_61_clk sg13g2_dfrbpq_2
X_3286_ _2873_ _2866_ _2872_ VPWR VGND sg13g2_xnor2_1
X_6074_ net835 _0258_ VPWR VGND sg13g2_buf_1
X_5025_ _1764_ VPWR _1773_ VGND _1756_ _1765_ sg13g2_o21ai_1
X_5927_ VGND VPWR net785 _2578_ _0173_ _2577_ sg13g2_a21oi_1
XFILLER_22_753 VPWR VGND sg13g2_fill_1
X_5858_ _2513_ net803 net895 VPWR VGND sg13g2_nand2b_1
X_4809_ net866 net862 net908 net1050 _1569_ VPWR VGND sg13g2_and4_1
XFILLER_10_959 VPWR VGND sg13g2_decap_8
X_5789_ net974 _2397_ _2445_ VPWR VGND sg13g2_and2_1
XFILLER_5_996 VPWR VGND sg13g2_decap_8
X_3140_ VGND VPWR _2728_ _2729_ _2731_ _2711_ sg13g2_a21oi_1
X_3071_ _2664_ net998 net936 VPWR VGND sg13g2_nand2_1
XFILLER_39_1028 VPWR VGND sg13g2_fill_1
X_3973_ _0766_ _0758_ _0765_ VPWR VGND sg13g2_nand2_1
X_5712_ net21 _2370_ _2373_ VPWR VGND sg13g2_xnor2_1
X_5643_ VGND VPWR _2312_ _2317_ _2320_ net411 sg13g2_a21oi_1
X_5574_ _2266_ mac2.sum_lvl2_ff\[33\] mac2.sum_lvl2_ff\[14\] VPWR VGND sg13g2_nand2_1
Xhold201 mac1.products_ff\[77\] VPWR VGND net241 sg13g2_dlygate4sd3_1
X_4525_ VGND VPWR _1252_ _1257_ _1298_ _1269_ sg13g2_a21oi_1
Xhold234 DP_2.matrix\[44\] VPWR VGND net274 sg13g2_dlygate4sd3_1
Xhold223 mac1.products_ff\[148\] VPWR VGND net263 sg13g2_dlygate4sd3_1
Xhold212 mac2.products_ff\[77\] VPWR VGND net252 sg13g2_dlygate4sd3_1
Xhold278 DP_4.matrix\[77\] VPWR VGND net318 sg13g2_dlygate4sd3_1
Xhold267 DP_3.matrix\[74\] VPWR VGND net307 sg13g2_dlygate4sd3_1
Xhold256 _0011_ VPWR VGND net296 sg13g2_dlygate4sd3_1
Xhold245 _2157_ VPWR VGND net285 sg13g2_dlygate4sd3_1
X_4456_ net841 net839 net895 net893 _1231_ VPWR VGND sg13g2_and4_1
X_3407_ _2990_ _2989_ _2986_ VPWR VGND sg13g2_nand2b_1
X_4387_ _1164_ _1128_ _1162_ _1163_ VPWR VGND sg13g2_and3_1
Xhold289 DP_4.matrix\[38\] VPWR VGND net329 sg13g2_dlygate4sd3_1
X_6126_ net1127 VGND VPWR _0166_ DP_3.matrix\[8\] clknet_leaf_36_clk sg13g2_dfrbpq_1
X_3338_ _2891_ _2923_ _2889_ _2924_ VPWR VGND sg13g2_nand3_1
X_3269_ _2857_ _2826_ _2855_ VPWR VGND sg13g2_xnor2_1
X_6057_ net897 _0233_ VPWR VGND sg13g2_buf_1
X_5008_ _1743_ VPWR _1757_ VGND _1741_ _1744_ sg13g2_o21ai_1
XFILLER_27_845 VPWR VGND sg13g2_decap_4
XFILLER_14_528 VPWR VGND sg13g2_fill_1
XFILLER_2_966 VPWR VGND sg13g2_decap_8
Xclkbuf_4_3_0_clk clknet_0_clk clknet_4_3_0_clk VPWR VGND sg13g2_buf_8
XFILLER_18_834 VPWR VGND sg13g2_decap_8
XFILLER_29_171 VPWR VGND sg13g2_fill_2
XFILLER_17_366 VPWR VGND sg13g2_fill_1
XFILLER_18_889 VPWR VGND sg13g2_decap_8
XFILLER_9_510 VPWR VGND sg13g2_fill_1
X_5290_ _2031_ net874 net812 VPWR VGND sg13g2_nand2_1
X_4310_ _1088_ _1087_ _0134_ VPWR VGND sg13g2_xor2_1
X_4241_ VGND VPWR _1019_ _1020_ _1022_ _1014_ sg13g2_a21oi_1
XFILLER_45_1021 VPWR VGND sg13g2_decap_8
X_4172_ _0934_ _0957_ _0959_ VPWR VGND sg13g2_and2_1
X_3123_ _2714_ net997 net935 VPWR VGND sg13g2_nand2_1
X_3054_ net946 net942 net999 net997 _2648_ VPWR VGND sg13g2_and4_1
X_3956_ _0748_ _0749_ _0718_ _0750_ VPWR VGND sg13g2_nand3_1
X_3887_ _0680_ _0681_ _0656_ _0683_ VPWR VGND sg13g2_nand3_1
X_5626_ net346 mac2.sum_lvl3_ff\[30\] _2306_ VPWR VGND sg13g2_xor2_1
X_5557_ mac2.sum_lvl2_ff\[30\] mac2.sum_lvl2_ff\[11\] _2252_ VPWR VGND sg13g2_nor2_1
X_5488_ _0018_ _2197_ _2198_ VPWR VGND sg13g2_xnor2_1
X_4508_ _1281_ net837 net1048 VPWR VGND sg13g2_nand2_2
X_4439_ VGND VPWR _1179_ _1185_ _1214_ _1187_ sg13g2_a21oi_1
X_6109_ net1090 VGND VPWR _0116_ mac1.products_ff\[73\] clknet_leaf_63_clk sg13g2_dfrbpq_1
XFILLER_27_642 VPWR VGND sg13g2_fill_1
XFILLER_27_664 VPWR VGND sg13g2_fill_1
XFILLER_41_155 VPWR VGND sg13g2_fill_2
XFILLER_23_881 VPWR VGND sg13g2_fill_1
XFILLER_2_752 VPWR VGND sg13g2_fill_1
XFILLER_49_211 VPWR VGND sg13g2_fill_2
XFILLER_2_68 VPWR VGND sg13g2_fill_2
XFILLER_46_973 VPWR VGND sg13g2_decap_8
XFILLER_45_472 VPWR VGND sg13g2_fill_2
X_4790_ _1515_ VPWR _1550_ VGND _1512_ _1516_ sg13g2_o21ai_1
X_3810_ _0611_ _0595_ _0612_ VPWR VGND sg13g2_xor2_1
XFILLER_14_881 VPWR VGND sg13g2_decap_8
X_3741_ net1031 net1027 net969 net966 _0546_ VPWR VGND sg13g2_and4_1
X_3672_ _0479_ _0438_ _0477_ VPWR VGND sg13g2_xnor2_1
X_6460_ net1134 VGND VPWR _0136_ mac2.products_ff\[76\] clknet_leaf_48_clk sg13g2_dfrbpq_1
X_6391_ net1071 VGND VPWR net477 mac1.sum_lvl3_ff\[3\] clknet_leaf_66_clk sg13g2_dfrbpq_1
X_5411_ _0001_ _2136_ _2137_ VPWR VGND sg13g2_xnor2_1
X_5342_ _2081_ net812 net1046 VPWR VGND sg13g2_nand2_1
XFILLER_49_0 VPWR VGND sg13g2_fill_1
XFILLER_5_590 VPWR VGND sg13g2_fill_2
X_5273_ _2015_ _1994_ _2014_ VPWR VGND sg13g2_xnor2_1
X_4224_ _1006_ _0997_ _1004_ VPWR VGND sg13g2_xnor2_1
X_4155_ _0942_ _0916_ _0943_ VPWR VGND sg13g2_xor2_1
X_3106_ _2696_ _2697_ _2679_ _2698_ VPWR VGND sg13g2_nand3_1
X_4086_ VGND VPWR _0876_ _0877_ _0842_ _0802_ sg13g2_a21oi_2
X_3037_ VPWR _2634_ net906 VGND sg13g2_inv_1
XFILLER_37_995 VPWR VGND sg13g2_decap_8
XFILLER_23_122 VPWR VGND sg13g2_fill_1
XFILLER_24_634 VPWR VGND sg13g2_fill_1
XFILLER_23_155 VPWR VGND sg13g2_fill_2
X_4988_ _1737_ _1730_ _0091_ VPWR VGND sg13g2_xor2_1
X_3939_ _0701_ VPWR _0733_ VGND _0699_ _0702_ sg13g2_o21ai_1
X_5609_ _2292_ net454 mac2.sum_lvl3_ff\[7\] VPWR VGND sg13g2_nand2_1
X_6589_ net1080 VGND VPWR net14 DP_3.I_range.out_data\[3\] clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_3_538 VPWR VGND sg13g2_fill_1
XFILLER_19_406 VPWR VGND sg13g2_fill_1
XFILLER_28_995 VPWR VGND sg13g2_decap_8
XFILLER_15_656 VPWR VGND sg13g2_fill_2
XFILLER_35_1020 VPWR VGND sg13g2_decap_8
XFILLER_11_840 VPWR VGND sg13g2_decap_8
Xinput16 uio_in[7] net16 VPWR VGND sg13g2_buf_1
XFILLER_7_877 VPWR VGND sg13g2_decap_8
XFILLER_6_365 VPWR VGND sg13g2_fill_1
XFILLER_19_951 VPWR VGND sg13g2_decap_8
XFILLER_37_225 VPWR VGND sg13g2_fill_1
X_5960_ _2600_ _2444_ _2463_ VPWR VGND sg13g2_xnor2_1
X_4911_ VGND VPWR _1668_ _1667_ _1655_ sg13g2_or2_1
X_5891_ VGND VPWR _2542_ _2543_ _2545_ _2544_ sg13g2_a21oi_1
XFILLER_34_976 VPWR VGND sg13g2_decap_8
X_4842_ _1601_ net858 net908 VPWR VGND sg13g2_nand2_1
XFILLER_21_615 VPWR VGND sg13g2_fill_1
XFILLER_20_136 VPWR VGND sg13g2_decap_4
X_4773_ _1510_ VPWR _1534_ VGND _1530_ _1532_ sg13g2_o21ai_1
X_3724_ _0529_ _0507_ _0530_ VPWR VGND sg13g2_nor2b_1
X_6512_ net1141 VGND VPWR net110 mac2.sum_lvl1_ff\[48\] clknet_leaf_42_clk sg13g2_dfrbpq_1
X_3655_ _0462_ _0445_ _0463_ VPWR VGND sg13g2_xor2_1
X_6443_ net1140 VGND VPWR _0146_ mac2.products_ff\[7\] clknet_leaf_41_clk sg13g2_dfrbpq_1
X_6374_ net1069 VGND VPWR net129 mac1.sum_lvl3_ff\[22\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3586_ _0395_ _0386_ _0393_ VPWR VGND sg13g2_xnor2_1
X_5325_ _2065_ _2025_ _2063_ VPWR VGND sg13g2_xnor2_1
X_5256_ VGND VPWR _1998_ _1997_ _1973_ sg13g2_or2_1
X_4207_ net850 net905 net847 net902 _0990_ VPWR VGND sg13g2_and4_1
X_5187_ _1931_ _1921_ _1929_ VPWR VGND sg13g2_xnor2_1
X_4138_ VGND VPWR _0881_ _0886_ _0927_ _0898_ sg13g2_a21oi_1
XFILLER_29_748 VPWR VGND sg13g2_decap_8
X_4069_ net954 net952 net1008 net1006 _0860_ VPWR VGND sg13g2_and4_1
XFILLER_43_217 VPWR VGND sg13g2_fill_2
XFILLER_25_954 VPWR VGND sg13g2_decap_8
XFILLER_40_957 VPWR VGND sg13g2_fill_1
XFILLER_11_169 VPWR VGND sg13g2_fill_1
Xfanout1103 net1106 net1103 VPWR VGND sg13g2_buf_8
Xfanout1114 net1115 net1114 VPWR VGND sg13g2_buf_8
Xfanout1147 net1148 net1147 VPWR VGND sg13g2_buf_8
Xfanout1136 net1137 net1136 VPWR VGND sg13g2_buf_8
Xfanout1125 net1130 net1125 VPWR VGND sg13g2_buf_8
XFILLER_16_910 VPWR VGND sg13g2_decap_8
XFILLER_15_431 VPWR VGND sg13g2_fill_2
XFILLER_16_987 VPWR VGND sg13g2_decap_8
XFILLER_30_456 VPWR VGND sg13g2_fill_2
XFILLER_8_45 VPWR VGND sg13g2_fill_1
XFILLER_6_162 VPWR VGND sg13g2_fill_1
X_3440_ VGND VPWR _3018_ _3013_ _3011_ sg13g2_or2_1
X_3371_ VGND VPWR _2893_ _2924_ _2956_ _2926_ sg13g2_a21oi_1
X_5110_ VGND VPWR _1852_ _1853_ _1856_ _1847_ sg13g2_a21oi_1
X_6090_ net1070 VGND VPWR _0071_ mac1.products_ff\[2\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_5041_ VGND VPWR _1785_ _1786_ _1789_ _1780_ sg13g2_a21oi_1
XFILLER_38_545 VPWR VGND sg13g2_fill_1
X_5943_ _2589_ net280 net787 VPWR VGND sg13g2_nand2b_1
X_5874_ _2522_ _2528_ _2529_ VPWR VGND sg13g2_nor2_1
XFILLER_22_924 VPWR VGND sg13g2_decap_8
X_4825_ _1584_ _1545_ _0148_ VPWR VGND sg13g2_xor2_1
X_4756_ _1517_ _1512_ _1516_ VPWR VGND sg13g2_xnor2_1
X_3707_ _0513_ _0487_ _0511_ VPWR VGND sg13g2_xnor2_1
X_4687_ _1448_ _1449_ _1439_ _1450_ VPWR VGND sg13g2_nand3_1
XFILLER_49_1008 VPWR VGND sg13g2_decap_8
X_3638_ _0412_ VPWR _0446_ VGND _0403_ _0413_ sg13g2_o21ai_1
X_6426_ net1060 VGND VPWR _0028_ mac1.total_sum\[6\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_3569_ VGND VPWR _0376_ _0377_ _0379_ _0346_ sg13g2_a21oi_1
X_6357_ net1102 VGND VPWR net61 mac2.sum_lvl1_ff\[73\] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_5308_ _2047_ _2046_ _2049_ VPWR VGND sg13g2_xor2_1
X_6288_ net1098 VGND VPWR net204 mac1.sum_lvl2_ff\[12\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_5239_ _1981_ _1969_ _1982_ VPWR VGND sg13g2_xor2_1
XFILLER_17_43 VPWR VGND sg13g2_fill_1
XFILLER_9_917 VPWR VGND sg13g2_decap_8
XFILLER_12_445 VPWR VGND sg13g2_fill_2
XFILLER_13_968 VPWR VGND sg13g2_decap_8
XFILLER_32_1012 VPWR VGND sg13g2_decap_8
XFILLER_8_449 VPWR VGND sg13g2_fill_1
XFILLER_48_821 VPWR VGND sg13g2_fill_2
XFILLER_48_810 VPWR VGND sg13g2_fill_2
XFILLER_0_861 VPWR VGND sg13g2_decap_8
Xhold5 mac2.products_ff\[82\] VPWR VGND net45 sg13g2_dlygate4sd3_1
XFILLER_48_876 VPWR VGND sg13g2_fill_1
XFILLER_48_898 VPWR VGND sg13g2_decap_8
XFILLER_31_732 VPWR VGND sg13g2_fill_1
X_4610_ _1376_ _1368_ _1375_ VPWR VGND sg13g2_nand2_1
XFILLER_12_990 VPWR VGND sg13g2_decap_8
X_5590_ net499 _2275_ _0056_ VPWR VGND sg13g2_xor2_1
XFILLER_8_983 VPWR VGND sg13g2_decap_8
X_4541_ _1313_ net836 net893 VPWR VGND sg13g2_nand2_1
X_4472_ VGND VPWR _1170_ _1212_ _1247_ _1211_ sg13g2_a21oi_1
Xhold427 _2151_ VPWR VGND net467 sg13g2_dlygate4sd3_1
Xhold416 _2299_ VPWR VGND net456 sg13g2_dlygate4sd3_1
Xhold405 _2283_ VPWR VGND net445 sg13g2_dlygate4sd3_1
X_6211_ net1124 VGND VPWR net421 DP_3.matrix\[4\] clknet_leaf_35_clk sg13g2_dfrbpq_2
X_3423_ _3005_ _3003_ _3004_ VPWR VGND sg13g2_xnor2_1
Xhold438 mac1.sum_lvl2_ff\[10\] VPWR VGND net478 sg13g2_dlygate4sd3_1
Xhold449 _2291_ VPWR VGND net489 sg13g2_dlygate4sd3_1
X_6142_ net1095 VGND VPWR net409 DP_1.matrix\[6\] clknet_leaf_8_clk sg13g2_dfrbpq_1
Xfanout907 DP_3.matrix\[36\] net907 VPWR VGND sg13g2_buf_1
Xfanout929 net426 net929 VPWR VGND sg13g2_buf_2
X_3354_ VGND VPWR _2939_ _2937_ _2913_ sg13g2_or2_1
Xfanout918 net387 net918 VPWR VGND sg13g2_buf_8
X_3285_ _2871_ _2867_ _2872_ VPWR VGND sg13g2_xor2_1
X_6073_ net837 _0257_ VPWR VGND sg13g2_buf_1
X_5024_ _1771_ _1751_ _0093_ VPWR VGND sg13g2_xor2_1
XFILLER_38_375 VPWR VGND sg13g2_fill_1
X_5926_ _2578_ _2416_ _2420_ VPWR VGND sg13g2_xnor2_1
X_5857_ _2512_ net279 net797 VPWR VGND sg13g2_nand2_1
X_4808_ _1568_ net861 net1049 VPWR VGND sg13g2_nand2_1
XFILLER_10_938 VPWR VGND sg13g2_decap_8
XFILLER_6_909 VPWR VGND sg13g2_decap_8
X_5788_ _2444_ net799 _2443_ net801 net931 VPWR VGND sg13g2_a22oi_1
X_4739_ _1471_ VPWR _1500_ VGND _1468_ _1472_ sg13g2_o21ai_1
X_6409_ net1084 VGND VPWR net115 mac2.sum_lvl3_ff\[25\] clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_0_157 VPWR VGND sg13g2_fill_1
XFILLER_48_139 VPWR VGND sg13g2_fill_2
XFILLER_28_20 VPWR VGND sg13g2_fill_1
XFILLER_28_75 VPWR VGND sg13g2_fill_1
XFILLER_44_301 VPWR VGND sg13g2_fill_1
XFILLER_5_975 VPWR VGND sg13g2_decap_8
X_3070_ _2649_ VPWR _2663_ VGND _2647_ _2650_ sg13g2_o21ai_1
XFILLER_39_1007 VPWR VGND sg13g2_decap_8
XFILLER_23_529 VPWR VGND sg13g2_fill_2
X_3972_ _0763_ _0759_ _0765_ VPWR VGND sg13g2_xor2_1
X_5711_ VPWR VGND _2372_ _2371_ _2363_ mac1.total_sum\[11\] _2373_ mac2.total_sum\[11\]
+ sg13g2_a221oi_1
X_5642_ _2319_ mac2.sum_lvl3_ff\[33\] net410 VPWR VGND sg13g2_xnor2_1
X_5573_ VGND VPWR _2261_ _2263_ _2265_ _2262_ sg13g2_a21oi_1
Xhold202 mac2.products_ff\[13\] VPWR VGND net242 sg13g2_dlygate4sd3_1
X_4524_ _1295_ _1283_ _1297_ VPWR VGND sg13g2_xor2_1
Xhold235 DP_3.matrix\[72\] VPWR VGND net275 sg13g2_dlygate4sd3_1
Xhold224 mac1.products_ff\[151\] VPWR VGND net264 sg13g2_dlygate4sd3_1
Xhold213 mac1.products_ff\[81\] VPWR VGND net253 sg13g2_dlygate4sd3_1
Xhold246 _0006_ VPWR VGND net286 sg13g2_dlygate4sd3_1
X_4455_ _1230_ net839 net893 VPWR VGND sg13g2_nand2_1
Xhold257 mac2.sum_lvl3_ff\[14\] VPWR VGND net297 sg13g2_dlygate4sd3_1
Xhold268 mac2.sum_lvl2_ff\[19\] VPWR VGND net308 sg13g2_dlygate4sd3_1
X_3406_ _2988_ _2962_ _2989_ VPWR VGND sg13g2_xor2_1
X_4386_ _1139_ VPWR _1163_ VGND _1159_ _1161_ sg13g2_o21ai_1
Xhold279 mac1.sum_lvl2_ff\[12\] VPWR VGND net319 sg13g2_dlygate4sd3_1
X_3337_ _2921_ _2899_ _2923_ VPWR VGND sg13g2_xor2_1
X_6125_ net1118 VGND VPWR _0165_ DP_2.matrix\[80\] clknet_leaf_58_clk sg13g2_dfrbpq_2
X_3268_ _2856_ _2826_ _2855_ VPWR VGND sg13g2_nand2_1
XFILLER_22_1022 VPWR VGND sg13g2_decap_8
X_6056_ net899 _0232_ VPWR VGND sg13g2_buf_1
X_3199_ _2788_ _2741_ _2787_ VPWR VGND sg13g2_xnor2_1
X_5007_ VPWR _1756_ _1755_ VGND sg13g2_inv_1
XFILLER_26_389 VPWR VGND sg13g2_fill_1
X_5909_ _2558_ _2562_ _2563_ VPWR VGND sg13g2_nor2b_1
XFILLER_2_945 VPWR VGND sg13g2_decap_8
XFILLER_18_868 VPWR VGND sg13g2_decap_8
XFILLER_17_356 VPWR VGND sg13g2_fill_1
XFILLER_41_860 VPWR VGND sg13g2_decap_8
XFILLER_13_584 VPWR VGND sg13g2_fill_1
XFILLER_40_392 VPWR VGND sg13g2_fill_1
XFILLER_45_1000 VPWR VGND sg13g2_decap_8
X_4240_ _1019_ _1020_ _1014_ _1021_ VPWR VGND sg13g2_nand3_1
X_4171_ _0120_ _0957_ _0958_ VPWR VGND sg13g2_xnor2_1
X_3122_ _2713_ net997 net933 VPWR VGND sg13g2_nand2_1
X_3053_ _2647_ net1001 net937 VPWR VGND sg13g2_nand2_1
XFILLER_17_890 VPWR VGND sg13g2_decap_8
X_3955_ _0724_ VPWR _0749_ VGND _0745_ _0747_ sg13g2_o21ai_1
XFILLER_32_871 VPWR VGND sg13g2_fill_1
X_3886_ _0680_ _0681_ _0682_ VPWR VGND sg13g2_and2_1
X_5625_ _2305_ net401 net346 VPWR VGND sg13g2_nand2_1
X_5556_ _0033_ _2249_ _2250_ VPWR VGND sg13g2_xnor2_1
X_5487_ _2198_ _2192_ _2194_ VPWR VGND sg13g2_nand2_1
X_4507_ _1280_ net1048 net839 net893 DP_4.matrix\[41\] VPWR VGND sg13g2_a22oi_1
X_4438_ _1213_ _1174_ _0137_ VPWR VGND sg13g2_xor2_1
X_4369_ _1146_ _1141_ _1145_ VPWR VGND sg13g2_xnor2_1
X_6108_ net1090 VGND VPWR _0078_ mac1.products_ff\[72\] clknet_leaf_63_clk sg13g2_dfrbpq_1
X_6039_ net955 _0207_ VPWR VGND sg13g2_buf_1
XFILLER_15_838 VPWR VGND sg13g2_decap_8
XFILLER_25_32 VPWR VGND sg13g2_fill_1
XFILLER_41_101 VPWR VGND sg13g2_fill_1
XFILLER_29_1017 VPWR VGND sg13g2_decap_8
XFILLER_29_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_245 VPWR VGND sg13g2_fill_2
XFILLER_49_278 VPWR VGND sg13g2_fill_1
XFILLER_49_267 VPWR VGND sg13g2_fill_2
XFILLER_46_952 VPWR VGND sg13g2_decap_8
XFILLER_18_687 VPWR VGND sg13g2_fill_1
XFILLER_14_860 VPWR VGND sg13g2_decap_8
X_3740_ _0545_ net1027 net966 VPWR VGND sg13g2_nand2_1
XFILLER_41_690 VPWR VGND sg13g2_fill_1
X_3671_ VGND VPWR _0478_ _0476_ _0439_ sg13g2_or2_1
X_6390_ net1069 VGND VPWR net391 mac1.sum_lvl3_ff\[2\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_5410_ _2138_ _2135_ _2137_ VPWR VGND sg13g2_nand2_1
X_5341_ _2080_ net874 net1042 VPWR VGND sg13g2_nand2_1
X_5272_ _2014_ _2003_ _2013_ VPWR VGND sg13g2_xnor2_1
X_4223_ _1005_ _0997_ _1004_ VPWR VGND sg13g2_nand2_1
X_4154_ _0942_ net949 net1007 VPWR VGND sg13g2_nand2_1
X_4085_ VGND VPWR _0799_ _0841_ _0876_ _0840_ sg13g2_a21oi_1
X_3105_ _2685_ VPWR _2697_ VGND _2693_ _2695_ sg13g2_o21ai_1
X_3036_ VPWR _2633_ DP_3.I_range.out_data\[5\] VGND sg13g2_inv_1
XFILLER_37_974 VPWR VGND sg13g2_decap_8
XFILLER_23_112 VPWR VGND sg13g2_fill_1
X_4987_ _1738_ _1730_ _1737_ VPWR VGND sg13g2_nand2_1
X_3938_ _0732_ _0726_ _0731_ VPWR VGND sg13g2_xnor2_1
X_3869_ _0663_ _0660_ _0665_ VPWR VGND sg13g2_xor2_1
Xclkbuf_4_2_0_clk clknet_0_clk clknet_4_2_0_clk VPWR VGND sg13g2_buf_8
X_6588_ net1080 VGND VPWR net13 DP_3.I_range.out_data\[2\] clknet_leaf_22_clk sg13g2_dfrbpq_2
X_5608_ _2290_ net489 _0060_ VPWR VGND sg13g2_nor2b_1
X_5539_ _2237_ VPWR _2238_ VGND _2231_ _2234_ sg13g2_o21ai_1
XFILLER_46_215 VPWR VGND sg13g2_fill_1
XFILLER_28_974 VPWR VGND sg13g2_decap_8
XFILLER_14_167 VPWR VGND sg13g2_fill_2
XFILLER_30_638 VPWR VGND sg13g2_fill_1
XFILLER_10_373 VPWR VGND sg13g2_fill_2
XFILLER_7_856 VPWR VGND sg13g2_decap_8
XFILLER_11_896 VPWR VGND sg13g2_decap_8
XFILLER_42_1025 VPWR VGND sg13g2_decap_4
XFILLER_38_716 VPWR VGND sg13g2_decap_4
XFILLER_19_930 VPWR VGND sg13g2_decap_8
XFILLER_46_760 VPWR VGND sg13g2_fill_2
X_4910_ _1665_ _1656_ _1667_ VPWR VGND sg13g2_xor2_1
X_5890_ net863 _2495_ _2544_ VPWR VGND sg13g2_nor2_1
X_4841_ _1600_ net914 net856 VPWR VGND sg13g2_nand2_1
XFILLER_20_104 VPWR VGND sg13g2_fill_1
XFILLER_20_126 VPWR VGND sg13g2_fill_2
XFILLER_21_649 VPWR VGND sg13g2_decap_8
X_4772_ _1510_ _1530_ _1532_ _1533_ VPWR VGND sg13g2_or3_1
X_3723_ _0529_ _0508_ _0528_ VPWR VGND sg13g2_xnor2_1
X_6511_ net1136 VGND VPWR net224 mac2.sum_lvl1_ff\[47\] clknet_leaf_43_clk sg13g2_dfrbpq_1
XFILLER_9_171 VPWR VGND sg13g2_fill_1
X_3654_ _0462_ _0446_ _0460_ VPWR VGND sg13g2_xnor2_1
X_6442_ net1139 VGND VPWR _0145_ mac2.products_ff\[6\] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_6373_ net1064 VGND VPWR net119 mac1.sum_lvl3_ff\[21\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3585_ _0394_ _0386_ _0393_ VPWR VGND sg13g2_nand2_1
X_5324_ _2025_ _2063_ _2064_ VPWR VGND sg13g2_nor2_1
X_5255_ _1997_ net821 net1046 VPWR VGND sg13g2_nand2_1
X_4206_ _0989_ net906 net842 VPWR VGND sg13g2_nand2_1
X_5186_ _1921_ _1929_ _1930_ VPWR VGND sg13g2_nor2_1
XFILLER_29_738 VPWR VGND sg13g2_fill_2
X_4137_ _0924_ _0912_ _0926_ VPWR VGND sg13g2_xor2_1
X_4068_ _0859_ net952 net1007 VPWR VGND sg13g2_nand2_1
XFILLER_24_421 VPWR VGND sg13g2_fill_2
XFILLER_25_933 VPWR VGND sg13g2_decap_8
XFILLER_24_487 VPWR VGND sg13g2_decap_8
XFILLER_4_859 VPWR VGND sg13g2_decap_8
Xfanout1104 net1106 net1104 VPWR VGND sg13g2_buf_8
Xfanout1115 net1130 net1115 VPWR VGND sg13g2_buf_8
Xfanout1137 net1138 net1137 VPWR VGND sg13g2_buf_8
Xfanout1126 net1128 net1126 VPWR VGND sg13g2_buf_8
Xfanout1148 rst_n net1148 VPWR VGND sg13g2_buf_8
XFILLER_19_215 VPWR VGND sg13g2_decap_4
XFILLER_16_966 VPWR VGND sg13g2_decap_8
XFILLER_43_774 VPWR VGND sg13g2_fill_2
XFILLER_30_413 VPWR VGND sg13g2_decap_4
XFILLER_8_57 VPWR VGND sg13g2_fill_1
X_3370_ _2953_ _2952_ _2955_ VPWR VGND sg13g2_xor2_1
XFILLER_3_881 VPWR VGND sg13g2_decap_8
X_5040_ _1785_ _1786_ _1780_ _1788_ VPWR VGND sg13g2_nand3_1
XFILLER_38_513 VPWR VGND sg13g2_fill_2
X_5942_ VGND VPWR net787 _2588_ _0178_ _2587_ sg13g2_a21oi_1
XFILLER_19_771 VPWR VGND sg13g2_fill_2
XFILLER_22_903 VPWR VGND sg13g2_decap_8
XFILLER_34_752 VPWR VGND sg13g2_fill_2
X_5873_ _2523_ VPWR _2528_ VGND net791 _2526_ sg13g2_o21ai_1
X_4824_ _1582_ _1583_ _1584_ VPWR VGND sg13g2_nor2b_1
X_4755_ _1516_ _1469_ _1514_ VPWR VGND sg13g2_xnor2_1
X_3706_ VGND VPWR _0512_ _0511_ _0487_ sg13g2_or2_1
X_4686_ _1446_ _1445_ _1440_ _1449_ VPWR VGND sg13g2_a21o_1
X_3637_ _0445_ _0435_ _0443_ VPWR VGND sg13g2_xnor2_1
X_6425_ net1060 VGND VPWR _0027_ mac1.total_sum\[5\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_3568_ _0376_ _0377_ _0346_ _0378_ VPWR VGND sg13g2_nand3_1
X_6356_ net1102 VGND VPWR net145 mac2.sum_lvl1_ff\[72\] clknet_leaf_24_clk sg13g2_dfrbpq_1
X_5307_ _2046_ _2047_ _2048_ VPWR VGND sg13g2_nor2_1
X_3499_ _0308_ _0309_ _0284_ _0311_ VPWR VGND sg13g2_nand3_1
X_6287_ net1120 VGND VPWR net226 mac1.sum_lvl2_ff\[11\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_5238_ _1979_ _1970_ _1981_ VPWR VGND sg13g2_xor2_1
X_5169_ _1911_ _1910_ _1912_ _1914_ VPWR VGND sg13g2_a21o_1
XFILLER_25_730 VPWR VGND sg13g2_decap_4
XFILLER_25_752 VPWR VGND sg13g2_decap_4
XFILLER_13_947 VPWR VGND sg13g2_decap_8
XFILLER_40_755 VPWR VGND sg13g2_fill_1
XFILLER_0_840 VPWR VGND sg13g2_decap_8
Xhold6 mac1.sum_lvl1_ff\[10\] VPWR VGND net46 sg13g2_dlygate4sd3_1
XFILLER_31_700 VPWR VGND sg13g2_decap_4
XFILLER_31_744 VPWR VGND sg13g2_fill_1
XFILLER_30_265 VPWR VGND sg13g2_fill_2
X_4540_ _1312_ net893 net834 VPWR VGND sg13g2_nand2_1
XFILLER_8_962 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_10_clk clknet_4_9_0_clk clknet_leaf_10_clk VPWR VGND sg13g2_buf_8
X_4471_ _1246_ _1245_ _1244_ VPWR VGND sg13g2_nand2b_1
Xhold406 _0058_ VPWR VGND net446 sg13g2_dlygate4sd3_1
Xhold417 _0062_ VPWR VGND net457 sg13g2_dlygate4sd3_1
X_3422_ _2990_ VPWR _3004_ VGND _2962_ _2988_ sg13g2_o21ai_1
Xhold439 _0001_ VPWR VGND net479 sg13g2_dlygate4sd3_1
X_6210_ net1120 VGND VPWR net246 mac1.sum_lvl1_ff\[10\] clknet_leaf_60_clk sg13g2_dfrbpq_1
Xhold428 _0004_ VPWR VGND net468 sg13g2_dlygate4sd3_1
X_6141_ net1071 VGND VPWR _0067_ mac1.products_ff\[139\] clknet_leaf_66_clk sg13g2_dfrbpq_1
Xfanout908 net909 net908 VPWR VGND sg13g2_buf_8
X_3353_ net993 net990 net928 net926 _2938_ VPWR VGND sg13g2_and4_1
Xfanout919 DP_3.matrix\[3\] net919 VPWR VGND sg13g2_buf_8
X_3284_ _2871_ _2830_ _2869_ VPWR VGND sg13g2_xnor2_1
X_6072_ net838 _0256_ VPWR VGND sg13g2_buf_1
X_5023_ VGND VPWR _1772_ _1771_ _1751_ sg13g2_or2_1
XFILLER_0_1022 VPWR VGND sg13g2_decap_8
X_5925_ net1038 net785 _2577_ VPWR VGND sg13g2_nor2_1
X_5856_ VGND VPWR _2511_ _2510_ _2485_ sg13g2_or2_1
XFILLER_16_1008 VPWR VGND sg13g2_decap_8
XFILLER_22_744 VPWR VGND sg13g2_decap_8
X_4807_ _1521_ VPWR _1567_ VGND _1519_ _1522_ sg13g2_o21ai_1
XFILLER_10_917 VPWR VGND sg13g2_decap_8
X_5787_ net971 DP_2.matrix\[41\] net809 _2443_ VPWR VGND sg13g2_mux2_1
X_4738_ _1488_ VPWR _1499_ VGND _1466_ _1489_ sg13g2_o21ai_1
X_4669_ _1430_ _1429_ _1432_ VPWR VGND sg13g2_xor2_1
X_6408_ net1084 VGND VPWR net97 mac2.sum_lvl3_ff\[24\] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_6339_ net1103 VGND VPWR net44 mac2.sum_lvl2_ff\[53\] clknet_leaf_26_clk sg13g2_dfrbpq_1
XFILLER_12_221 VPWR VGND sg13g2_fill_2
XFILLER_12_232 VPWR VGND sg13g2_fill_1
XFILLER_40_541 VPWR VGND sg13g2_decap_4
XFILLER_5_954 VPWR VGND sg13g2_decap_8
XFILLER_4_442 VPWR VGND sg13g2_fill_2
XFILLER_5_47 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_59_clk clknet_4_8_0_clk clknet_leaf_59_clk VPWR VGND sg13g2_buf_8
XFILLER_35_302 VPWR VGND sg13g2_fill_1
X_3971_ _0759_ _0763_ _0764_ VPWR VGND sg13g2_nor2_1
X_5710_ _2362_ _2366_ _2372_ VPWR VGND sg13g2_nor2_1
X_5641_ _2317_ _2318_ _0051_ VPWR VGND sg13g2_and2_1
X_5572_ _0036_ _2261_ _2264_ VPWR VGND sg13g2_xnor2_1
X_4523_ VGND VPWR _1296_ _1295_ _1283_ sg13g2_or2_1
Xhold203 mac1.sum_lvl1_ff\[80\] VPWR VGND net243 sg13g2_dlygate4sd3_1
Xhold214 mac1.sum_lvl1_ff\[76\] VPWR VGND net254 sg13g2_dlygate4sd3_1
Xhold225 mac1.sum_lvl3_ff\[0\] VPWR VGND net265 sg13g2_dlygate4sd3_1
Xhold236 DP_3.matrix\[79\] VPWR VGND net276 sg13g2_dlygate4sd3_1
Xhold247 mac1.sum_lvl2_ff\[19\] VPWR VGND net287 sg13g2_dlygate4sd3_1
X_4454_ _1229_ net897 DP_4.matrix\[41\] VPWR VGND sg13g2_nand2_1
Xhold258 _2325_ VPWR VGND net298 sg13g2_dlygate4sd3_1
Xhold269 _0039_ VPWR VGND net309 sg13g2_dlygate4sd3_1
X_3405_ _2988_ net929 net1054 VPWR VGND sg13g2_nand2_1
X_4385_ _1139_ _1159_ _1161_ _1162_ VPWR VGND sg13g2_or3_1
X_6124_ net1089 VGND VPWR _0164_ DP_2.matrix\[44\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_3336_ _2921_ _2899_ _2922_ VPWR VGND sg13g2_nor2b_1
X_6055_ net900 _0231_ VPWR VGND sg13g2_buf_1
X_3267_ _2854_ _2837_ _2855_ VPWR VGND sg13g2_xor2_1
XFILLER_22_1001 VPWR VGND sg13g2_decap_8
X_5006_ _1752_ _1754_ _1755_ VPWR VGND sg13g2_nor2_1
X_3198_ _2787_ _2778_ _2785_ VPWR VGND sg13g2_xnor2_1
X_5908_ _2559_ VPWR _2562_ VGND net794 _2561_ sg13g2_o21ai_1
X_5839_ _2494_ net905 net795 VPWR VGND sg13g2_nand2b_1
XFILLER_10_769 VPWR VGND sg13g2_fill_2
XFILLER_2_924 VPWR VGND sg13g2_decap_8
XFILLER_7_1017 VPWR VGND sg13g2_decap_8
XFILLER_7_1028 VPWR VGND sg13g2_fill_1
XFILLER_18_814 VPWR VGND sg13g2_decap_8
XFILLER_9_501 VPWR VGND sg13g2_decap_8
XFILLER_41_883 VPWR VGND sg13g2_fill_2
X_4170_ VGND VPWR _0934_ _0937_ _0958_ _0933_ sg13g2_a21oi_1
X_3121_ _2712_ net1000 net930 VPWR VGND sg13g2_nand2_1
XFILLER_49_994 VPWR VGND sg13g2_decap_8
X_3052_ VGND VPWR _2646_ _2641_ _2639_ sg13g2_or2_1
X_3954_ _0724_ _0745_ _0747_ _0748_ VPWR VGND sg13g2_or3_1
X_3885_ _0679_ _0678_ _0640_ _0681_ VPWR VGND sg13g2_a21o_1
X_5624_ _2304_ _2301_ _2303_ VPWR VGND sg13g2_nand2_1
X_5555_ _2251_ _2248_ _2250_ VPWR VGND sg13g2_nand2_1
X_5486_ _2197_ _2196_ _2195_ VPWR VGND sg13g2_nand2b_1
X_4506_ _1265_ _1260_ _1267_ _1279_ VPWR VGND sg13g2_a21o_1
X_4437_ _1211_ _1212_ _1213_ VPWR VGND sg13g2_nor2b_1
X_6107_ net1088 VGND VPWR _0077_ mac1.products_ff\[71\] clknet_leaf_64_clk sg13g2_dfrbpq_1
X_4368_ _1145_ _1098_ _1143_ VPWR VGND sg13g2_xnor2_1
X_3319_ _2905_ _2879_ _2903_ VPWR VGND sg13g2_xnor2_1
X_4299_ _1075_ _1074_ _1069_ _1078_ VPWR VGND sg13g2_a21o_1
X_6038_ net957 _0206_ VPWR VGND sg13g2_buf_1
XFILLER_1_231 VPWR VGND sg13g2_decap_4
XFILLER_1_220 VPWR VGND sg13g2_fill_2
XFILLER_38_909 VPWR VGND sg13g2_decap_4
XFILLER_33_614 VPWR VGND sg13g2_fill_1
XFILLER_12_1011 VPWR VGND sg13g2_decap_8
X_3670_ _0477_ net1032 net969 VPWR VGND sg13g2_nand2_1
X_5340_ _2059_ VPWR _2079_ VGND _2031_ _2057_ sg13g2_o21ai_1
X_5271_ _2013_ _2004_ _2011_ VPWR VGND sg13g2_xnor2_1
XFILLER_5_592 VPWR VGND sg13g2_fill_1
X_4222_ _1002_ _1003_ _1004_ VPWR VGND sg13g2_nor2b_1
X_4153_ _0941_ net1007 net947 VPWR VGND sg13g2_nand2_1
X_3104_ _2685_ _2693_ _2695_ _2696_ VPWR VGND sg13g2_or3_1
X_4084_ _0875_ _0874_ _0873_ VPWR VGND sg13g2_nand2b_1
XFILLER_28_419 VPWR VGND sg13g2_fill_1
X_3035_ VPWR DP_1.Q_range.data_plus_4\[6\] net8 VGND sg13g2_inv_1
X_4986_ _1735_ _1736_ _1737_ VPWR VGND sg13g2_nor2b_1
X_3937_ _0731_ _0693_ _0728_ VPWR VGND sg13g2_xnor2_1
XFILLER_23_157 VPWR VGND sg13g2_fill_1
XFILLER_32_680 VPWR VGND sg13g2_fill_2
X_3868_ _0664_ _0663_ _0660_ VPWR VGND sg13g2_nand2b_1
X_6587_ net1075 VGND VPWR DP_1.Q_range.data_plus_4\[6\] DP_1.Q_range.out_data\[5\]
+ clknet_leaf_5_clk sg13g2_dfrbpq_1
X_3799_ _0602_ _0578_ _0601_ VPWR VGND sg13g2_xnor2_1
X_5607_ net488 VPWR _2291_ VGND _2285_ _2289_ sg13g2_o21ai_1
X_5538_ mac2.sum_lvl2_ff\[7\] mac2.sum_lvl2_ff\[26\] _2237_ VPWR VGND sg13g2_xor2_1
X_5469_ mac1.sum_lvl3_ff\[28\] mac1.sum_lvl3_ff\[8\] _2183_ VPWR VGND sg13g2_and2_1
XFILLER_47_739 VPWR VGND sg13g2_fill_2
XFILLER_28_953 VPWR VGND sg13g2_decap_8
XFILLER_27_452 VPWR VGND sg13g2_decap_8
XFILLER_43_934 VPWR VGND sg13g2_fill_2
XFILLER_15_658 VPWR VGND sg13g2_fill_1
XFILLER_23_691 VPWR VGND sg13g2_decap_8
XFILLER_7_802 VPWR VGND sg13g2_decap_4
XFILLER_11_875 VPWR VGND sg13g2_decap_8
XFILLER_7_835 VPWR VGND sg13g2_decap_8
XFILLER_42_1004 VPWR VGND sg13g2_decap_8
XFILLER_18_452 VPWR VGND sg13g2_fill_1
XFILLER_19_986 VPWR VGND sg13g2_decap_8
XFILLER_18_496 VPWR VGND sg13g2_fill_1
X_4840_ VGND VPWR net864 net908 _1599_ _1568_ sg13g2_a21oi_1
X_6510_ net1136 VGND VPWR net245 mac2.sum_lvl1_ff\[46\] clknet_leaf_50_clk sg13g2_dfrbpq_1
X_4771_ VGND VPWR _1528_ _1529_ _1532_ _1511_ sg13g2_a21oi_1
X_3722_ _0528_ _0517_ _0527_ VPWR VGND sg13g2_xnor2_1
XFILLER_9_194 VPWR VGND sg13g2_decap_4
X_3653_ _0461_ _0446_ _0460_ VPWR VGND sg13g2_nand2_1
X_6441_ net1127 VGND VPWR _0138_ mac2.products_ff\[5\] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_6372_ net1062 VGND VPWR net170 mac1.sum_lvl3_ff\[20\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_5323_ _2063_ _2054_ _2062_ VPWR VGND sg13g2_xnor2_1
X_3584_ _0391_ _0387_ _0393_ VPWR VGND sg13g2_xor2_1
X_5254_ _1996_ net816 net874 VPWR VGND sg13g2_nand2_1
X_5185_ _1929_ _1922_ _1928_ VPWR VGND sg13g2_xnor2_1
X_4205_ _0987_ _0988_ _0080_ VPWR VGND sg13g2_nor2_1
X_4136_ VGND VPWR _0925_ _0924_ _0912_ sg13g2_or2_1
XFILLER_29_728 VPWR VGND sg13g2_fill_1
X_4067_ _0858_ net1010 net951 VPWR VGND sg13g2_nand2_1
XFILLER_25_912 VPWR VGND sg13g2_decap_8
XFILLER_36_260 VPWR VGND sg13g2_fill_2
XFILLER_11_105 VPWR VGND sg13g2_fill_2
XFILLER_19_1028 VPWR VGND sg13g2_fill_1
XFILLER_25_989 VPWR VGND sg13g2_decap_8
X_4969_ VGND VPWR _1692_ _1715_ _1723_ _1717_ sg13g2_a21oi_1
XFILLER_11_116 VPWR VGND sg13g2_fill_2
XFILLER_4_838 VPWR VGND sg13g2_decap_8
Xfanout1105 net1106 net1105 VPWR VGND sg13g2_buf_8
Xfanout1116 net1119 net1116 VPWR VGND sg13g2_buf_8
Xfanout1138 net1147 net1138 VPWR VGND sg13g2_buf_8
Xfanout1127 net1128 net1127 VPWR VGND sg13g2_buf_8
XFILLER_15_433 VPWR VGND sg13g2_fill_1
XFILLER_16_945 VPWR VGND sg13g2_decap_8
XFILLER_30_436 VPWR VGND sg13g2_fill_2
XFILLER_30_458 VPWR VGND sg13g2_fill_1
XFILLER_11_672 VPWR VGND sg13g2_fill_1
XFILLER_6_131 VPWR VGND sg13g2_fill_2
XFILLER_3_860 VPWR VGND sg13g2_decap_8
XFILLER_38_503 VPWR VGND sg13g2_fill_2
Xclkbuf_4_1_0_clk clknet_0_clk clknet_4_1_0_clk VPWR VGND sg13g2_buf_8
X_5941_ _2588_ _2429_ _2431_ VPWR VGND sg13g2_xnor2_1
XFILLER_19_794 VPWR VGND sg13g2_fill_2
X_5872_ VGND VPWR net273 net797 _2527_ _2526_ sg13g2_a21oi_1
XFILLER_22_959 VPWR VGND sg13g2_decap_8
X_4823_ _1583_ _1546_ _1581_ VPWR VGND sg13g2_nand2_1
X_4754_ VGND VPWR _1515_ _1513_ _1470_ sg13g2_or2_1
XFILLER_21_458 VPWR VGND sg13g2_fill_1
X_3705_ _0511_ net975 net1058 VPWR VGND sg13g2_nand2_1
XFILLER_30_992 VPWR VGND sg13g2_decap_8
X_4685_ _1445_ _1446_ _1440_ _1448_ VPWR VGND sg13g2_nand3_1
X_3636_ _0435_ _0443_ _0444_ VPWR VGND sg13g2_nor2_1
X_6424_ net1060 VGND VPWR _0026_ mac1.total_sum\[4\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_3567_ _0352_ VPWR _0377_ VGND _0373_ _0375_ sg13g2_o21ai_1
X_6355_ net1089 VGND VPWR net264 mac1.sum_lvl1_ff\[87\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_5306_ VGND VPWR _1994_ _2014_ _2047_ _2016_ sg13g2_a21oi_1
X_6286_ net1120 VGND VPWR net46 mac1.sum_lvl2_ff\[10\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_5237_ _1980_ _1970_ _1979_ VPWR VGND sg13g2_nand2b_1
X_3498_ _0308_ _0309_ _0310_ VPWR VGND sg13g2_and2_1
XFILLER_25_1010 VPWR VGND sg13g2_decap_8
X_5168_ _1911_ _1912_ _1910_ _1913_ VPWR VGND sg13g2_nand3_1
X_5099_ _1845_ _1807_ _1842_ VPWR VGND sg13g2_xnor2_1
X_4119_ _0894_ _0889_ _0896_ _0908_ VPWR VGND sg13g2_a21o_1
XFILLER_16_219 VPWR VGND sg13g2_fill_2
XFILLER_13_926 VPWR VGND sg13g2_decap_8
XFILLER_12_469 VPWR VGND sg13g2_decap_4
XFILLER_21_992 VPWR VGND sg13g2_decap_8
XFILLER_20_491 VPWR VGND sg13g2_decap_4
XFILLER_48_812 VPWR VGND sg13g2_fill_1
XFILLER_48_823 VPWR VGND sg13g2_fill_1
XFILLER_0_896 VPWR VGND sg13g2_decap_8
Xhold7 mac2.sum_lvl1_ff\[78\] VPWR VGND net47 sg13g2_dlygate4sd3_1
XFILLER_16_775 VPWR VGND sg13g2_fill_1
XFILLER_16_797 VPWR VGND sg13g2_decap_8
XFILLER_8_941 VPWR VGND sg13g2_decap_8
Xhold407 DP_3.matrix\[5\] VPWR VGND net447 sg13g2_dlygate4sd3_1
Xhold418 mac1.sum_lvl2_ff\[27\] VPWR VGND net458 sg13g2_dlygate4sd3_1
X_4470_ _1209_ _1243_ _1207_ _1245_ VPWR VGND sg13g2_nand3_1
X_3421_ _3002_ _2987_ _3003_ VPWR VGND sg13g2_xor2_1
Xhold429 mac2.sum_lvl2_ff\[5\] VPWR VGND net469 sg13g2_dlygate4sd3_1
X_3352_ _2937_ net990 net926 VPWR VGND sg13g2_nand2_1
X_6140_ net1094 VGND VPWR net283 DP_1.matrix\[5\] clknet_leaf_8_clk sg13g2_dfrbpq_2
Xfanout909 net910 net909 VPWR VGND sg13g2_buf_8
X_3283_ VGND VPWR _2870_ _2868_ _2831_ sg13g2_or2_1
X_6071_ net841 _0255_ VPWR VGND sg13g2_buf_1
XFILLER_38_300 VPWR VGND sg13g2_fill_2
X_5022_ _1769_ _1768_ _1771_ VPWR VGND sg13g2_xor2_1
XFILLER_17_0 VPWR VGND sg13g2_fill_2
XFILLER_0_1001 VPWR VGND sg13g2_decap_8
X_5924_ net786 net1040 _0172_ VPWR VGND sg13g2_xor2_1
X_5855_ VGND VPWR _2510_ _2509_ _2505_ sg13g2_or2_1
X_4806_ _1566_ _1561_ _1565_ VPWR VGND sg13g2_xnor2_1
XFILLER_22_778 VPWR VGND sg13g2_fill_2
X_5786_ VGND VPWR net784 _2441_ _2442_ _2437_ sg13g2_a21oi_1
X_4737_ _1497_ _1496_ _0146_ VPWR VGND sg13g2_xor2_1
X_4668_ _1431_ _1429_ VPWR VGND _1430_ sg13g2_nand2b_2
X_3619_ _0425_ _0424_ _0426_ _0428_ VPWR VGND sg13g2_a21o_1
X_6407_ net1100 VGND VPWR net76 mac2.sum_lvl3_ff\[23\] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_4599_ _1366_ _1358_ _1365_ VPWR VGND sg13g2_nand2_1
X_6338_ net1084 VGND VPWR net194 mac2.sum_lvl2_ff\[52\] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_6269_ net1115 VGND VPWR net241 mac1.sum_lvl1_ff\[45\] clknet_leaf_59_clk sg13g2_dfrbpq_1
XFILLER_44_314 VPWR VGND sg13g2_fill_2
XFILLER_44_21 VPWR VGND sg13g2_fill_1
XFILLER_5_933 VPWR VGND sg13g2_decap_8
X_3970_ VGND VPWR _0763_ _0762_ _0761_ sg13g2_or2_1
X_5640_ net531 _2314_ _2316_ _2318_ VPWR VGND sg13g2_or3_1
X_5571_ _2264_ _2263_ _2262_ VPWR VGND sg13g2_nand2b_1
X_4522_ _1293_ _1284_ _1295_ VPWR VGND sg13g2_xor2_1
Xhold204 mac1.sum_lvl1_ff\[79\] VPWR VGND net244 sg13g2_dlygate4sd3_1
Xhold215 mac1.sum_lvl1_ff\[40\] VPWR VGND net255 sg13g2_dlygate4sd3_1
Xhold226 _0016_ VPWR VGND net266 sg13g2_dlygate4sd3_1
X_4453_ VGND VPWR net844 net891 _1228_ _1197_ sg13g2_a21oi_1
Xhold237 DP_3.matrix\[77\] VPWR VGND net277 sg13g2_dlygate4sd3_1
Xhold248 _0007_ VPWR VGND net288 sg13g2_dlygate4sd3_1
X_3404_ _2987_ net927 net1054 VPWR VGND sg13g2_nand2_1
Xhold259 _0053_ VPWR VGND net299 sg13g2_dlygate4sd3_1
X_4384_ VGND VPWR _1157_ _1158_ _1161_ _1140_ sg13g2_a21oi_1
X_3335_ _2921_ _2900_ _2920_ VPWR VGND sg13g2_xnor2_1
X_6123_ net1094 VGND VPWR _0163_ DP_2.matrix\[8\] clknet_leaf_10_clk sg13g2_dfrbpq_2
X_3266_ _2854_ _2838_ _2852_ VPWR VGND sg13g2_xnor2_1
X_6054_ net902 _0230_ VPWR VGND sg13g2_buf_1
X_5005_ net889 net886 net820 net818 _1754_ VPWR VGND sg13g2_and4_1
X_3197_ _2786_ _2778_ _2785_ VPWR VGND sg13g2_nand2_1
X_5907_ _2560_ VPWR _2561_ VGND net855 net804 sg13g2_o21ai_1
X_5838_ _2493_ _2490_ _2492_ VPWR VGND sg13g2_nand2_1
X_5769_ net1033 net1015 net810 _2426_ VPWR VGND sg13g2_mux2_1
XFILLER_2_903 VPWR VGND sg13g2_decap_8
XFILLER_44_122 VPWR VGND sg13g2_fill_2
XFILLER_18_848 VPWR VGND sg13g2_decap_4
XFILLER_33_807 VPWR VGND sg13g2_fill_2
XFILLER_44_199 VPWR VGND sg13g2_fill_2
XFILLER_32_339 VPWR VGND sg13g2_fill_1
X_3120_ _2694_ VPWR _2711_ VGND _2685_ _2695_ sg13g2_o21ai_1
XFILLER_1_991 VPWR VGND sg13g2_decap_8
XFILLER_49_973 VPWR VGND sg13g2_decap_8
X_3051_ _2645_ net1003 DP_2.matrix\[75\] VPWR VGND sg13g2_nand2_1
X_3953_ VGND VPWR _0743_ _0744_ _0747_ _0725_ sg13g2_a21oi_1
X_3884_ _0678_ _0679_ _0640_ _0680_ VPWR VGND sg13g2_nand3_1
X_5623_ _0063_ _2300_ net316 VPWR VGND sg13g2_xnor2_1
X_5554_ _2245_ _2243_ _2244_ _2250_ VPWR VGND sg13g2_a21o_2
X_5485_ _2196_ mac1.sum_lvl3_ff\[31\] mac1.sum_lvl3_ff\[11\] VPWR VGND sg13g2_nand2_1
X_4505_ _0129_ _1277_ _1278_ VPWR VGND sg13g2_xnor2_1
X_4436_ _1212_ _1175_ _1210_ VPWR VGND sg13g2_nand2_1
X_4367_ VGND VPWR _1144_ _1142_ _1099_ sg13g2_or2_1
X_6106_ net1069 VGND VPWR _0076_ mac1.products_ff\[70\] clknet_leaf_67_clk sg13g2_dfrbpq_1
X_3318_ VGND VPWR _2904_ _2903_ _2879_ sg13g2_or2_1
X_4298_ _1074_ _1075_ _1069_ _1077_ VPWR VGND sg13g2_nand3_1
X_6037_ net960 _0205_ VPWR VGND sg13g2_buf_1
X_3249_ _2837_ _2827_ _2835_ VPWR VGND sg13g2_xnor2_1
XFILLER_41_147 VPWR VGND sg13g2_fill_2
XFILLER_41_99 VPWR VGND sg13g2_fill_2
XFILLER_46_987 VPWR VGND sg13g2_decap_8
XFILLER_18_678 VPWR VGND sg13g2_fill_1
XFILLER_14_895 VPWR VGND sg13g2_decap_8
X_5270_ _2011_ _2004_ _2012_ VPWR VGND sg13g2_nor2b_1
X_4221_ _0998_ VPWR _1003_ VGND _0999_ _1001_ sg13g2_o21ai_1
X_4152_ _0940_ net1010 net1052 VPWR VGND sg13g2_nand2_1
X_3103_ VGND VPWR _2691_ _2692_ _2695_ _2686_ sg13g2_a21oi_1
X_4083_ _0838_ _0872_ _0836_ _0874_ VPWR VGND sg13g2_nand3_1
X_3034_ VPWR DP_3.Q_range.data_plus_4\[6\] net12 VGND sg13g2_inv_1
XFILLER_36_475 VPWR VGND sg13g2_fill_2
X_4985_ _1732_ VPWR _1736_ VGND _1733_ _1734_ sg13g2_o21ai_1
X_3936_ _0693_ _0728_ _0730_ VPWR VGND sg13g2_and2_1
X_3867_ _0662_ _0639_ _0663_ VPWR VGND sg13g2_xor2_1
XFILLER_20_887 VPWR VGND sg13g2_decap_8
X_6586_ net1075 VGND VPWR net7 DP_1.Q_range.out_data\[4\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_3798_ _0599_ _0593_ _0601_ VPWR VGND sg13g2_xor2_1
X_5606_ _2285_ net488 _2289_ _2290_ VPWR VGND sg13g2_nor3_1
X_5537_ _2236_ mac2.sum_lvl2_ff\[26\] mac2.sum_lvl2_ff\[7\] VPWR VGND sg13g2_nand2_1
X_5468_ _2181_ _2182_ _0029_ VPWR VGND sg13g2_and2_1
X_5399_ _2125_ net393 _2123_ _2129_ VPWR VGND sg13g2_nand3_1
X_4419_ _1195_ _1190_ _1194_ VPWR VGND sg13g2_xnor2_1
XFILLER_43_979 VPWR VGND sg13g2_decap_8
XFILLER_15_637 VPWR VGND sg13g2_fill_2
XFILLER_14_169 VPWR VGND sg13g2_fill_1
XFILLER_11_854 VPWR VGND sg13g2_decap_8
XFILLER_19_965 VPWR VGND sg13g2_decap_8
XFILLER_46_784 VPWR VGND sg13g2_fill_2
XFILLER_45_272 VPWR VGND sg13g2_fill_1
XFILLER_18_486 VPWR VGND sg13g2_fill_2
XFILLER_21_629 VPWR VGND sg13g2_fill_2
XFILLER_33_456 VPWR VGND sg13g2_fill_1
X_4770_ _1528_ _1529_ _1511_ _1531_ VPWR VGND sg13g2_nand3_1
XFILLER_42_990 VPWR VGND sg13g2_decap_8
XFILLER_9_140 VPWR VGND sg13g2_fill_1
X_3721_ _0527_ _0518_ _0525_ VPWR VGND sg13g2_xnor2_1
X_3652_ _0459_ _0452_ _0460_ VPWR VGND sg13g2_xor2_1
X_6440_ net1126 VGND VPWR _0088_ mac2.products_ff\[4\] clknet_leaf_33_clk sg13g2_dfrbpq_1
X_3583_ _0387_ _0391_ _0392_ VPWR VGND sg13g2_nor2_1
X_6371_ net1101 VGND VPWR net172 mac2.sum_lvl1_ff\[87\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_5322_ _2062_ _2026_ _2060_ VPWR VGND sg13g2_xnor2_1
XFILLER_47_0 VPWR VGND sg13g2_fill_2
X_5253_ _1978_ _1971_ _1941_ _1995_ VPWR VGND sg13g2_a21o_1
X_5184_ _1928_ _1923_ _1926_ VPWR VGND sg13g2_xnor2_1
X_4204_ _0988_ net847 net906 net905 net850 VPWR VGND sg13g2_a22oi_1
X_4135_ _0922_ _0913_ _0924_ VPWR VGND sg13g2_xor2_1
XFILLER_3_1021 VPWR VGND sg13g2_decap_8
X_4066_ VGND VPWR net960 net1006 _0857_ _0826_ sg13g2_a21oi_1
XFILLER_25_902 VPWR VGND sg13g2_fill_1
XFILLER_19_1007 VPWR VGND sg13g2_decap_8
XFILLER_25_968 VPWR VGND sg13g2_decap_8
X_4968_ _1720_ VPWR _1722_ VGND _1705_ _1718_ sg13g2_o21ai_1
X_4899_ _1636_ VPWR _1656_ VGND _1634_ _1637_ sg13g2_o21ai_1
X_3919_ _0714_ _0690_ _0713_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_662 VPWR VGND sg13g2_fill_2
X_6569_ net1061 VGND VPWR net481 mac2.total_sum\[1\] clknet_leaf_4_clk sg13g2_dfrbpq_1
Xfanout1117 net1119 net1117 VPWR VGND sg13g2_buf_8
Xfanout1106 net1107 net1106 VPWR VGND sg13g2_buf_8
Xfanout1128 net1129 net1128 VPWR VGND sg13g2_buf_8
Xfanout1139 net1146 net1139 VPWR VGND sg13g2_buf_8
XFILLER_19_228 VPWR VGND sg13g2_fill_2
XFILLER_16_924 VPWR VGND sg13g2_decap_8
XFILLER_27_283 VPWR VGND sg13g2_fill_1
XFILLER_43_798 VPWR VGND sg13g2_fill_2
XFILLER_6_176 VPWR VGND sg13g2_fill_2
X_5940_ net1029 net787 _2587_ VPWR VGND sg13g2_nor2_1
XFILLER_18_261 VPWR VGND sg13g2_fill_1
XFILLER_19_773 VPWR VGND sg13g2_fill_1
XFILLER_46_581 VPWR VGND sg13g2_fill_2
X_5871_ net794 _2524_ _2525_ _2526_ VPWR VGND sg13g2_nor3_1
XFILLER_34_754 VPWR VGND sg13g2_fill_1
XFILLER_22_938 VPWR VGND sg13g2_decap_8
X_4822_ _1546_ _1581_ _1582_ VPWR VGND sg13g2_nor2_1
X_4753_ _1514_ net859 net915 VPWR VGND sg13g2_nand2_1
X_3704_ _0510_ net971 net1027 VPWR VGND sg13g2_nand2_1
XFILLER_30_971 VPWR VGND sg13g2_decap_8
X_6423_ net1061 VGND VPWR net443 mac1.total_sum\[3\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_4684_ _1447_ _1440_ _1445_ _1446_ VPWR VGND sg13g2_and3_1
X_3635_ _0443_ _0436_ _0442_ VPWR VGND sg13g2_xnor2_1
XFILLER_1_809 VPWR VGND sg13g2_decap_8
X_3566_ _0352_ _0373_ _0375_ _0376_ VPWR VGND sg13g2_or3_1
X_6354_ net1067 VGND VPWR net223 mac1.sum_lvl1_ff\[86\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_5305_ _2044_ _2023_ _2046_ VPWR VGND sg13g2_xor2_1
X_3497_ _0307_ _0306_ _0268_ _0309_ VPWR VGND sg13g2_a21o_1
X_6285_ net1114 VGND VPWR net182 mac1.sum_lvl2_ff\[9\] clknet_leaf_59_clk sg13g2_dfrbpq_1
X_5236_ _1979_ _1971_ _1978_ VPWR VGND sg13g2_xnor2_1
X_5167_ _1864_ VPWR _1912_ VGND _1803_ _1865_ sg13g2_o21ai_1
X_5098_ _1807_ _1842_ _1844_ VPWR VGND sg13g2_and2_1
X_4118_ _0118_ _0906_ _0907_ VPWR VGND sg13g2_xnor2_1
X_4049_ _0841_ _0804_ _0839_ VPWR VGND sg13g2_nand2_1
XFILLER_13_905 VPWR VGND sg13g2_decap_8
XFILLER_33_23 VPWR VGND sg13g2_fill_2
XFILLER_21_971 VPWR VGND sg13g2_decap_8
XFILLER_32_1026 VPWR VGND sg13g2_fill_2
XFILLER_0_875 VPWR VGND sg13g2_decap_8
Xhold8 mac1.sum_lvl1_ff\[77\] VPWR VGND net48 sg13g2_dlygate4sd3_1
XFILLER_15_220 VPWR VGND sg13g2_fill_1
XFILLER_8_920 VPWR VGND sg13g2_decap_8
XFILLER_8_997 VPWR VGND sg13g2_decap_8
XFILLER_7_485 VPWR VGND sg13g2_fill_2
Xhold408 DP_1.matrix\[37\] VPWR VGND net448 sg13g2_dlygate4sd3_1
X_3420_ _3002_ net988 net1051 VPWR VGND sg13g2_nand2_1
Xhold419 _0015_ VPWR VGND net459 sg13g2_dlygate4sd3_1
X_3351_ _2936_ net994 net1051 VPWR VGND sg13g2_nand2_1
X_3282_ _2869_ net994 net929 VPWR VGND sg13g2_nand2_1
X_6070_ net842 _0254_ VPWR VGND sg13g2_buf_1
X_5021_ _1768_ _1769_ _1770_ VPWR VGND sg13g2_nor2b_2
X_5923_ VGND VPWR _2572_ _2573_ _0169_ _2576_ sg13g2_a21oi_1
XFILLER_34_540 VPWR VGND sg13g2_fill_2
X_5854_ VGND VPWR net879 net797 _2509_ _2508_ sg13g2_a21oi_1
XFILLER_21_201 VPWR VGND sg13g2_decap_4
X_4805_ _1565_ _1513_ _1562_ VPWR VGND sg13g2_xnor2_1
X_5785_ _2438_ VPWR _2441_ VGND _2439_ _2440_ sg13g2_o21ai_1
XFILLER_30_790 VPWR VGND sg13g2_decap_4
X_4736_ _1498_ _1496_ _1497_ VPWR VGND sg13g2_nand2_1
X_4667_ _1430_ net925 net855 VPWR VGND sg13g2_nand2_1
X_3618_ _0425_ _0426_ _0424_ _0427_ VPWR VGND sg13g2_nand3_1
X_6406_ net1101 VGND VPWR net195 mac2.sum_lvl3_ff\[22\] clknet_leaf_29_clk sg13g2_dfrbpq_1
X_6337_ net1081 VGND VPWR net202 mac2.sum_lvl2_ff\[51\] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_4598_ _1363_ _1364_ _1365_ VPWR VGND sg13g2_nor2b_1
X_3549_ _0359_ _0321_ _0356_ VPWR VGND sg13g2_xnor2_1
X_6268_ net1110 VGND VPWR net175 mac1.sum_lvl1_ff\[44\] clknet_leaf_57_clk sg13g2_dfrbpq_1
X_5219_ _1962_ net878 net811 VPWR VGND sg13g2_nand2_1
X_6199_ net1112 VGND VPWR _0216_ DP_2.matrix\[76\] clknet_leaf_57_clk sg13g2_dfrbpq_2
XFILLER_29_389 VPWR VGND sg13g2_fill_2
XFILLER_44_66 VPWR VGND sg13g2_fill_2
XFILLER_12_223 VPWR VGND sg13g2_fill_1
XFILLER_8_205 VPWR VGND sg13g2_fill_2
XFILLER_5_912 VPWR VGND sg13g2_decap_8
XFILLER_5_27 VPWR VGND sg13g2_fill_1
XFILLER_4_433 VPWR VGND sg13g2_fill_1
Xclkbuf_4_0_0_clk clknet_0_clk clknet_4_0_0_clk VPWR VGND sg13g2_buf_8
XFILLER_5_989 VPWR VGND sg13g2_decap_8
XFILLER_4_444 VPWR VGND sg13g2_fill_1
XFILLER_36_838 VPWR VGND sg13g2_fill_2
XFILLER_44_860 VPWR VGND sg13g2_fill_2
X_5570_ VGND VPWR _2263_ mac2.sum_lvl2_ff\[13\] mac2.sum_lvl2_ff\[32\] sg13g2_or2_1
X_4521_ _1293_ _1284_ _1294_ VPWR VGND sg13g2_nor2b_1
Xhold205 mac2.products_ff\[78\] VPWR VGND net245 sg13g2_dlygate4sd3_1
X_4452_ _1201_ VPWR _1227_ VGND _1195_ _1202_ sg13g2_o21ai_1
Xhold216 mac2.sum_lvl1_ff\[11\] VPWR VGND net256 sg13g2_dlygate4sd3_1
Xhold238 DP_4.matrix\[80\] VPWR VGND net278 sg13g2_dlygate4sd3_1
Xhold227 mac1.sum_lvl2_ff\[0\] VPWR VGND net267 sg13g2_dlygate4sd3_1
X_3403_ _2986_ net990 net1051 VPWR VGND sg13g2_nand2_1
Xhold249 mac1.sum_lvl3_ff\[15\] VPWR VGND net289 sg13g2_dlygate4sd3_1
X_4383_ _1157_ _1158_ _1140_ _1160_ VPWR VGND sg13g2_nand3_1
X_3334_ _2920_ _2909_ _2919_ VPWR VGND sg13g2_xnor2_1
X_6122_ net1135 VGND VPWR _0162_ DP_1.matrix\[80\] clknet_leaf_48_clk sg13g2_dfrbpq_2
X_3265_ _2853_ _2838_ _2852_ VPWR VGND sg13g2_nand2_1
X_6053_ net905 _0229_ VPWR VGND sg13g2_buf_1
X_5004_ _1753_ net886 net818 VPWR VGND sg13g2_nand2_1
X_3196_ _2783_ _2779_ _2785_ VPWR VGND sg13g2_xor2_1
X_5906_ _2560_ net803 net835 VPWR VGND sg13g2_nand2b_1
XFILLER_41_329 VPWR VGND sg13g2_fill_1
X_5837_ _2491_ VPWR _2492_ VGND net924 net805 sg13g2_o21ai_1
X_5768_ _2425_ _2412_ _2424_ VPWR VGND sg13g2_nand2_1
X_4719_ _1476_ VPWR _1481_ VGND _1477_ _1479_ sg13g2_o21ai_1
X_5699_ _2358_ _2356_ _2357_ _2363_ VPWR VGND sg13g2_a21o_1
XFILLER_2_959 VPWR VGND sg13g2_decap_8
XFILLER_29_186 VPWR VGND sg13g2_fill_1
XFILLER_41_874 VPWR VGND sg13g2_fill_1
XFILLER_45_1014 VPWR VGND sg13g2_decap_8
XFILLER_1_970 VPWR VGND sg13g2_decap_8
XFILLER_49_952 VPWR VGND sg13g2_decap_8
X_3050_ _2643_ _2636_ _0066_ VPWR VGND sg13g2_xor2_1
X_3952_ _0743_ _0744_ _0725_ _0746_ VPWR VGND sg13g2_nand3_1
X_3883_ _0677_ _0676_ _0659_ _0679_ VPWR VGND sg13g2_a21o_1
X_5622_ _2302_ VPWR _2303_ VGND _2296_ _2298_ sg13g2_o21ai_1
X_5553_ VPWR _2249_ _2248_ VGND sg13g2_inv_1
X_4504_ _1244_ _1249_ _1278_ VPWR VGND sg13g2_nor2_1
X_5484_ mac1.sum_lvl3_ff\[31\] mac1.sum_lvl3_ff\[11\] _2195_ VPWR VGND sg13g2_nor2_1
X_4435_ _1175_ _1210_ _1211_ VPWR VGND sg13g2_nor2_1
X_4366_ _1143_ net840 net897 VPWR VGND sg13g2_nand2_1
X_6105_ net1063 VGND VPWR _0075_ mac1.products_ff\[69\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3317_ _2903_ net934 net1054 VPWR VGND sg13g2_nand2_1
X_4297_ _1076_ _1069_ _1074_ _1075_ VPWR VGND sg13g2_and3_1
X_6036_ net964 _0204_ VPWR VGND sg13g2_buf_1
X_3248_ _2827_ _2835_ _2836_ VPWR VGND sg13g2_nor2_1
X_3179_ _2744_ VPWR _2769_ VGND _2765_ _2767_ sg13g2_o21ai_1
XFILLER_39_473 VPWR VGND sg13g2_fill_1
XFILLER_27_657 VPWR VGND sg13g2_fill_2
XFILLER_22_362 VPWR VGND sg13g2_fill_2
XFILLER_41_67 VPWR VGND sg13g2_fill_2
XFILLER_1_222 VPWR VGND sg13g2_fill_1
XFILLER_46_966 VPWR VGND sg13g2_decap_8
XFILLER_17_145 VPWR VGND sg13g2_fill_1
XFILLER_18_646 VPWR VGND sg13g2_fill_2
XFILLER_14_874 VPWR VGND sg13g2_decap_8
X_4220_ _0998_ _0999_ _1001_ _1002_ VPWR VGND sg13g2_nor3_1
X_4151_ _0918_ VPWR _0939_ VGND _0915_ _0919_ sg13g2_o21ai_1
X_3102_ _2691_ _2692_ _2686_ _2694_ VPWR VGND sg13g2_nand3_1
X_4082_ VGND VPWR _0836_ _0838_ _0873_ _0872_ sg13g2_a21oi_1
X_3033_ VPWR DP_3.I_range.data_plus_4\[6\] net16 VGND sg13g2_inv_1
XFILLER_37_988 VPWR VGND sg13g2_decap_8
X_4984_ _1732_ _1733_ _1734_ _1735_ VPWR VGND sg13g2_nor3_1
X_3935_ VGND VPWR _0729_ _0727_ _0694_ sg13g2_or2_1
X_3866_ _0662_ net1020 net955 VPWR VGND sg13g2_nand2_1
X_5605_ VPWR VGND _2283_ _2282_ _2281_ mac2.sum_lvl3_ff\[25\] _2289_ net359 sg13g2_a221oi_1
X_6585_ net1075 VGND VPWR net6 DP_1.Q_range.out_data\[3\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_3797_ _0600_ _0593_ _0599_ VPWR VGND sg13g2_nand2_1
X_5536_ _2234_ net549 _0044_ VPWR VGND sg13g2_nor2b_2
X_5467_ _2174_ _2177_ _2180_ _2182_ VPWR VGND sg13g2_or3_1
X_4418_ _1194_ _1142_ _1191_ VPWR VGND sg13g2_xnor2_1
X_5398_ VGND VPWR _2123_ _2125_ _2128_ net393 sg13g2_a21oi_1
X_4349_ _1127_ _1125_ _1126_ VPWR VGND sg13g2_nand2_1
X_6019_ net278 _0171_ VPWR VGND sg13g2_buf_1
XFILLER_14_104 VPWR VGND sg13g2_fill_1
XFILLER_28_988 VPWR VGND sg13g2_decap_8
XFILLER_42_402 VPWR VGND sg13g2_fill_2
XFILLER_35_1013 VPWR VGND sg13g2_decap_8
XFILLER_11_833 VPWR VGND sg13g2_decap_8
XFILLER_6_314 VPWR VGND sg13g2_fill_2
XFILLER_7_0 VPWR VGND sg13g2_fill_1
Xfanout890 net275 net890 VPWR VGND sg13g2_buf_1
XFILLER_46_730 VPWR VGND sg13g2_fill_2
XFILLER_19_944 VPWR VGND sg13g2_decap_8
X_3720_ _0525_ _0518_ _0526_ VPWR VGND sg13g2_nor2b_1
Xclkbuf_leaf_40_clk clknet_4_15_0_clk clknet_leaf_40_clk VPWR VGND sg13g2_buf_8
X_3651_ _0459_ _0453_ _0457_ VPWR VGND sg13g2_xnor2_1
X_3582_ VGND VPWR _0391_ _0390_ _0389_ sg13g2_or2_1
X_6370_ net1085 VGND VPWR net233 mac2.sum_lvl1_ff\[86\] clknet_leaf_20_clk sg13g2_dfrbpq_1
X_5321_ _2026_ _2060_ _2061_ VPWR VGND sg13g2_nor2b_1
XFILLER_6_881 VPWR VGND sg13g2_decap_8
X_5252_ _1980_ VPWR _1994_ VGND _1969_ _1981_ sg13g2_o21ai_1
X_5183_ _1927_ _1926_ _1923_ VPWR VGND sg13g2_nand2b_1
X_4203_ _0987_ net905 net847 _0079_ VPWR VGND sg13g2_and3_2
XFILLER_3_82 VPWR VGND sg13g2_fill_2
X_4134_ _0922_ _0913_ _0923_ VPWR VGND sg13g2_nor2b_1
XFILLER_3_1000 VPWR VGND sg13g2_decap_8
X_4065_ _0830_ VPWR _0856_ VGND _0824_ _0831_ sg13g2_o21ai_1
XFILLER_36_262 VPWR VGND sg13g2_fill_1
XFILLER_25_947 VPWR VGND sg13g2_decap_8
X_4967_ _1720_ _1721_ _0143_ VPWR VGND sg13g2_and2_1
X_4898_ _1655_ _1654_ _1652_ VPWR VGND sg13g2_nand2b_1
X_3918_ _0713_ _0710_ _0712_ VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_31_clk clknet_4_12_0_clk clknet_leaf_31_clk VPWR VGND sg13g2_buf_8
X_3849_ net961 net1017 net965 _0646_ VPWR VGND net1014 sg13g2_nand4_1
X_6568_ net1061 VGND VPWR net326 mac2.total_sum\[0\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_5519_ VGND VPWR _2219_ _2221_ _2222_ _2220_ sg13g2_a21oi_1
X_6499_ net1145 VGND VPWR net70 mac2.sum_lvl1_ff\[15\] clknet_leaf_38_clk sg13g2_dfrbpq_1
Xfanout1107 net1108 net1107 VPWR VGND sg13g2_buf_8
Xfanout1118 net1119 net1118 VPWR VGND sg13g2_buf_8
Xfanout1129 net1130 net1129 VPWR VGND sg13g2_buf_8
XFILLER_47_44 VPWR VGND sg13g2_fill_1
XFILLER_16_903 VPWR VGND sg13g2_decap_8
XFILLER_28_796 VPWR VGND sg13g2_fill_1
XFILLER_8_27 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_22_clk clknet_4_5_0_clk clknet_leaf_22_clk VPWR VGND sg13g2_buf_8
XFILLER_6_133 VPWR VGND sg13g2_fill_1
XFILLER_3_895 VPWR VGND sg13g2_decap_8
XFILLER_46_560 VPWR VGND sg13g2_fill_1
XFILLER_19_796 VPWR VGND sg13g2_fill_1
XFILLER_34_744 VPWR VGND sg13g2_fill_2
X_5870_ net1047 net807 _2525_ VPWR VGND sg13g2_nor2_1
XFILLER_22_917 VPWR VGND sg13g2_decap_8
X_4821_ _1581_ _1547_ _1579_ VPWR VGND sg13g2_xnor2_1
X_4752_ _1513_ net857 net914 VPWR VGND sg13g2_nand2_2
XFILLER_21_449 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_13_clk clknet_4_6_0_clk clknet_leaf_13_clk VPWR VGND sg13g2_buf_8
X_4683_ _1441_ VPWR _1446_ VGND _1442_ _1444_ sg13g2_o21ai_1
X_3703_ _0492_ _0485_ _0455_ _0509_ VPWR VGND sg13g2_a21o_1
X_6422_ net1061 VGND VPWR net383 mac1.total_sum\[2\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_3634_ _0442_ _0437_ _0440_ VPWR VGND sg13g2_xnor2_1
X_3565_ VGND VPWR _0371_ _0372_ _0375_ _0353_ sg13g2_a21oi_1
X_6353_ net1073 VGND VPWR net192 mac1.sum_lvl1_ff\[85\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_5304_ _2044_ _2023_ _2045_ VPWR VGND sg13g2_nor2b_1
X_3496_ _0306_ _0307_ _0268_ _0308_ VPWR VGND sg13g2_nand3_1
X_6284_ net1114 VGND VPWR net156 mac1.sum_lvl2_ff\[8\] clknet_leaf_59_clk sg13g2_dfrbpq_1
X_5235_ _1976_ _1977_ _1978_ VPWR VGND sg13g2_nor2b_1
X_5166_ _1837_ VPWR _1911_ VGND _1907_ _1909_ sg13g2_o21ai_1
X_5097_ VGND VPWR _1843_ _1841_ _1808_ sg13g2_or2_1
X_4117_ _0873_ _0878_ _0907_ VPWR VGND sg13g2_nor2_1
X_4048_ _0804_ _0839_ _0840_ VPWR VGND sg13g2_nor2_1
XFILLER_25_711 VPWR VGND sg13g2_fill_2
X_5999_ _2624_ VPWR _0247_ VGND net790 _2623_ sg13g2_o21ai_1
XFILLER_21_950 VPWR VGND sg13g2_decap_8
XFILLER_40_747 VPWR VGND sg13g2_fill_1
XFILLER_32_1005 VPWR VGND sg13g2_decap_8
XFILLER_3_158 VPWR VGND sg13g2_fill_1
XFILLER_0_854 VPWR VGND sg13g2_decap_8
Xhold9 mac2.products_ff\[68\] VPWR VGND net49 sg13g2_dlygate4sd3_1
XFILLER_48_847 VPWR VGND sg13g2_decap_4
XFILLER_47_335 VPWR VGND sg13g2_fill_2
XFILLER_28_593 VPWR VGND sg13g2_fill_2
XFILLER_43_574 VPWR VGND sg13g2_fill_1
XFILLER_31_714 VPWR VGND sg13g2_fill_2
XFILLER_12_983 VPWR VGND sg13g2_decap_8
XFILLER_7_442 VPWR VGND sg13g2_fill_2
XFILLER_8_976 VPWR VGND sg13g2_decap_8
Xhold409 _0617_ VPWR VGND net449 sg13g2_dlygate4sd3_1
XFILLER_48_1012 VPWR VGND sg13g2_decap_8
X_3350_ _2904_ VPWR _2935_ VGND _2902_ _2905_ sg13g2_o21ai_1
X_5020_ _1748_ VPWR _1769_ VGND _1739_ _1749_ sg13g2_o21ai_1
X_3281_ _2868_ net994 net926 VPWR VGND sg13g2_nand2_1
XFILLER_31_4 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_2_clk clknet_4_0_0_clk clknet_leaf_2_clk VPWR VGND sg13g2_buf_8
XFILLER_17_2 VPWR VGND sg13g2_fill_1
X_5922_ _2573_ _2575_ _2576_ VPWR VGND sg13g2_nor2_1
X_5853_ net794 _2506_ _2507_ _2508_ VPWR VGND sg13g2_nor3_1
XFILLER_22_725 VPWR VGND sg13g2_decap_8
X_4804_ _1513_ _1562_ _1564_ VPWR VGND sg13g2_and2_1
X_5784_ net799 VPWR _2440_ VGND net1052 _2397_ sg13g2_o21ai_1
XFILLER_22_758 VPWR VGND sg13g2_fill_2
XFILLER_21_279 VPWR VGND sg13g2_fill_2
X_4735_ _1459_ _1458_ _1457_ _1497_ VPWR VGND sg13g2_a21o_2
XFILLER_9_92 VPWR VGND sg13g2_fill_2
X_4666_ _1406_ VPWR _1429_ VGND _1381_ _1404_ sg13g2_o21ai_1
X_3617_ _0378_ VPWR _0426_ VGND _0317_ _0379_ sg13g2_o21ai_1
X_6405_ net1101 VGND VPWR net123 mac2.sum_lvl3_ff\[21\] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_4597_ _1360_ VPWR _1364_ VGND _1361_ _1362_ sg13g2_o21ai_1
X_3548_ _0321_ _0356_ _0358_ VPWR VGND sg13g2_and2_1
X_6336_ net1076 VGND VPWR net94 mac2.sum_lvl2_ff\[50\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_3479_ _0290_ _3031_ _0291_ VPWR VGND sg13g2_xor2_1
X_6267_ net1092 VGND VPWR net146 mac1.sum_lvl1_ff\[43\] clknet_leaf_63_clk sg13g2_dfrbpq_1
X_5218_ _1961_ net885 net1042 VPWR VGND sg13g2_nand2_1
X_6198_ net1110 VGND VPWR net149 mac1.sum_lvl1_ff\[6\] clknet_leaf_56_clk sg13g2_dfrbpq_1
X_5149_ _1894_ net1045 net831 net870 net826 VPWR VGND sg13g2_a22oi_1
XFILLER_44_316 VPWR VGND sg13g2_fill_1
XFILLER_44_12 VPWR VGND sg13g2_fill_1
XFILLER_8_217 VPWR VGND sg13g2_decap_4
XFILLER_40_588 VPWR VGND sg13g2_fill_2
XFILLER_21_780 VPWR VGND sg13g2_decap_4
XFILLER_5_968 VPWR VGND sg13g2_decap_8
XFILLER_44_850 VPWR VGND sg13g2_fill_1
X_4520_ _1293_ _1285_ _1292_ VPWR VGND sg13g2_xnor2_1
Xhold206 mac1.products_ff\[10\] VPWR VGND net246 sg13g2_dlygate4sd3_1
X_4451_ _1224_ _1216_ _1226_ VPWR VGND sg13g2_xor2_1
Xhold217 mac2.sum_lvl1_ff\[10\] VPWR VGND net257 sg13g2_dlygate4sd3_1
Xhold239 DP_3.matrix\[78\] VPWR VGND net279 sg13g2_dlygate4sd3_1
Xhold228 _0000_ VPWR VGND net268 sg13g2_dlygate4sd3_1
X_3402_ _2965_ VPWR _2985_ VGND _2937_ _2963_ sg13g2_o21ai_1
X_6121_ net1073 VGND VPWR _0161_ DP_1.matrix\[44\] clknet_leaf_2_clk sg13g2_dfrbpq_2
X_4382_ _1159_ _1140_ _1157_ _1158_ VPWR VGND sg13g2_and3_1
X_3333_ _2919_ _2910_ _2917_ VPWR VGND sg13g2_xnor2_1
X_3264_ _2851_ _2844_ _2852_ VPWR VGND sg13g2_xor2_1
X_6052_ net906 _0228_ VPWR VGND sg13g2_buf_1
XFILLER_39_611 VPWR VGND sg13g2_fill_1
XFILLER_22_1015 VPWR VGND sg13g2_decap_8
X_5003_ _1752_ net818 net889 net820 net886 VPWR VGND sg13g2_a22oi_1
X_3195_ _2779_ _2783_ _2784_ VPWR VGND sg13g2_nor2_1
X_5905_ _2559_ DP_4.matrix\[78\] net797 VPWR VGND sg13g2_nand2_1
X_5836_ VGND VPWR _2634_ net805 _2491_ net795 sg13g2_a21oi_1
XFILLER_10_739 VPWR VGND sg13g2_decap_4
X_5767_ _2423_ _2421_ _2424_ VPWR VGND sg13g2_nor2b_1
X_5698_ VPWR _2362_ _2361_ VGND sg13g2_inv_1
X_4718_ _1476_ _1477_ _1479_ _1480_ VPWR VGND sg13g2_or3_1
X_4649_ _1409_ _1410_ _1412_ _1413_ VPWR VGND sg13g2_or3_1
XFILLER_2_938 VPWR VGND sg13g2_decap_8
X_6319_ net1137 VGND VPWR net102 mac1.sum_lvl2_ff\[49\] clknet_leaf_49_clk sg13g2_dfrbpq_1
XFILLER_45_669 VPWR VGND sg13g2_fill_1
XFILLER_4_231 VPWR VGND sg13g2_fill_2
XFILLER_5_787 VPWR VGND sg13g2_fill_1
XFILLER_49_931 VPWR VGND sg13g2_decap_8
X_3951_ _0745_ _0725_ _0743_ _0744_ VPWR VGND sg13g2_and3_1
XFILLER_17_883 VPWR VGND sg13g2_decap_8
XFILLER_32_831 VPWR VGND sg13g2_decap_4
X_3882_ _0676_ _0677_ _0659_ _0678_ VPWR VGND sg13g2_nand3_1
XFILLER_32_886 VPWR VGND sg13g2_fill_2
X_5621_ net315 mac2.sum_lvl3_ff\[29\] _2302_ VPWR VGND sg13g2_xor2_1
X_5552_ mac2.sum_lvl2_ff\[10\] mac2.sum_lvl2_ff\[29\] _2248_ VPWR VGND sg13g2_xor2_1
X_4503_ _1275_ _1276_ _1277_ VPWR VGND sg13g2_nor2_1
X_5483_ net522 _2191_ _0017_ VPWR VGND sg13g2_xor2_1
X_4434_ _1210_ _1176_ _1208_ VPWR VGND sg13g2_xnor2_1
X_4365_ _1142_ net839 net897 VPWR VGND sg13g2_nand2_2
X_6104_ net1070 VGND VPWR _0074_ mac1.products_ff\[68\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3316_ _2902_ net930 net990 VPWR VGND sg13g2_nand2_1
X_6035_ net987 _0195_ VPWR VGND sg13g2_buf_1
X_4296_ _1070_ VPWR _1075_ VGND _1071_ _1073_ sg13g2_o21ai_1
X_3247_ _2835_ _2828_ _2834_ VPWR VGND sg13g2_xnor2_1
X_3178_ _2744_ _2765_ _2767_ _2768_ VPWR VGND sg13g2_or3_1
XFILLER_41_149 VPWR VGND sg13g2_fill_1
X_5819_ DP_3.I_range.out_data\[2\] DP_3.I_range.out_data\[3\] _2633_ DP_3.I_range.out_data\[4\]
+ _2474_ VPWR VGND sg13g2_nor4_1
XFILLER_41_35 VPWR VGND sg13g2_fill_1
XFILLER_18_625 VPWR VGND sg13g2_fill_2
XFILLER_18_658 VPWR VGND sg13g2_decap_4
XFILLER_17_168 VPWR VGND sg13g2_fill_1
XFILLER_14_853 VPWR VGND sg13g2_decap_8
XFILLER_12_1025 VPWR VGND sg13g2_decap_4
X_4150_ _0921_ _0914_ _0923_ _0938_ VPWR VGND sg13g2_a21o_1
X_3101_ _2693_ _2686_ _2691_ _2692_ VPWR VGND sg13g2_and3_1
X_4081_ _0870_ _0843_ _0872_ VPWR VGND sg13g2_xor2_1
X_3032_ VPWR DP_1.I_range.data_plus_4\[6\] net4 VGND sg13g2_inv_1
X_4983_ _1734_ net884 net831 net826 net887 VPWR VGND sg13g2_a22oi_1
X_3934_ _0728_ net954 net1013 VPWR VGND sg13g2_nand2_1
XFILLER_32_650 VPWR VGND sg13g2_fill_1
X_3865_ _0661_ net1019 net952 VPWR VGND sg13g2_nand2_1
X_5604_ _2288_ net487 mac2.sum_lvl3_ff\[6\] VPWR VGND sg13g2_xnor2_1
X_6584_ net1076 VGND VPWR net5 DP_1.Q_range.out_data\[2\] clknet_leaf_4_clk sg13g2_dfrbpq_2
X_3796_ _0599_ _0594_ _0597_ VPWR VGND sg13g2_xnor2_1
X_5535_ _2232_ VPWR _2235_ VGND _2229_ _2233_ sg13g2_o21ai_1
X_5466_ _2180_ VPWR _2181_ VGND _2174_ _2177_ sg13g2_o21ai_1
X_4417_ _1142_ _1191_ _1193_ VPWR VGND sg13g2_and2_1
X_5397_ _2127_ mac1.sum_lvl2_ff\[27\] net392 VPWR VGND sg13g2_xnor2_1
X_4348_ _1088_ _1087_ _1086_ _1126_ VPWR VGND sg13g2_a21o_2
XFILLER_47_709 VPWR VGND sg13g2_fill_1
X_4279_ _1035_ VPWR _1058_ VGND _1010_ _1033_ sg13g2_o21ai_1
XFILLER_28_923 VPWR VGND sg13g2_fill_2
X_6018_ net1043 _0170_ VPWR VGND sg13g2_buf_1
XFILLER_28_967 VPWR VGND sg13g2_decap_8
XFILLER_27_466 VPWR VGND sg13g2_fill_2
XFILLER_7_849 VPWR VGND sg13g2_decap_8
XFILLER_11_889 VPWR VGND sg13g2_decap_8
XFILLER_42_1018 VPWR VGND sg13g2_decap_8
Xfanout880 net881 net880 VPWR VGND sg13g2_buf_8
XFILLER_19_923 VPWR VGND sg13g2_decap_8
Xfanout891 net892 net891 VPWR VGND sg13g2_buf_2
XFILLER_46_742 VPWR VGND sg13g2_fill_1
XFILLER_18_422 VPWR VGND sg13g2_fill_2
XFILLER_45_252 VPWR VGND sg13g2_fill_2
XFILLER_33_403 VPWR VGND sg13g2_decap_4
XFILLER_18_488 VPWR VGND sg13g2_fill_1
X_3650_ _0458_ _0453_ _0457_ VPWR VGND sg13g2_nand2_1
X_3581_ _0390_ net967 net1039 net970 net1037 VPWR VGND sg13g2_a22oi_1
X_5320_ _2060_ _2055_ _2058_ VPWR VGND sg13g2_xnor2_1
XFILLER_6_860 VPWR VGND sg13g2_decap_8
X_5251_ _1966_ _1960_ _1968_ _1993_ VPWR VGND sg13g2_a21o_1
X_4202_ _2634_ _2635_ _0079_ VPWR VGND sg13g2_nor2_1
X_5182_ _1925_ _1874_ _1926_ VPWR VGND sg13g2_xor2_1
X_4133_ _0922_ _0914_ _0921_ VPWR VGND sg13g2_xnor2_1
X_4064_ _0853_ _0845_ _0855_ VPWR VGND sg13g2_xor2_1
XFILLER_25_926 VPWR VGND sg13g2_decap_8
X_4966_ _1702_ _1704_ _1719_ _1721_ VPWR VGND sg13g2_or3_1
XFILLER_33_981 VPWR VGND sg13g2_decap_8
X_4897_ VGND VPWR _1654_ _1653_ _1601_ sg13g2_or2_1
X_3917_ _0709_ _0708_ _0691_ _0712_ VPWR VGND sg13g2_a21o_1
X_3848_ net965 net961 net1016 net1013 _0645_ VPWR VGND sg13g2_and4_1
XFILLER_20_664 VPWR VGND sg13g2_fill_1
XFILLER_20_697 VPWR VGND sg13g2_fill_1
X_3779_ _0582_ VPWR _0583_ VGND _0557_ _0559_ sg13g2_o21ai_1
X_6567_ net1129 VGND VPWR net486 mac2.sum_lvl3_ff\[15\] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_5518_ net351 _2219_ _0040_ VPWR VGND sg13g2_xor2_1
X_6498_ net1145 VGND VPWR net130 mac2.sum_lvl1_ff\[14\] clknet_leaf_38_clk sg13g2_dfrbpq_1
X_5449_ net442 _2165_ _0025_ VPWR VGND sg13g2_xor2_1
Xfanout1108 net1148 net1108 VPWR VGND sg13g2_buf_8
Xfanout1119 net1130 net1119 VPWR VGND sg13g2_buf_8
XFILLER_47_506 VPWR VGND sg13g2_fill_2
XFILLER_19_219 VPWR VGND sg13g2_fill_2
XFILLER_43_701 VPWR VGND sg13g2_fill_2
XFILLER_43_745 VPWR VGND sg13g2_fill_2
XFILLER_16_959 VPWR VGND sg13g2_decap_8
XFILLER_42_200 VPWR VGND sg13g2_fill_2
XFILLER_30_417 VPWR VGND sg13g2_fill_2
XFILLER_11_686 VPWR VGND sg13g2_fill_1
XFILLER_6_178 VPWR VGND sg13g2_fill_1
XFILLER_3_874 VPWR VGND sg13g2_decap_8
XFILLER_2_395 VPWR VGND sg13g2_fill_2
XFILLER_46_550 VPWR VGND sg13g2_fill_1
XFILLER_46_583 VPWR VGND sg13g2_fill_1
X_4820_ _1580_ _1547_ _1579_ VPWR VGND sg13g2_nand2b_1
XFILLER_15_981 VPWR VGND sg13g2_decap_8
X_4751_ _1512_ net919 net856 VPWR VGND sg13g2_nand2_1
X_3702_ _0494_ VPWR _0508_ VGND _0483_ _0495_ sg13g2_o21ai_1
X_4682_ _1441_ _1442_ _1444_ _1445_ VPWR VGND sg13g2_or3_1
X_6421_ net1061 VGND VPWR net293 mac1.total_sum\[1\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_3633_ _0441_ _0440_ _0437_ VPWR VGND sg13g2_nand2b_1
X_3564_ _0371_ _0372_ _0353_ _0374_ VPWR VGND sg13g2_nand3_1
X_6352_ net1073 VGND VPWR net263 mac1.sum_lvl1_ff\[84\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_5303_ _2042_ _2041_ _2044_ VPWR VGND sg13g2_xor2_1
X_3495_ _0305_ _0304_ _0287_ _0307_ VPWR VGND sg13g2_a21o_1
X_6283_ net1114 VGND VPWR net168 mac1.sum_lvl2_ff\[7\] clknet_leaf_57_clk sg13g2_dfrbpq_1
X_5234_ _1972_ VPWR _1977_ VGND _1974_ _1975_ sg13g2_o21ai_1
X_5165_ _1837_ _1907_ _1909_ _1910_ VPWR VGND sg13g2_or3_1
XFILLER_25_1024 VPWR VGND sg13g2_decap_4
X_4116_ _0904_ _0905_ _0906_ VPWR VGND sg13g2_nor2_1
X_5096_ _1842_ net820 net877 VPWR VGND sg13g2_nand2_1
X_4047_ _0839_ _0805_ _0837_ VPWR VGND sg13g2_xnor2_1
XFILLER_37_561 VPWR VGND sg13g2_fill_1
XFILLER_25_745 VPWR VGND sg13g2_decap_8
X_5998_ _2624_ net859 net790 VPWR VGND sg13g2_nand2_1
XFILLER_25_778 VPWR VGND sg13g2_decap_4
XFILLER_33_25 VPWR VGND sg13g2_fill_1
X_4949_ _1704_ _1697_ _1703_ VPWR VGND sg13g2_nand2_1
XFILLER_32_1028 VPWR VGND sg13g2_fill_1
XFILLER_3_137 VPWR VGND sg13g2_fill_2
XFILLER_0_833 VPWR VGND sg13g2_decap_8
XFILLER_48_859 VPWR VGND sg13g2_fill_1
XFILLER_16_701 VPWR VGND sg13g2_fill_1
XFILLER_16_723 VPWR VGND sg13g2_fill_2
XFILLER_15_244 VPWR VGND sg13g2_fill_2
XFILLER_12_962 VPWR VGND sg13g2_decap_8
XFILLER_8_955 VPWR VGND sg13g2_decap_8
XFILLER_11_483 VPWR VGND sg13g2_fill_2
X_3280_ _2867_ net998 net1051 VPWR VGND sg13g2_nand2_1
XFILLER_24_4 VPWR VGND sg13g2_fill_1
X_5921_ _2574_ VPWR _2575_ VGND net791 _2571_ sg13g2_o21ai_1
XFILLER_0_1015 VPWR VGND sg13g2_decap_8
XFILLER_34_542 VPWR VGND sg13g2_fill_1
X_5852_ net898 net807 _2507_ VPWR VGND sg13g2_nor2_1
X_4803_ VGND VPWR _1563_ _1562_ _1513_ sg13g2_or2_1
X_5783_ net1053 net809 _2439_ VPWR VGND sg13g2_nor2_1
XFILLER_22_737 VPWR VGND sg13g2_decap_8
X_4734_ _1495_ _1431_ _1496_ VPWR VGND sg13g2_xor2_1
X_4665_ _1428_ _1420_ _1422_ VPWR VGND sg13g2_nand2_1
X_3616_ _0351_ VPWR _0425_ VGND _0421_ _0423_ sg13g2_o21ai_1
X_6404_ net1102 VGND VPWR net116 mac2.sum_lvl3_ff\[20\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_4596_ _1360_ _1361_ _1362_ _1363_ VPWR VGND sg13g2_nor3_1
X_3547_ VGND VPWR _0357_ _0355_ _0322_ sg13g2_or2_1
X_6335_ net1077 VGND VPWR net69 mac2.sum_lvl2_ff\[49\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_6266_ net1092 VGND VPWR net189 mac1.sum_lvl1_ff\[42\] clknet_leaf_63_clk sg13g2_dfrbpq_1
X_3478_ _0290_ net1037 net974 VPWR VGND sg13g2_nand2_1
X_5217_ _1935_ VPWR _1960_ VGND _1933_ _1936_ sg13g2_o21ai_1
X_6197_ net1117 VGND VPWR _0215_ DP_2.matrix\[75\] clknet_leaf_53_clk sg13g2_dfrbpq_2
X_5148_ net827 net870 net831 _1893_ VPWR VGND net1045 sg13g2_nand4_1
X_5079_ _1823_ _1822_ _1805_ _1826_ VPWR VGND sg13g2_a21o_1
XFILLER_25_575 VPWR VGND sg13g2_fill_1
XFILLER_40_534 VPWR VGND sg13g2_decap_8
XFILLER_40_545 VPWR VGND sg13g2_fill_1
XFILLER_8_207 VPWR VGND sg13g2_fill_1
XFILLER_5_947 VPWR VGND sg13g2_decap_8
XFILLER_18_91 VPWR VGND sg13g2_fill_2
XFILLER_44_862 VPWR VGND sg13g2_fill_1
XFILLER_15_1023 VPWR VGND sg13g2_decap_4
X_4450_ _1224_ _1216_ _1225_ VPWR VGND sg13g2_nor2b_1
Xhold207 mac2.sum_lvl1_ff\[8\] VPWR VGND net247 sg13g2_dlygate4sd3_1
Xhold229 DP_4.matrix\[76\] VPWR VGND net269 sg13g2_dlygate4sd3_1
X_3401_ _2968_ _2960_ _2967_ _2984_ VPWR VGND sg13g2_a21o_1
X_4381_ _1146_ VPWR _1158_ VGND _1154_ _1156_ sg13g2_o21ai_1
Xhold218 mac2.products_ff\[149\] VPWR VGND net258 sg13g2_dlygate4sd3_1
X_6120_ net1095 VGND VPWR _0160_ DP_1.matrix\[8\] clknet_leaf_61_clk sg13g2_dfrbpq_1
X_3332_ _2917_ _2910_ _2918_ VPWR VGND sg13g2_nor2b_1
X_6051_ net926 _0219_ VPWR VGND sg13g2_buf_1
X_3263_ _2851_ _2845_ _2849_ VPWR VGND sg13g2_xnor2_1
X_3194_ VGND VPWR _2783_ _2782_ _2781_ sg13g2_or2_1
X_5002_ _0092_ _1738_ _1750_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_328 VPWR VGND sg13g2_fill_2
X_5904_ _2558_ _2533_ _2557_ VPWR VGND sg13g2_nand2b_1
X_5835_ _2490_ net275 net798 VPWR VGND sg13g2_nand2_1
X_5766_ _2423_ net800 _2422_ net801 net999 VPWR VGND sg13g2_a22oi_1
XFILLER_22_589 VPWR VGND sg13g2_fill_1
X_5697_ mac2.total_sum\[10\] mac1.total_sum\[10\] _2361_ VPWR VGND sg13g2_xor2_1
X_4717_ _1479_ net909 net867 net911 net864 VPWR VGND sg13g2_a22oi_1
X_4648_ _1412_ net915 net868 net916 net865 VPWR VGND sg13g2_a22oi_1
XFILLER_2_917 VPWR VGND sg13g2_decap_8
X_4579_ _1349_ _1333_ _0132_ VPWR VGND sg13g2_xor2_1
X_6318_ net1133 VGND VPWR net109 mac1.sum_lvl2_ff\[48\] clknet_leaf_49_clk sg13g2_dfrbpq_1
X_6249_ net1139 VGND VPWR _0257_ DP_4.matrix\[41\] clknet_leaf_44_clk sg13g2_dfrbpq_2
XFILLER_18_807 VPWR VGND sg13g2_decap_8
XFILLER_17_339 VPWR VGND sg13g2_fill_1
XFILLER_25_361 VPWR VGND sg13g2_fill_1
XFILLER_38_1023 VPWR VGND sg13g2_decap_4
XFILLER_13_545 VPWR VGND sg13g2_fill_2
XFILLER_20_70 VPWR VGND sg13g2_fill_1
XFILLER_49_910 VPWR VGND sg13g2_decap_8
XFILLER_49_987 VPWR VGND sg13g2_decap_8
Xhold90 mac2.products_ff\[14\] VPWR VGND net130 sg13g2_dlygate4sd3_1
X_3950_ _0732_ VPWR _0744_ VGND _0740_ _0742_ sg13g2_o21ai_1
XFILLER_17_862 VPWR VGND sg13g2_decap_8
XFILLER_44_681 VPWR VGND sg13g2_fill_1
XFILLER_32_821 VPWR VGND sg13g2_fill_2
X_3881_ _0665_ VPWR _0677_ VGND _0673_ _0675_ sg13g2_o21ai_1
XFILLER_31_320 VPWR VGND sg13g2_fill_1
X_5620_ _2301_ mac2.sum_lvl3_ff\[29\] net315 VPWR VGND sg13g2_nand2_1
X_5551_ _2247_ mac2.sum_lvl2_ff\[29\] mac2.sum_lvl2_ff\[10\] VPWR VGND sg13g2_nand2_1
X_4502_ VGND VPWR _1240_ _1242_ _1276_ _1273_ sg13g2_a21oi_1
X_5482_ _2194_ _2191_ _2193_ VPWR VGND sg13g2_nand2_1
X_4433_ _1209_ _1176_ _1208_ VPWR VGND sg13g2_nand2b_1
X_4364_ _1141_ net901 net837 VPWR VGND sg13g2_nand2_1
X_3315_ _2884_ _2877_ _2847_ _2901_ VPWR VGND sg13g2_a21o_1
X_4295_ _1070_ _1071_ _1073_ _1074_ VPWR VGND sg13g2_or3_1
X_6103_ net1084 VGND VPWR _0111_ mac1.products_ff\[15\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_6_1021 VPWR VGND sg13g2_decap_8
X_6034_ net989 _0194_ VPWR VGND sg13g2_buf_1
X_3246_ _2834_ _2829_ _2832_ VPWR VGND sg13g2_xnor2_1
X_3177_ VGND VPWR _2763_ _2764_ _2767_ _2745_ sg13g2_a21oi_1
XFILLER_39_486 VPWR VGND sg13g2_fill_1
XFILLER_27_659 VPWR VGND sg13g2_fill_1
X_5818_ DP_3.Q_range.out_data\[2\] net505 _2472_ _2473_ VPWR VGND sg13g2_nor3_1
X_5749_ VGND VPWR net787 _2405_ _2406_ _2394_ sg13g2_a21oi_1
XFILLER_41_69 VPWR VGND sg13g2_fill_1
XFILLER_17_136 VPWR VGND sg13g2_fill_1
XFILLER_18_648 VPWR VGND sg13g2_fill_1
XFILLER_41_651 VPWR VGND sg13g2_fill_2
XFILLER_12_1004 VPWR VGND sg13g2_decap_8
X_3100_ _2687_ VPWR _2692_ VGND _2688_ _2690_ sg13g2_o21ai_1
X_4080_ _0871_ _0870_ _0843_ VPWR VGND sg13g2_nand2b_1
XFILLER_49_784 VPWR VGND sg13g2_fill_2
X_4982_ net830 net887 net825 net884 _1733_ VPWR VGND sg13g2_and4_1
X_3933_ _0727_ net1014 net952 VPWR VGND sg13g2_nand2_1
X_3864_ _0660_ net1023 net951 VPWR VGND sg13g2_nand2_1
XFILLER_31_150 VPWR VGND sg13g2_fill_2
XFILLER_20_846 VPWR VGND sg13g2_decap_4
XFILLER_32_695 VPWR VGND sg13g2_fill_2
X_5603_ net487 mac2.sum_lvl3_ff\[6\] _2287_ VPWR VGND sg13g2_and2_1
X_3795_ _0598_ _0597_ _0594_ VPWR VGND sg13g2_nand2b_1
X_6583_ net1074 VGND VPWR net439 mac2.total_sum\[15\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_5534_ _2229_ _2232_ _2233_ _2234_ VPWR VGND sg13g2_nor3_2
X_5465_ mac1.sum_lvl3_ff\[7\] mac1.sum_lvl3_ff\[27\] _2180_ VPWR VGND sg13g2_xor2_1
X_4416_ VGND VPWR _1192_ _1191_ _1142_ sg13g2_or2_1
X_5396_ net537 _2126_ _0013_ VPWR VGND sg13g2_and2_1
X_4347_ _1124_ _1060_ _1125_ VPWR VGND sg13g2_xor2_1
X_4278_ _1057_ _1049_ _1051_ VPWR VGND sg13g2_nand2_1
X_6017_ net273 _0168_ VPWR VGND sg13g2_buf_1
X_3229_ _2770_ VPWR _2818_ VGND _2709_ _2771_ sg13g2_o21ai_1
XFILLER_42_404 VPWR VGND sg13g2_fill_1
XFILLER_14_128 VPWR VGND sg13g2_fill_2
XFILLER_7_806 VPWR VGND sg13g2_fill_2
XFILLER_6_316 VPWR VGND sg13g2_fill_1
XFILLER_11_868 VPWR VGND sg13g2_decap_8
Xhold390 _0020_ VPWR VGND net430 sg13g2_dlygate4sd3_1
Xfanout870 net872 net870 VPWR VGND sg13g2_buf_8
Xfanout881 net882 net881 VPWR VGND sg13g2_buf_1
XFILLER_19_902 VPWR VGND sg13g2_decap_8
Xfanout892 net893 net892 VPWR VGND sg13g2_buf_1
XFILLER_45_220 VPWR VGND sg13g2_fill_2
XFILLER_18_445 VPWR VGND sg13g2_decap_8
XFILLER_19_979 VPWR VGND sg13g2_decap_8
XFILLER_13_194 VPWR VGND sg13g2_fill_1
XFILLER_41_481 VPWR VGND sg13g2_fill_2
XFILLER_9_198 VPWR VGND sg13g2_fill_2
X_3580_ net1039 net1037 net970 net967 _0389_ VPWR VGND sg13g2_and4_1
XFILLER_42_90 VPWR VGND sg13g2_fill_1
X_5250_ _1991_ _1989_ _0150_ VPWR VGND sg13g2_xor2_1
X_4201_ _0122_ _0979_ _0986_ VPWR VGND sg13g2_xnor2_1
X_5181_ _1925_ net881 net814 VPWR VGND sg13g2_nand2_1
X_4132_ _0921_ _0915_ _0920_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_84 VPWR VGND sg13g2_fill_1
X_4063_ _0853_ _0845_ _0854_ VPWR VGND sg13g2_nor2b_1
XFILLER_24_404 VPWR VGND sg13g2_fill_2
X_4965_ _1719_ VPWR _1720_ VGND _1702_ _1704_ sg13g2_o21ai_1
XFILLER_36_297 VPWR VGND sg13g2_fill_2
X_3916_ VGND VPWR _0708_ _0709_ _0711_ _0691_ sg13g2_a21oi_1
X_4896_ _1653_ DP_4.matrix\[5\] net1049 VPWR VGND sg13g2_nand2_2
X_3847_ _0644_ net1018 net957 VPWR VGND sg13g2_nand2_1
XFILLER_22_27 VPWR VGND sg13g2_fill_1
X_3778_ _0581_ _0567_ _0582_ VPWR VGND sg13g2_xor2_1
X_6566_ net1084 VGND VPWR _0037_ mac2.sum_lvl3_ff\[14\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_5517_ net350 mac2.sum_lvl2_ff\[21\] _2221_ VPWR VGND sg13g2_xor2_1
X_6497_ net1142 VGND VPWR net242 mac2.sum_lvl1_ff\[13\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_5448_ _2167_ mac1.sum_lvl3_ff\[23\] net441 VPWR VGND sg13g2_xnor2_1
Xfanout1109 net1113 net1109 VPWR VGND sg13g2_buf_8
X_5379_ mac1.sum_lvl2_ff\[23\] net340 _2113_ VPWR VGND sg13g2_and2_1
XFILLER_16_938 VPWR VGND sg13g2_decap_8
XFILLER_15_448 VPWR VGND sg13g2_fill_1
XFILLER_15_459 VPWR VGND sg13g2_decap_4
XFILLER_24_982 VPWR VGND sg13g2_decap_8
XFILLER_23_481 VPWR VGND sg13g2_fill_2
XFILLER_3_853 VPWR VGND sg13g2_decap_8
XFILLER_26_8 VPWR VGND sg13g2_fill_1
XFILLER_18_220 VPWR VGND sg13g2_fill_1
XFILLER_15_960 VPWR VGND sg13g2_decap_8
X_4750_ _1483_ VPWR _1511_ VGND _1474_ _1484_ sg13g2_o21ai_1
X_3701_ _0480_ _0474_ _0482_ _0507_ VPWR VGND sg13g2_a21o_1
X_4681_ _1444_ net913 net867 net914 net864 VPWR VGND sg13g2_a22oi_1
X_6420_ net1061 VGND VPWR net266 mac1.total_sum\[0\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_3632_ _0439_ _0388_ _0440_ VPWR VGND sg13g2_xor2_1
XFILLER_30_985 VPWR VGND sg13g2_decap_8
X_6351_ net1133 VGND VPWR net57 mac1.sum_lvl1_ff\[83\] clknet_leaf_49_clk sg13g2_dfrbpq_1
X_5302_ _2042_ _2041_ _2043_ VPWR VGND sg13g2_nor2b_1
X_3563_ _0373_ _0353_ _0371_ _0372_ VPWR VGND sg13g2_and3_1
XFILLER_45_0 VPWR VGND sg13g2_fill_2
X_3494_ _0304_ _0305_ _0287_ _0306_ VPWR VGND sg13g2_nand3_1
X_6282_ net1111 VGND VPWR net73 mac1.sum_lvl2_ff\[6\] clknet_leaf_56_clk sg13g2_dfrbpq_1
X_5233_ _1972_ _1974_ _1975_ _1976_ VPWR VGND sg13g2_nor3_1
X_5164_ VGND VPWR _1905_ _1906_ _1909_ _1871_ sg13g2_a21oi_1
XFILLER_25_1003 VPWR VGND sg13g2_decap_8
X_4115_ VGND VPWR _0869_ _0871_ _0905_ _0902_ sg13g2_a21oi_1
X_5095_ _1841_ net877 net818 VPWR VGND sg13g2_nand2_1
X_4046_ _0838_ _0805_ _0837_ VPWR VGND sg13g2_nand2b_1
XFILLER_25_713 VPWR VGND sg13g2_fill_1
X_5997_ _2551_ _2537_ _2623_ VPWR VGND sg13g2_xor2_1
XFILLER_13_919 VPWR VGND sg13g2_decap_8
X_4948_ _1703_ _1676_ _1698_ VPWR VGND sg13g2_nand2_1
X_4879_ _1637_ _1590_ _1635_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_451 VPWR VGND sg13g2_fill_1
XFILLER_20_484 VPWR VGND sg13g2_decap_8
XFILLER_21_985 VPWR VGND sg13g2_decap_8
X_6549_ net1076 VGND VPWR net2 DP_1.I_range.out_data\[3\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_0_812 VPWR VGND sg13g2_decap_8
XFILLER_0_889 VPWR VGND sg13g2_decap_8
XFILLER_16_746 VPWR VGND sg13g2_fill_2
XFILLER_31_716 VPWR VGND sg13g2_fill_1
XFILLER_12_941 VPWR VGND sg13g2_decap_8
XFILLER_31_738 VPWR VGND sg13g2_fill_1
XFILLER_8_934 VPWR VGND sg13g2_decap_8
XFILLER_7_411 VPWR VGND sg13g2_fill_1
XFILLER_23_70 VPWR VGND sg13g2_fill_1
XFILLER_7_444 VPWR VGND sg13g2_fill_1
X_5920_ _2574_ net1044 net791 VPWR VGND sg13g2_nand2_1
X_5851_ net916 net804 _2506_ VPWR VGND sg13g2_nor2_1
X_4802_ _1562_ net860 net911 VPWR VGND sg13g2_nand2_1
X_5782_ _2438_ net386 net802 VPWR VGND sg13g2_nand2_1
XFILLER_21_237 VPWR VGND sg13g2_fill_2
X_4733_ _1495_ _1492_ _1494_ VPWR VGND sg13g2_nand2_1
XFILLER_30_771 VPWR VGND sg13g2_fill_1
X_6403_ net1096 VGND VPWR net286 mac1.sum_lvl3_ff\[15\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_4664_ _0138_ _1400_ _1427_ VPWR VGND sg13g2_xnor2_1
X_3615_ _0351_ _0421_ _0423_ _0424_ VPWR VGND sg13g2_or3_1
X_4595_ _1362_ net920 net869 net863 net923 VPWR VGND sg13g2_a22oi_1
X_3546_ _0356_ net974 net1032 VPWR VGND sg13g2_nand2_1
X_6334_ net1077 VGND VPWR net106 mac2.sum_lvl2_ff\[48\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_6265_ net1092 VGND VPWR net237 mac1.sum_lvl1_ff\[41\] clknet_leaf_62_clk sg13g2_dfrbpq_1
X_5216_ _1927_ VPWR _1959_ VGND _1874_ _1925_ sg13g2_o21ai_1
X_3477_ _0289_ net1037 net972 VPWR VGND sg13g2_nand2_1
X_6196_ net1131 VGND VPWR _0214_ DP_2.matrix\[74\] clknet_leaf_52_clk sg13g2_dfrbpq_1
X_5147_ net831 net826 net870 net1045 _1892_ VPWR VGND sg13g2_and4_1
X_5078_ VGND VPWR _1822_ _1823_ _1825_ _1805_ sg13g2_a21oi_1
X_4029_ VGND VPWR _0821_ _0820_ _0771_ sg13g2_or2_1
XFILLER_40_524 VPWR VGND sg13g2_fill_1
XFILLER_5_926 VPWR VGND sg13g2_decap_8
XFILLER_47_112 VPWR VGND sg13g2_fill_2
XFILLER_36_819 VPWR VGND sg13g2_fill_2
XFILLER_16_565 VPWR VGND sg13g2_fill_1
XFILLER_15_1002 VPWR VGND sg13g2_decap_8
XFILLER_7_241 VPWR VGND sg13g2_fill_1
XFILLER_8_775 VPWR VGND sg13g2_fill_2
Xhold208 mac1.sum_lvl1_ff\[84\] VPWR VGND net248 sg13g2_dlygate4sd3_1
X_3400_ VGND VPWR _2959_ _2973_ _2983_ _2972_ sg13g2_a21oi_1
X_4380_ _1146_ _1154_ _1156_ _1157_ VPWR VGND sg13g2_or3_1
Xhold219 mac2.sum_lvl1_ff\[9\] VPWR VGND net259 sg13g2_dlygate4sd3_1
X_3331_ _2917_ _2911_ _2916_ VPWR VGND sg13g2_xnor2_1
XFILLER_4_992 VPWR VGND sg13g2_decap_8
X_6050_ net929 _0218_ VPWR VGND sg13g2_buf_1
X_3262_ _2850_ _2845_ _2849_ VPWR VGND sg13g2_nand2_1
X_3193_ _2782_ net927 net1000 net929 net998 VPWR VGND sg13g2_a22oi_1
X_5001_ _1751_ _1750_ _1738_ VPWR VGND sg13g2_nand2b_1
X_5903_ _2557_ _2556_ _2552_ VPWR VGND sg13g2_nand2b_1
X_5834_ _2488_ VPWR _2489_ VGND net795 _2487_ sg13g2_o21ai_1
X_5765_ net1036 net1020 net809 _2422_ VPWR VGND sg13g2_mux2_1
X_5696_ _2360_ mac1.total_sum\[10\] mac2.total_sum\[10\] VPWR VGND sg13g2_nand2_1
X_4716_ net864 net911 DP_4.matrix\[0\] _1478_ VPWR VGND net909 sg13g2_nand4_1
X_4647_ net865 net916 net868 _1411_ VPWR VGND net915 sg13g2_nand4_1
X_6317_ net1138 VGND VPWR net138 mac1.sum_lvl2_ff\[47\] clknet_leaf_51_clk sg13g2_dfrbpq_1
X_4578_ _1347_ _1334_ _1349_ VPWR VGND sg13g2_xor2_1
X_3529_ _0337_ _0336_ _0319_ _0340_ VPWR VGND sg13g2_a21o_1
X_6248_ net1139 VGND VPWR _0256_ DP_4.matrix\[40\] clknet_leaf_45_clk sg13g2_dfrbpq_1
X_6179_ net1094 VGND VPWR net378 DP_2.matrix\[7\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_45_627 VPWR VGND sg13g2_fill_1
XFILLER_44_104 VPWR VGND sg13g2_fill_1
XFILLER_38_1002 VPWR VGND sg13g2_decap_8
XFILLER_41_833 VPWR VGND sg13g2_fill_1
XFILLER_4_266 VPWR VGND sg13g2_fill_2
XFILLER_45_1028 VPWR VGND sg13g2_fill_1
XFILLER_1_984 VPWR VGND sg13g2_decap_8
XFILLER_49_966 VPWR VGND sg13g2_decap_8
Xhold80 mac1.products_ff\[71\] VPWR VGND net120 sg13g2_dlygate4sd3_1
Xhold91 mac2.products_ff\[74\] VPWR VGND net131 sg13g2_dlygate4sd3_1
XFILLER_17_841 VPWR VGND sg13g2_decap_8
X_3880_ _0665_ _0673_ _0675_ _0676_ VPWR VGND sg13g2_or3_1
XFILLER_32_877 VPWR VGND sg13g2_fill_2
X_5550_ _0047_ _2243_ _2246_ VPWR VGND sg13g2_xnor2_1
X_5481_ net521 mac1.sum_lvl3_ff\[30\] _2193_ VPWR VGND sg13g2_xor2_1
X_4501_ VPWR _1275_ _1274_ VGND sg13g2_inv_1
X_4432_ _1208_ _1177_ _1206_ VPWR VGND sg13g2_xnor2_1
X_4363_ _1112_ VPWR _1140_ VGND _1103_ _1113_ sg13g2_o21ai_1
X_3314_ _2886_ VPWR _2900_ VGND _2875_ _2887_ sg13g2_o21ai_1
X_4294_ _1073_ net894 net848 net896 net844 VPWR VGND sg13g2_a22oi_1
X_6102_ net1097 VGND VPWR _0110_ mac1.products_ff\[14\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_6_1000 VPWR VGND sg13g2_decap_8
X_3245_ _2833_ _2832_ _2829_ VPWR VGND sg13g2_nand2b_1
X_6033_ net991 _0193_ VPWR VGND sg13g2_buf_1
X_3176_ _2763_ _2764_ _2745_ _2766_ VPWR VGND sg13g2_nand3_1
XFILLER_27_605 VPWR VGND sg13g2_fill_1
XFILLER_27_627 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_61_clk clknet_4_3_0_clk clknet_leaf_61_clk VPWR VGND sg13g2_buf_8
X_5817_ _2472_ DP_3.Q_range.out_data\[3\] DP_3.Q_range.out_data\[5\] VPWR VGND sg13g2_nand2_1
X_5748_ _2399_ VPWR _2405_ VGND _2403_ _2404_ sg13g2_o21ai_1
X_5679_ _2342_ _2345_ _2346_ _2347_ VPWR VGND sg13g2_nor3_1
XFILLER_18_627 VPWR VGND sg13g2_fill_1
XFILLER_45_446 VPWR VGND sg13g2_fill_2
XFILLER_17_126 VPWR VGND sg13g2_fill_2
XFILLER_26_693 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_52_clk clknet_4_10_0_clk clknet_leaf_52_clk VPWR VGND sg13g2_buf_8
XFILLER_14_888 VPWR VGND sg13g2_decap_8
XFILLER_9_347 VPWR VGND sg13g2_fill_2
XFILLER_1_781 VPWR VGND sg13g2_decap_8
X_4981_ _1732_ net890 net822 VPWR VGND sg13g2_nand2_1
X_3932_ _0726_ net1019 DP_2.matrix\[41\] VPWR VGND sg13g2_nand2_1
XFILLER_16_170 VPWR VGND sg13g2_fill_2
XFILLER_16_192 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_43_clk clknet_4_11_0_clk clknet_leaf_43_clk VPWR VGND sg13g2_buf_8
X_3863_ _0650_ VPWR _0659_ VGND _0642_ _0651_ sg13g2_o21ai_1
X_5602_ _0059_ _2284_ net360 VPWR VGND sg13g2_xnor2_1
X_6582_ net1066 VGND VPWR net299 mac2.total_sum\[14\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_3794_ _0596_ _0570_ _0597_ VPWR VGND sg13g2_xor2_1
X_5533_ VPWR VGND _2227_ _2226_ _2225_ mac2.sum_lvl2_ff\[24\] _2233_ mac2.sum_lvl2_ff\[5\]
+ sg13g2_a221oi_1
X_5464_ _2179_ mac1.sum_lvl3_ff\[27\] mac1.sum_lvl3_ff\[7\] VPWR VGND sg13g2_nand2_1
X_5395_ _2118_ _2121_ net536 _2126_ VPWR VGND sg13g2_or3_1
X_4415_ _1191_ net841 net895 VPWR VGND sg13g2_nand2_1
X_4346_ _1124_ _1121_ _1123_ VPWR VGND sg13g2_nand2_1
XFILLER_28_1023 VPWR VGND sg13g2_decap_4
X_4277_ _0127_ _1029_ _1056_ VPWR VGND sg13g2_xnor2_1
X_3228_ _2743_ VPWR _2817_ VGND _2813_ _2815_ sg13g2_o21ai_1
X_6016_ net1047 _0167_ VPWR VGND sg13g2_buf_1
X_3159_ VGND VPWR _2749_ _2747_ _2714_ sg13g2_or2_1
XFILLER_27_446 VPWR VGND sg13g2_fill_1
XFILLER_27_468 VPWR VGND sg13g2_fill_1
XFILLER_36_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_34_clk clknet_4_15_0_clk clknet_leaf_34_clk VPWR VGND sg13g2_buf_8
XFILLER_23_663 VPWR VGND sg13g2_decap_4
XFILLER_35_1027 VPWR VGND sg13g2_fill_2
XFILLER_11_847 VPWR VGND sg13g2_decap_8
XFILLER_6_339 VPWR VGND sg13g2_fill_1
Xhold380 DP_3.matrix\[4\] VPWR VGND net420 sg13g2_dlygate4sd3_1
Xhold391 DP_2.matrix\[39\] VPWR VGND net431 sg13g2_dlygate4sd3_1
XFILLER_2_567 VPWR VGND sg13g2_fill_1
Xfanout860 DP_4.matrix\[3\] net860 VPWR VGND sg13g2_buf_1
Xfanout882 net301 net882 VPWR VGND sg13g2_buf_2
Xfanout871 net872 net871 VPWR VGND sg13g2_buf_1
Xfanout893 net529 net893 VPWR VGND sg13g2_buf_8
XFILLER_18_424 VPWR VGND sg13g2_fill_1
XFILLER_19_958 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_25_clk clknet_4_13_0_clk clknet_leaf_25_clk VPWR VGND sg13g2_buf_8
XFILLER_42_983 VPWR VGND sg13g2_decap_8
XFILLER_9_188 VPWR VGND sg13g2_fill_2
XFILLER_6_895 VPWR VGND sg13g2_decap_8
XFILLER_5_361 VPWR VGND sg13g2_fill_2
X_4200_ _0986_ _0980_ _0985_ VPWR VGND sg13g2_xnor2_1
X_5180_ _1924_ net882 net811 VPWR VGND sg13g2_nand2_1
X_4131_ _0917_ _0919_ _0920_ VPWR VGND sg13g2_nor2_1
X_4062_ _0853_ _0846_ _0852_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_1014 VPWR VGND sg13g2_decap_8
XFILLER_36_232 VPWR VGND sg13g2_fill_1
XFILLER_18_980 VPWR VGND sg13g2_decap_8
X_4964_ _1718_ _1705_ _1719_ VPWR VGND sg13g2_xor2_1
Xclkbuf_leaf_16_clk clknet_4_4_0_clk clknet_leaf_16_clk VPWR VGND sg13g2_buf_8
X_3915_ _0708_ _0709_ _0691_ _0710_ VPWR VGND sg13g2_nand3_1
X_4895_ _1652_ net1049 net858 net908 net856 VPWR VGND sg13g2_a22oi_1
X_3846_ _0629_ VPWR _0643_ VGND _0627_ _0630_ sg13g2_o21ai_1
X_3777_ _0579_ _0554_ _0581_ VPWR VGND sg13g2_xor2_1
X_6565_ net1084 VGND VPWR _0036_ mac2.sum_lvl3_ff\[13\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_5516_ mac2.sum_lvl2_ff\[21\] net350 _2220_ VPWR VGND sg13g2_and2_1
X_6496_ net1142 VGND VPWR net225 mac2.sum_lvl1_ff\[12\] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_5447_ _2166_ mac1.sum_lvl3_ff\[23\] mac1.sum_lvl3_ff\[3\] VPWR VGND sg13g2_nand2_1
X_5378_ _2110_ VPWR _2112_ VGND _2109_ _2111_ sg13g2_o21ai_1
X_4329_ net844 net894 net848 _1107_ VPWR VGND net891 sg13g2_nand4_1
XFILLER_47_508 VPWR VGND sg13g2_fill_1
XFILLER_16_917 VPWR VGND sg13g2_decap_8
XFILLER_28_744 VPWR VGND sg13g2_decap_4
XFILLER_28_777 VPWR VGND sg13g2_fill_2
XFILLER_43_703 VPWR VGND sg13g2_fill_1
XFILLER_42_202 VPWR VGND sg13g2_fill_1
XFILLER_24_961 VPWR VGND sg13g2_decap_8
XFILLER_23_460 VPWR VGND sg13g2_fill_1
XFILLER_3_832 VPWR VGND sg13g2_decap_8
XFILLER_18_1022 VPWR VGND sg13g2_decap_8
X_3700_ _0505_ _0503_ _0106_ VPWR VGND sg13g2_xor2_1
XFILLER_30_964 VPWR VGND sg13g2_decap_8
X_4680_ net864 net914 net867 _1443_ VPWR VGND net913 sg13g2_nand4_1
X_3631_ _0439_ net1035 net970 VPWR VGND sg13g2_nand2_1
X_3562_ _0360_ VPWR _0372_ VGND _0368_ _0370_ sg13g2_o21ai_1
X_6350_ net1133 VGND VPWR net155 mac1.sum_lvl1_ff\[82\] clknet_leaf_48_clk sg13g2_dfrbpq_1
X_5301_ VGND VPWR _2002_ _2013_ _2042_ _2001_ sg13g2_a21oi_1
X_3493_ _0293_ VPWR _0305_ VGND _0301_ _0303_ sg13g2_o21ai_1
X_6281_ net1109 VGND VPWR net127 mac1.sum_lvl2_ff\[5\] clknet_leaf_55_clk sg13g2_dfrbpq_1
X_5232_ _1975_ net871 net821 net874 net819 VPWR VGND sg13g2_a22oi_1
Xclkbuf_leaf_5_clk clknet_4_1_0_clk clknet_leaf_5_clk VPWR VGND sg13g2_buf_8
X_5163_ _1905_ _1906_ _1871_ _1908_ VPWR VGND sg13g2_nand3_1
X_4114_ VPWR _0904_ _0903_ VGND sg13g2_inv_1
X_5094_ _1840_ net883 net816 VPWR VGND sg13g2_nand2_1
X_4045_ _0837_ _0806_ _0835_ VPWR VGND sg13g2_xnor2_1
X_5996_ _2622_ VPWR _0246_ VGND net789 _2621_ sg13g2_o21ai_1
XFILLER_40_728 VPWR VGND sg13g2_fill_2
X_4947_ VPWR VGND _1648_ _1701_ _1679_ _1619_ _1702_ _1678_ sg13g2_a221oi_1
X_4878_ VGND VPWR _1636_ _1635_ _1590_ sg13g2_or2_1
XFILLER_20_430 VPWR VGND sg13g2_fill_2
XFILLER_21_964 VPWR VGND sg13g2_decap_8
XFILLER_32_1019 VPWR VGND sg13g2_decap_8
X_3829_ _0627_ net1022 net957 VPWR VGND sg13g2_nand2_1
X_6548_ net1076 VGND VPWR net1 DP_1.I_range.out_data\[2\] clknet_leaf_4_clk sg13g2_dfrbpq_2
X_6479_ net1079 VGND VPWR _0151_ mac2.products_ff\[147\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_0_868 VPWR VGND sg13g2_decap_8
XFILLER_12_920 VPWR VGND sg13g2_decap_8
XFILLER_8_913 VPWR VGND sg13g2_decap_8
XFILLER_11_441 VPWR VGND sg13g2_fill_1
XFILLER_12_997 VPWR VGND sg13g2_decap_8
XFILLER_11_485 VPWR VGND sg13g2_fill_1
XFILLER_48_1026 VPWR VGND sg13g2_fill_2
XFILLER_39_839 VPWR VGND sg13g2_fill_2
X_5850_ _2505_ _2489_ _2504_ VPWR VGND sg13g2_nand2_1
X_4801_ _1561_ net917 net856 VPWR VGND sg13g2_nand2_1
X_5781_ net1053 net784 _2437_ VPWR VGND sg13g2_nor2_1
X_4732_ _1491_ _1490_ _1460_ _1494_ VPWR VGND sg13g2_a21o_1
XFILLER_30_761 VPWR VGND sg13g2_fill_2
X_4663_ _1424_ _1398_ _1427_ VPWR VGND sg13g2_xor2_1
X_3614_ VGND VPWR _0419_ _0420_ _0423_ _0385_ sg13g2_a21oi_1
X_6402_ net1083 VGND VPWR net305 mac1.sum_lvl3_ff\[14\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_30_794 VPWR VGND sg13g2_fill_1
X_4594_ net869 net923 net863 net920 _1361_ VPWR VGND sg13g2_and4_1
X_3545_ _0355_ net1032 net972 VPWR VGND sg13g2_nand2_1
X_6333_ net1078 VGND VPWR net51 mac2.sum_lvl2_ff\[47\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_3476_ _0288_ net1040 DP_2.matrix\[5\] VPWR VGND sg13g2_nand2_1
X_6264_ net1092 VGND VPWR net72 mac1.sum_lvl1_ff\[40\] clknet_leaf_62_clk sg13g2_dfrbpq_1
X_5215_ _1947_ VPWR _1958_ VGND _1931_ _1948_ sg13g2_o21ai_1
X_6195_ net1109 VGND VPWR net86 mac1.sum_lvl1_ff\[5\] clknet_leaf_55_clk sg13g2_dfrbpq_1
Xclkbuf_4_15_0_clk clknet_0_clk clknet_4_15_0_clk VPWR VGND sg13g2_buf_8
X_5146_ _1891_ net822 net873 VPWR VGND sg13g2_nand2_1
X_5077_ _1822_ _1823_ _1805_ _1824_ VPWR VGND sg13g2_nand3_1
X_4028_ _0820_ net954 net1008 VPWR VGND sg13g2_nand2_1
XFILLER_38_872 VPWR VGND sg13g2_fill_1
XFILLER_44_37 VPWR VGND sg13g2_fill_2
X_5979_ _2612_ _2505_ _2509_ VPWR VGND sg13g2_xnor2_1
XFILLER_5_905 VPWR VGND sg13g2_decap_8
XFILLER_18_93 VPWR VGND sg13g2_fill_1
XFILLER_7_231 VPWR VGND sg13g2_fill_2
Xhold209 mac2.products_ff\[5\] VPWR VGND net249 sg13g2_dlygate4sd3_1
XFILLER_4_971 VPWR VGND sg13g2_decap_8
X_3330_ _2915_ _2912_ _2916_ VPWR VGND sg13g2_xor2_1
XFILLER_3_481 VPWR VGND sg13g2_fill_1
X_3261_ _2847_ _2848_ _2849_ VPWR VGND sg13g2_nor2_1
X_5000_ _1749_ _1739_ _1750_ VPWR VGND sg13g2_xor2_1
X_3192_ net1001 net998 net929 net926 _2781_ VPWR VGND sg13g2_and4_1
XFILLER_39_669 VPWR VGND sg13g2_fill_2
XFILLER_35_842 VPWR VGND sg13g2_fill_1
X_5902_ _2553_ VPWR _2556_ VGND net794 _2555_ sg13g2_o21ai_1
X_5833_ net806 net795 net882 _2488_ VPWR VGND sg13g2_nand3_1
X_5764_ _2416_ _2420_ _2421_ VPWR VGND sg13g2_and2_1
X_5695_ net18 _2356_ _2359_ VPWR VGND sg13g2_xnor2_1
X_4715_ net867 net864 net911 net909 _1477_ VPWR VGND sg13g2_and4_1
X_4646_ net868 net865 net916 net915 _1410_ VPWR VGND sg13g2_and4_1
X_4577_ _1334_ _1347_ _1348_ VPWR VGND sg13g2_nor2_1
X_6316_ net1111 VGND VPWR net243 mac1.sum_lvl2_ff\[46\] clknet_leaf_54_clk sg13g2_dfrbpq_1
X_3528_ VGND VPWR _0336_ _0337_ _0339_ _0319_ sg13g2_a21oi_1
X_3459_ _0272_ net1037 net976 VPWR VGND sg13g2_nand2_1
X_6247_ net1129 VGND VPWR _0255_ DP_4.matrix\[39\] clknet_leaf_45_clk sg13g2_dfrbpq_1
X_6178_ net1094 VGND VPWR net417 DP_2.matrix\[6\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_5129_ _1874_ net884 net811 VPWR VGND sg13g2_nand2_1
XFILLER_45_606 VPWR VGND sg13g2_fill_2
XFILLER_41_801 VPWR VGND sg13g2_fill_2
XFILLER_13_547 VPWR VGND sg13g2_fill_1
XFILLER_41_867 VPWR VGND sg13g2_decap_8
XFILLER_45_1007 VPWR VGND sg13g2_decap_8
XFILLER_1_963 VPWR VGND sg13g2_decap_8
XFILLER_0_473 VPWR VGND sg13g2_fill_2
XFILLER_49_945 VPWR VGND sg13g2_decap_8
Xhold70 mac2.products_ff\[80\] VPWR VGND net110 sg13g2_dlygate4sd3_1
Xhold92 mac2.sum_lvl1_ff\[49\] VPWR VGND net132 sg13g2_dlygate4sd3_1
Xhold81 mac2.products_ff\[145\] VPWR VGND net121 sg13g2_dlygate4sd3_1
XFILLER_45_80 VPWR VGND sg13g2_fill_2
XFILLER_17_897 VPWR VGND sg13g2_decap_8
X_5480_ _2192_ net525 net521 VPWR VGND sg13g2_nand2_1
X_4500_ _1242_ _1273_ _1240_ _1274_ VPWR VGND sg13g2_nand3_1
X_4431_ _1207_ _1177_ _1206_ VPWR VGND sg13g2_nand2_1
X_4362_ _1139_ _1092_ _1138_ VPWR VGND sg13g2_xnor2_1
X_3313_ _2872_ _2866_ _2874_ _2899_ VPWR VGND sg13g2_a21o_1
X_4293_ net844 net896 net848 _1072_ VPWR VGND net894 sg13g2_nand4_1
X_6101_ net1098 VGND VPWR _0109_ mac1.products_ff\[13\] clknet_leaf_29_clk sg13g2_dfrbpq_1
X_6032_ net994 _0192_ VPWR VGND sg13g2_buf_1
X_3244_ _2831_ _2780_ _2832_ VPWR VGND sg13g2_xor2_1
X_3175_ _2765_ _2745_ _2763_ _2764_ VPWR VGND sg13g2_and3_1
Xfanout1090 net1093 net1090 VPWR VGND sg13g2_buf_8
XFILLER_35_694 VPWR VGND sg13g2_fill_1
XFILLER_10_506 VPWR VGND sg13g2_decap_8
X_5816_ _2441_ _2442_ _2471_ _0163_ VPWR VGND sg13g2_mux2_1
X_5747_ net799 VPWR _2404_ VGND DP_1.matrix\[44\] net808 sg13g2_o21ai_1
X_5678_ VPWR VGND _2340_ _2339_ _2338_ mac1.total_sum\[5\] _2346_ mac2.total_sum\[5\]
+ sg13g2_a221oi_1
X_4629_ _1391_ _1390_ _1385_ _1394_ VPWR VGND sg13g2_a21o_1
XFILLER_46_904 VPWR VGND sg13g2_fill_2
XFILLER_46_959 VPWR VGND sg13g2_decap_8
XFILLER_25_160 VPWR VGND sg13g2_fill_1
XFILLER_26_683 VPWR VGND sg13g2_decap_4
XFILLER_14_867 VPWR VGND sg13g2_decap_8
XFILLER_41_653 VPWR VGND sg13g2_fill_1
XFILLER_9_326 VPWR VGND sg13g2_fill_2
XFILLER_15_94 VPWR VGND sg13g2_fill_1
XFILLER_0_270 VPWR VGND sg13g2_decap_8
XFILLER_49_786 VPWR VGND sg13g2_fill_1
X_4980_ _1730_ _1731_ _0090_ VPWR VGND sg13g2_nor2_1
X_3931_ _0707_ _0697_ _0705_ _0725_ VPWR VGND sg13g2_a21o_1
XFILLER_17_694 VPWR VGND sg13g2_decap_4
X_3862_ _0657_ _0637_ _0078_ VPWR VGND sg13g2_xor2_1
XFILLER_31_152 VPWR VGND sg13g2_fill_1
XFILLER_32_664 VPWR VGND sg13g2_fill_2
X_5601_ net359 mac2.sum_lvl3_ff\[25\] _2286_ VPWR VGND sg13g2_xor2_1
X_6581_ net1066 VGND VPWR net413 mac2.total_sum\[13\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_32_697 VPWR VGND sg13g2_fill_1
X_3793_ _0596_ net969 net1058 VPWR VGND sg13g2_nand2_1
X_5532_ _2232_ mac2.sum_lvl2_ff\[25\] mac2.sum_lvl2_ff\[6\] VPWR VGND sg13g2_xnor2_1
XFILLER_9_882 VPWR VGND sg13g2_decap_8
X_5463_ _2177_ net534 _0028_ VPWR VGND sg13g2_nor2b_2
X_5394_ net536 VPWR _2125_ VGND _2118_ _2121_ sg13g2_o21ai_1
X_4414_ _1190_ net899 DP_4.matrix\[41\] VPWR VGND sg13g2_nand2_1
X_4345_ _1120_ _1119_ _1089_ _1123_ VPWR VGND sg13g2_a21o_1
XFILLER_28_1002 VPWR VGND sg13g2_decap_8
X_4276_ _1053_ _1027_ _1056_ VPWR VGND sg13g2_xor2_1
X_3227_ _2743_ _2813_ _2815_ _2816_ VPWR VGND sg13g2_or3_1
X_6015_ net1051 _0165_ VPWR VGND sg13g2_buf_1
X_3158_ _2748_ net934 net995 VPWR VGND sg13g2_nand2_1
X_3089_ _2681_ net998 net933 VPWR VGND sg13g2_nand2_1
XFILLER_35_1006 VPWR VGND sg13g2_decap_8
XFILLER_11_826 VPWR VGND sg13g2_decap_8
XFILLER_22_174 VPWR VGND sg13g2_decap_4
XFILLER_2_513 VPWR VGND sg13g2_fill_1
Xhold381 _0224_ VPWR VGND net421 sg13g2_dlygate4sd3_1
Xhold370 mac2.sum_lvl3_ff\[13\] VPWR VGND net410 sg13g2_dlygate4sd3_1
Xhold392 mac2.sum_lvl2_ff\[3\] VPWR VGND net432 sg13g2_dlygate4sd3_1
Xfanout861 net379 net861 VPWR VGND sg13g2_buf_8
Xfanout850 net343 net850 VPWR VGND sg13g2_buf_8
Xfanout872 DP_3.matrix\[79\] net872 VPWR VGND sg13g2_buf_2
Xfanout883 net884 net883 VPWR VGND sg13g2_buf_8
Xfanout894 net895 net894 VPWR VGND sg13g2_buf_2
XFILLER_18_403 VPWR VGND sg13g2_fill_1
XFILLER_19_937 VPWR VGND sg13g2_decap_8
XFILLER_45_222 VPWR VGND sg13g2_fill_1
XFILLER_41_461 VPWR VGND sg13g2_fill_2
XFILLER_41_483 VPWR VGND sg13g2_fill_1
XFILLER_6_874 VPWR VGND sg13g2_decap_8
X_4130_ _0919_ net947 net1010 net949 net1008 VPWR VGND sg13g2_a22oi_1
XFILLER_49_550 VPWR VGND sg13g2_fill_2
X_4061_ _0851_ _0847_ _0852_ VPWR VGND sg13g2_xor2_1
XFILLER_37_767 VPWR VGND sg13g2_fill_1
XFILLER_24_406 VPWR VGND sg13g2_fill_1
XFILLER_37_789 VPWR VGND sg13g2_fill_1
X_4963_ _1716_ _1706_ _1718_ VPWR VGND sg13g2_xor2_1
XFILLER_36_299 VPWR VGND sg13g2_fill_1
X_3914_ _0707_ _0706_ _0697_ _0709_ VPWR VGND sg13g2_a21o_1
X_4894_ _1638_ _1633_ _1640_ _1651_ VPWR VGND sg13g2_a21o_1
XFILLER_33_995 VPWR VGND sg13g2_decap_8
X_3845_ VPWR _0642_ _0641_ VGND sg13g2_inv_1
X_3776_ _0554_ _0579_ _0580_ VPWR VGND sg13g2_nor2_1
X_6564_ net1082 VGND VPWR _0035_ mac2.sum_lvl3_ff\[12\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_5515_ _2216_ VPWR _2219_ VGND _2215_ _2217_ sg13g2_o21ai_1
X_6495_ net1142 VGND VPWR net84 mac2.sum_lvl1_ff\[11\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_5446_ VGND VPWR _2162_ _2164_ _2165_ _2163_ sg13g2_a21oi_1
X_5377_ net476 _2109_ _0009_ VPWR VGND sg13g2_xor2_1
X_4328_ net849 net844 net894 net891 _1106_ VPWR VGND sg13g2_and4_1
X_4259_ net849 net846 net898 net896 _1039_ VPWR VGND sg13g2_and4_1
XFILLER_41_1021 VPWR VGND sg13g2_decap_8
XFILLER_24_940 VPWR VGND sg13g2_decap_8
XFILLER_10_144 VPWR VGND sg13g2_fill_1
XFILLER_3_811 VPWR VGND sg13g2_decap_8
XFILLER_3_888 VPWR VGND sg13g2_decap_8
XFILLER_38_509 VPWR VGND sg13g2_decap_4
XFILLER_19_701 VPWR VGND sg13g2_fill_1
XFILLER_18_288 VPWR VGND sg13g2_fill_1
XFILLER_18_1001 VPWR VGND sg13g2_decap_8
XFILLER_14_461 VPWR VGND sg13g2_fill_2
XFILLER_15_995 VPWR VGND sg13g2_decap_8
XFILLER_30_932 VPWR VGND sg13g2_decap_4
X_3630_ _0438_ net1035 net967 VPWR VGND sg13g2_nand2_1
X_3561_ _0360_ _0368_ _0370_ _0371_ VPWR VGND sg13g2_or3_1
X_5300_ _2039_ _2027_ _2041_ VPWR VGND sg13g2_xor2_1
X_3492_ _0293_ _0301_ _0303_ _0304_ VPWR VGND sg13g2_or3_1
X_6280_ net1109 VGND VPWR net88 mac1.sum_lvl2_ff\[4\] clknet_leaf_55_clk sg13g2_dfrbpq_1
X_5231_ net821 net818 net874 net871 _1974_ VPWR VGND sg13g2_and4_1
XFILLER_45_2 VPWR VGND sg13g2_fill_1
X_5162_ _1907_ _1871_ _1905_ _1906_ VPWR VGND sg13g2_and3_1
X_5093_ _1821_ _1811_ _1819_ _1839_ VPWR VGND sg13g2_a21o_1
X_4113_ _0871_ _0902_ _0869_ _0903_ VPWR VGND sg13g2_nand3_1
X_4044_ _0836_ _0806_ _0835_ VPWR VGND sg13g2_nand2_1
X_5995_ _2622_ net861 net789 VPWR VGND sg13g2_nand2_1
XFILLER_24_258 VPWR VGND sg13g2_fill_1
X_4946_ _1701_ _1677_ _1699_ VPWR VGND sg13g2_nand2_1
X_4877_ _1635_ net914 net854 VPWR VGND sg13g2_nand2_1
XFILLER_21_943 VPWR VGND sg13g2_decap_8
X_3828_ VGND VPWR _0626_ _0621_ _0619_ sg13g2_or2_1
X_6547_ net1145 VGND VPWR net75 mac2.sum_lvl2_ff\[34\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_3759_ VGND VPWR _0501_ _0532_ _0564_ _0534_ sg13g2_a21oi_1
X_6478_ net1079 VGND VPWR _0150_ mac2.products_ff\[146\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_5429_ _2153_ mac1.sum_lvl2_ff\[33\] mac1.sum_lvl2_ff\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_0_847 VPWR VGND sg13g2_decap_8
XFILLER_43_512 VPWR VGND sg13g2_fill_1
XFILLER_16_748 VPWR VGND sg13g2_fill_1
XFILLER_28_586 VPWR VGND sg13g2_fill_1
XFILLER_12_976 VPWR VGND sg13g2_decap_8
XFILLER_8_969 VPWR VGND sg13g2_decap_8
XFILLER_48_1005 VPWR VGND sg13g2_decap_8
XFILLER_2_151 VPWR VGND sg13g2_fill_1
X_4800_ _1526_ VPWR _1560_ VGND _1517_ _1527_ sg13g2_o21ai_1
X_5780_ _2405_ _2406_ _2436_ _0160_ VPWR VGND sg13g2_mux2_1
X_4731_ VGND VPWR _1490_ _1491_ _1493_ _1460_ sg13g2_a21oi_1
X_4662_ VGND VPWR _1422_ _1423_ _1426_ _1398_ sg13g2_a21oi_1
X_3613_ _0419_ _0420_ _0385_ _0422_ VPWR VGND sg13g2_nand3_1
X_6401_ net1083 VGND VPWR net468 mac1.sum_lvl3_ff\[13\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_31_1020 VPWR VGND sg13g2_decap_8
X_4593_ _1360_ net924 net861 VPWR VGND sg13g2_nand2_1
X_3544_ _0354_ net1036 DP_2.matrix\[5\] VPWR VGND sg13g2_nand2_1
X_6332_ net1077 VGND VPWR net64 mac2.sum_lvl2_ff\[46\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_3475_ _0278_ VPWR _0287_ VGND _0270_ _0279_ sg13g2_o21ai_1
X_6263_ net1088 VGND VPWR net120 mac1.sum_lvl1_ff\[39\] clknet_leaf_64_clk sg13g2_dfrbpq_1
X_5214_ VGND VPWR _1922_ _1928_ _1957_ _1930_ sg13g2_a21oi_1
X_6194_ net1131 VGND VPWR _0213_ DP_2.matrix\[73\] clknet_leaf_53_clk sg13g2_dfrbpq_1
X_5145_ _1850_ VPWR _1890_ VGND _1848_ _1851_ sg13g2_o21ai_1
X_5076_ _1821_ _1820_ _1811_ _1823_ VPWR VGND sg13g2_a21o_1
X_4027_ _0819_ net1013 net951 VPWR VGND sg13g2_nand2_1
X_5978_ _2611_ net916 net793 VPWR VGND sg13g2_nand2_1
X_4929_ _1685_ net855 net908 VPWR VGND sg13g2_nand2_1
XFILLER_21_784 VPWR VGND sg13g2_fill_1
XFILLER_44_832 VPWR VGND sg13g2_decap_4
XFILLER_28_394 VPWR VGND sg13g2_fill_2
XFILLER_8_722 VPWR VGND sg13g2_fill_2
XFILLER_8_777 VPWR VGND sg13g2_fill_1
XFILLER_4_950 VPWR VGND sg13g2_decap_8
X_3260_ _2848_ net1055 net938 net987 net936 VPWR VGND sg13g2_a22oi_1
X_3191_ _2780_ net998 net926 VPWR VGND sg13g2_nand2_1
XFILLER_22_1008 VPWR VGND sg13g2_decap_8
XFILLER_39_637 VPWR VGND sg13g2_fill_2
X_5901_ _2554_ VPWR _2555_ VGND net857 net804 sg13g2_o21ai_1
XFILLER_35_832 VPWR VGND sg13g2_decap_4
X_5832_ VGND VPWR net918 net806 _2487_ _2486_ sg13g2_a21oi_1
X_5763_ VGND VPWR _2417_ _2418_ _2420_ _2419_ sg13g2_a21oi_1
X_4714_ _1476_ net861 net914 VPWR VGND sg13g2_nand2_1
X_5694_ _2359_ _2358_ _2357_ VPWR VGND sg13g2_nand2b_1
X_4645_ _1409_ net862 net919 VPWR VGND sg13g2_nand2_1
X_4576_ _1345_ _1335_ _1347_ VPWR VGND sg13g2_xor2_1
X_3527_ _0336_ _0337_ _0319_ _0338_ VPWR VGND sg13g2_nand3_1
X_6315_ net1132 VGND VPWR net244 mac1.sum_lvl2_ff\[45\] clknet_leaf_51_clk sg13g2_dfrbpq_1
X_3458_ _3021_ VPWR _0271_ VGND _3019_ _3022_ sg13g2_o21ai_1
X_6246_ net1120 VGND VPWR _0254_ DP_4.matrix\[38\] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_3389_ _2971_ _2946_ _2973_ VPWR VGND sg13g2_xor2_1
X_6177_ net1118 VGND VPWR _0100_ mac1.products_ff\[151\] clknet_leaf_47_clk sg13g2_dfrbpq_2
X_5128_ _1873_ net889 net1042 VPWR VGND sg13g2_nand2_1
X_5059_ _1806_ net886 net816 VPWR VGND sg13g2_nand2_1
XFILLER_38_670 VPWR VGND sg13g2_fill_1
XFILLER_25_331 VPWR VGND sg13g2_fill_1
XFILLER_25_375 VPWR VGND sg13g2_fill_2
XFILLER_26_898 VPWR VGND sg13g2_decap_4
XFILLER_9_508 VPWR VGND sg13g2_fill_2
XFILLER_5_769 VPWR VGND sg13g2_fill_2
XFILLER_1_942 VPWR VGND sg13g2_decap_8
XFILLER_49_924 VPWR VGND sg13g2_decap_8
XFILLER_0_452 VPWR VGND sg13g2_decap_8
XFILLER_29_71 VPWR VGND sg13g2_fill_1
Xhold71 mac2.sum_lvl1_ff\[47\] VPWR VGND net111 sg13g2_dlygate4sd3_1
Xhold82 mac2.sum_lvl1_ff\[37\] VPWR VGND net122 sg13g2_dlygate4sd3_1
Xhold60 mac2.sum_lvl1_ff\[0\] VPWR VGND net100 sg13g2_dlygate4sd3_1
Xhold93 mac2.products_ff\[4\] VPWR VGND net133 sg13g2_dlygate4sd3_1
XFILLER_17_876 VPWR VGND sg13g2_decap_8
XFILLER_32_835 VPWR VGND sg13g2_fill_1
Xclkbuf_4_14_0_clk clknet_0_clk clknet_4_14_0_clk VPWR VGND sg13g2_buf_8
XFILLER_12_592 VPWR VGND sg13g2_fill_2
X_4430_ _1205_ _1188_ _1206_ VPWR VGND sg13g2_xor2_1
X_4361_ _1138_ _1129_ _1136_ VPWR VGND sg13g2_xnor2_1
X_6100_ net1098 VGND VPWR _0108_ mac1.products_ff\[12\] clknet_leaf_29_clk sg13g2_dfrbpq_1
X_3312_ _2897_ _2895_ _0095_ VPWR VGND sg13g2_xor2_1
X_4292_ net848 net844 net896 net894 _1071_ VPWR VGND sg13g2_and4_1
X_6031_ net997 _0191_ VPWR VGND sg13g2_buf_1
X_3243_ _2831_ net996 net928 VPWR VGND sg13g2_nand2_1
X_3174_ _2752_ VPWR _2764_ VGND _2760_ _2762_ sg13g2_o21ai_1
Xfanout1091 net1093 net1091 VPWR VGND sg13g2_buf_8
XFILLER_13_0 VPWR VGND sg13g2_fill_1
Xfanout1080 net1086 net1080 VPWR VGND sg13g2_buf_8
XFILLER_27_629 VPWR VGND sg13g2_fill_1
X_5815_ net784 VPWR _2471_ VGND _2468_ _2470_ sg13g2_o21ai_1
X_5746_ net1059 net810 _2403_ VPWR VGND sg13g2_nor2_1
X_5677_ _2345_ mac1.total_sum\[6\] mac2.total_sum\[6\] VPWR VGND sg13g2_xnor2_1
X_4628_ VGND VPWR _1390_ _1391_ _1393_ _1385_ sg13g2_a21oi_1
X_4559_ _1305_ _1328_ _1330_ VPWR VGND sg13g2_and2_1
X_6229_ net1104 VGND VPWR _0237_ DP_3.matrix\[73\] clknet_leaf_26_clk sg13g2_dfrbpq_1
Xheichips25_template_40 VPWR VGND uio_oe[7] sg13g2_tiehi
XFILLER_45_448 VPWR VGND sg13g2_fill_1
XFILLER_14_846 VPWR VGND sg13g2_decap_8
XFILLER_9_349 VPWR VGND sg13g2_fill_1
XFILLER_12_1018 VPWR VGND sg13g2_decap_8
XFILLER_37_905 VPWR VGND sg13g2_fill_2
X_3930_ _0724_ _0719_ _0722_ VPWR VGND sg13g2_xnor2_1
XFILLER_45_993 VPWR VGND sg13g2_decap_8
X_3861_ VGND VPWR _0658_ _0657_ _0637_ sg13g2_or2_1
XFILLER_16_194 VPWR VGND sg13g2_fill_1
XFILLER_20_816 VPWR VGND sg13g2_fill_2
XFILLER_32_676 VPWR VGND sg13g2_decap_4
X_3792_ _0595_ net966 net1058 VPWR VGND sg13g2_nand2_1
X_6580_ net1066 VGND VPWR _0051_ mac2.total_sum\[12\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_5600_ mac2.sum_lvl3_ff\[25\] net359 _2285_ VPWR VGND sg13g2_nor2_1
XFILLER_9_861 VPWR VGND sg13g2_decap_8
X_5531_ mac2.sum_lvl2_ff\[25\] mac2.sum_lvl2_ff\[6\] _2231_ VPWR VGND sg13g2_and2_1
X_5462_ net533 VPWR _2178_ VGND _2172_ _2176_ sg13g2_o21ai_1
X_5393_ net535 mac1.sum_lvl2_ff\[26\] _2124_ VPWR VGND sg13g2_xor2_1
X_4413_ _1155_ VPWR _1189_ VGND _1146_ _1156_ sg13g2_o21ai_1
X_4344_ VGND VPWR _1119_ _1120_ _1122_ _1089_ sg13g2_a21oi_1
X_6014_ net274 _0164_ VPWR VGND sg13g2_buf_1
X_4275_ VGND VPWR _1051_ _1052_ _1055_ _1027_ sg13g2_a21oi_1
X_3226_ VGND VPWR _2811_ _2812_ _2815_ _2777_ sg13g2_a21oi_1
X_3157_ _2747_ net995 net933 VPWR VGND sg13g2_nand2_1
XFILLER_27_404 VPWR VGND sg13g2_fill_1
XFILLER_27_459 VPWR VGND sg13g2_decap_8
X_3088_ _2680_ net1003 net930 VPWR VGND sg13g2_nand2_1
XFILLER_23_698 VPWR VGND sg13g2_decap_4
XFILLER_10_337 VPWR VGND sg13g2_fill_1
X_5729_ _2386_ DP_1.I_range.out_data\[2\] DP_1.Q_range.out_data\[2\] VPWR VGND sg13g2_nand2_1
Xhold360 DP_2.matrix\[41\] VPWR VGND net400 sg13g2_dlygate4sd3_1
Xhold371 _2319_ VPWR VGND net411 sg13g2_dlygate4sd3_1
Xhold393 _2224_ VPWR VGND net433 sg13g2_dlygate4sd3_1
Xhold382 DP_3.matrix\[1\] VPWR VGND net422 sg13g2_dlygate4sd3_1
Xfanout851 net853 net851 VPWR VGND sg13g2_buf_8
Xfanout840 net398 net840 VPWR VGND sg13g2_buf_8
Xfanout873 net874 net873 VPWR VGND sg13g2_buf_8
Xfanout862 DP_4.matrix\[2\] net862 VPWR VGND sg13g2_buf_1
Xfanout884 net885 net884 VPWR VGND sg13g2_buf_1
XFILLER_19_916 VPWR VGND sg13g2_decap_8
Xfanout895 net539 net895 VPWR VGND sg13g2_buf_8
XFILLER_27_993 VPWR VGND sg13g2_decap_8
XFILLER_41_495 VPWR VGND sg13g2_fill_2
XFILLER_10_882 VPWR VGND sg13g2_decap_8
XFILLER_6_853 VPWR VGND sg13g2_decap_8
XFILLER_5_352 VPWR VGND sg13g2_fill_1
X_4060_ _0851_ _0810_ _0849_ VPWR VGND sg13g2_xnor2_1
XFILLER_49_562 VPWR VGND sg13g2_fill_2
XFILLER_25_919 VPWR VGND sg13g2_decap_8
X_4962_ _1716_ _1706_ _1717_ VPWR VGND sg13g2_nor2b_1
X_3913_ _0706_ _0707_ _0697_ _0708_ VPWR VGND sg13g2_nand3_1
XFILLER_33_974 VPWR VGND sg13g2_decap_8
X_4893_ _1650_ _1649_ _0140_ VPWR VGND sg13g2_xor2_1
X_3844_ _0638_ _0640_ _0641_ VPWR VGND sg13g2_nor2_1
X_6563_ net1077 VGND VPWR _0034_ mac2.sum_lvl3_ff\[11\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_3775_ _0579_ _0539_ _0577_ VPWR VGND sg13g2_xnor2_1
XFILLER_9_691 VPWR VGND sg13g2_fill_1
X_5514_ _0039_ _2215_ _2218_ VPWR VGND sg13g2_xnor2_1
X_6494_ net1142 VGND VPWR net80 mac2.sum_lvl1_ff\[10\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_5445_ net382 _2162_ _0024_ VPWR VGND sg13g2_xor2_1
X_5376_ _2111_ mac1.sum_lvl2_ff\[22\] net475 VPWR VGND sg13g2_xnor2_1
X_4327_ _1105_ net842 net896 VPWR VGND sg13g2_nand2_1
X_4258_ _1038_ net843 net901 VPWR VGND sg13g2_nand2_1
XFILLER_41_1000 VPWR VGND sg13g2_decap_8
X_3209_ net944 net939 net986 net1054 _2798_ VPWR VGND sg13g2_and4_1
X_4189_ _0974_ _0964_ _0976_ VPWR VGND sg13g2_xor2_1
XFILLER_28_735 VPWR VGND sg13g2_decap_4
XFILLER_28_779 VPWR VGND sg13g2_fill_1
XFILLER_42_237 VPWR VGND sg13g2_fill_1
XFILLER_23_451 VPWR VGND sg13g2_decap_8
XFILLER_24_996 VPWR VGND sg13g2_decap_8
XFILLER_11_657 VPWR VGND sg13g2_fill_2
XFILLER_3_867 VPWR VGND sg13g2_decap_8
Xhold190 mac1.products_ff\[80\] VPWR VGND net230 sg13g2_dlygate4sd3_1
XFILLER_46_576 VPWR VGND sg13g2_fill_1
XFILLER_15_974 VPWR VGND sg13g2_decap_8
XFILLER_14_484 VPWR VGND sg13g2_fill_2
XFILLER_30_999 VPWR VGND sg13g2_decap_8
X_3560_ VGND VPWR _0366_ _0367_ _0370_ _0361_ sg13g2_a21oi_1
X_5230_ _1973_ net819 net871 VPWR VGND sg13g2_nand2_1
X_3491_ VGND VPWR _0299_ _0300_ _0303_ _0294_ sg13g2_a21oi_1
X_5161_ _1882_ VPWR _1906_ VGND _1902_ _1904_ sg13g2_o21ai_1
X_5092_ _1838_ _1833_ _1836_ VPWR VGND sg13g2_xnor2_1
X_4112_ _0900_ _0879_ _0902_ VPWR VGND sg13g2_xor2_1
XFILLER_25_1017 VPWR VGND sg13g2_decap_8
XFILLER_25_1028 VPWR VGND sg13g2_fill_1
X_4043_ _0834_ _0817_ _0835_ VPWR VGND sg13g2_xor2_1
X_5994_ _2550_ _2546_ _2621_ VPWR VGND sg13g2_xor2_1
XFILLER_25_738 VPWR VGND sg13g2_decap_8
X_4945_ _0142_ _1699_ _1700_ VPWR VGND sg13g2_xnor2_1
XFILLER_21_922 VPWR VGND sg13g2_decap_8
X_4876_ _1634_ net919 net1044 VPWR VGND sg13g2_nand2_1
X_3827_ _0625_ net1023 net954 VPWR VGND sg13g2_nand2_1
XFILLER_21_999 VPWR VGND sg13g2_decap_8
X_3758_ _0561_ _0560_ _0563_ VPWR VGND sg13g2_xor2_1
X_6546_ net1142 VGND VPWR net141 mac2.sum_lvl2_ff\[33\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_3689_ _0495_ _0483_ _0496_ VPWR VGND sg13g2_xor2_1
X_6477_ net1075 VGND VPWR _0159_ mac2.products_ff\[145\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_5428_ VGND VPWR _2148_ _2150_ _2152_ _2149_ sg13g2_a21oi_1
X_5359_ _2097_ net872 net1042 VPWR VGND sg13g2_nand2_1
XFILLER_0_826 VPWR VGND sg13g2_decap_8
XFILLER_28_532 VPWR VGND sg13g2_fill_1
XFILLER_15_226 VPWR VGND sg13g2_fill_2
XFILLER_12_955 VPWR VGND sg13g2_decap_8
XFILLER_30_229 VPWR VGND sg13g2_fill_1
XFILLER_8_948 VPWR VGND sg13g2_decap_8
XFILLER_48_1028 VPWR VGND sg13g2_fill_1
XFILLER_48_92 VPWR VGND sg13g2_fill_2
XFILLER_0_1008 VPWR VGND sg13g2_decap_8
X_4730_ _1490_ _1491_ _1460_ _1492_ VPWR VGND sg13g2_nand3_1
X_4661_ _1422_ _1423_ _1398_ _1425_ VPWR VGND sg13g2_nand3_1
X_3612_ _0421_ _0385_ _0419_ _0420_ VPWR VGND sg13g2_and3_1
X_6400_ net1083 VGND VPWR net321 mac1.sum_lvl3_ff\[12\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_6331_ net1078 VGND VPWR net93 mac2.sum_lvl2_ff\[45\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_4592_ _1358_ _1359_ _0085_ VPWR VGND sg13g2_nor2_1
X_3543_ _0335_ _0325_ _0333_ _0353_ VPWR VGND sg13g2_a21o_1
X_3474_ _0285_ _3029_ _0073_ VPWR VGND sg13g2_xor2_1
X_6262_ net1069 VGND VPWR net54 mac1.sum_lvl1_ff\[38\] clknet_leaf_67_clk sg13g2_dfrbpq_1
X_6193_ net1131 VGND VPWR _0212_ DP_2.matrix\[72\] clknet_leaf_53_clk sg13g2_dfrbpq_1
XFILLER_9_1022 VPWR VGND sg13g2_decap_8
X_5213_ _1956_ _1917_ _0159_ VPWR VGND sg13g2_xor2_1
X_5144_ _1889_ _1884_ _1888_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_18 VPWR VGND sg13g2_fill_2
XFILLER_29_307 VPWR VGND sg13g2_fill_2
X_5075_ _1820_ _1821_ _1811_ _1822_ VPWR VGND sg13g2_nand3_1
XFILLER_38_830 VPWR VGND sg13g2_decap_4
X_4026_ _0784_ VPWR _0818_ VGND _0775_ _0785_ sg13g2_o21ai_1
X_5977_ _2610_ VPWR _0223_ VGND net790 _2609_ sg13g2_o21ai_1
XFILLER_40_505 VPWR VGND sg13g2_fill_2
X_4928_ _1684_ net909 net851 VPWR VGND sg13g2_nand2_1
XFILLER_21_741 VPWR VGND sg13g2_decap_8
XFILLER_21_752 VPWR VGND sg13g2_fill_2
X_4859_ VGND VPWR _1541_ _1583_ _1618_ _1582_ sg13g2_a21oi_1
X_6529_ net1144 VGND VPWR net250 mac2.sum_lvl2_ff\[13\] clknet_leaf_41_clk sg13g2_dfrbpq_1
XFILLER_0_612 VPWR VGND sg13g2_fill_1
XFILLER_28_384 VPWR VGND sg13g2_fill_2
XFILLER_8_701 VPWR VGND sg13g2_fill_1
XFILLER_15_1016 VPWR VGND sg13g2_decap_8
XFILLER_15_1027 VPWR VGND sg13g2_fill_2
XFILLER_34_94 VPWR VGND sg13g2_fill_1
XFILLER_7_233 VPWR VGND sg13g2_fill_1
XFILLER_3_450 VPWR VGND sg13g2_fill_2
X_3190_ _2779_ net1004 net1051 VPWR VGND sg13g2_nand2_1
XFILLER_39_605 VPWR VGND sg13g2_fill_1
X_5900_ _2554_ net803 net838 VPWR VGND sg13g2_nand2b_1
XFILLER_34_343 VPWR VGND sg13g2_fill_2
XFILLER_35_855 VPWR VGND sg13g2_decap_8
XFILLER_34_376 VPWR VGND sg13g2_fill_1
X_5831_ net900 net805 _2486_ VPWR VGND sg13g2_and2_1
X_5762_ net1038 _2417_ _2419_ VPWR VGND sg13g2_nor2_1
X_4713_ _1443_ VPWR _1475_ VGND _1441_ _1444_ sg13g2_o21ai_1
X_5693_ VGND VPWR _2358_ mac2.total_sum\[9\] mac1.total_sum\[9\] sg13g2_or2_1
X_4644_ _1388_ VPWR _1408_ VGND _1386_ _1389_ sg13g2_o21ai_1
X_4575_ _1345_ _1335_ _1346_ VPWR VGND sg13g2_nor2b_1
X_6314_ net1131 VGND VPWR net159 mac1.sum_lvl2_ff\[44\] clknet_leaf_52_clk sg13g2_dfrbpq_1
X_3526_ _0335_ _0334_ _0325_ _0337_ VPWR VGND sg13g2_a21o_1
X_6245_ net1105 VGND VPWR _0253_ DP_4.matrix\[37\] clknet_leaf_32_clk sg13g2_dfrbpq_2
X_3457_ VPWR _0270_ _0269_ VGND sg13g2_inv_1
X_6176_ net1089 VGND VPWR _0201_ DP_2.matrix\[5\] clknet_leaf_61_clk sg13g2_dfrbpq_2
X_3388_ _2946_ _2971_ _2972_ VPWR VGND sg13g2_nor2_1
X_5127_ _1843_ VPWR _1872_ VGND _1840_ _1844_ sg13g2_o21ai_1
XFILLER_45_608 VPWR VGND sg13g2_fill_1
X_5058_ _1788_ VPWR _1805_ VGND _1779_ _1789_ sg13g2_o21ai_1
X_4009_ _0754_ _0755_ _0799_ _0800_ _0802_ VPWR VGND sg13g2_and4_1
Xclkbuf_leaf_64_clk clknet_4_2_0_clk clknet_leaf_64_clk VPWR VGND sg13g2_buf_8
XFILLER_38_1016 VPWR VGND sg13g2_decap_8
XFILLER_38_1027 VPWR VGND sg13g2_fill_2
XFILLER_41_803 VPWR VGND sg13g2_fill_1
XFILLER_1_921 VPWR VGND sg13g2_decap_8
XFILLER_20_63 VPWR VGND sg13g2_fill_2
XFILLER_49_903 VPWR VGND sg13g2_decap_8
Xhold50 mac1.products_ff\[143\] VPWR VGND net90 sg13g2_dlygate4sd3_1
XFILLER_1_998 VPWR VGND sg13g2_decap_8
XFILLER_21_1020 VPWR VGND sg13g2_decap_8
Xhold61 mac2.sum_lvl2_ff\[48\] VPWR VGND net101 sg13g2_dlygate4sd3_1
Xhold72 mac2.sum_lvl1_ff\[77\] VPWR VGND net112 sg13g2_dlygate4sd3_1
Xhold83 mac2.sum_lvl2_ff\[39\] VPWR VGND net123 sg13g2_dlygate4sd3_1
XFILLER_17_811 VPWR VGND sg13g2_decap_8
Xhold94 mac1.products_ff\[11\] VPWR VGND net134 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_55_clk clknet_4_8_0_clk clknet_leaf_55_clk VPWR VGND sg13g2_buf_8
XFILLER_16_332 VPWR VGND sg13g2_fill_2
XFILLER_17_855 VPWR VGND sg13g2_decap_8
XFILLER_31_357 VPWR VGND sg13g2_fill_2
XFILLER_12_582 VPWR VGND sg13g2_fill_1
XFILLER_6_76 VPWR VGND sg13g2_fill_2
X_4360_ _1137_ _1129_ _1136_ VPWR VGND sg13g2_nand2_1
XFILLER_6_87 VPWR VGND sg13g2_fill_2
X_3311_ _2895_ _2897_ _2898_ VPWR VGND sg13g2_nor2_1
X_4291_ _1070_ net843 net898 VPWR VGND sg13g2_nand2_1
X_6030_ net998 _0190_ VPWR VGND sg13g2_buf_1
X_3242_ _2830_ net996 net927 VPWR VGND sg13g2_nand2_1
X_3173_ _2752_ _2760_ _2762_ _2763_ VPWR VGND sg13g2_or3_1
XFILLER_6_1014 VPWR VGND sg13g2_decap_8
Xfanout1092 net1093 net1092 VPWR VGND sg13g2_buf_8
Xfanout1070 net1072 net1070 VPWR VGND sg13g2_buf_8
Xfanout1081 net1082 net1081 VPWR VGND sg13g2_buf_8
XFILLER_48_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_46_clk clknet_4_9_0_clk clknet_leaf_46_clk VPWR VGND sg13g2_buf_8
XFILLER_35_630 VPWR VGND sg13g2_fill_1
X_5814_ _2470_ net800 _2469_ net802 DP_2.matrix\[79\] VPWR VGND sg13g2_a22oi_1
X_5745_ _2402_ _2395_ _2400_ VPWR VGND sg13g2_xnor2_1
X_5676_ mac1.total_sum\[6\] mac2.total_sum\[6\] _2344_ VPWR VGND sg13g2_and2_1
X_4627_ _1390_ _1391_ _1385_ _1392_ VPWR VGND sg13g2_nand3_1
X_4558_ _0131_ _1328_ _1329_ VPWR VGND sg13g2_xnor2_1
X_3509_ _0320_ net1039 DP_2.matrix\[5\] VPWR VGND sg13g2_nand2_1
X_4489_ VGND VPWR _1263_ _1262_ _1219_ sg13g2_or2_1
XFILLER_44_1020 VPWR VGND sg13g2_decap_8
X_6228_ net1100 VGND VPWR _0236_ DP_3.matrix\[72\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_6159_ net1132 VGND VPWR _0104_ mac1.products_ff\[145\] clknet_leaf_51_clk sg13g2_dfrbpq_1
XFILLER_46_906 VPWR VGND sg13g2_fill_1
XFILLER_17_107 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_37_clk clknet_4_13_0_clk clknet_leaf_37_clk VPWR VGND sg13g2_buf_8
XFILLER_26_652 VPWR VGND sg13g2_decap_4
XFILLER_22_880 VPWR VGND sg13g2_fill_2
XFILLER_31_73 VPWR VGND sg13g2_fill_2
XFILLER_49_711 VPWR VGND sg13g2_fill_1
XFILLER_1_795 VPWR VGND sg13g2_decap_8
XFILLER_49_799 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_28_clk clknet_4_7_0_clk clknet_leaf_28_clk VPWR VGND sg13g2_buf_8
XFILLER_45_972 VPWR VGND sg13g2_decap_8
X_3860_ _0655_ _0654_ _0657_ VPWR VGND sg13g2_xor2_1
XFILLER_32_666 VPWR VGND sg13g2_fill_1
X_3791_ _0594_ net1027 DP_2.matrix\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_13_891 VPWR VGND sg13g2_decap_8
X_5530_ _0043_ _2228_ net470 VPWR VGND sg13g2_xnor2_1
X_5461_ _2172_ _2175_ _2176_ _2177_ VPWR VGND sg13g2_nor3_1
X_4412_ _1188_ _1178_ _1186_ VPWR VGND sg13g2_xnor2_1
X_5392_ _2123_ mac1.sum_lvl2_ff\[26\] mac1.sum_lvl2_ff\[7\] VPWR VGND sg13g2_nand2_1
X_4343_ _1119_ _1120_ _1089_ _1121_ VPWR VGND sg13g2_nand3_1
X_4274_ _1051_ _1052_ _1027_ _1054_ VPWR VGND sg13g2_nand3_1
X_3225_ _2811_ _2812_ _2777_ _2814_ VPWR VGND sg13g2_nand3_1
X_6013_ net1054 _0162_ VPWR VGND sg13g2_buf_1
XFILLER_39_243 VPWR VGND sg13g2_fill_2
X_3156_ _2746_ net998 net930 VPWR VGND sg13g2_nand2_1
X_3087_ _2670_ VPWR _2679_ VGND _2662_ _2671_ sg13g2_o21ai_1
Xclkbuf_leaf_19_clk clknet_4_4_0_clk clknet_leaf_19_clk VPWR VGND sg13g2_buf_8
XFILLER_23_622 VPWR VGND sg13g2_decap_4
XFILLER_36_994 VPWR VGND sg13g2_decap_8
X_3989_ _0777_ VPWR _0782_ VGND _0778_ _0780_ sg13g2_o21ai_1
X_5728_ _2384_ VPWR _2385_ VGND DP_1.I_range.out_data\[3\] DP_1.Q_range.out_data\[5\]
+ sg13g2_o21ai_1
X_5659_ net26 _2328_ _2331_ VPWR VGND sg13g2_xnor2_1
Xhold350 _2108_ VPWR VGND net390 sg13g2_dlygate4sd3_1
Xhold361 mac2.sum_lvl3_ff\[30\] VPWR VGND net401 sg13g2_dlygate4sd3_1
Xhold372 _2320_ VPWR VGND net412 sg13g2_dlygate4sd3_1
Xhold394 _0041_ VPWR VGND net434 sg13g2_dlygate4sd3_1
Xhold383 _0221_ VPWR VGND net423 sg13g2_dlygate4sd3_1
Xfanout852 net853 net852 VPWR VGND sg13g2_buf_1
Xfanout841 net398 net841 VPWR VGND sg13g2_buf_1
Xfanout830 net831 net830 VPWR VGND sg13g2_buf_1
Xfanout874 DP_3.matrix\[78\] net874 VPWR VGND sg13g2_buf_8
Xfanout885 net307 net885 VPWR VGND sg13g2_buf_2
Xclkbuf_4_13_0_clk clknet_0_clk clknet_4_13_0_clk VPWR VGND sg13g2_buf_8
Xfanout863 net866 net863 VPWR VGND sg13g2_buf_8
XFILLER_45_202 VPWR VGND sg13g2_fill_2
Xfanout896 DP_3.matrix\[41\] net896 VPWR VGND sg13g2_buf_8
XFILLER_18_438 VPWR VGND sg13g2_decap_8
XFILLER_27_972 VPWR VGND sg13g2_decap_8
XFILLER_13_132 VPWR VGND sg13g2_fill_1
XFILLER_42_997 VPWR VGND sg13g2_decap_8
XFILLER_10_861 VPWR VGND sg13g2_decap_8
XFILLER_9_169 VPWR VGND sg13g2_fill_2
XFILLER_6_832 VPWR VGND sg13g2_decap_8
XFILLER_3_1028 VPWR VGND sg13g2_fill_1
XFILLER_36_213 VPWR VGND sg13g2_fill_1
X_4961_ _1716_ _1692_ _1715_ VPWR VGND sg13g2_xnor2_1
XFILLER_18_994 VPWR VGND sg13g2_decap_8
X_3912_ _0704_ _0703_ _0698_ _0707_ VPWR VGND sg13g2_a21o_1
X_4892_ _1615_ _1620_ _1650_ VPWR VGND sg13g2_nor2_1
X_3843_ net1024 DP_1.matrix\[37\] net955 net953 _0640_ VPWR VGND sg13g2_and4_1
X_6562_ net1067 VGND VPWR _0033_ mac2.sum_lvl3_ff\[10\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_3774_ _0539_ _0577_ _0578_ VPWR VGND sg13g2_nor2_1
X_5513_ mac2.sum_lvl2_ff\[1\] mac2.sum_lvl2_ff\[20\] _2218_ VPWR VGND sg13g2_xor2_1
X_6493_ net1140 VGND VPWR net83 mac2.sum_lvl1_ff\[9\] clknet_leaf_40_clk sg13g2_dfrbpq_1
X_5444_ net381 mac1.sum_lvl3_ff\[22\] _2164_ VPWR VGND sg13g2_xor2_1
Xclkbuf_leaf_8_clk clknet_4_3_0_clk clknet_leaf_8_clk VPWR VGND sg13g2_buf_8
X_5375_ _2110_ mac1.sum_lvl2_ff\[22\] mac1.sum_lvl2_ff\[3\] VPWR VGND sg13g2_nand2_1
X_4326_ _1072_ VPWR _1104_ VGND _1070_ _1073_ sg13g2_o21ai_1
X_4257_ _1017_ VPWR _1037_ VGND _1015_ _1018_ sg13g2_o21ai_1
X_3208_ _2797_ net936 net989 VPWR VGND sg13g2_nand2_1
X_4188_ _0974_ _0964_ _0975_ VPWR VGND sg13g2_nor2b_1
X_3139_ _2728_ _2729_ _2711_ _2730_ VPWR VGND sg13g2_nand3_1
XFILLER_28_758 VPWR VGND sg13g2_fill_2
XFILLER_24_975 VPWR VGND sg13g2_decap_8
XFILLER_3_846 VPWR VGND sg13g2_decap_8
Xhold180 mac2.products_ff\[1\] VPWR VGND net220 sg13g2_dlygate4sd3_1
Xhold191 mac2.sum_lvl1_ff\[41\] VPWR VGND net231 sg13g2_dlygate4sd3_1
XFILLER_46_500 VPWR VGND sg13g2_fill_1
XFILLER_19_714 VPWR VGND sg13g2_fill_1
XFILLER_19_725 VPWR VGND sg13g2_decap_4
XFILLER_15_953 VPWR VGND sg13g2_decap_8
XFILLER_30_901 VPWR VGND sg13g2_fill_1
XFILLER_30_978 VPWR VGND sg13g2_decap_8
X_3490_ _0299_ _0300_ _0294_ _0302_ VPWR VGND sg13g2_nand3_1
X_5160_ _1882_ _1902_ _1904_ _1905_ VPWR VGND sg13g2_or3_1
X_4111_ _0900_ _0879_ _0901_ VPWR VGND sg13g2_nor2b_1
X_5091_ _1837_ _1833_ _1836_ VPWR VGND sg13g2_nand2_1
X_4042_ _0834_ _0818_ _0832_ VPWR VGND sg13g2_xnor2_1
X_5993_ _2620_ VPWR _0245_ VGND net789 _2619_ sg13g2_o21ai_1
XFILLER_37_577 VPWR VGND sg13g2_fill_2
X_4944_ VGND VPWR _1677_ _1680_ _1700_ _1676_ sg13g2_a21oi_1
XFILLER_21_901 VPWR VGND sg13g2_decap_8
X_4875_ VGND VPWR _1633_ _1604_ _1602_ sg13g2_or2_1
X_3826_ _0623_ _0616_ _0076_ VPWR VGND sg13g2_xor2_1
XFILLER_21_978 VPWR VGND sg13g2_decap_8
X_3757_ _0560_ _0561_ _0562_ VPWR VGND sg13g2_nor2_1
X_6545_ net1142 VGND VPWR net132 mac2.sum_lvl2_ff\[32\] clknet_leaf_41_clk sg13g2_dfrbpq_1
X_3688_ _0493_ _0484_ _0495_ VPWR VGND sg13g2_xor2_1
X_6476_ net1075 VGND VPWR _0158_ mac2.products_ff\[144\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_0_805 VPWR VGND sg13g2_decap_8
X_5427_ _0004_ _2148_ net467 VPWR VGND sg13g2_xnor2_1
X_5358_ _2084_ VPWR _2096_ VGND _2056_ _2082_ sg13g2_o21ai_1
X_4309_ _1054_ VPWR _1088_ VGND _1029_ _1055_ sg13g2_o21ai_1
X_5289_ _2030_ net879 net1042 VPWR VGND sg13g2_nand2_1
XFILLER_28_555 VPWR VGND sg13g2_fill_1
XFILLER_12_934 VPWR VGND sg13g2_decap_8
XFILLER_8_927 VPWR VGND sg13g2_decap_8
XFILLER_23_41 VPWR VGND sg13g2_fill_2
XFILLER_11_477 VPWR VGND sg13g2_fill_1
XFILLER_3_0 VPWR VGND sg13g2_fill_1
XFILLER_39_809 VPWR VGND sg13g2_decap_4
XFILLER_46_374 VPWR VGND sg13g2_fill_1
X_4660_ _1422_ _1423_ _1424_ VPWR VGND sg13g2_and2_1
X_3611_ _0396_ VPWR _0420_ VGND _0416_ _0418_ sg13g2_o21ai_1
X_6330_ net1081 VGND VPWR net47 mac2.sum_lvl2_ff\[44\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_4591_ _1359_ net863 net924 net923 net869 VPWR VGND sg13g2_a22oi_1
XFILLER_7_982 VPWR VGND sg13g2_decap_8
X_3542_ _0352_ _0347_ _0350_ VPWR VGND sg13g2_xnor2_1
X_6261_ net1063 VGND VPWR net217 mac1.sum_lvl1_ff\[37\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3473_ VGND VPWR _0286_ _0285_ _3029_ sg13g2_or2_1
X_5212_ _1954_ _1955_ _1956_ VPWR VGND sg13g2_nor2b_2
X_6192_ net1109 VGND VPWR net183 mac1.sum_lvl1_ff\[4\] clknet_leaf_55_clk sg13g2_dfrbpq_1
XFILLER_9_1001 VPWR VGND sg13g2_decap_8
X_5143_ _1888_ _1841_ _1886_ VPWR VGND sg13g2_xnor2_1
X_5074_ _1818_ _1817_ _1812_ _1821_ VPWR VGND sg13g2_a21o_1
X_4025_ _0817_ _0807_ _0815_ VPWR VGND sg13g2_xnor2_1
XFILLER_37_385 VPWR VGND sg13g2_fill_2
XFILLER_13_709 VPWR VGND sg13g2_decap_8
X_5976_ _2610_ net918 net790 VPWR VGND sg13g2_nand2_1
X_4927_ _1683_ net915 net1044 VPWR VGND sg13g2_nand2_1
X_4858_ _1617_ _1616_ _1615_ VPWR VGND sg13g2_nand2b_1
X_3809_ _0611_ net1026 net1053 VPWR VGND sg13g2_nand2_1
XFILLER_5_919 VPWR VGND sg13g2_decap_8
X_4789_ _1503_ _1506_ _1549_ VPWR VGND sg13g2_nor2_1
X_6528_ net1143 VGND VPWR net251 mac2.sum_lvl2_ff\[12\] clknet_leaf_42_clk sg13g2_dfrbpq_1
X_6459_ net1134 VGND VPWR _0135_ mac2.products_ff\[75\] clknet_leaf_48_clk sg13g2_dfrbpq_1
XFILLER_47_105 VPWR VGND sg13g2_fill_2
XFILLER_29_875 VPWR VGND sg13g2_fill_2
XFILLER_29_886 VPWR VGND sg13g2_fill_2
XFILLER_28_396 VPWR VGND sg13g2_fill_1
XFILLER_43_377 VPWR VGND sg13g2_fill_2
XFILLER_4_985 VPWR VGND sg13g2_decap_8
XFILLER_46_193 VPWR VGND sg13g2_fill_1
X_5830_ VGND VPWR net277 net797 _2485_ _2484_ sg13g2_a21oi_1
X_5761_ _2418_ net799 net1022 net808 net1002 VPWR VGND sg13g2_a22oi_1
X_4712_ _1474_ _1468_ _1473_ VPWR VGND sg13g2_xnor2_1
X_5692_ mac1.total_sum\[9\] mac2.total_sum\[9\] _2357_ VPWR VGND sg13g2_and2_1
X_4643_ _1405_ _1402_ _1407_ VPWR VGND sg13g2_xor2_1
X_4574_ _1345_ _1320_ _1344_ VPWR VGND sg13g2_xnor2_1
X_6313_ net1131 VGND VPWR net48 mac1.sum_lvl2_ff\[43\] clknet_leaf_53_clk sg13g2_dfrbpq_1
X_3525_ _0334_ _0335_ _0325_ _0336_ VPWR VGND sg13g2_nand3_1
X_6244_ net1121 VGND VPWR _0252_ DP_4.matrix\[36\] clknet_leaf_32_clk sg13g2_dfrbpq_2
X_3456_ _3030_ _0268_ _0269_ VPWR VGND sg13g2_nor2_1
X_6175_ net1094 VGND VPWR _0200_ DP_2.matrix\[4\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_3387_ _2971_ _2931_ _2969_ VPWR VGND sg13g2_xnor2_1
X_5126_ _1860_ VPWR _1871_ VGND _1838_ _1861_ sg13g2_o21ai_1
X_5057_ _1802_ _1801_ _1804_ VPWR VGND sg13g2_xor2_1
X_4008_ _0801_ _0799_ _0800_ VPWR VGND sg13g2_nand2_1
X_5959_ net971 net783 _2599_ VPWR VGND sg13g2_nor2_1
XFILLER_25_377 VPWR VGND sg13g2_fill_1
XFILLER_1_900 VPWR VGND sg13g2_decap_8
XFILLER_1_977 VPWR VGND sg13g2_decap_8
XFILLER_49_959 VPWR VGND sg13g2_decap_8
Xhold40 mac2.products_ff\[10\] VPWR VGND net80 sg13g2_dlygate4sd3_1
Xhold51 mac1.products_ff\[136\] VPWR VGND net91 sg13g2_dlygate4sd3_1
Xhold62 mac1.sum_lvl1_ff\[83\] VPWR VGND net102 sg13g2_dlygate4sd3_1
Xhold73 mac2.sum_lvl2_ff\[44\] VPWR VGND net113 sg13g2_dlygate4sd3_1
Xhold95 mac1.products_ff\[141\] VPWR VGND net135 sg13g2_dlygate4sd3_1
Xhold84 mac1.products_ff\[78\] VPWR VGND net124 sg13g2_dlygate4sd3_1
XFILLER_43_130 VPWR VGND sg13g2_fill_2
XFILLER_43_141 VPWR VGND sg13g2_fill_1
X_3310_ VGND VPWR _2896_ _2897_ _2862_ _2822_ sg13g2_a21oi_2
X_4290_ _1040_ VPWR _1069_ VGND _1038_ _1041_ sg13g2_o21ai_1
X_3241_ _2829_ net1000 net1051 VPWR VGND sg13g2_nand2_1
X_3172_ VGND VPWR _2758_ _2759_ _2762_ _2753_ sg13g2_a21oi_1
Xfanout1071 net1072 net1071 VPWR VGND sg13g2_buf_8
Xfanout1060 net1068 net1060 VPWR VGND sg13g2_buf_8
Xfanout1082 net1085 net1082 VPWR VGND sg13g2_buf_8
XFILLER_48_970 VPWR VGND sg13g2_decap_8
Xfanout1093 net1095 net1093 VPWR VGND sg13g2_buf_8
X_5813_ net968 net948 _2396_ _2469_ VPWR VGND sg13g2_mux2_1
XFILLER_23_826 VPWR VGND sg13g2_fill_1
X_5744_ _2400_ _2395_ _2401_ VPWR VGND sg13g2_xor2_1
X_5675_ net30 _2341_ _2343_ VPWR VGND sg13g2_xnor2_1
X_4626_ _1386_ VPWR _1391_ VGND _1387_ _1389_ sg13g2_o21ai_1
Xhold510 DP_2.matrix\[75\] VPWR VGND net550 sg13g2_dlygate4sd3_1
X_4557_ VGND VPWR _1305_ _1308_ _1329_ _1304_ sg13g2_a21oi_1
X_3508_ _0302_ VPWR _0319_ VGND _0293_ _0303_ sg13g2_o21ai_1
X_4488_ _1262_ net897 net836 VPWR VGND sg13g2_nand2_2
X_3439_ _3017_ net1040 net974 VPWR VGND sg13g2_nand2_1
X_6227_ net1129 VGND VPWR _0235_ DP_3.matrix\[43\] clknet_leaf_34_clk sg13g2_dfrbpq_1
X_6158_ net1116 VGND VPWR _0189_ DP_1.matrix\[73\] clknet_leaf_54_clk sg13g2_dfrbpq_1
X_5109_ _1852_ _1853_ _1847_ _1855_ VPWR VGND sg13g2_nand3_1
X_6089_ net1063 VGND VPWR _0070_ mac1.products_ff\[1\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_26_675 VPWR VGND sg13g2_fill_1
XFILLER_40_100 VPWR VGND sg13g2_fill_2
XFILLER_40_144 VPWR VGND sg13g2_fill_2
Xoutput30 net30 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_1_774 VPWR VGND sg13g2_decap_8
XFILLER_49_745 VPWR VGND sg13g2_fill_2
XFILLER_16_152 VPWR VGND sg13g2_fill_2
XFILLER_13_870 VPWR VGND sg13g2_decap_8
XFILLER_20_818 VPWR VGND sg13g2_fill_1
X_3790_ _0573_ VPWR _0593_ VGND _0545_ _0571_ sg13g2_o21ai_1
XFILLER_9_841 VPWR VGND sg13g2_decap_4
XFILLER_9_896 VPWR VGND sg13g2_decap_8
X_5460_ VPWR VGND _2170_ _2169_ _2168_ mac1.sum_lvl3_ff\[25\] _2176_ mac1.sum_lvl3_ff\[5\]
+ sg13g2_a221oi_1
X_4411_ _1178_ _1186_ _1187_ VPWR VGND sg13g2_nor2_1
X_5391_ _2121_ net463 _0012_ VPWR VGND sg13g2_nor2b_1
X_4342_ _1095_ VPWR _1120_ VGND _1116_ _1118_ sg13g2_o21ai_1
XFILLER_28_1016 VPWR VGND sg13g2_decap_8
X_4273_ _1051_ _1052_ _1053_ VPWR VGND sg13g2_and2_1
XFILLER_28_1027 VPWR VGND sg13g2_fill_2
X_3224_ _2813_ _2777_ _2811_ _2812_ VPWR VGND sg13g2_and3_1
X_6012_ net1056 _0161_ VPWR VGND sg13g2_buf_1
.ends

