* NGSPICE file created from heichips25_template.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

.subckt heichips25_template VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
XFILLER_39_244 VPWR VGND sg13g2_fill_2
XFILLER_28_918 VPWR VGND sg13g2_decap_8
XFILLER_39_288 VPWR VGND sg13g2_decap_8
XFILLER_36_995 VPWR VGND sg13g2_decap_8
XFILLER_23_656 VPWR VGND sg13g2_decap_8
XFILLER_35_1009 VPWR VGND sg13g2_decap_8
XFILLER_10_306 VPWR VGND sg13g2_decap_8
XFILLER_22_166 VPWR VGND sg13g2_fill_2
XFILLER_22_177 VPWR VGND sg13g2_decap_8
XFILLER_7_7 VPWR VGND sg13g2_decap_8
XFILLER_2_516 VPWR VGND sg13g2_decap_8
XFILLER_46_715 VPWR VGND sg13g2_decap_8
XFILLER_18_428 VPWR VGND sg13g2_decap_8
X_501_ net57 VGND VPWR _123_ DP_3.matrix\[129\] clknet_5_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_27_973 VPWR VGND sg13g2_decap_8
X_432_ net133 _126_ VPWR VGND sg13g2_buf_1
XFILLER_14_612 VPWR VGND sg13g2_decap_8
XFILLER_26_63 VPWR VGND sg13g2_decap_8
XFILLER_26_483 VPWR VGND sg13g2_decap_8
XFILLER_42_976 VPWR VGND sg13g2_decap_8
XFILLER_13_144 VPWR VGND sg13g2_decap_8
XFILLER_14_667 VPWR VGND sg13g2_decap_8
X_363_ _214_ net47 net120 VPWR VGND sg13g2_nand2_1
X_294_ mac2.sum_lvl1_ff\[17\] mac2.sum_lvl1_ff\[25\] _173_ VPWR VGND sg13g2_xor2_1
XFILLER_10_895 VPWR VGND sg13g2_decap_8
XFILLER_6_866 VPWR VGND sg13g2_decap_8
XFILLER_5_365 VPWR VGND sg13g2_fill_2
XFILLER_49_531 VPWR VGND sg13g2_decap_8
XFILLER_3_67 VPWR VGND sg13g2_decap_8
XFILLER_36_225 VPWR VGND sg13g2_decap_8
XFILLER_18_940 VPWR VGND sg13g2_decap_8
XFILLER_33_954 VPWR VGND sg13g2_decap_8
XFILLER_9_660 VPWR VGND sg13g2_decap_8
XFILLER_8_170 VPWR VGND sg13g2_decap_8
XFILLER_28_715 VPWR VGND sg13g2_decap_8
XFILLER_41_1024 VPWR VGND sg13g2_decap_4
XFILLER_27_214 VPWR VGND sg13g2_decap_8
XFILLER_43_707 VPWR VGND sg13g2_decap_8
XFILLER_24_943 VPWR VGND sg13g2_decap_8
XFILLER_36_792 VPWR VGND sg13g2_decap_8
XFILLER_10_114 VPWR VGND sg13g2_decap_8
XFILLER_11_648 VPWR VGND sg13g2_decap_8
XFILLER_23_486 VPWR VGND sg13g2_decap_8
XFILLER_3_803 VPWR VGND sg13g2_decap_8
XFILLER_12_87 VPWR VGND sg13g2_decap_8
XFILLER_5_4 VPWR VGND sg13g2_fill_2
XFILLER_2_335 VPWR VGND sg13g2_decap_8
XFILLER_46_512 VPWR VGND sg13g2_decap_8
XFILLER_46_589 VPWR VGND sg13g2_decap_8
XFILLER_27_770 VPWR VGND sg13g2_decap_8
XFILLER_33_217 VPWR VGND sg13g2_fill_1
XFILLER_34_729 VPWR VGND sg13g2_decap_8
XFILLER_26_291 VPWR VGND sg13g2_decap_8
X_415_ net82 _109_ VPWR VGND sg13g2_buf_1
XFILLER_42_773 VPWR VGND sg13g2_decap_8
XFILLER_15_965 VPWR VGND sg13g2_decap_8
XFILLER_14_475 VPWR VGND sg13g2_decap_4
X_346_ _203_ _202_ _051_ VPWR VGND sg13g2_xor2_1
XFILLER_41_272 VPWR VGND sg13g2_decap_8
XFILLER_30_968 VPWR VGND sg13g2_decap_8
X_277_ _003_ _162_ _163_ VPWR VGND sg13g2_xnor2_1
XFILLER_10_692 VPWR VGND sg13g2_decap_8
XFILLER_6_663 VPWR VGND sg13g2_decap_8
XFILLER_5_184 VPWR VGND sg13g2_decap_8
XFILLER_49_350 VPWR VGND sg13g2_decap_8
XFILLER_37_567 VPWR VGND sg13g2_decap_8
XFILLER_33_751 VPWR VGND sg13g2_decap_8
XFILLER_20_423 VPWR VGND sg13g2_fill_2
XFILLER_21_946 VPWR VGND sg13g2_decap_8
XFILLER_32_272 VPWR VGND sg13g2_decap_8
XFILLER_20_434 VPWR VGND sg13g2_decap_8
Xclkbuf_4_12_0_clk clknet_0_clk clknet_4_12_0_clk VPWR VGND sg13g2_buf_8
XFILLER_9_490 VPWR VGND sg13g2_decap_8
XFILLER_28_501 VPWR VGND sg13g2_decap_4
XFILLER_43_504 VPWR VGND sg13g2_decap_8
XFILLER_15_206 VPWR VGND sg13g2_decap_8
XFILLER_28_589 VPWR VGND sg13g2_decap_8
XFILLER_24_740 VPWR VGND sg13g2_decap_8
XFILLER_30_209 VPWR VGND sg13g2_fill_1
XFILLER_11_456 VPWR VGND sg13g2_decap_8
XFILLER_12_957 VPWR VGND sg13g2_decap_8
XFILLER_23_86 VPWR VGND sg13g2_decap_8
XFILLER_3_600 VPWR VGND sg13g2_decap_8
XFILLER_3_677 VPWR VGND sg13g2_decap_8
XFILLER_2_187 VPWR VGND sg13g2_fill_1
XFILLER_47_821 VPWR VGND sg13g2_decap_8
XFILLER_46_342 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_47_898 VPWR VGND sg13g2_decap_8
XFILLER_46_364 VPWR VGND sg13g2_decap_4
XFILLER_19_567 VPWR VGND sg13g2_decap_8
XFILLER_34_526 VPWR VGND sg13g2_decap_8
XFILLER_46_386 VPWR VGND sg13g2_decap_8
XFILLER_9_11 VPWR VGND sg13g2_decap_8
XFILLER_15_762 VPWR VGND sg13g2_decap_8
XFILLER_42_570 VPWR VGND sg13g2_decap_8
XFILLER_14_261 VPWR VGND sg13g2_decap_8
XFILLER_30_765 VPWR VGND sg13g2_decap_8
X_329_ _192_ net136 net85 VPWR VGND sg13g2_nand2_1
XFILLER_31_1023 VPWR VGND sg13g2_decap_4
XFILLER_7_961 VPWR VGND sg13g2_decap_8
XFILLER_6_460 VPWR VGND sg13g2_decap_8
XFILLER_9_1024 VPWR VGND sg13g2_decap_4
XFILLER_29_0 VPWR VGND sg13g2_decap_8
XFILLER_38_810 VPWR VGND sg13g2_decap_8
XFILLER_37_342 VPWR VGND sg13g2_decap_8
XFILLER_38_887 VPWR VGND sg13g2_decap_8
XFILLER_20_231 VPWR VGND sg13g2_decap_8
XFILLER_21_743 VPWR VGND sg13g2_decap_8
XFILLER_48_618 VPWR VGND sg13g2_decap_8
XFILLER_0_658 VPWR VGND sg13g2_decap_8
XFILLER_47_139 VPWR VGND sg13g2_decap_8
XFILLER_29_854 VPWR VGND sg13g2_decap_8
XFILLER_28_364 VPWR VGND sg13g2_decap_8
XFILLER_44_857 VPWR VGND sg13g2_decap_8
XFILLER_18_97 VPWR VGND sg13g2_decap_8
XFILLER_43_345 VPWR VGND sg13g2_decap_8
XFILLER_12_754 VPWR VGND sg13g2_decap_8
XFILLER_15_1007 VPWR VGND sg13g2_decap_8
XFILLER_8_747 VPWR VGND sg13g2_decap_8
XFILLER_7_202 VPWR VGND sg13g2_decap_8
XFILLER_11_286 VPWR VGND sg13g2_decap_8
XFILLER_7_279 VPWR VGND sg13g2_decap_8
XFILLER_4_986 VPWR VGND sg13g2_decap_8
XFILLER_38_139 VPWR VGND sg13g2_decap_4
XFILLER_35_813 VPWR VGND sg13g2_decap_8
XFILLER_47_695 VPWR VGND sg13g2_decap_8
XFILLER_46_183 VPWR VGND sg13g2_decap_8
XFILLER_34_389 VPWR VGND sg13g2_decap_8
XFILLER_30_562 VPWR VGND sg13g2_decap_8
XFILLER_26_824 VPWR VGND sg13g2_decap_8
XFILLER_38_684 VPWR VGND sg13g2_decap_8
XFILLER_25_378 VPWR VGND sg13g2_decap_8
XFILLER_34_890 VPWR VGND sg13g2_decap_8
XFILLER_40_304 VPWR VGND sg13g2_decap_8
XFILLER_41_849 VPWR VGND sg13g2_decap_8
XFILLER_20_32 VPWR VGND sg13g2_decap_8
XFILLER_1_934 VPWR VGND sg13g2_decap_8
XFILLER_49_916 VPWR VGND sg13g2_decap_8
XFILLER_0_455 VPWR VGND sg13g2_decap_8
XFILLER_48_415 VPWR VGND sg13g2_decap_8
Xhold30 DP_4.matrix\[33\] VPWR VGND net54 sg13g2_dlygate4sd3_1
Xhold41 DP_2.matrix\[65\] VPWR VGND net91 sg13g2_dlygate4sd3_1
Xhold74 DP_4.matrix\[128\] VPWR VGND net124 sg13g2_dlygate4sd3_1
Xhold52 mac1.sum_lvl1_ff\[16\] VPWR VGND net102 sg13g2_dlygate4sd3_1
Xhold63 mac2.products_ff\[112\] VPWR VGND net113 sg13g2_dlygate4sd3_1
Xhold96 DP_3.matrix\[0\] VPWR VGND net146 sg13g2_dlygate4sd3_1
Xhold85 DP_2.matrix\[16\] VPWR VGND net135 sg13g2_dlygate4sd3_1
XFILLER_29_651 VPWR VGND sg13g2_decap_8
XFILLER_16_323 VPWR VGND sg13g2_decap_8
XFILLER_17_824 VPWR VGND sg13g2_decap_8
XFILLER_28_183 VPWR VGND sg13g2_decap_8
XFILLER_45_73 VPWR VGND sg13g2_decap_8
XFILLER_44_654 VPWR VGND sg13g2_decap_8
XFILLER_43_142 VPWR VGND sg13g2_decap_8
X_594_ net63 VGND VPWR _041_ mac2.products_ff\[97\] clknet_5_3__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_827 VPWR VGND sg13g2_decap_8
XFILLER_31_337 VPWR VGND sg13g2_decap_8
XFILLER_8_500 VPWR VGND sg13g2_fill_2
XFILLER_12_573 VPWR VGND sg13g2_fill_2
XFILLER_12_584 VPWR VGND sg13g2_decap_8
XFILLER_8_566 VPWR VGND sg13g2_decap_8
XFILLER_6_67 VPWR VGND sg13g2_decap_8
XFILLER_4_783 VPWR VGND sg13g2_decap_8
XFILLER_3_271 VPWR VGND sg13g2_decap_8
XFILLER_6_1027 VPWR VGND sg13g2_fill_2
XFILLER_20_4 VPWR VGND sg13g2_decap_8
XFILLER_39_459 VPWR VGND sg13g2_fill_2
XFILLER_48_982 VPWR VGND sg13g2_decap_8
XFILLER_47_492 VPWR VGND sg13g2_decap_8
XFILLER_35_610 VPWR VGND sg13g2_decap_8
XFILLER_23_838 VPWR VGND sg13g2_decap_8
XFILLER_34_175 VPWR VGND sg13g2_decap_8
XFILLER_35_687 VPWR VGND sg13g2_decap_8
XFILLER_22_337 VPWR VGND sg13g2_decap_8
XFILLER_44_1011 VPWR VGND sg13g2_decap_8
Xheichips25_template_10 VPWR VGND uio_out[5] sg13g2_tielo
Xheichips25_template_21 VPWR VGND uio_oe[4] sg13g2_tiehi
XFILLER_26_621 VPWR VGND sg13g2_decap_8
XFILLER_38_481 VPWR VGND sg13g2_fill_1
XFILLER_14_849 VPWR VGND sg13g2_decap_8
XFILLER_15_32 VPWR VGND sg13g2_decap_8
XFILLER_25_153 VPWR VGND sg13g2_decap_8
XFILLER_26_698 VPWR VGND sg13g2_decap_8
XFILLER_41_646 VPWR VGND sg13g2_decap_8
XFILLER_9_308 VPWR VGND sg13g2_decap_8
XFILLER_40_167 VPWR VGND sg13g2_decap_8
XFILLER_31_42 VPWR VGND sg13g2_decap_8
XFILLER_1_731 VPWR VGND sg13g2_decap_8
XFILLER_49_713 VPWR VGND sg13g2_decap_8
XFILLER_0_252 VPWR VGND sg13g2_decap_8
XFILLER_48_234 VPWR VGND sg13g2_decap_8
XFILLER_48_267 VPWR VGND sg13g2_decap_8
XFILLER_45_941 VPWR VGND sg13g2_decap_8
XFILLER_44_451 VPWR VGND sg13g2_decap_8
X_577_ net57 VGND VPWR net28 mac2.sum_lvl1_ff\[32\] clknet_5_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_698 VPWR VGND sg13g2_decap_8
XFILLER_32_624 VPWR VGND sg13g2_decap_8
XFILLER_31_112 VPWR VGND sg13g2_decap_4
XFILLER_8_330 VPWR VGND sg13g2_decap_8
XFILLER_9_842 VPWR VGND sg13g2_decap_8
XFILLER_13_893 VPWR VGND sg13g2_decap_8
XFILLER_8_352 VPWR VGND sg13g2_decap_8
Xclkbuf_5_17__f_clk clknet_4_8_0_clk clknet_5_17__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_4_580 VPWR VGND sg13g2_decap_8
XFILLER_39_267 VPWR VGND sg13g2_decap_4
XFILLER_27_429 VPWR VGND sg13g2_decap_8
XFILLER_36_974 VPWR VGND sg13g2_decap_8
XFILLER_35_484 VPWR VGND sg13g2_decap_8
XFILLER_23_635 VPWR VGND sg13g2_decap_8
XFILLER_22_145 VPWR VGND sg13g2_decap_8
XFILLER_22_156 VPWR VGND sg13g2_fill_2
XFILLER_18_407 VPWR VGND sg13g2_decap_8
X_500_ net57 VGND VPWR _122_ DP_3.matrix\[128\] clknet_5_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_248 VPWR VGND sg13g2_fill_2
XFILLER_26_440 VPWR VGND sg13g2_decap_8
XFILLER_27_952 VPWR VGND sg13g2_decap_8
X_431_ net51 _125_ VPWR VGND sg13g2_buf_1
XFILLER_42_955 VPWR VGND sg13g2_decap_8
XFILLER_14_646 VPWR VGND sg13g2_decap_8
X_362_ _213_ _212_ _061_ VPWR VGND sg13g2_xor2_1
XFILLER_9_138 VPWR VGND sg13g2_decap_8
X_293_ _172_ net186 net105 VPWR VGND sg13g2_nand2_1
XFILLER_42_74 VPWR VGND sg13g2_decap_8
XFILLER_6_845 VPWR VGND sg13g2_decap_8
XFILLER_10_874 VPWR VGND sg13g2_decap_8
XFILLER_5_344 VPWR VGND sg13g2_decap_8
XFILLER_3_46 VPWR VGND sg13g2_decap_8
XFILLER_49_510 VPWR VGND sg13g2_decap_8
XFILLER_49_587 VPWR VGND sg13g2_decap_8
XFILLER_37_749 VPWR VGND sg13g2_decap_8
XFILLER_18_996 VPWR VGND sg13g2_decap_8
XFILLER_33_933 VPWR VGND sg13g2_decap_8
XFILLER_20_649 VPWR VGND sg13g2_decap_8
XFILLER_32_498 VPWR VGND sg13g2_decap_8
XFILLER_13_690 VPWR VGND sg13g2_decap_8
XFILLER_41_1003 VPWR VGND sg13g2_decap_8
XFILLER_24_922 VPWR VGND sg13g2_decap_8
XFILLER_36_771 VPWR VGND sg13g2_decap_8
XFILLER_23_465 VPWR VGND sg13g2_decap_8
XFILLER_24_999 VPWR VGND sg13g2_decap_8
XFILLER_12_11 VPWR VGND sg13g2_decap_8
XFILLER_12_66 VPWR VGND sg13g2_decap_8
XFILLER_2_314 VPWR VGND sg13g2_decap_8
XFILLER_3_859 VPWR VGND sg13g2_decap_8
XFILLER_18_204 VPWR VGND sg13g2_decap_8
XFILLER_19_749 VPWR VGND sg13g2_decap_8
XFILLER_46_568 VPWR VGND sg13g2_decap_8
XFILLER_34_708 VPWR VGND sg13g2_decap_8
XFILLER_37_63 VPWR VGND sg13g2_decap_8
XFILLER_37_74 VPWR VGND sg13g2_fill_1
X_414_ net161 _108_ VPWR VGND sg13g2_buf_1
XFILLER_15_944 VPWR VGND sg13g2_decap_8
XFILLER_42_752 VPWR VGND sg13g2_decap_8
XFILLER_14_454 VPWR VGND sg13g2_decap_8
XFILLER_41_251 VPWR VGND sg13g2_decap_8
X_345_ _203_ net131 net91 VPWR VGND sg13g2_nand2_1
XFILLER_30_947 VPWR VGND sg13g2_decap_8
X_276_ mac1.products_ff\[49\] mac1.products_ff\[33\] _163_ VPWR VGND sg13g2_xor2_1
XFILLER_10_671 VPWR VGND sg13g2_decap_8
XFILLER_6_642 VPWR VGND sg13g2_decap_8
XFILLER_5_163 VPWR VGND sg13g2_decap_8
XFILLER_49_384 VPWR VGND sg13g2_decap_8
XFILLER_37_546 VPWR VGND sg13g2_decap_8
XFILLER_18_793 VPWR VGND sg13g2_decap_8
XFILLER_24_229 VPWR VGND sg13g2_decap_8
XFILLER_33_730 VPWR VGND sg13g2_decap_8
XFILLER_20_402 VPWR VGND sg13g2_decap_8
XFILLER_21_925 VPWR VGND sg13g2_decap_8
XFILLER_16_719 VPWR VGND sg13g2_decap_8
XFILLER_28_568 VPWR VGND sg13g2_decap_8
XFILLER_15_229 VPWR VGND sg13g2_fill_1
XFILLER_12_936 VPWR VGND sg13g2_decap_8
XFILLER_24_796 VPWR VGND sg13g2_decap_8
XFILLER_8_929 VPWR VGND sg13g2_decap_8
XFILLER_11_435 VPWR VGND sg13g2_decap_8
XFILLER_23_65 VPWR VGND sg13g2_decap_8
XFILLER_3_656 VPWR VGND sg13g2_decap_8
XFILLER_24_1020 VPWR VGND sg13g2_decap_8
XFILLER_47_800 VPWR VGND sg13g2_decap_8
XFILLER_48_84 VPWR VGND sg13g2_decap_4
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_19_546 VPWR VGND sg13g2_decap_8
XFILLER_47_877 VPWR VGND sg13g2_decap_8
XFILLER_34_505 VPWR VGND sg13g2_decap_8
XFILLER_15_741 VPWR VGND sg13g2_decap_8
XFILLER_30_744 VPWR VGND sg13g2_decap_8
X_328_ _191_ _190_ _039_ VPWR VGND sg13g2_xor2_1
XFILLER_9_89 VPWR VGND sg13g2_decap_8
XFILLER_31_1002 VPWR VGND sg13g2_decap_8
XFILLER_7_940 VPWR VGND sg13g2_decap_8
XFILLER_11_991 VPWR VGND sg13g2_decap_8
X_259_ _154_ net173 net102 VPWR VGND sg13g2_nand2_1
XFILLER_9_1003 VPWR VGND sg13g2_decap_8
XFILLER_37_321 VPWR VGND sg13g2_decap_8
XFILLER_38_866 VPWR VGND sg13g2_decap_8
XFILLER_37_398 VPWR VGND sg13g2_decap_8
XFILLER_21_722 VPWR VGND sg13g2_decap_8
XFILLER_21_799 VPWR VGND sg13g2_decap_8
XFILLER_20_287 VPWR VGND sg13g2_decap_8
XFILLER_4_409 VPWR VGND sg13g2_decap_8
XFILLER_0_637 VPWR VGND sg13g2_decap_8
XFILLER_47_118 VPWR VGND sg13g2_decap_8
XFILLER_18_32 VPWR VGND sg13g2_fill_1
XFILLER_29_833 VPWR VGND sg13g2_decap_8
XFILLER_18_76 VPWR VGND sg13g2_fill_1
XFILLER_44_836 VPWR VGND sg13g2_decap_8
XFILLER_43_324 VPWR VGND sg13g2_decap_8
XFILLER_16_538 VPWR VGND sg13g2_decap_8
XFILLER_24_560 VPWR VGND sg13g2_decap_8
XFILLER_31_519 VPWR VGND sg13g2_decap_8
XFILLER_12_733 VPWR VGND sg13g2_decap_8
XFILLER_34_97 VPWR VGND sg13g2_fill_2
XFILLER_8_726 VPWR VGND sg13g2_decap_8
XFILLER_11_265 VPWR VGND sg13g2_decap_8
XFILLER_7_258 VPWR VGND sg13g2_decap_8
XFILLER_4_965 VPWR VGND sg13g2_decap_8
XFILLER_3_497 VPWR VGND sg13g2_fill_2
XFILLER_38_118 VPWR VGND sg13g2_decap_8
XFILLER_47_674 VPWR VGND sg13g2_decap_8
Xclkbuf_4_11_0_clk clknet_0_clk clknet_4_11_0_clk VPWR VGND sg13g2_buf_8
XFILLER_46_162 VPWR VGND sg13g2_decap_8
XFILLER_19_376 VPWR VGND sg13g2_decap_8
XFILLER_34_324 VPWR VGND sg13g2_decap_8
XFILLER_35_869 VPWR VGND sg13g2_decap_8
XFILLER_30_541 VPWR VGND sg13g2_decap_8
XFILLER_41_0 VPWR VGND sg13g2_decap_8
XFILLER_29_129 VPWR VGND sg13g2_decap_8
XFILLER_26_803 VPWR VGND sg13g2_decap_8
XFILLER_37_140 VPWR VGND sg13g2_decap_8
XFILLER_38_663 VPWR VGND sg13g2_decap_8
XFILLER_25_313 VPWR VGND sg13g2_decap_4
XFILLER_25_357 VPWR VGND sg13g2_decap_8
XFILLER_37_195 VPWR VGND sg13g2_decap_8
XFILLER_41_828 VPWR VGND sg13g2_decap_8
XFILLER_40_327 VPWR VGND sg13g2_decap_8
XFILLER_5_729 VPWR VGND sg13g2_decap_8
XFILLER_20_11 VPWR VGND sg13g2_decap_8
XFILLER_1_913 VPWR VGND sg13g2_decap_8
XFILLER_20_88 VPWR VGND sg13g2_decap_8
XFILLER_0_434 VPWR VGND sg13g2_decap_8
Xhold31 DP_2.matrix\[1\] VPWR VGND net55 sg13g2_dlygate4sd3_1
XFILLER_29_42 VPWR VGND sg13g2_decap_8
Xhold20 DP_4.matrix\[65\] VPWR VGND net44 sg13g2_dlygate4sd3_1
Xhold42 DP_1.matrix\[33\] VPWR VGND net92 sg13g2_dlygate4sd3_1
Xhold53 _010_ VPWR VGND net103 sg13g2_dlygate4sd3_1
Xhold64 _023_ VPWR VGND net114 sg13g2_dlygate4sd3_1
XFILLER_29_630 VPWR VGND sg13g2_decap_8
XFILLER_17_803 VPWR VGND sg13g2_decap_8
Xhold75 DP_3.matrix\[112\] VPWR VGND net125 sg13g2_dlygate4sd3_1
XFILLER_21_1023 VPWR VGND sg13g2_decap_4
Xhold86 DP_4.matrix\[96\] VPWR VGND net136 sg13g2_dlygate4sd3_1
Xhold97 mac2.products_ff\[0\] VPWR VGND net147 sg13g2_dlygate4sd3_1
XFILLER_44_633 VPWR VGND sg13g2_decap_8
XFILLER_16_302 VPWR VGND sg13g2_decap_8
XFILLER_28_162 VPWR VGND sg13g2_decap_8
XFILLER_45_63 VPWR VGND sg13g2_decap_4
XFILLER_45_52 VPWR VGND sg13g2_fill_2
XFILLER_43_121 VPWR VGND sg13g2_decap_8
X_593_ net64 VGND VPWR _040_ mac2.products_ff\[96\] clknet_5_9__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_806 VPWR VGND sg13g2_decap_8
XFILLER_16_379 VPWR VGND sg13g2_decap_8
XFILLER_24_390 VPWR VGND sg13g2_decap_8
XFILLER_8_545 VPWR VGND sg13g2_decap_8
XFILLER_40_894 VPWR VGND sg13g2_decap_8
XFILLER_6_35 VPWR VGND sg13g2_decap_4
XFILLER_4_762 VPWR VGND sg13g2_decap_8
XFILLER_3_250 VPWR VGND sg13g2_decap_8
XFILLER_6_1006 VPWR VGND sg13g2_decap_8
XFILLER_13_4 VPWR VGND sg13g2_decap_8
XFILLER_39_438 VPWR VGND sg13g2_decap_8
XFILLER_48_961 VPWR VGND sg13g2_decap_8
XFILLER_47_471 VPWR VGND sg13g2_decap_8
XFILLER_19_151 VPWR VGND sg13g2_decap_4
XFILLER_19_173 VPWR VGND sg13g2_fill_2
XFILLER_35_666 VPWR VGND sg13g2_decap_8
XFILLER_16_880 VPWR VGND sg13g2_decap_8
XFILLER_22_316 VPWR VGND sg13g2_decap_8
XFILLER_23_817 VPWR VGND sg13g2_decap_8
XFILLER_34_154 VPWR VGND sg13g2_decap_8
XFILLER_30_382 VPWR VGND sg13g2_decap_8
XFILLER_31_883 VPWR VGND sg13g2_decap_8
Xheichips25_template_11 VPWR VGND uio_out[6] sg13g2_tielo
Xheichips25_template_22 VPWR VGND uio_oe[5] sg13g2_tiehi
XFILLER_26_600 VPWR VGND sg13g2_decap_8
XFILLER_25_132 VPWR VGND sg13g2_decap_8
XFILLER_14_828 VPWR VGND sg13g2_decap_8
XFILLER_15_11 VPWR VGND sg13g2_decap_8
XFILLER_26_677 VPWR VGND sg13g2_decap_8
XFILLER_41_625 VPWR VGND sg13g2_decap_8
XFILLER_40_102 VPWR VGND sg13g2_decap_8
XFILLER_40_146 VPWR VGND sg13g2_decap_8
XFILLER_31_21 VPWR VGND sg13g2_decap_8
XFILLER_31_98 VPWR VGND sg13g2_decap_8
XFILLER_1_710 VPWR VGND sg13g2_decap_8
XFILLER_0_231 VPWR VGND sg13g2_decap_8
XFILLER_1_787 VPWR VGND sg13g2_decap_8
XFILLER_49_769 VPWR VGND sg13g2_decap_8
XFILLER_36_408 VPWR VGND sg13g2_fill_2
XFILLER_45_920 VPWR VGND sg13g2_decap_8
XFILLER_44_430 VPWR VGND sg13g2_decap_8
XFILLER_45_997 VPWR VGND sg13g2_decap_8
XFILLER_16_165 VPWR VGND sg13g2_decap_4
XFILLER_17_677 VPWR VGND sg13g2_decap_8
X_576_ net67 VGND VPWR net181 mac2.sum_lvl1_ff\[25\] clknet_5_6__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_603 VPWR VGND sg13g2_decap_8
XFILLER_13_872 VPWR VGND sg13g2_decap_8
XFILLER_9_821 VPWR VGND sg13g2_decap_8
XFILLER_40_691 VPWR VGND sg13g2_decap_8
XFILLER_9_898 VPWR VGND sg13g2_decap_8
XFILLER_39_202 VPWR VGND sg13g2_fill_1
XFILLER_27_408 VPWR VGND sg13g2_decap_8
XFILLER_47_290 VPWR VGND sg13g2_decap_8
XFILLER_36_953 VPWR VGND sg13g2_decap_8
XFILLER_23_614 VPWR VGND sg13g2_decap_8
XFILLER_35_463 VPWR VGND sg13g2_decap_8
XFILLER_22_124 VPWR VGND sg13g2_decap_8
XFILLER_11_809 VPWR VGND sg13g2_decap_8
XFILLER_31_680 VPWR VGND sg13g2_decap_8
XFILLER_45_227 VPWR VGND sg13g2_decap_8
Xclkbuf_5_23__f_clk clknet_4_11_0_clk clknet_5_23__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_26_32 VPWR VGND sg13g2_decap_8
XFILLER_27_931 VPWR VGND sg13g2_decap_8
X_430_ net143 _124_ VPWR VGND sg13g2_buf_1
XFILLER_41_400 VPWR VGND sg13g2_decap_8
XFILLER_42_934 VPWR VGND sg13g2_decap_8
XFILLER_13_124 VPWR VGND sg13g2_decap_4
XFILLER_26_98 VPWR VGND sg13g2_decap_8
X_361_ _213_ net141 net44 VPWR VGND sg13g2_nand2_1
XFILLER_42_42 VPWR VGND sg13g2_decap_8
XFILLER_9_117 VPWR VGND sg13g2_decap_8
X_292_ net152 mac2.sum_lvl2_ff\[4\] _029_ VPWR VGND sg13g2_xor2_1
XFILLER_41_499 VPWR VGND sg13g2_decap_8
XFILLER_10_853 VPWR VGND sg13g2_decap_8
XFILLER_6_824 VPWR VGND sg13g2_decap_8
XFILLER_5_323 VPWR VGND sg13g2_decap_8
XFILLER_5_367 VPWR VGND sg13g2_fill_1
XFILLER_3_25 VPWR VGND sg13g2_decap_8
XFILLER_1_584 VPWR VGND sg13g2_decap_8
XFILLER_49_566 VPWR VGND sg13g2_decap_8
XFILLER_37_728 VPWR VGND sg13g2_decap_8
XFILLER_18_975 VPWR VGND sg13g2_decap_8
XFILLER_33_912 VPWR VGND sg13g2_decap_8
XFILLER_45_794 VPWR VGND sg13g2_decap_8
XFILLER_17_485 VPWR VGND sg13g2_fill_1
X_559_ net61 VGND VPWR net31 mac1.sum_lvl3_ff\[2\] clknet_5_16__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_444 VPWR VGND sg13g2_decap_8
XFILLER_33_989 VPWR VGND sg13g2_decap_8
XFILLER_20_628 VPWR VGND sg13g2_decap_8
XFILLER_12_190 VPWR VGND sg13g2_decap_8
XFILLER_9_695 VPWR VGND sg13g2_decap_8
XFILLER_5_890 VPWR VGND sg13g2_decap_8
XFILLER_27_249 VPWR VGND sg13g2_decap_8
XFILLER_42_219 VPWR VGND sg13g2_fill_1
XFILLER_24_901 VPWR VGND sg13g2_decap_8
XFILLER_36_750 VPWR VGND sg13g2_decap_8
XFILLER_23_444 VPWR VGND sg13g2_decap_8
XFILLER_24_978 VPWR VGND sg13g2_decap_8
XFILLER_10_149 VPWR VGND sg13g2_decap_8
XFILLER_12_34 VPWR VGND sg13g2_fill_2
XFILLER_12_45 VPWR VGND sg13g2_decap_8
XFILLER_3_838 VPWR VGND sg13g2_decap_8
XFILLER_5_6 VPWR VGND sg13g2_fill_1
Xhold150 _026_ VPWR VGND net200 sg13g2_dlygate4sd3_1
XFILLER_19_728 VPWR VGND sg13g2_decap_8
XFILLER_46_547 VPWR VGND sg13g2_decap_8
XFILLER_18_249 VPWR VGND sg13g2_decap_8
XFILLER_42_731 VPWR VGND sg13g2_decap_8
XFILLER_15_923 VPWR VGND sg13g2_decap_8
X_413_ net45 _107_ VPWR VGND sg13g2_buf_1
XFILLER_18_1017 VPWR VGND sg13g2_decap_8
XFILLER_18_1028 VPWR VGND sg13g2_fill_1
XFILLER_41_230 VPWR VGND sg13g2_decap_8
XFILLER_14_488 VPWR VGND sg13g2_decap_8
XFILLER_14_499 VPWR VGND sg13g2_fill_2
XFILLER_30_926 VPWR VGND sg13g2_decap_8
X_344_ _202_ net101 net157 VPWR VGND sg13g2_nand2_1
X_275_ _162_ net182 net109 VPWR VGND sg13g2_nand2_1
XFILLER_10_650 VPWR VGND sg13g2_decap_8
XFILLER_6_621 VPWR VGND sg13g2_decap_8
XFILLER_5_142 VPWR VGND sg13g2_decap_8
XFILLER_45_7 VPWR VGND sg13g2_decap_8
XFILLER_6_698 VPWR VGND sg13g2_decap_8
XFILLER_2_893 VPWR VGND sg13g2_decap_8
XFILLER_1_381 VPWR VGND sg13g2_decap_8
XFILLER_37_525 VPWR VGND sg13g2_decap_8
XFILLER_18_772 VPWR VGND sg13g2_decap_8
XFILLER_45_591 VPWR VGND sg13g2_decap_8
XFILLER_17_293 VPWR VGND sg13g2_decap_8
XFILLER_21_904 VPWR VGND sg13g2_decap_8
XFILLER_33_786 VPWR VGND sg13g2_decap_8
XFILLER_20_469 VPWR VGND sg13g2_fill_1
XFILLER_0_819 VPWR VGND sg13g2_decap_8
XFILLER_28_547 VPWR VGND sg13g2_decap_8
XFILLER_43_539 VPWR VGND sg13g2_decap_8
XFILLER_11_414 VPWR VGND sg13g2_decap_8
XFILLER_12_915 VPWR VGND sg13g2_decap_8
XFILLER_23_11 VPWR VGND sg13g2_decap_4
XFILLER_24_775 VPWR VGND sg13g2_decap_8
XFILLER_8_908 VPWR VGND sg13g2_decap_8
XFILLER_23_44 VPWR VGND sg13g2_decap_8
XFILLER_7_429 VPWR VGND sg13g2_decap_8
XFILLER_20_992 VPWR VGND sg13g2_decap_8
XFILLER_3_635 VPWR VGND sg13g2_decap_8
XFILLER_48_63 VPWR VGND sg13g2_decap_8
XFILLER_47_856 VPWR VGND sg13g2_decap_8
XFILLER_19_525 VPWR VGND sg13g2_decap_8
XFILLER_15_720 VPWR VGND sg13g2_decap_8
XFILLER_14_230 VPWR VGND sg13g2_decap_4
XFILLER_15_797 VPWR VGND sg13g2_decap_8
XFILLER_30_723 VPWR VGND sg13g2_decap_8
X_327_ _191_ net138 net50 VPWR VGND sg13g2_nand2_1
XFILLER_14_296 VPWR VGND sg13g2_decap_8
XFILLER_11_970 VPWR VGND sg13g2_decap_8
X_258_ net115 mac1.sum_lvl2_ff\[4\] _012_ VPWR VGND sg13g2_xor2_1
XFILLER_7_996 VPWR VGND sg13g2_decap_8
XFILLER_2_690 VPWR VGND sg13g2_decap_8
XFILLER_49_182 VPWR VGND sg13g2_decap_8
XFILLER_38_845 VPWR VGND sg13g2_decap_8
XFILLER_25_517 VPWR VGND sg13g2_decap_8
XFILLER_37_377 VPWR VGND sg13g2_decap_8
XFILLER_18_591 VPWR VGND sg13g2_decap_8
XFILLER_40_509 VPWR VGND sg13g2_decap_8
XFILLER_21_701 VPWR VGND sg13g2_decap_8
XFILLER_33_583 VPWR VGND sg13g2_decap_8
XFILLER_20_266 VPWR VGND sg13g2_decap_8
XFILLER_21_778 VPWR VGND sg13g2_decap_8
XFILLER_47_1010 VPWR VGND sg13g2_decap_8
XFILLER_0_616 VPWR VGND sg13g2_decap_8
XFILLER_29_812 VPWR VGND sg13g2_decap_8
XFILLER_18_11 VPWR VGND sg13g2_decap_8
XFILLER_44_815 VPWR VGND sg13g2_decap_8
XFILLER_28_344 VPWR VGND sg13g2_decap_4
XFILLER_29_889 VPWR VGND sg13g2_decap_8
XFILLER_43_303 VPWR VGND sg13g2_decap_8
XFILLER_16_517 VPWR VGND sg13g2_decap_8
XFILLER_28_399 VPWR VGND sg13g2_decap_8
XFILLER_34_21 VPWR VGND sg13g2_decap_4
XFILLER_12_712 VPWR VGND sg13g2_decap_8
XFILLER_34_76 VPWR VGND sg13g2_decap_8
XFILLER_8_705 VPWR VGND sg13g2_decap_8
XFILLER_11_244 VPWR VGND sg13g2_decap_8
XFILLER_12_789 VPWR VGND sg13g2_decap_8
XFILLER_7_237 VPWR VGND sg13g2_decap_8
XFILLER_4_944 VPWR VGND sg13g2_decap_8
XFILLER_3_410 VPWR VGND sg13g2_fill_1
XFILLER_3_454 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_47_653 VPWR VGND sg13g2_decap_8
XFILLER_46_141 VPWR VGND sg13g2_decap_8
XFILLER_19_333 VPWR VGND sg13g2_decap_8
XFILLER_19_355 VPWR VGND sg13g2_decap_8
XFILLER_34_303 VPWR VGND sg13g2_decap_8
XFILLER_35_848 VPWR VGND sg13g2_decap_8
XFILLER_15_594 VPWR VGND sg13g2_decap_8
XFILLER_30_520 VPWR VGND sg13g2_decap_8
XFILLER_30_597 VPWR VGND sg13g2_decap_8
XFILLER_7_793 VPWR VGND sg13g2_decap_8
XFILLER_6_281 VPWR VGND sg13g2_decap_8
XFILLER_34_0 VPWR VGND sg13g2_decap_8
XFILLER_29_108 VPWR VGND sg13g2_decap_8
Xclkbuf_5_4__f_clk clknet_4_2_0_clk clknet_5_4__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_38_642 VPWR VGND sg13g2_decap_8
XFILLER_1_91 VPWR VGND sg13g2_decap_8
XFILLER_26_859 VPWR VGND sg13g2_decap_8
XFILLER_41_807 VPWR VGND sg13g2_decap_8
XFILLER_33_391 VPWR VGND sg13g2_decap_8
XFILLER_5_708 VPWR VGND sg13g2_decap_8
XFILLER_4_218 VPWR VGND sg13g2_decap_8
XFILLER_20_67 VPWR VGND sg13g2_decap_8
XFILLER_0_413 VPWR VGND sg13g2_decap_8
XFILLER_1_969 VPWR VGND sg13g2_decap_8
Xhold32 DP_3.matrix\[17\] VPWR VGND net82 sg13g2_dlygate4sd3_1
Xhold10 mac1.sum_lvl1_ff\[32\] VPWR VGND net34 sg13g2_dlygate4sd3_1
Xhold21 DP_3.matrix\[1\] VPWR VGND net45 sg13g2_dlygate4sd3_1
Xhold54 DP_1.matrix\[129\] VPWR VGND net104 sg13g2_dlygate4sd3_1
Xhold65 mac1.sum_lvl2_ff\[0\] VPWR VGND net115 sg13g2_dlygate4sd3_1
XFILLER_21_1002 VPWR VGND sg13g2_decap_8
XFILLER_29_87 VPWR VGND sg13g2_decap_8
Xhold43 DP_3.matrix\[65\] VPWR VGND net93 sg13g2_dlygate4sd3_1
Xhold76 mac1.products_ff\[16\] VPWR VGND net126 sg13g2_dlygate4sd3_1
Xhold87 DP_3.matrix\[96\] VPWR VGND net137 sg13g2_dlygate4sd3_1
Xhold98 _017_ VPWR VGND net148 sg13g2_dlygate4sd3_1
XFILLER_44_612 VPWR VGND sg13g2_decap_8
XFILLER_29_686 VPWR VGND sg13g2_decap_8
X_592_ net80 VGND VPWR _045_ mac2.products_ff\[1\] clknet_5_30__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_42 VPWR VGND sg13g2_fill_2
XFILLER_16_358 VPWR VGND sg13g2_decap_8
XFILLER_17_859 VPWR VGND sg13g2_decap_8
XFILLER_44_689 VPWR VGND sg13g2_decap_8
XFILLER_31_306 VPWR VGND sg13g2_decap_8
XFILLER_31_317 VPWR VGND sg13g2_fill_2
XFILLER_43_199 VPWR VGND sg13g2_decap_8
XFILLER_25_881 VPWR VGND sg13g2_decap_8
XFILLER_12_564 VPWR VGND sg13g2_decap_4
XFILLER_40_873 VPWR VGND sg13g2_decap_8
XFILLER_4_741 VPWR VGND sg13g2_decap_8
XFILLER_48_940 VPWR VGND sg13g2_decap_8
XFILLER_0_980 VPWR VGND sg13g2_decap_8
XFILLER_47_450 VPWR VGND sg13g2_decap_8
XFILLER_19_130 VPWR VGND sg13g2_decap_8
XFILLER_34_133 VPWR VGND sg13g2_decap_8
XFILLER_35_645 VPWR VGND sg13g2_decap_8
XFILLER_15_391 VPWR VGND sg13g2_decap_8
XFILLER_31_862 VPWR VGND sg13g2_decap_8
XFILLER_7_590 VPWR VGND sg13g2_decap_8
Xheichips25_template_12 VPWR VGND uio_out[7] sg13g2_tielo
XFILLER_45_409 VPWR VGND sg13g2_decap_8
Xheichips25_template_23 VPWR VGND uio_oe[6] sg13g2_tiehi
XFILLER_38_450 VPWR VGND sg13g2_decap_8
XFILLER_39_984 VPWR VGND sg13g2_decap_8
XFILLER_26_656 VPWR VGND sg13g2_decap_8
XFILLER_14_807 VPWR VGND sg13g2_decap_8
XFILLER_41_604 VPWR VGND sg13g2_decap_8
XFILLER_25_188 VPWR VGND sg13g2_decap_8
XFILLER_40_125 VPWR VGND sg13g2_decap_8
XFILLER_15_67 VPWR VGND sg13g2_decap_8
XFILLER_21_361 VPWR VGND sg13g2_fill_1
XFILLER_22_884 VPWR VGND sg13g2_decap_8
XFILLER_5_527 VPWR VGND sg13g2_decap_8
Xclkbuf_4_10_0_clk clknet_0_clk clknet_4_10_0_clk VPWR VGND sg13g2_buf_8
XFILLER_31_77 VPWR VGND sg13g2_decap_8
XFILLER_0_210 VPWR VGND sg13g2_decap_8
XFILLER_1_766 VPWR VGND sg13g2_decap_8
XFILLER_49_748 VPWR VGND sg13g2_decap_8
XFILLER_0_287 VPWR VGND sg13g2_decap_8
XFILLER_17_656 VPWR VGND sg13g2_decap_8
XFILLER_29_483 VPWR VGND sg13g2_decap_8
XFILLER_45_976 VPWR VGND sg13g2_decap_8
XFILLER_16_144 VPWR VGND sg13g2_decap_8
X_575_ net67 VGND VPWR net114 mac2.sum_lvl1_ff\[24\] clknet_5_9__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_486 VPWR VGND sg13g2_decap_8
XFILLER_9_800 VPWR VGND sg13g2_decap_8
XFILLER_13_851 VPWR VGND sg13g2_decap_8
XFILLER_31_136 VPWR VGND sg13g2_decap_8
XFILLER_32_659 VPWR VGND sg13g2_decap_8
XFILLER_12_361 VPWR VGND sg13g2_decap_8
XFILLER_40_670 VPWR VGND sg13g2_decap_8
XFILLER_9_877 VPWR VGND sg13g2_decap_8
XFILLER_8_387 VPWR VGND sg13g2_decap_8
XFILLER_36_932 VPWR VGND sg13g2_decap_8
XFILLER_35_442 VPWR VGND sg13g2_decap_8
XFILLER_11_1012 VPWR VGND sg13g2_decap_8
XFILLER_46_729 VPWR VGND sg13g2_decap_8
XFILLER_27_910 VPWR VGND sg13g2_decap_8
XFILLER_39_781 VPWR VGND sg13g2_decap_8
XFILLER_26_11 VPWR VGND sg13g2_decap_8
XFILLER_42_913 VPWR VGND sg13g2_decap_8
XFILLER_27_987 VPWR VGND sg13g2_decap_8
XFILLER_13_103 VPWR VGND sg13g2_decap_8
XFILLER_14_626 VPWR VGND sg13g2_decap_4
XFILLER_26_77 VPWR VGND sg13g2_decap_8
XFILLER_26_497 VPWR VGND sg13g2_decap_8
X_360_ _212_ net134 net93 VPWR VGND sg13g2_nand2_1
XFILLER_41_423 VPWR VGND sg13g2_decap_8
XFILLER_41_434 VPWR VGND sg13g2_fill_2
XFILLER_42_21 VPWR VGND sg13g2_decap_8
X_291_ _030_ _170_ _171_ VPWR VGND sg13g2_xnor2_1
XFILLER_41_478 VPWR VGND sg13g2_decap_8
XFILLER_6_803 VPWR VGND sg13g2_decap_8
XFILLER_10_832 VPWR VGND sg13g2_decap_8
XFILLER_22_681 VPWR VGND sg13g2_decap_8
XFILLER_1_563 VPWR VGND sg13g2_decap_8
XFILLER_49_545 VPWR VGND sg13g2_decap_8
XFILLER_37_707 VPWR VGND sg13g2_decap_8
XFILLER_17_431 VPWR VGND sg13g2_decap_8
XFILLER_18_954 VPWR VGND sg13g2_decap_8
XFILLER_36_239 VPWR VGND sg13g2_decap_8
XFILLER_45_773 VPWR VGND sg13g2_decap_8
XFILLER_44_283 VPWR VGND sg13g2_decap_8
X_558_ net69 VGND VPWR net204 mac1.sum_lvl3_ff\[1\] clknet_5_18__leaf_clk sg13g2_dfrbpq_2
XFILLER_32_423 VPWR VGND sg13g2_decap_8
XFILLER_20_607 VPWR VGND sg13g2_decap_8
XFILLER_33_968 VPWR VGND sg13g2_decap_8
X_489_ net76 VGND VPWR _111_ DP_3.matrix\[33\] clknet_5_14__leaf_clk sg13g2_dfrbpq_1
XFILLER_34_1023 VPWR VGND sg13g2_decap_4
XFILLER_9_674 VPWR VGND sg13g2_decap_8
XFILLER_8_184 VPWR VGND sg13g2_decap_8
XFILLER_28_729 VPWR VGND sg13g2_decap_8
XFILLER_27_228 VPWR VGND sg13g2_decap_8
XFILLER_24_957 VPWR VGND sg13g2_decap_8
XFILLER_10_128 VPWR VGND sg13g2_decap_8
XFILLER_3_817 VPWR VGND sg13g2_decap_8
Xhold151 mac2.products_ff\[16\] VPWR VGND net201 sg13g2_dlygate4sd3_1
Xhold140 _005_ VPWR VGND net190 sg13g2_dlygate4sd3_1
XFILLER_2_349 VPWR VGND sg13g2_decap_8
XFILLER_19_707 VPWR VGND sg13g2_decap_8
XFILLER_37_21 VPWR VGND sg13g2_fill_1
XFILLER_46_526 VPWR VGND sg13g2_decap_8
XFILLER_15_902 VPWR VGND sg13g2_decap_8
XFILLER_42_710 VPWR VGND sg13g2_decap_8
XFILLER_27_784 VPWR VGND sg13g2_decap_8
X_412_ net146 _106_ VPWR VGND sg13g2_buf_1
XFILLER_15_979 VPWR VGND sg13g2_decap_8
XFILLER_30_905 VPWR VGND sg13g2_decap_8
XFILLER_42_787 VPWR VGND sg13g2_decap_8
X_343_ _201_ _200_ _049_ VPWR VGND sg13g2_xor2_1
X_274_ net97 mac1.products_ff\[80\] _004_ VPWR VGND sg13g2_xor2_1
XFILLER_41_286 VPWR VGND sg13g2_decap_8
XFILLER_6_600 VPWR VGND sg13g2_decap_8
XFILLER_5_121 VPWR VGND sg13g2_decap_8
XFILLER_6_677 VPWR VGND sg13g2_decap_8
XFILLER_5_198 VPWR VGND sg13g2_decap_8
XFILLER_2_872 VPWR VGND sg13g2_decap_8
XFILLER_1_360 VPWR VGND sg13g2_decap_8
XFILLER_38_7 VPWR VGND sg13g2_decap_8
XFILLER_49_364 VPWR VGND sg13g2_decap_8
XFILLER_37_504 VPWR VGND sg13g2_decap_8
XFILLER_18_751 VPWR VGND sg13g2_decap_8
XFILLER_45_570 VPWR VGND sg13g2_decap_8
XFILLER_17_272 VPWR VGND sg13g2_fill_1
XFILLER_33_765 VPWR VGND sg13g2_decap_8
XFILLER_32_242 VPWR VGND sg13g2_fill_2
XFILLER_20_448 VPWR VGND sg13g2_decap_8
XFILLER_32_286 VPWR VGND sg13g2_decap_4
XFILLER_28_526 VPWR VGND sg13g2_decap_8
XFILLER_43_518 VPWR VGND sg13g2_decap_8
XFILLER_24_754 VPWR VGND sg13g2_decap_8
XFILLER_23_253 VPWR VGND sg13g2_decap_8
XFILLER_23_297 VPWR VGND sg13g2_decap_8
XFILLER_20_971 VPWR VGND sg13g2_decap_8
XFILLER_3_614 VPWR VGND sg13g2_decap_8
XFILLER_2_102 VPWR VGND sg13g2_decap_8
XFILLER_3_4 VPWR VGND sg13g2_decap_8
XFILLER_2_157 VPWR VGND sg13g2_decap_8
XFILLER_2_168 VPWR VGND sg13g2_fill_1
XFILLER_2_179 VPWR VGND sg13g2_fill_2
XFILLER_48_42 VPWR VGND sg13g2_decap_8
XFILLER_19_504 VPWR VGND sg13g2_decap_8
XFILLER_47_835 VPWR VGND sg13g2_decap_8
XFILLER_46_356 VPWR VGND sg13g2_decap_4
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_27_581 VPWR VGND sg13g2_decap_8
XFILLER_9_36 VPWR VGND sg13g2_fill_2
XFILLER_9_25 VPWR VGND sg13g2_decap_8
XFILLER_14_242 VPWR VGND sg13g2_fill_2
XFILLER_15_776 VPWR VGND sg13g2_decap_8
XFILLER_30_702 VPWR VGND sg13g2_decap_8
X_326_ _190_ net144 net52 VPWR VGND sg13g2_nand2_1
XFILLER_42_584 VPWR VGND sg13g2_decap_8
XFILLER_14_275 VPWR VGND sg13g2_decap_8
XFILLER_30_779 VPWR VGND sg13g2_decap_8
X_257_ _013_ _152_ _153_ VPWR VGND sg13g2_xnor2_1
XFILLER_7_975 VPWR VGND sg13g2_decap_8
XFILLER_6_474 VPWR VGND sg13g2_fill_2
XFILLER_49_161 VPWR VGND sg13g2_decap_8
XFILLER_38_824 VPWR VGND sg13g2_decap_8
XFILLER_37_356 VPWR VGND sg13g2_decap_8
XFILLER_46_890 VPWR VGND sg13g2_decap_8
XFILLER_33_562 VPWR VGND sg13g2_decap_8
XFILLER_20_245 VPWR VGND sg13g2_decap_8
XFILLER_21_757 VPWR VGND sg13g2_decap_8
XFILLER_28_323 VPWR VGND sg13g2_decap_8
XFILLER_29_868 VPWR VGND sg13g2_decap_8
XFILLER_28_378 VPWR VGND sg13g2_decap_8
XFILLER_43_359 VPWR VGND sg13g2_decap_8
XFILLER_34_55 VPWR VGND sg13g2_decap_8
XFILLER_12_768 VPWR VGND sg13g2_decap_8
XFILLER_7_216 VPWR VGND sg13g2_decap_8
XFILLER_4_923 VPWR VGND sg13g2_decap_8
XFILLER_3_433 VPWR VGND sg13g2_decap_8
XFILLER_47_632 VPWR VGND sg13g2_decap_8
XFILLER_19_312 VPWR VGND sg13g2_decap_8
XFILLER_46_120 VPWR VGND sg13g2_decap_8
XFILLER_35_827 VPWR VGND sg13g2_decap_8
XFILLER_28_890 VPWR VGND sg13g2_decap_8
XFILLER_15_540 VPWR VGND sg13g2_decap_4
XFILLER_43_882 VPWR VGND sg13g2_decap_8
XFILLER_30_576 VPWR VGND sg13g2_decap_8
X_309_ _180_ net184 net117 VPWR VGND sg13g2_nand2_1
XFILLER_7_772 VPWR VGND sg13g2_decap_8
XFILLER_6_260 VPWR VGND sg13g2_decap_8
XFILLER_27_0 VPWR VGND sg13g2_decap_8
XFILLER_38_621 VPWR VGND sg13g2_decap_8
XFILLER_1_70 VPWR VGND sg13g2_decap_8
XFILLER_26_838 VPWR VGND sg13g2_decap_8
XFILLER_38_698 VPWR VGND sg13g2_decap_8
XFILLER_21_532 VPWR VGND sg13g2_decap_8
XFILLER_14_1010 VPWR VGND sg13g2_decap_8
XFILLER_20_46 VPWR VGND sg13g2_decap_8
XFILLER_1_948 VPWR VGND sg13g2_decap_8
Xhold11 mac1.products_ff\[128\] VPWR VGND net35 sg13g2_dlygate4sd3_1
XFILLER_0_469 VPWR VGND sg13g2_decap_8
Xhold22 DP_1.matrix\[1\] VPWR VGND net46 sg13g2_dlygate4sd3_1
XFILLER_48_429 VPWR VGND sg13g2_decap_8
Xhold33 DP_4.matrix\[129\] VPWR VGND net83 sg13g2_dlygate4sd3_1
Xhold44 DP_4.matrix\[97\] VPWR VGND net94 sg13g2_dlygate4sd3_1
XFILLER_29_66 VPWR VGND sg13g2_decap_8
Xhold55 mac2.sum_lvl1_ff\[16\] VPWR VGND net105 sg13g2_dlygate4sd3_1
Xhold88 DP_3.matrix\[80\] VPWR VGND net138 sg13g2_dlygate4sd3_1
Xhold99 DP_3.matrix\[48\] VPWR VGND net149 sg13g2_dlygate4sd3_1
Xhold66 _012_ VPWR VGND net116 sg13g2_dlygate4sd3_1
Xhold77 _000_ VPWR VGND net127 sg13g2_dlygate4sd3_1
XFILLER_29_665 VPWR VGND sg13g2_decap_8
XFILLER_45_21 VPWR VGND sg13g2_decap_8
XFILLER_17_838 VPWR VGND sg13g2_decap_8
X_591_ net79 VGND VPWR _044_ mac2.products_ff\[0\] clknet_5_27__leaf_clk sg13g2_dfrbpq_1
XFILLER_16_337 VPWR VGND sg13g2_decap_8
XFILLER_28_197 VPWR VGND sg13g2_decap_8
XFILLER_45_87 VPWR VGND sg13g2_fill_2
XFILLER_44_668 VPWR VGND sg13g2_decap_8
XFILLER_25_860 VPWR VGND sg13g2_decap_8
XFILLER_12_543 VPWR VGND sg13g2_decap_8
XFILLER_40_852 VPWR VGND sg13g2_decap_8
XFILLER_12_598 VPWR VGND sg13g2_decap_4
XFILLER_4_720 VPWR VGND sg13g2_decap_8
XFILLER_4_797 VPWR VGND sg13g2_decap_8
XFILLER_3_285 VPWR VGND sg13g2_decap_8
XFILLER_48_996 VPWR VGND sg13g2_decap_8
XFILLER_35_624 VPWR VGND sg13g2_decap_8
XFILLER_34_112 VPWR VGND sg13g2_decap_8
XFILLER_15_370 VPWR VGND sg13g2_decap_8
XFILLER_34_189 VPWR VGND sg13g2_decap_8
XFILLER_31_841 VPWR VGND sg13g2_decap_8
XFILLER_44_1025 VPWR VGND sg13g2_decap_4
Xheichips25_template_13 VPWR VGND uo_out[4] sg13g2_tielo
Xheichips25_template_24 VPWR VGND uio_oe[7] sg13g2_tiehi
XFILLER_39_963 VPWR VGND sg13g2_decap_8
XFILLER_25_101 VPWR VGND sg13g2_decap_8
XFILLER_26_635 VPWR VGND sg13g2_decap_8
XFILLER_25_167 VPWR VGND sg13g2_decap_8
XFILLER_15_46 VPWR VGND sg13g2_decap_8
XFILLER_22_863 VPWR VGND sg13g2_decap_8
XFILLER_5_506 VPWR VGND sg13g2_decap_8
XFILLER_31_56 VPWR VGND sg13g2_decap_8
XFILLER_1_745 VPWR VGND sg13g2_decap_8
XFILLER_49_727 VPWR VGND sg13g2_decap_8
XFILLER_0_266 VPWR VGND sg13g2_decap_8
XFILLER_48_248 VPWR VGND sg13g2_fill_2
XFILLER_29_462 VPWR VGND sg13g2_decap_8
XFILLER_45_955 VPWR VGND sg13g2_decap_8
XFILLER_16_123 VPWR VGND sg13g2_decap_8
XFILLER_17_635 VPWR VGND sg13g2_decap_8
XFILLER_44_465 VPWR VGND sg13g2_decap_8
X_574_ net76 VGND VPWR _065_ mac2.products_ff\[49\] clknet_5_12__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_638 VPWR VGND sg13g2_decap_8
XFILLER_13_830 VPWR VGND sg13g2_decap_8
XFILLER_12_340 VPWR VGND sg13g2_decap_8
XFILLER_9_856 VPWR VGND sg13g2_decap_8
XFILLER_8_366 VPWR VGND sg13g2_decap_8
XFILLER_4_594 VPWR VGND sg13g2_decap_8
XFILLER_28_1009 VPWR VGND sg13g2_decap_8
XFILLER_39_237 VPWR VGND sg13g2_decap_8
XFILLER_36_911 VPWR VGND sg13g2_decap_8
XFILLER_48_793 VPWR VGND sg13g2_decap_8
XFILLER_35_421 VPWR VGND sg13g2_decap_8
XFILLER_36_988 VPWR VGND sg13g2_decap_8
XFILLER_35_498 VPWR VGND sg13g2_decap_8
XFILLER_23_649 VPWR VGND sg13g2_decap_8
XFILLER_7_91 VPWR VGND sg13g2_fill_2
XFILLER_46_708 VPWR VGND sg13g2_decap_8
XFILLER_39_760 VPWR VGND sg13g2_decap_8
XFILLER_14_605 VPWR VGND sg13g2_decap_8
XFILLER_26_56 VPWR VGND sg13g2_decap_8
XFILLER_26_454 VPWR VGND sg13g2_fill_2
XFILLER_27_966 VPWR VGND sg13g2_decap_8
XFILLER_42_969 VPWR VGND sg13g2_decap_8
XFILLER_13_137 VPWR VGND sg13g2_decap_8
X_290_ mac2.sum_lvl2_ff\[1\] mac2.sum_lvl2_ff\[5\] _171_ VPWR VGND sg13g2_xor2_1
XFILLER_10_811 VPWR VGND sg13g2_decap_8
XFILLER_22_660 VPWR VGND sg13g2_decap_8
XFILLER_10_888 VPWR VGND sg13g2_decap_8
XFILLER_6_859 VPWR VGND sg13g2_decap_8
XFILLER_5_358 VPWR VGND sg13g2_decap_8
XFILLER_1_542 VPWR VGND sg13g2_decap_8
XFILLER_49_524 VPWR VGND sg13g2_decap_8
XFILLER_17_410 VPWR VGND sg13g2_decap_8
XFILLER_18_933 VPWR VGND sg13g2_decap_8
XFILLER_36_218 VPWR VGND sg13g2_decap_8
XFILLER_45_752 VPWR VGND sg13g2_decap_8
XFILLER_44_262 VPWR VGND sg13g2_decap_8
X_557_ net69 VGND VPWR net116 mac1.sum_lvl3_ff\[0\] clknet_5_18__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_402 VPWR VGND sg13g2_decap_8
XFILLER_33_947 VPWR VGND sg13g2_decap_8
X_488_ net76 VGND VPWR _110_ DP_3.matrix\[32\] clknet_5_15__leaf_clk sg13g2_dfrbpq_1
XFILLER_34_1002 VPWR VGND sg13g2_decap_8
XFILLER_9_653 VPWR VGND sg13g2_decap_8
XFILLER_8_163 VPWR VGND sg13g2_decap_8
XFILLER_41_1017 VPWR VGND sg13g2_decap_8
XFILLER_41_1028 VPWR VGND sg13g2_fill_1
XFILLER_28_708 VPWR VGND sg13g2_decap_8
XFILLER_48_590 VPWR VGND sg13g2_decap_8
XFILLER_23_413 VPWR VGND sg13g2_decap_4
XFILLER_24_936 VPWR VGND sg13g2_decap_8
XFILLER_36_785 VPWR VGND sg13g2_decap_8
XFILLER_10_107 VPWR VGND sg13g2_decap_8
XFILLER_23_479 VPWR VGND sg13g2_decap_8
XFILLER_12_25 VPWR VGND sg13g2_fill_1
XFILLER_2_328 VPWR VGND sg13g2_decap_8
Xhold141 mac1.sum_lvl1_ff\[8\] VPWR VGND net191 sg13g2_dlygate4sd3_1
Xhold130 mac2.products_ff\[96\] VPWR VGND net180 sg13g2_dlygate4sd3_1
Xhold152 _018_ VPWR VGND net202 sg13g2_dlygate4sd3_1
XFILLER_46_505 VPWR VGND sg13g2_decap_8
XFILLER_27_763 VPWR VGND sg13g2_decap_8
X_411_ net96 _105_ VPWR VGND sg13g2_buf_1
XFILLER_14_413 VPWR VGND sg13g2_decap_4
XFILLER_15_958 VPWR VGND sg13g2_decap_8
XFILLER_26_284 VPWR VGND sg13g2_decap_8
XFILLER_42_766 VPWR VGND sg13g2_decap_8
XFILLER_14_468 VPWR VGND sg13g2_decap_8
X_342_ _201_ net162 net84 VPWR VGND sg13g2_nand2_1
XFILLER_41_265 VPWR VGND sg13g2_decap_8
X_273_ _005_ _160_ net189 VPWR VGND sg13g2_xnor2_1
XFILLER_10_685 VPWR VGND sg13g2_decap_8
XFILLER_5_100 VPWR VGND sg13g2_decap_8
XFILLER_6_656 VPWR VGND sg13g2_decap_8
XFILLER_5_177 VPWR VGND sg13g2_decap_8
XFILLER_2_851 VPWR VGND sg13g2_decap_8
XFILLER_49_343 VPWR VGND sg13g2_decap_8
XFILLER_49_398 VPWR VGND sg13g2_decap_8
XFILLER_18_730 VPWR VGND sg13g2_decap_8
XFILLER_17_251 VPWR VGND sg13g2_decap_8
XFILLER_33_744 VPWR VGND sg13g2_decap_8
XFILLER_21_939 VPWR VGND sg13g2_decap_8
XFILLER_32_265 VPWR VGND sg13g2_decap_8
XFILLER_20_416 VPWR VGND sg13g2_decap_8
XFILLER_4_92 VPWR VGND sg13g2_decap_8
XFILLER_28_505 VPWR VGND sg13g2_fill_1
XFILLER_23_232 VPWR VGND sg13g2_decap_8
XFILLER_24_733 VPWR VGND sg13g2_decap_8
XFILLER_36_582 VPWR VGND sg13g2_decap_8
XFILLER_11_449 VPWR VGND sg13g2_decap_8
XFILLER_20_950 VPWR VGND sg13g2_decap_8
XFILLER_23_79 VPWR VGND sg13g2_decap_8
XFILLER_48_21 VPWR VGND sg13g2_decap_8
XFILLER_47_814 VPWR VGND sg13g2_decap_8
XFILLER_46_335 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_46_368 VPWR VGND sg13g2_fill_1
XFILLER_27_560 VPWR VGND sg13g2_decap_8
XFILLER_34_519 VPWR VGND sg13g2_decap_8
XFILLER_15_755 VPWR VGND sg13g2_decap_8
XFILLER_42_563 VPWR VGND sg13g2_decap_8
XFILLER_14_254 VPWR VGND sg13g2_decap_8
X_325_ _148_ _146_ _147_ net4 VPWR VGND sg13g2_a21o_2
XFILLER_30_758 VPWR VGND sg13g2_decap_8
Xfanout80 net81 net80 VPWR VGND sg13g2_buf_8
X_256_ mac1.sum_lvl2_ff\[1\] mac1.sum_lvl2_ff\[5\] _153_ VPWR VGND sg13g2_xor2_1
XFILLER_31_1016 VPWR VGND sg13g2_decap_8
XFILLER_31_1027 VPWR VGND sg13g2_fill_2
XFILLER_10_493 VPWR VGND sg13g2_decap_8
XFILLER_7_954 VPWR VGND sg13g2_decap_8
XFILLER_9_1017 VPWR VGND sg13g2_decap_8
XFILLER_9_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_140 VPWR VGND sg13g2_decap_8
XFILLER_38_803 VPWR VGND sg13g2_decap_8
XFILLER_37_302 VPWR VGND sg13g2_fill_2
XFILLER_37_335 VPWR VGND sg13g2_decap_8
XFILLER_33_541 VPWR VGND sg13g2_decap_8
XFILLER_20_224 VPWR VGND sg13g2_decap_8
XFILLER_21_736 VPWR VGND sg13g2_decap_8
XFILLER_9_280 VPWR VGND sg13g2_fill_1
XFILLER_28_302 VPWR VGND sg13g2_decap_8
XFILLER_29_847 VPWR VGND sg13g2_decap_8
XFILLER_43_338 VPWR VGND sg13g2_decap_8
XFILLER_24_530 VPWR VGND sg13g2_decap_8
XFILLER_36_390 VPWR VGND sg13g2_decap_8
XFILLER_12_747 VPWR VGND sg13g2_decap_8
XFILLER_11_279 VPWR VGND sg13g2_decap_8
Xclkload0 VPWR clkload0/Y clknet_5_7__leaf_clk VGND sg13g2_inv_1
XFILLER_4_902 VPWR VGND sg13g2_decap_8
XFILLER_3_401 VPWR VGND sg13g2_fill_1
XFILLER_4_979 VPWR VGND sg13g2_decap_8
Xclkbuf_5_29__f_clk clknet_4_14_0_clk clknet_5_29__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_47_611 VPWR VGND sg13g2_decap_8
XFILLER_35_806 VPWR VGND sg13g2_decap_8
XFILLER_47_688 VPWR VGND sg13g2_decap_8
XFILLER_46_176 VPWR VGND sg13g2_decap_8
XFILLER_46_198 VPWR VGND sg13g2_fill_2
XFILLER_34_338 VPWR VGND sg13g2_fill_1
XFILLER_43_861 VPWR VGND sg13g2_decap_8
XFILLER_42_371 VPWR VGND sg13g2_decap_8
XFILLER_30_555 VPWR VGND sg13g2_decap_8
X_308_ mac2.products_ff\[80\] net111 _021_ VPWR VGND sg13g2_xor2_1
X_239_ net133 net161 _068_ VPWR VGND sg13g2_and2_1
XFILLER_7_751 VPWR VGND sg13g2_decap_8
XFILLER_38_600 VPWR VGND sg13g2_decap_8
XFILLER_26_817 VPWR VGND sg13g2_decap_8
XFILLER_38_677 VPWR VGND sg13g2_decap_8
XFILLER_34_883 VPWR VGND sg13g2_decap_8
XFILLER_21_577 VPWR VGND sg13g2_decap_4
XFILLER_20_25 VPWR VGND sg13g2_decap_8
XFILLER_1_927 VPWR VGND sg13g2_decap_8
XFILLER_49_909 VPWR VGND sg13g2_decap_8
XFILLER_48_408 VPWR VGND sg13g2_decap_8
Xhold12 mac2.sum_lvl2_ff\[8\] VPWR VGND net36 sg13g2_dlygate4sd3_1
XFILLER_0_448 VPWR VGND sg13g2_decap_8
Xhold23 DP_1.matrix\[113\] VPWR VGND net47 sg13g2_dlygate4sd3_1
Xhold45 DP_2.matrix\[97\] VPWR VGND net95 sg13g2_dlygate4sd3_1
Xhold56 _027_ VPWR VGND net106 sg13g2_dlygate4sd3_1
Xhold34 DP_2.matrix\[81\] VPWR VGND net84 sg13g2_dlygate4sd3_1
Xhold89 DP_4.matrix\[32\] VPWR VGND net139 sg13g2_dlygate4sd3_1
Xhold78 DP_1.matrix\[16\] VPWR VGND net128 sg13g2_dlygate4sd3_1
XFILLER_28_121 VPWR VGND sg13g2_decap_8
XFILLER_29_644 VPWR VGND sg13g2_decap_8
Xhold67 mac2.products_ff\[32\] VPWR VGND net117 sg13g2_dlygate4sd3_1
X_590_ net58 VGND VPWR net25 mac2.sum_lvl2_ff\[9\] clknet_5_6__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_817 VPWR VGND sg13g2_decap_8
XFILLER_44_647 VPWR VGND sg13g2_decap_8
XFILLER_16_316 VPWR VGND sg13g2_decap_8
XFILLER_28_176 VPWR VGND sg13g2_decap_8
XFILLER_43_135 VPWR VGND sg13g2_decap_8
XFILLER_12_522 VPWR VGND sg13g2_decap_8
XFILLER_40_831 VPWR VGND sg13g2_decap_8
XFILLER_8_515 VPWR VGND sg13g2_fill_2
XFILLER_8_559 VPWR VGND sg13g2_decap_8
XFILLER_4_776 VPWR VGND sg13g2_decap_8
XFILLER_3_264 VPWR VGND sg13g2_decap_8
XFILLER_48_975 VPWR VGND sg13g2_decap_8
XFILLER_35_603 VPWR VGND sg13g2_decap_8
XFILLER_47_485 VPWR VGND sg13g2_decap_8
XFILLER_19_198 VPWR VGND sg13g2_fill_2
XFILLER_16_894 VPWR VGND sg13g2_decap_8
XFILLER_31_820 VPWR VGND sg13g2_decap_8
XFILLER_34_168 VPWR VGND sg13g2_decap_8
XFILLER_37_1022 VPWR VGND sg13g2_decap_8
XFILLER_31_897 VPWR VGND sg13g2_decap_8
XFILLER_30_396 VPWR VGND sg13g2_decap_8
XFILLER_44_1004 VPWR VGND sg13g2_decap_8
Xclkbuf_5_12__f_clk clknet_4_6_0_clk clknet_5_12__leaf_clk VPWR VGND sg13g2_buf_8
Xheichips25_template_14 VPWR VGND uo_out[5] sg13g2_tielo
XFILLER_39_942 VPWR VGND sg13g2_decap_8
XFILLER_26_614 VPWR VGND sg13g2_decap_8
XFILLER_25_146 VPWR VGND sg13g2_decap_8
XFILLER_15_25 VPWR VGND sg13g2_decap_8
XFILLER_34_680 VPWR VGND sg13g2_decap_8
XFILLER_41_639 VPWR VGND sg13g2_decap_8
XFILLER_22_842 VPWR VGND sg13g2_decap_8
XFILLER_31_35 VPWR VGND sg13g2_decap_8
XFILLER_1_724 VPWR VGND sg13g2_decap_8
XFILLER_49_706 VPWR VGND sg13g2_decap_8
XFILLER_0_245 VPWR VGND sg13g2_decap_8
XFILLER_48_227 VPWR VGND sg13g2_decap_8
XFILLER_29_441 VPWR VGND sg13g2_decap_8
XFILLER_45_934 VPWR VGND sg13g2_decap_8
XFILLER_44_444 VPWR VGND sg13g2_decap_8
X_573_ net76 VGND VPWR _064_ mac2.products_ff\[48\] clknet_5_12__leaf_clk sg13g2_dfrbpq_1
XFILLER_31_105 VPWR VGND sg13g2_decap_8
XFILLER_32_617 VPWR VGND sg13g2_decap_8
XFILLER_9_835 VPWR VGND sg13g2_decap_8
XFILLER_13_886 VPWR VGND sg13g2_decap_8
XFILLER_8_323 VPWR VGND sg13g2_decap_8
XFILLER_4_573 VPWR VGND sg13g2_decap_8
XFILLER_48_772 VPWR VGND sg13g2_decap_8
XFILLER_11_4 VPWR VGND sg13g2_decap_8
XFILLER_36_967 VPWR VGND sg13g2_decap_8
XFILLER_23_628 VPWR VGND sg13g2_decap_8
XFILLER_35_477 VPWR VGND sg13g2_decap_8
XFILLER_16_691 VPWR VGND sg13g2_decap_8
XFILLER_22_138 VPWR VGND sg13g2_decap_8
XFILLER_31_694 VPWR VGND sg13g2_decap_8
XFILLER_7_70 VPWR VGND sg13g2_decap_8
XFILLER_45_208 VPWR VGND sg13g2_decap_8
XFILLER_27_945 VPWR VGND sg13g2_decap_8
XFILLER_26_46 VPWR VGND sg13g2_decap_4
XFILLER_26_433 VPWR VGND sg13g2_decap_8
XFILLER_42_948 VPWR VGND sg13g2_decap_8
XFILLER_14_639 VPWR VGND sg13g2_decap_8
XFILLER_42_56 VPWR VGND sg13g2_decap_4
XFILLER_10_867 VPWR VGND sg13g2_decap_8
XFILLER_21_182 VPWR VGND sg13g2_decap_8
XFILLER_6_838 VPWR VGND sg13g2_decap_8
XFILLER_5_337 VPWR VGND sg13g2_decap_8
XFILLER_1_521 VPWR VGND sg13g2_decap_8
XFILLER_49_503 VPWR VGND sg13g2_decap_8
XFILLER_3_39 VPWR VGND sg13g2_decap_8
XFILLER_1_598 VPWR VGND sg13g2_decap_8
XFILLER_18_912 VPWR VGND sg13g2_decap_8
XFILLER_45_731 VPWR VGND sg13g2_decap_8
XFILLER_44_241 VPWR VGND sg13g2_decap_8
X_556_ net56 VGND VPWR net169 mac1.total_sum\[2\] clknet_5_18__leaf_clk sg13g2_dfrbpq_1
XFILLER_18_989 VPWR VGND sg13g2_decap_8
XFILLER_33_926 VPWR VGND sg13g2_decap_8
X_487_ net79 VGND VPWR _109_ DP_3.matrix\[17\] clknet_5_26__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_458 VPWR VGND sg13g2_decap_4
XFILLER_9_632 VPWR VGND sg13g2_decap_8
XFILLER_13_683 VPWR VGND sg13g2_decap_8
XFILLER_4_381 VPWR VGND sg13g2_decap_8
XFILLER_36_764 VPWR VGND sg13g2_decap_8
XFILLER_24_915 VPWR VGND sg13g2_decap_8
XFILLER_35_263 VPWR VGND sg13g2_fill_2
XFILLER_23_458 VPWR VGND sg13g2_decap_8
XFILLER_32_981 VPWR VGND sg13g2_decap_8
XFILLER_12_59 VPWR VGND sg13g2_decap_8
Xhold153 mac1.sum_lvl2_ff\[4\] VPWR VGND net203 sg13g2_dlygate4sd3_1
Xhold142 _009_ VPWR VGND net192 sg13g2_dlygate4sd3_1
Xhold120 mac2.sum_lvl3_ff\[1\] VPWR VGND net170 sg13g2_dlygate4sd3_1
Xhold131 _024_ VPWR VGND net181 sg13g2_dlygate4sd3_1
XFILLER_2_1012 VPWR VGND sg13g2_decap_8
XFILLER_37_56 VPWR VGND sg13g2_decap_8
XFILLER_27_742 VPWR VGND sg13g2_decap_8
X_410_ net150 _104_ VPWR VGND sg13g2_buf_1
XFILLER_15_937 VPWR VGND sg13g2_decap_8
XFILLER_26_252 VPWR VGND sg13g2_decap_8
XFILLER_42_745 VPWR VGND sg13g2_decap_8
XFILLER_14_447 VPWR VGND sg13g2_decap_8
X_341_ _200_ net89 net158 VPWR VGND sg13g2_nand2_1
XFILLER_41_244 VPWR VGND sg13g2_decap_8
XFILLER_23_992 VPWR VGND sg13g2_decap_8
X_272_ net188 mac1.products_ff\[81\] _161_ VPWR VGND sg13g2_xor2_1
XFILLER_10_664 VPWR VGND sg13g2_decap_8
XFILLER_6_635 VPWR VGND sg13g2_decap_8
XFILLER_5_156 VPWR VGND sg13g2_decap_8
XFILLER_2_830 VPWR VGND sg13g2_decap_8
XFILLER_49_322 VPWR VGND sg13g2_decap_8
XFILLER_1_395 VPWR VGND sg13g2_decap_8
XFILLER_37_539 VPWR VGND sg13g2_decap_8
XFILLER_17_230 VPWR VGND sg13g2_decap_8
XFILLER_18_786 VPWR VGND sg13g2_decap_8
XFILLER_32_200 VPWR VGND sg13g2_decap_8
XFILLER_33_723 VPWR VGND sg13g2_decap_8
X_539_ net60 VGND VPWR _063_ mac1.products_ff\[113\] clknet_5_24__leaf_clk sg13g2_dfrbpq_1
XFILLER_21_918 VPWR VGND sg13g2_decap_8
XFILLER_32_244 VPWR VGND sg13g2_fill_1
XFILLER_9_473 VPWR VGND sg13g2_decap_4
XFILLER_4_71 VPWR VGND sg13g2_decap_8
XFILLER_24_712 VPWR VGND sg13g2_decap_8
XFILLER_36_561 VPWR VGND sg13g2_decap_8
XFILLER_23_211 VPWR VGND sg13g2_decap_8
XFILLER_12_929 VPWR VGND sg13g2_decap_8
XFILLER_24_789 VPWR VGND sg13g2_decap_8
XFILLER_11_428 VPWR VGND sg13g2_decap_8
XFILLER_17_1020 VPWR VGND sg13g2_decap_8
XFILLER_23_58 VPWR VGND sg13g2_decap_8
XFILLER_3_649 VPWR VGND sg13g2_decap_8
XFILLER_24_1013 VPWR VGND sg13g2_decap_8
XFILLER_48_88 VPWR VGND sg13g2_fill_2
XFILLER_48_77 VPWR VGND sg13g2_decap_8
XFILLER_46_303 VPWR VGND sg13g2_decap_4
XFILLER_19_539 VPWR VGND sg13g2_decap_8
XFILLER_15_734 VPWR VGND sg13g2_decap_8
XFILLER_42_542 VPWR VGND sg13g2_decap_8
XFILLER_14_244 VPWR VGND sg13g2_fill_1
X_324_ _189_ _188_ _037_ VPWR VGND sg13g2_xor2_1
XFILLER_9_38 VPWR VGND sg13g2_fill_1
XFILLER_30_737 VPWR VGND sg13g2_decap_8
X_255_ _152_ net203 net115 VPWR VGND sg13g2_nand2_1
Xfanout70 net75 net70 VPWR VGND sg13g2_buf_8
Xfanout81 rst_n net81 VPWR VGND sg13g2_buf_8
XFILLER_7_933 VPWR VGND sg13g2_decap_8
XFILLER_11_984 VPWR VGND sg13g2_decap_8
XFILLER_6_432 VPWR VGND sg13g2_fill_1
XFILLER_6_421 VPWR VGND sg13g2_decap_8
XFILLER_43_7 VPWR VGND sg13g2_decap_8
XFILLER_1_192 VPWR VGND sg13g2_decap_8
XFILLER_37_314 VPWR VGND sg13g2_decap_8
XFILLER_49_196 VPWR VGND sg13g2_decap_8
XFILLER_38_859 VPWR VGND sg13g2_decap_8
XFILLER_18_561 VPWR VGND sg13g2_decap_8
XFILLER_33_520 VPWR VGND sg13g2_decap_8
XFILLER_21_715 VPWR VGND sg13g2_decap_8
XFILLER_33_597 VPWR VGND sg13g2_decap_8
XFILLER_47_1024 VPWR VGND sg13g2_decap_4
XFILLER_18_25 VPWR VGND sg13g2_decap_8
XFILLER_29_826 VPWR VGND sg13g2_decap_8
XFILLER_44_829 VPWR VGND sg13g2_decap_8
XFILLER_43_317 VPWR VGND sg13g2_decap_8
XFILLER_18_69 VPWR VGND sg13g2_decap_8
XFILLER_34_35 VPWR VGND sg13g2_fill_2
XFILLER_11_214 VPWR VGND sg13g2_decap_8
XFILLER_12_726 VPWR VGND sg13g2_decap_8
XFILLER_8_719 VPWR VGND sg13g2_decap_8
Xclkload1 VPWR clkload1/Y clknet_5_11__leaf_clk VGND sg13g2_inv_1
XFILLER_11_258 VPWR VGND sg13g2_decap_8
XFILLER_4_958 VPWR VGND sg13g2_decap_8
XFILLER_3_468 VPWR VGND sg13g2_fill_2
XFILLER_47_667 VPWR VGND sg13g2_decap_8
XFILLER_46_155 VPWR VGND sg13g2_decap_8
XFILLER_19_369 VPWR VGND sg13g2_decap_8
XFILLER_34_317 VPWR VGND sg13g2_decap_8
XFILLER_43_840 VPWR VGND sg13g2_decap_8
XFILLER_42_350 VPWR VGND sg13g2_decap_8
XFILLER_42_394 VPWR VGND sg13g2_decap_8
XFILLER_30_534 VPWR VGND sg13g2_decap_8
X_307_ _022_ _178_ net176 VPWR VGND sg13g2_xnor2_1
X_238_ net139 net163 _066_ VPWR VGND sg13g2_and2_1
XFILLER_7_730 VPWR VGND sg13g2_decap_8
XFILLER_11_781 VPWR VGND sg13g2_decap_8
XFILLER_6_295 VPWR VGND sg13g2_decap_8
XFILLER_37_133 VPWR VGND sg13g2_decap_8
XFILLER_38_656 VPWR VGND sg13g2_decap_8
XFILLER_25_306 VPWR VGND sg13g2_decap_8
XFILLER_37_188 VPWR VGND sg13g2_decap_8
XFILLER_18_391 VPWR VGND sg13g2_fill_1
XFILLER_34_862 VPWR VGND sg13g2_decap_8
XFILLER_33_361 VPWR VGND sg13g2_fill_2
XFILLER_1_906 VPWR VGND sg13g2_decap_8
XFILLER_0_427 VPWR VGND sg13g2_decap_8
Xhold13 mac1.products_ff\[96\] VPWR VGND net37 sg13g2_dlygate4sd3_1
XFILLER_29_35 VPWR VGND sg13g2_fill_2
Xhold46 DP_2.matrix\[129\] VPWR VGND net96 sg13g2_dlygate4sd3_1
Xhold35 DP_3.matrix\[97\] VPWR VGND net85 sg13g2_dlygate4sd3_1
Xhold24 DP_1.matrix\[97\] VPWR VGND net48 sg13g2_dlygate4sd3_1
Xhold57 mac2.sum_lvl3_ff\[2\] VPWR VGND net107 sg13g2_dlygate4sd3_1
Xhold79 mac1.sum_lvl1_ff\[0\] VPWR VGND net129 sg13g2_dlygate4sd3_1
XFILLER_21_1016 VPWR VGND sg13g2_decap_8
XFILLER_21_1027 VPWR VGND sg13g2_fill_2
XFILLER_28_100 VPWR VGND sg13g2_decap_8
XFILLER_29_623 VPWR VGND sg13g2_decap_8
Xhold68 _019_ VPWR VGND net118 sg13g2_dlygate4sd3_1
XFILLER_44_626 VPWR VGND sg13g2_decap_8
XFILLER_45_89 VPWR VGND sg13g2_fill_1
XFILLER_45_67 VPWR VGND sg13g2_fill_2
XFILLER_25_895 VPWR VGND sg13g2_decap_8
XFILLER_40_810 VPWR VGND sg13g2_decap_8
XFILLER_24_383 VPWR VGND sg13g2_decap_8
XFILLER_40_887 VPWR VGND sg13g2_decap_8
XFILLER_6_39 VPWR VGND sg13g2_fill_1
XFILLER_6_28 VPWR VGND sg13g2_decap_8
XFILLER_4_755 VPWR VGND sg13g2_decap_8
XFILLER_3_243 VPWR VGND sg13g2_decap_8
XFILLER_48_954 VPWR VGND sg13g2_decap_8
XFILLER_0_994 VPWR VGND sg13g2_decap_8
XFILLER_47_464 VPWR VGND sg13g2_decap_8
XFILLER_19_144 VPWR VGND sg13g2_decap_8
XFILLER_19_155 VPWR VGND sg13g2_fill_1
XFILLER_34_147 VPWR VGND sg13g2_decap_8
XFILLER_35_659 VPWR VGND sg13g2_decap_8
XFILLER_37_1001 VPWR VGND sg13g2_decap_8
XFILLER_16_873 VPWR VGND sg13g2_decap_8
XFILLER_22_309 VPWR VGND sg13g2_decap_8
XFILLER_42_191 VPWR VGND sg13g2_decap_8
XFILLER_30_342 VPWR VGND sg13g2_decap_8
XFILLER_31_876 VPWR VGND sg13g2_decap_8
XFILLER_30_375 VPWR VGND sg13g2_decap_8
XFILLER_32_0 VPWR VGND sg13g2_decap_8
XFILLER_39_921 VPWR VGND sg13g2_decap_8
Xheichips25_template_15 VPWR VGND uo_out[6] sg13g2_tielo
XFILLER_39_998 VPWR VGND sg13g2_decap_8
XFILLER_25_125 VPWR VGND sg13g2_decap_8
XFILLER_41_618 VPWR VGND sg13g2_decap_8
XFILLER_22_821 VPWR VGND sg13g2_decap_8
XFILLER_40_139 VPWR VGND sg13g2_decap_8
XFILLER_21_342 VPWR VGND sg13g2_fill_2
XFILLER_22_898 VPWR VGND sg13g2_decap_8
XFILLER_31_14 VPWR VGND sg13g2_decap_8
XFILLER_1_703 VPWR VGND sg13g2_decap_8
XFILLER_0_224 VPWR VGND sg13g2_decap_8
XFILLER_29_420 VPWR VGND sg13g2_decap_8
XFILLER_45_913 VPWR VGND sg13g2_decap_8
XFILLER_44_423 VPWR VGND sg13g2_decap_8
XFILLER_29_497 VPWR VGND sg13g2_decap_8
X_572_ net65 VGND VPWR net177 mac2.sum_lvl1_ff\[17\] clknet_5_9__leaf_clk sg13g2_dfrbpq_1
XFILLER_16_158 VPWR VGND sg13g2_decap_8
XFILLER_25_692 VPWR VGND sg13g2_decap_8
XFILLER_8_302 VPWR VGND sg13g2_decap_8
XFILLER_9_814 VPWR VGND sg13g2_decap_8
XFILLER_13_865 VPWR VGND sg13g2_decap_8
XFILLER_12_375 VPWR VGND sg13g2_fill_2
XFILLER_40_684 VPWR VGND sg13g2_decap_8
XFILLER_4_552 VPWR VGND sg13g2_decap_8
XFILLER_0_791 VPWR VGND sg13g2_decap_8
XFILLER_48_751 VPWR VGND sg13g2_decap_8
XFILLER_47_283 VPWR VGND sg13g2_decap_8
XFILLER_36_946 VPWR VGND sg13g2_decap_8
XFILLER_35_456 VPWR VGND sg13g2_decap_8
XFILLER_16_670 VPWR VGND sg13g2_decap_8
XFILLER_23_607 VPWR VGND sg13g2_decap_8
XFILLER_44_990 VPWR VGND sg13g2_decap_8
XFILLER_22_117 VPWR VGND sg13g2_decap_8
XFILLER_31_673 VPWR VGND sg13g2_decap_8
XFILLER_8_880 VPWR VGND sg13g2_decap_8
XFILLER_11_1026 VPWR VGND sg13g2_fill_2
XFILLER_7_93 VPWR VGND sg13g2_fill_1
XFILLER_27_924 VPWR VGND sg13g2_decap_8
XFILLER_39_795 VPWR VGND sg13g2_decap_8
XFILLER_26_25 VPWR VGND sg13g2_decap_8
XFILLER_42_927 VPWR VGND sg13g2_decap_8
XFILLER_13_117 VPWR VGND sg13g2_decap_8
XFILLER_42_35 VPWR VGND sg13g2_decap_8
XFILLER_22_695 VPWR VGND sg13g2_decap_8
XFILLER_6_817 VPWR VGND sg13g2_decap_8
XFILLER_10_846 VPWR VGND sg13g2_decap_8
XFILLER_5_316 VPWR VGND sg13g2_decap_8
XFILLER_1_500 VPWR VGND sg13g2_decap_8
XFILLER_3_18 VPWR VGND sg13g2_decap_8
XFILLER_1_577 VPWR VGND sg13g2_decap_8
XFILLER_27_1022 VPWR VGND sg13g2_decap_8
XFILLER_49_559 VPWR VGND sg13g2_decap_8
XFILLER_45_710 VPWR VGND sg13g2_decap_8
XFILLER_29_272 VPWR VGND sg13g2_decap_8
XFILLER_44_220 VPWR VGND sg13g2_decap_8
XFILLER_17_445 VPWR VGND sg13g2_fill_1
XFILLER_18_968 VPWR VGND sg13g2_decap_8
XFILLER_33_905 VPWR VGND sg13g2_decap_8
XFILLER_45_787 VPWR VGND sg13g2_decap_8
X_555_ net56 VGND VPWR net206 mac1.total_sum\[1\] clknet_5_16__leaf_clk sg13g2_dfrbpq_1
X_486_ net79 VGND VPWR _108_ DP_3.matrix\[16\] clknet_5_27__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_297 VPWR VGND sg13g2_decap_8
XFILLER_32_437 VPWR VGND sg13g2_decap_8
XFILLER_9_611 VPWR VGND sg13g2_decap_8
XFILLER_13_662 VPWR VGND sg13g2_decap_8
XFILLER_40_481 VPWR VGND sg13g2_decap_8
XFILLER_41_982 VPWR VGND sg13g2_decap_8
XFILLER_12_183 VPWR VGND sg13g2_decap_8
XFILLER_9_688 VPWR VGND sg13g2_decap_8
XFILLER_8_198 VPWR VGND sg13g2_decap_8
XFILLER_5_883 VPWR VGND sg13g2_decap_8
XFILLER_4_360 VPWR VGND sg13g2_decap_8
XFILLER_36_743 VPWR VGND sg13g2_decap_8
XFILLER_35_242 VPWR VGND sg13g2_decap_8
XFILLER_32_960 VPWR VGND sg13g2_decap_8
Xhold110 DP_1.matrix\[32\] VPWR VGND net160 sg13g2_dlygate4sd3_1
Xhold132 mac1.products_ff\[32\] VPWR VGND net182 sg13g2_dlygate4sd3_1
Xhold121 _183_ VPWR VGND net171 sg13g2_dlygate4sd3_1
Xhold143 mac1.products_ff\[97\] VPWR VGND net193 sg13g2_dlygate4sd3_1
Xhold154 _013_ VPWR VGND net204 sg13g2_dlygate4sd3_1
XFILLER_27_721 VPWR VGND sg13g2_decap_8
XFILLER_26_231 VPWR VGND sg13g2_decap_8
XFILLER_39_592 VPWR VGND sg13g2_decap_8
XFILLER_15_916 VPWR VGND sg13g2_decap_8
XFILLER_42_724 VPWR VGND sg13g2_decap_8
X_340_ _199_ _198_ _047_ VPWR VGND sg13g2_xor2_1
XFILLER_27_798 VPWR VGND sg13g2_decap_8
XFILLER_41_223 VPWR VGND sg13g2_decap_8
XFILLER_30_919 VPWR VGND sg13g2_decap_8
XFILLER_23_971 VPWR VGND sg13g2_decap_8
X_271_ _160_ mac1.products_ff\[80\] net97 VPWR VGND sg13g2_nand2_1
XFILLER_10_643 VPWR VGND sg13g2_decap_8
XFILLER_6_614 VPWR VGND sg13g2_decap_8
XFILLER_5_135 VPWR VGND sg13g2_decap_8
XFILLER_49_301 VPWR VGND sg13g2_decap_8
XFILLER_2_886 VPWR VGND sg13g2_decap_8
XFILLER_1_374 VPWR VGND sg13g2_decap_8
XFILLER_37_518 VPWR VGND sg13g2_decap_8
XFILLER_18_765 VPWR VGND sg13g2_decap_8
XFILLER_33_702 VPWR VGND sg13g2_decap_8
XFILLER_45_584 VPWR VGND sg13g2_decap_8
XFILLER_17_286 VPWR VGND sg13g2_decap_8
X_538_ net62 VGND VPWR _062_ mac1.products_ff\[112\] clknet_5_7__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_779 VPWR VGND sg13g2_decap_8
XFILLER_14_982 VPWR VGND sg13g2_decap_8
X_469_ net74 VGND VPWR _091_ DP_2.matrix\[17\] clknet_5_22__leaf_clk sg13g2_dfrbpq_1
XFILLER_9_452 VPWR VGND sg13g2_decap_8
XFILLER_13_492 VPWR VGND sg13g2_decap_8
XFILLER_5_680 VPWR VGND sg13g2_decap_8
XFILLER_4_190 VPWR VGND sg13g2_decap_8
XFILLER_4_50 VPWR VGND sg13g2_decap_8
XFILLER_36_540 VPWR VGND sg13g2_decap_8
XFILLER_12_908 VPWR VGND sg13g2_decap_8
XFILLER_24_768 VPWR VGND sg13g2_decap_8
XFILLER_11_407 VPWR VGND sg13g2_decap_8
XFILLER_23_15 VPWR VGND sg13g2_fill_2
XFILLER_23_267 VPWR VGND sg13g2_decap_4
XFILLER_20_985 VPWR VGND sg13g2_decap_8
XFILLER_3_628 VPWR VGND sg13g2_decap_8
XFILLER_2_116 VPWR VGND sg13g2_decap_4
XFILLER_48_56 VPWR VGND sg13g2_decap_8
XFILLER_19_518 VPWR VGND sg13g2_decap_8
XFILLER_47_849 VPWR VGND sg13g2_decap_8
XFILLER_42_521 VPWR VGND sg13g2_decap_8
XFILLER_15_713 VPWR VGND sg13g2_decap_8
XFILLER_27_595 VPWR VGND sg13g2_decap_8
XFILLER_14_223 VPWR VGND sg13g2_decap_8
XFILLER_42_598 VPWR VGND sg13g2_decap_8
X_323_ _189_ net142 net83 VPWR VGND sg13g2_nand2_1
XFILLER_14_289 VPWR VGND sg13g2_decap_8
XFILLER_30_716 VPWR VGND sg13g2_decap_8
Xfanout71 net74 net71 VPWR VGND sg13g2_buf_8
Xfanout60 net61 net60 VPWR VGND sg13g2_buf_8
X_254_ net126 mac1.products_ff\[0\] _000_ VPWR VGND sg13g2_xor2_1
XFILLER_7_912 VPWR VGND sg13g2_decap_8
XFILLER_11_963 VPWR VGND sg13g2_decap_8
XFILLER_13_81 VPWR VGND sg13g2_decap_8
XFILLER_7_989 VPWR VGND sg13g2_decap_8
XFILLER_2_683 VPWR VGND sg13g2_decap_8
XFILLER_36_7 VPWR VGND sg13g2_decap_8
XFILLER_1_171 VPWR VGND sg13g2_decap_8
XFILLER_49_175 VPWR VGND sg13g2_decap_8
XFILLER_37_304 VPWR VGND sg13g2_fill_1
XFILLER_38_838 VPWR VGND sg13g2_decap_8
XFILLER_18_540 VPWR VGND sg13g2_decap_4
XFILLER_45_381 VPWR VGND sg13g2_decap_8
XFILLER_33_576 VPWR VGND sg13g2_decap_8
XFILLER_20_259 VPWR VGND sg13g2_decap_8
XFILLER_9_271 VPWR VGND sg13g2_decap_8
XFILLER_47_1003 VPWR VGND sg13g2_decap_8
XFILLER_0_609 VPWR VGND sg13g2_decap_8
XFILLER_29_805 VPWR VGND sg13g2_decap_8
XFILLER_18_37 VPWR VGND sg13g2_fill_2
XFILLER_28_337 VPWR VGND sg13g2_fill_2
XFILLER_28_348 VPWR VGND sg13g2_fill_2
XFILLER_44_808 VPWR VGND sg13g2_decap_8
XFILLER_37_882 VPWR VGND sg13g2_decap_8
XFILLER_34_14 VPWR VGND sg13g2_decap_8
XFILLER_34_25 VPWR VGND sg13g2_fill_2
XFILLER_12_705 VPWR VGND sg13g2_decap_8
XFILLER_34_69 VPWR VGND sg13g2_decap_8
XFILLER_11_237 VPWR VGND sg13g2_decap_8
Xclkload2 clknet_5_12__leaf_clk clkload2/X VPWR VGND sg13g2_buf_1
XFILLER_20_782 VPWR VGND sg13g2_decap_8
XFILLER_4_937 VPWR VGND sg13g2_decap_8
XFILLER_3_447 VPWR VGND sg13g2_decap_8
XFILLER_47_646 VPWR VGND sg13g2_decap_8
XFILLER_19_326 VPWR VGND sg13g2_decap_8
XFILLER_46_134 VPWR VGND sg13g2_decap_8
XFILLER_43_896 VPWR VGND sg13g2_decap_8
XFILLER_15_587 VPWR VGND sg13g2_decap_8
XFILLER_30_513 VPWR VGND sg13g2_decap_8
X_306_ net175 mac2.products_ff\[65\] _179_ VPWR VGND sg13g2_xor2_1
XFILLER_11_760 VPWR VGND sg13g2_decap_8
X_237_ net145 net149 _064_ VPWR VGND sg13g2_and2_1
XFILLER_7_786 VPWR VGND sg13g2_decap_8
XFILLER_6_274 VPWR VGND sg13g2_decap_8
XFILLER_3_992 VPWR VGND sg13g2_decap_8
XFILLER_38_635 VPWR VGND sg13g2_decap_8
XFILLER_1_84 VPWR VGND sg13g2_decap_8
XFILLER_19_882 VPWR VGND sg13g2_decap_8
XFILLER_34_841 VPWR VGND sg13g2_decap_8
XFILLER_33_384 VPWR VGND sg13g2_decap_8
XFILLER_14_1024 VPWR VGND sg13g2_decap_4
XFILLER_0_406 VPWR VGND sg13g2_decap_8
Xhold14 _006_ VPWR VGND net38 sg13g2_dlygate4sd3_1
XFILLER_29_14 VPWR VGND sg13g2_fill_1
Xhold36 DP_1.matrix\[49\] VPWR VGND net86 sg13g2_dlygate4sd3_1
Xhold25 DP_2.matrix\[17\] VPWR VGND net49 sg13g2_dlygate4sd3_1
Xhold47 mac1.products_ff\[64\] VPWR VGND net97 sg13g2_dlygate4sd3_1
XFILLER_29_602 VPWR VGND sg13g2_decap_8
Xhold69 DP_1.matrix\[128\] VPWR VGND net119 sg13g2_dlygate4sd3_1
Xhold58 _032_ VPWR VGND net108 sg13g2_dlygate4sd3_1
XFILLER_44_605 VPWR VGND sg13g2_decap_8
XFILLER_29_679 VPWR VGND sg13g2_decap_8
XFILLER_45_35 VPWR VGND sg13g2_decap_8
XFILLER_24_351 VPWR VGND sg13g2_decap_4
XFILLER_25_874 VPWR VGND sg13g2_decap_8
XFILLER_8_517 VPWR VGND sg13g2_fill_1
XFILLER_12_557 VPWR VGND sg13g2_decap_8
XFILLER_40_866 VPWR VGND sg13g2_decap_8
XFILLER_4_734 VPWR VGND sg13g2_decap_8
XFILLER_3_222 VPWR VGND sg13g2_decap_8
XFILLER_10_93 VPWR VGND sg13g2_decap_8
XFILLER_3_299 VPWR VGND sg13g2_decap_8
XFILLER_0_973 VPWR VGND sg13g2_decap_8
XFILLER_48_933 VPWR VGND sg13g2_decap_8
XFILLER_19_123 VPWR VGND sg13g2_decap_8
XFILLER_47_443 VPWR VGND sg13g2_decap_8
XFILLER_35_638 VPWR VGND sg13g2_decap_8
XFILLER_16_852 VPWR VGND sg13g2_decap_8
XFILLER_34_126 VPWR VGND sg13g2_decap_8
XFILLER_43_693 VPWR VGND sg13g2_decap_8
XFILLER_42_170 VPWR VGND sg13g2_decap_8
XFILLER_15_384 VPWR VGND sg13g2_decap_8
XFILLER_31_855 VPWR VGND sg13g2_decap_8
XFILLER_7_583 VPWR VGND sg13g2_decap_8
XFILLER_39_900 VPWR VGND sg13g2_decap_8
Xheichips25_template_16 VPWR VGND uo_out[7] sg13g2_tielo
XFILLER_38_443 VPWR VGND sg13g2_decap_8
XFILLER_39_977 VPWR VGND sg13g2_decap_8
XFILLER_25_115 VPWR VGND sg13g2_fill_2
XFILLER_26_649 VPWR VGND sg13g2_decap_8
XFILLER_22_800 VPWR VGND sg13g2_decap_8
XFILLER_21_321 VPWR VGND sg13g2_decap_8
XFILLER_33_170 VPWR VGND sg13g2_decap_8
XFILLER_40_118 VPWR VGND sg13g2_decap_8
XFILLER_21_332 VPWR VGND sg13g2_fill_2
XFILLER_21_354 VPWR VGND sg13g2_decap_8
XFILLER_22_877 VPWR VGND sg13g2_decap_8
XFILLER_21_398 VPWR VGND sg13g2_decap_8
XFILLER_0_203 VPWR VGND sg13g2_decap_8
XFILLER_1_759 VPWR VGND sg13g2_decap_8
XFILLER_29_476 VPWR VGND sg13g2_decap_8
X_571_ net65 VGND VPWR net112 mac2.sum_lvl1_ff\[16\] clknet_5_9__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_969 VPWR VGND sg13g2_decap_8
XFILLER_16_137 VPWR VGND sg13g2_decap_8
XFILLER_17_649 VPWR VGND sg13g2_decap_8
XFILLER_44_479 VPWR VGND sg13g2_decap_8
XFILLER_25_671 VPWR VGND sg13g2_decap_8
XFILLER_13_844 VPWR VGND sg13g2_decap_8
XFILLER_31_129 VPWR VGND sg13g2_decap_8
XFILLER_12_354 VPWR VGND sg13g2_decap_8
XFILLER_24_192 VPWR VGND sg13g2_decap_8
XFILLER_40_663 VPWR VGND sg13g2_decap_8
XFILLER_48_730 VPWR VGND sg13g2_decap_8
XFILLER_0_770 VPWR VGND sg13g2_decap_8
XFILLER_36_925 VPWR VGND sg13g2_decap_8
XFILLER_35_435 VPWR VGND sg13g2_decap_8
XFILLER_43_490 VPWR VGND sg13g2_decap_8
XFILLER_31_652 VPWR VGND sg13g2_decap_8
XFILLER_30_140 VPWR VGND sg13g2_decap_8
XFILLER_11_1005 VPWR VGND sg13g2_decap_8
XFILLER_27_903 VPWR VGND sg13g2_decap_8
XFILLER_38_251 VPWR VGND sg13g2_decap_4
XFILLER_39_774 VPWR VGND sg13g2_decap_8
XFILLER_42_906 VPWR VGND sg13g2_decap_8
XFILLER_14_619 VPWR VGND sg13g2_decap_8
XFILLER_41_416 VPWR VGND sg13g2_decap_8
XFILLER_42_14 VPWR VGND sg13g2_decap_8
XFILLER_10_825 VPWR VGND sg13g2_decap_8
XFILLER_22_674 VPWR VGND sg13g2_decap_8
XFILLER_27_1001 VPWR VGND sg13g2_decap_8
XFILLER_1_556 VPWR VGND sg13g2_decap_8
XFILLER_49_538 VPWR VGND sg13g2_decap_8
XFILLER_29_251 VPWR VGND sg13g2_decap_8
XFILLER_17_424 VPWR VGND sg13g2_decap_8
XFILLER_18_947 VPWR VGND sg13g2_decap_8
XFILLER_45_766 VPWR VGND sg13g2_decap_8
X_554_ net56 VGND VPWR net166 mac1.total_sum\[0\] clknet_5_5__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_276 VPWR VGND sg13g2_decap_8
XFILLER_32_416 VPWR VGND sg13g2_decap_8
X_485_ net78 VGND VPWR _107_ DP_3.matrix\[1\] clknet_5_31__leaf_clk sg13g2_dfrbpq_1
XFILLER_13_641 VPWR VGND sg13g2_decap_8
XFILLER_41_961 VPWR VGND sg13g2_decap_8
XFILLER_12_162 VPWR VGND sg13g2_decap_8
XFILLER_34_1016 VPWR VGND sg13g2_decap_8
XFILLER_34_1027 VPWR VGND sg13g2_fill_2
XFILLER_40_460 VPWR VGND sg13g2_decap_8
XFILLER_9_667 VPWR VGND sg13g2_decap_8
XFILLER_8_177 VPWR VGND sg13g2_decap_8
XFILLER_5_862 VPWR VGND sg13g2_decap_8
XFILLER_35_221 VPWR VGND sg13g2_decap_8
XFILLER_36_722 VPWR VGND sg13g2_decap_8
XFILLER_35_265 VPWR VGND sg13g2_fill_1
XFILLER_36_799 VPWR VGND sg13g2_decap_8
XFILLER_31_460 VPWR VGND sg13g2_fill_1
Xhold100 DP_2.matrix\[128\] VPWR VGND net150 sg13g2_dlygate4sd3_1
Xhold111 DP_3.matrix\[16\] VPWR VGND net161 sg13g2_dlygate4sd3_1
Xhold133 _003_ VPWR VGND net183 sg13g2_dlygate4sd3_1
Xhold122 _031_ VPWR VGND net172 sg13g2_dlygate4sd3_1
Xhold144 _159_ VPWR VGND net194 sg13g2_dlygate4sd3_1
Xhold155 mac1.sum_lvl3_ff\[2\] VPWR VGND net205 sg13g2_dlygate4sd3_1
XFILLER_37_14 VPWR VGND sg13g2_decap_8
XFILLER_46_519 VPWR VGND sg13g2_decap_8
XFILLER_27_700 VPWR VGND sg13g2_decap_8
XFILLER_39_571 VPWR VGND sg13g2_decap_8
XFILLER_26_210 VPWR VGND sg13g2_fill_1
XFILLER_42_703 VPWR VGND sg13g2_decap_8
XFILLER_27_777 VPWR VGND sg13g2_decap_8
XFILLER_26_298 VPWR VGND sg13g2_decap_8
XFILLER_41_202 VPWR VGND sg13g2_decap_8
XFILLER_23_950 VPWR VGND sg13g2_decap_8
X_270_ net37 mac1.products_ff\[112\] _006_ VPWR VGND sg13g2_xor2_1
XFILLER_41_279 VPWR VGND sg13g2_decap_8
XFILLER_10_622 VPWR VGND sg13g2_decap_8
XFILLER_22_493 VPWR VGND sg13g2_decap_8
XFILLER_10_699 VPWR VGND sg13g2_decap_8
XFILLER_5_114 VPWR VGND sg13g2_decap_8
XFILLER_2_865 VPWR VGND sg13g2_decap_8
XFILLER_1_353 VPWR VGND sg13g2_decap_8
XFILLER_49_357 VPWR VGND sg13g2_decap_8
XFILLER_40_1020 VPWR VGND sg13g2_decap_8
XFILLER_18_744 VPWR VGND sg13g2_decap_8
XFILLER_45_563 VPWR VGND sg13g2_decap_8
X_537_ net61 VGND VPWR net27 mac1.sum_lvl1_ff\[33\] clknet_5_5__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_265 VPWR VGND sg13g2_decap_8
XFILLER_32_235 VPWR VGND sg13g2_decap_8
XFILLER_33_758 VPWR VGND sg13g2_decap_8
XFILLER_14_961 VPWR VGND sg13g2_decap_8
X_468_ net73 VGND VPWR _090_ DP_2.matrix\[16\] clknet_5_29__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_279 VPWR VGND sg13g2_decap_8
XFILLER_9_431 VPWR VGND sg13g2_decap_8
X_399_ net53 _093_ VPWR VGND sg13g2_buf_1
XFILLER_13_471 VPWR VGND sg13g2_decap_8
XFILLER_40_290 VPWR VGND sg13g2_decap_8
XFILLER_9_497 VPWR VGND sg13g2_fill_2
XFILLER_28_519 VPWR VGND sg13g2_decap_8
XFILLER_36_596 VPWR VGND sg13g2_decap_8
XFILLER_23_246 VPWR VGND sg13g2_decap_8
XFILLER_24_747 VPWR VGND sg13g2_decap_8
XFILLER_23_279 VPWR VGND sg13g2_fill_2
Xclkbuf_5_18__f_clk clknet_4_9_0_clk clknet_5_18__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_20_964 VPWR VGND sg13g2_decap_8
XFILLER_3_607 VPWR VGND sg13g2_decap_8
XFILLER_48_35 VPWR VGND sg13g2_decap_8
XFILLER_47_828 VPWR VGND sg13g2_decap_8
XFILLER_46_349 VPWR VGND sg13g2_decap_8
XFILLER_42_500 VPWR VGND sg13g2_decap_8
XFILLER_14_202 VPWR VGND sg13g2_decap_8
XFILLER_27_574 VPWR VGND sg13g2_decap_8
XFILLER_9_18 VPWR VGND sg13g2_decap_8
XFILLER_15_769 VPWR VGND sg13g2_decap_8
XFILLER_42_577 VPWR VGND sg13g2_decap_8
X_322_ _188_ net124 net87 VPWR VGND sg13g2_nand2_1
XFILLER_14_268 VPWR VGND sg13g2_decap_8
XFILLER_11_942 VPWR VGND sg13g2_decap_8
Xfanout61 net62 net61 VPWR VGND sg13g2_buf_8
Xfanout72 net74 net72 VPWR VGND sg13g2_buf_8
X_253_ _001_ _150_ _151_ VPWR VGND sg13g2_xnor2_1
XFILLER_6_401 VPWR VGND sg13g2_fill_2
XFILLER_13_60 VPWR VGND sg13g2_decap_8
XFILLER_7_968 VPWR VGND sg13g2_decap_8
XFILLER_6_467 VPWR VGND sg13g2_decap_8
XFILLER_1_150 VPWR VGND sg13g2_decap_8
XFILLER_2_662 VPWR VGND sg13g2_decap_8
XFILLER_29_7 VPWR VGND sg13g2_decap_8
XFILLER_49_154 VPWR VGND sg13g2_decap_8
XFILLER_38_817 VPWR VGND sg13g2_decap_8
XFILLER_37_349 VPWR VGND sg13g2_decap_8
XFILLER_46_883 VPWR VGND sg13g2_decap_8
XFILLER_33_555 VPWR VGND sg13g2_decap_8
XFILLER_20_238 VPWR VGND sg13g2_decap_8
XFILLER_28_316 VPWR VGND sg13g2_decap_8
XFILLER_37_861 VPWR VGND sg13g2_decap_8
XFILLER_24_544 VPWR VGND sg13g2_decap_8
Xclkload3 VPWR clkload3/Y clknet_5_15__leaf_clk VGND sg13g2_inv_1
XFILLER_7_209 VPWR VGND sg13g2_decap_8
XFILLER_20_761 VPWR VGND sg13g2_decap_8
XFILLER_4_916 VPWR VGND sg13g2_decap_8
XFILLER_8_1020 VPWR VGND sg13g2_decap_8
XFILLER_19_305 VPWR VGND sg13g2_decap_8
XFILLER_47_625 VPWR VGND sg13g2_decap_8
XFILLER_15_511 VPWR VGND sg13g2_decap_8
XFILLER_28_883 VPWR VGND sg13g2_decap_8
XFILLER_15_533 VPWR VGND sg13g2_decap_8
XFILLER_15_544 VPWR VGND sg13g2_fill_2
XFILLER_43_875 VPWR VGND sg13g2_decap_8
X_305_ _178_ net111 mac2.products_ff\[80\] VPWR VGND sg13g2_nand2_1
XFILLER_30_569 VPWR VGND sg13g2_decap_8
X_236_ net159 net120 _062_ VPWR VGND sg13g2_and2_1
XFILLER_7_765 VPWR VGND sg13g2_decap_8
XFILLER_6_253 VPWR VGND sg13g2_decap_8
XFILLER_3_971 VPWR VGND sg13g2_decap_8
XFILLER_38_614 VPWR VGND sg13g2_decap_8
XFILLER_37_102 VPWR VGND sg13g2_decap_8
XFILLER_1_63 VPWR VGND sg13g2_decap_8
XFILLER_19_861 VPWR VGND sg13g2_decap_8
XFILLER_46_680 VPWR VGND sg13g2_decap_8
XFILLER_34_820 VPWR VGND sg13g2_decap_8
XFILLER_33_363 VPWR VGND sg13g2_fill_1
XFILLER_21_525 VPWR VGND sg13g2_decap_8
XFILLER_34_897 VPWR VGND sg13g2_decap_8
XFILLER_14_1003 VPWR VGND sg13g2_decap_8
XFILLER_20_39 VPWR VGND sg13g2_decap_8
Xhold26 DP_4.matrix\[81\] VPWR VGND net50 sg13g2_dlygate4sd3_1
Xhold15 DP_4.matrix\[17\] VPWR VGND net39 sg13g2_dlygate4sd3_1
Xhold37 DP_3.matrix\[129\] VPWR VGND net87 sg13g2_dlygate4sd3_1
XFILLER_29_37 VPWR VGND sg13g2_fill_1
XFILLER_29_59 VPWR VGND sg13g2_decap_8
Xhold59 mac1.products_ff\[48\] VPWR VGND net109 sg13g2_dlygate4sd3_1
Xhold48 _004_ VPWR VGND net98 sg13g2_dlygate4sd3_1
XFILLER_29_658 VPWR VGND sg13g2_decap_8
XFILLER_45_14 VPWR VGND sg13g2_decap_8
XFILLER_25_853 VPWR VGND sg13g2_decap_8
XFILLER_12_536 VPWR VGND sg13g2_decap_8
XFILLER_40_845 VPWR VGND sg13g2_decap_8
XFILLER_4_713 VPWR VGND sg13g2_decap_8
XFILLER_10_72 VPWR VGND sg13g2_decap_8
XFILLER_3_278 VPWR VGND sg13g2_decap_8
XFILLER_48_912 VPWR VGND sg13g2_decap_8
XFILLER_0_952 VPWR VGND sg13g2_decap_8
XFILLER_47_422 VPWR VGND sg13g2_decap_8
XFILLER_19_102 VPWR VGND sg13g2_decap_8
XFILLER_48_989 VPWR VGND sg13g2_decap_8
XFILLER_19_81 VPWR VGND sg13g2_decap_8
XFILLER_47_499 VPWR VGND sg13g2_decap_8
XFILLER_35_617 VPWR VGND sg13g2_decap_8
XFILLER_16_831 VPWR VGND sg13g2_decap_8
XFILLER_28_680 VPWR VGND sg13g2_decap_8
XFILLER_43_672 VPWR VGND sg13g2_decap_8
XFILLER_31_834 VPWR VGND sg13g2_decap_8
XFILLER_7_562 VPWR VGND sg13g2_decap_8
XFILLER_44_1018 VPWR VGND sg13g2_decap_8
Xheichips25_template_17 VPWR VGND uio_oe[0] sg13g2_tiehi
XFILLER_38_422 VPWR VGND sg13g2_decap_8
XFILLER_39_956 VPWR VGND sg13g2_decap_8
XFILLER_26_628 VPWR VGND sg13g2_decap_8
XFILLER_38_477 VPWR VGND sg13g2_decap_4
XFILLER_15_39 VPWR VGND sg13g2_decap_8
XFILLER_18_190 VPWR VGND sg13g2_decap_8
XFILLER_21_300 VPWR VGND sg13g2_decap_8
XFILLER_34_694 VPWR VGND sg13g2_decap_8
XFILLER_21_344 VPWR VGND sg13g2_fill_1
XFILLER_22_856 VPWR VGND sg13g2_decap_8
XFILLER_31_49 VPWR VGND sg13g2_decap_8
XFILLER_1_738 VPWR VGND sg13g2_decap_8
XFILLER_0_259 VPWR VGND sg13g2_decap_8
XFILLER_5_1023 VPWR VGND sg13g2_decap_4
XFILLER_29_411 VPWR VGND sg13g2_fill_1
XFILLER_29_455 VPWR VGND sg13g2_decap_8
X_570_ net57 VGND VPWR _037_ mac2.products_ff\[129\] clknet_5_2__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_606 VPWR VGND sg13g2_fill_2
XFILLER_45_948 VPWR VGND sg13g2_decap_8
XFILLER_44_458 VPWR VGND sg13g2_decap_8
XFILLER_25_650 VPWR VGND sg13g2_decap_8
XFILLER_13_823 VPWR VGND sg13g2_decap_8
XFILLER_24_171 VPWR VGND sg13g2_decap_8
XFILLER_12_333 VPWR VGND sg13g2_decap_8
XFILLER_40_642 VPWR VGND sg13g2_decap_8
XFILLER_8_337 VPWR VGND sg13g2_fill_2
XFILLER_9_849 VPWR VGND sg13g2_decap_8
XFILLER_12_377 VPWR VGND sg13g2_fill_1
XFILLER_8_359 VPWR VGND sg13g2_decap_8
XFILLER_4_587 VPWR VGND sg13g2_decap_8
XFILLER_36_904 VPWR VGND sg13g2_decap_8
XFILLER_48_786 VPWR VGND sg13g2_decap_8
XFILLER_43_480 VPWR VGND sg13g2_fill_1
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
XFILLER_31_631 VPWR VGND sg13g2_decap_8
XFILLER_11_1028 VPWR VGND sg13g2_fill_1
XFILLER_7_84 VPWR VGND sg13g2_decap_8
XFILLER_39_753 VPWR VGND sg13g2_decap_8
XFILLER_26_403 VPWR VGND sg13g2_decap_4
XFILLER_26_447 VPWR VGND sg13g2_decap_8
XFILLER_27_959 VPWR VGND sg13g2_decap_8
XFILLER_35_981 VPWR VGND sg13g2_decap_8
XFILLER_22_653 VPWR VGND sg13g2_decap_8
XFILLER_34_491 VPWR VGND sg13g2_decap_8
XFILLER_10_804 VPWR VGND sg13g2_decap_8
XFILLER_21_141 VPWR VGND sg13g2_decap_8
XFILLER_1_535 VPWR VGND sg13g2_decap_8
XFILLER_49_517 VPWR VGND sg13g2_decap_8
XFILLER_29_230 VPWR VGND sg13g2_decap_8
XFILLER_17_403 VPWR VGND sg13g2_decap_8
XFILLER_18_926 VPWR VGND sg13g2_decap_8
XFILLER_45_745 VPWR VGND sg13g2_decap_8
XFILLER_29_296 VPWR VGND sg13g2_decap_8
XFILLER_44_255 VPWR VGND sg13g2_decap_8
X_553_ net75 VGND VPWR _047_ mac1.products_ff\[97\] clknet_5_25__leaf_clk sg13g2_dfrbpq_1
X_484_ net78 VGND VPWR _106_ DP_3.matrix\[0\] clknet_5_31__leaf_clk sg13g2_dfrbpq_1
XFILLER_26_992 VPWR VGND sg13g2_decap_8
XFILLER_41_940 VPWR VGND sg13g2_decap_8
XFILLER_9_646 VPWR VGND sg13g2_decap_8
XFILLER_13_697 VPWR VGND sg13g2_decap_8
XFILLER_8_156 VPWR VGND sg13g2_decap_8
XFILLER_32_81 VPWR VGND sg13g2_decap_8
XFILLER_5_841 VPWR VGND sg13g2_decap_8
XFILLER_4_395 VPWR VGND sg13g2_decap_8
XFILLER_36_701 VPWR VGND sg13g2_decap_8
XFILLER_48_583 VPWR VGND sg13g2_decap_8
XFILLER_35_200 VPWR VGND sg13g2_decap_8
XFILLER_24_929 VPWR VGND sg13g2_decap_8
XFILLER_36_778 VPWR VGND sg13g2_decap_8
XFILLER_17_992 VPWR VGND sg13g2_decap_8
XFILLER_23_406 VPWR VGND sg13g2_decap_8
XFILLER_32_995 VPWR VGND sg13g2_decap_8
XFILLER_12_18 VPWR VGND sg13g2_decap_8
Xhold101 DP_1.matrix\[96\] VPWR VGND net151 sg13g2_dlygate4sd3_1
Xhold123 mac1.sum_lvl1_ff\[24\] VPWR VGND net173 sg13g2_dlygate4sd3_1
Xhold112 DP_1.matrix\[80\] VPWR VGND net162 sg13g2_dlygate4sd3_1
Xhold134 mac2.products_ff\[48\] VPWR VGND net184 sg13g2_dlygate4sd3_1
Xhold156 _016_ VPWR VGND net206 sg13g2_dlygate4sd3_1
Xhold145 _007_ VPWR VGND net195 sg13g2_dlygate4sd3_1
XFILLER_39_550 VPWR VGND sg13g2_decap_8
XFILLER_2_1026 VPWR VGND sg13g2_fill_2
XFILLER_27_756 VPWR VGND sg13g2_decap_8
XFILLER_14_406 VPWR VGND sg13g2_decap_8
XFILLER_26_266 VPWR VGND sg13g2_fill_2
XFILLER_26_277 VPWR VGND sg13g2_decap_8
XFILLER_42_759 VPWR VGND sg13g2_decap_8
XFILLER_10_601 VPWR VGND sg13g2_decap_8
XFILLER_41_258 VPWR VGND sg13g2_decap_8
XFILLER_22_472 VPWR VGND sg13g2_decap_8
XFILLER_10_678 VPWR VGND sg13g2_decap_8
XFILLER_6_649 VPWR VGND sg13g2_decap_8
XFILLER_2_844 VPWR VGND sg13g2_decap_8
XFILLER_1_332 VPWR VGND sg13g2_decap_8
XFILLER_49_336 VPWR VGND sg13g2_decap_8
XFILLER_18_723 VPWR VGND sg13g2_decap_8
XFILLER_45_542 VPWR VGND sg13g2_decap_8
XFILLER_17_244 VPWR VGND sg13g2_decap_8
X_536_ net61 VGND VPWR net35 mac1.sum_lvl1_ff\[32\] clknet_5_5__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_214 VPWR VGND sg13g2_decap_4
XFILLER_33_737 VPWR VGND sg13g2_decap_8
XFILLER_14_940 VPWR VGND sg13g2_decap_8
XFILLER_9_410 VPWR VGND sg13g2_decap_8
X_467_ net72 VGND VPWR _089_ DP_2.matrix\[1\] clknet_5_23__leaf_clk sg13g2_dfrbpq_1
XFILLER_20_409 VPWR VGND sg13g2_decap_8
XFILLER_32_258 VPWR VGND sg13g2_decap_8
XFILLER_43_91 VPWR VGND sg13g2_decap_8
X_398_ net123 _092_ VPWR VGND sg13g2_buf_1
XFILLER_4_85 VPWR VGND sg13g2_decap_8
XFILLER_49_881 VPWR VGND sg13g2_decap_8
XFILLER_24_726 VPWR VGND sg13g2_decap_8
XFILLER_36_575 VPWR VGND sg13g2_decap_8
XFILLER_23_225 VPWR VGND sg13g2_decap_8
XFILLER_20_943 VPWR VGND sg13g2_decap_8
XFILLER_32_792 VPWR VGND sg13g2_decap_8
XFILLER_48_14 VPWR VGND sg13g2_decap_8
XFILLER_24_1027 VPWR VGND sg13g2_fill_2
XFILLER_47_807 VPWR VGND sg13g2_decap_8
XFILLER_27_553 VPWR VGND sg13g2_decap_8
XFILLER_42_556 VPWR VGND sg13g2_decap_8
XFILLER_15_748 VPWR VGND sg13g2_decap_8
X_321_ _187_ _186_ _035_ VPWR VGND sg13g2_xor2_1
XFILLER_11_921 VPWR VGND sg13g2_decap_8
X_252_ mac1.products_ff\[17\] mac1.products_ff\[1\] _151_ VPWR VGND sg13g2_xor2_1
Xfanout73 net74 net73 VPWR VGND sg13g2_buf_8
Xfanout62 rst_n net62 VPWR VGND sg13g2_buf_8
XFILLER_31_1009 VPWR VGND sg13g2_decap_8
XFILLER_10_486 VPWR VGND sg13g2_decap_8
XFILLER_7_947 VPWR VGND sg13g2_decap_8
XFILLER_11_998 VPWR VGND sg13g2_decap_8
XFILLER_2_641 VPWR VGND sg13g2_decap_8
XFILLER_49_133 VPWR VGND sg13g2_decap_8
XFILLER_37_328 VPWR VGND sg13g2_decap_8
XFILLER_46_862 VPWR VGND sg13g2_decap_8
Xclkbuf_5_24__f_clk clknet_4_12_0_clk clknet_5_24__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_33_534 VPWR VGND sg13g2_decap_8
X_519_ net57 VGND VPWR _141_ DP_4.matrix\[129\] clknet_5_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_21_729 VPWR VGND sg13g2_decap_8
XFILLER_20_217 VPWR VGND sg13g2_decap_8
XFILLER_48_0 VPWR VGND sg13g2_decap_8
XFILLER_18_39 VPWR VGND sg13g2_fill_1
XFILLER_28_339 VPWR VGND sg13g2_fill_1
XFILLER_37_840 VPWR VGND sg13g2_decap_8
XFILLER_24_523 VPWR VGND sg13g2_decap_8
XFILLER_36_383 VPWR VGND sg13g2_decap_8
XFILLER_24_567 VPWR VGND sg13g2_fill_2
Xclkload4 clknet_5_17__leaf_clk clkload4/X VPWR VGND sg13g2_buf_1
XFILLER_20_740 VPWR VGND sg13g2_decap_8
XFILLER_47_604 VPWR VGND sg13g2_decap_8
XFILLER_46_169 VPWR VGND sg13g2_decap_8
XFILLER_28_862 VPWR VGND sg13g2_decap_8
XFILLER_43_854 VPWR VGND sg13g2_decap_8
XFILLER_42_364 VPWR VGND sg13g2_decap_8
X_304_ net113 mac2.products_ff\[96\] _023_ VPWR VGND sg13g2_xor2_1
XFILLER_30_548 VPWR VGND sg13g2_decap_8
X_235_ net134 net141 _060_ VPWR VGND sg13g2_and2_1
XFILLER_10_261 VPWR VGND sg13g2_fill_2
XFILLER_10_250 VPWR VGND sg13g2_decap_8
XFILLER_7_744 VPWR VGND sg13g2_decap_8
XFILLER_6_232 VPWR VGND sg13g2_decap_8
XFILLER_11_795 VPWR VGND sg13g2_decap_8
XFILLER_40_81 VPWR VGND sg13g2_decap_8
XFILLER_3_950 VPWR VGND sg13g2_decap_8
XFILLER_41_7 VPWR VGND sg13g2_decap_8
XFILLER_1_42 VPWR VGND sg13g2_decap_8
XFILLER_19_840 VPWR VGND sg13g2_decap_8
XFILLER_37_147 VPWR VGND sg13g2_fill_2
XFILLER_45_180 VPWR VGND sg13g2_decap_8
XFILLER_33_320 VPWR VGND sg13g2_decap_8
XFILLER_34_876 VPWR VGND sg13g2_decap_8
XFILLER_20_18 VPWR VGND sg13g2_decap_8
Xhold38 DP_2.matrix\[113\] VPWR VGND net88 sg13g2_dlygate4sd3_1
Xhold16 DP_1.matrix\[17\] VPWR VGND net40 sg13g2_dlygate4sd3_1
XFILLER_29_49 VPWR VGND sg13g2_fill_1
Xhold27 DP_4.matrix\[1\] VPWR VGND net51 sg13g2_dlygate4sd3_1
Xhold49 DP_3.matrix\[33\] VPWR VGND net99 sg13g2_dlygate4sd3_1
XFILLER_28_114 VPWR VGND sg13g2_decap_8
XFILLER_29_637 VPWR VGND sg13g2_decap_8
XFILLER_16_309 VPWR VGND sg13g2_decap_8
XFILLER_28_169 VPWR VGND sg13g2_decap_8
XFILLER_45_48 VPWR VGND sg13g2_decap_4
XFILLER_43_128 VPWR VGND sg13g2_decap_8
XFILLER_25_832 VPWR VGND sg13g2_decap_8
XFILLER_36_180 VPWR VGND sg13g2_decap_8
XFILLER_12_515 VPWR VGND sg13g2_decap_8
XFILLER_24_397 VPWR VGND sg13g2_decap_8
XFILLER_40_824 VPWR VGND sg13g2_decap_8
XFILLER_10_51 VPWR VGND sg13g2_decap_8
XFILLER_4_769 VPWR VGND sg13g2_decap_8
XFILLER_3_257 VPWR VGND sg13g2_decap_8
XFILLER_0_931 VPWR VGND sg13g2_decap_8
XFILLER_47_401 VPWR VGND sg13g2_decap_8
XFILLER_48_968 VPWR VGND sg13g2_decap_8
XFILLER_19_60 VPWR VGND sg13g2_decap_8
XFILLER_47_478 VPWR VGND sg13g2_decap_8
XFILLER_16_810 VPWR VGND sg13g2_decap_8
XFILLER_27_180 VPWR VGND sg13g2_decap_8
XFILLER_43_651 VPWR VGND sg13g2_decap_8
XFILLER_15_342 VPWR VGND sg13g2_decap_8
XFILLER_37_1015 VPWR VGND sg13g2_decap_8
XFILLER_16_887 VPWR VGND sg13g2_decap_8
XFILLER_31_813 VPWR VGND sg13g2_decap_8
XFILLER_30_389 VPWR VGND sg13g2_decap_8
XFILLER_7_541 VPWR VGND sg13g2_decap_8
Xheichips25_template_18 VPWR VGND uio_oe[1] sg13g2_tiehi
XFILLER_39_935 VPWR VGND sg13g2_decap_8
XFILLER_26_607 VPWR VGND sg13g2_decap_8
XFILLER_25_139 VPWR VGND sg13g2_decap_8
XFILLER_15_18 VPWR VGND sg13g2_decap_8
XFILLER_22_835 VPWR VGND sg13g2_decap_8
XFILLER_34_673 VPWR VGND sg13g2_decap_8
XFILLER_31_28 VPWR VGND sg13g2_decap_8
XFILLER_1_717 VPWR VGND sg13g2_decap_8
XFILLER_0_238 VPWR VGND sg13g2_decap_8
XFILLER_5_1002 VPWR VGND sg13g2_decap_8
XFILLER_29_434 VPWR VGND sg13g2_decap_8
XFILLER_45_927 VPWR VGND sg13g2_decap_8
XFILLER_44_437 VPWR VGND sg13g2_decap_8
XFILLER_13_802 VPWR VGND sg13g2_decap_8
XFILLER_12_312 VPWR VGND sg13g2_decap_8
XFILLER_24_150 VPWR VGND sg13g2_decap_8
XFILLER_40_621 VPWR VGND sg13g2_decap_8
XFILLER_8_316 VPWR VGND sg13g2_decap_8
XFILLER_9_828 VPWR VGND sg13g2_decap_8
XFILLER_13_879 VPWR VGND sg13g2_decap_8
XFILLER_21_890 VPWR VGND sg13g2_decap_8
XFILLER_40_698 VPWR VGND sg13g2_decap_8
XFILLER_4_533 VPWR VGND sg13g2_fill_1
XFILLER_21_72 VPWR VGND sg13g2_decap_8
XFILLER_4_566 VPWR VGND sg13g2_decap_8
XFILLER_48_765 VPWR VGND sg13g2_decap_8
XFILLER_47_297 VPWR VGND sg13g2_decap_8
XFILLER_16_684 VPWR VGND sg13g2_decap_8
XFILLER_31_610 VPWR VGND sg13g2_decap_8
XFILLER_15_172 VPWR VGND sg13g2_decap_8
XFILLER_31_687 VPWR VGND sg13g2_decap_8
XFILLER_7_63 VPWR VGND sg13g2_decap_8
XFILLER_8_894 VPWR VGND sg13g2_decap_8
XFILLER_7_371 VPWR VGND sg13g2_decap_8
XFILLER_30_0 VPWR VGND sg13g2_decap_8
XFILLER_39_732 VPWR VGND sg13g2_decap_8
XFILLER_26_39 VPWR VGND sg13g2_decap_8
XFILLER_26_426 VPWR VGND sg13g2_decap_8
XFILLER_27_938 VPWR VGND sg13g2_decap_8
XFILLER_35_960 VPWR VGND sg13g2_decap_8
XFILLER_34_470 VPWR VGND sg13g2_decap_8
XFILLER_41_407 VPWR VGND sg13g2_fill_1
XFILLER_21_120 VPWR VGND sg13g2_decap_8
XFILLER_22_632 VPWR VGND sg13g2_decap_8
XFILLER_42_49 VPWR VGND sg13g2_decap_8
XFILLER_21_175 VPWR VGND sg13g2_decap_8
XFILLER_1_514 VPWR VGND sg13g2_decap_8
Xclkbuf_5_5__f_clk clknet_4_2_0_clk clknet_5_5__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_18_905 VPWR VGND sg13g2_decap_8
XFILLER_45_724 VPWR VGND sg13g2_decap_8
XFILLER_44_234 VPWR VGND sg13g2_decap_8
X_552_ net75 VGND VPWR _046_ mac1.products_ff\[96\] clknet_5_25__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_919 VPWR VGND sg13g2_decap_8
X_483_ net59 VGND VPWR _105_ DP_2.matrix\[129\] clknet_5_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_26_971 VPWR VGND sg13g2_decap_8
XFILLER_16_83 VPWR VGND sg13g2_decap_4
XFILLER_9_625 VPWR VGND sg13g2_decap_8
XFILLER_8_102 VPWR VGND sg13g2_decap_8
XFILLER_13_676 VPWR VGND sg13g2_decap_8
XFILLER_40_451 VPWR VGND sg13g2_decap_4
XFILLER_40_495 VPWR VGND sg13g2_decap_8
XFILLER_41_996 VPWR VGND sg13g2_decap_8
XFILLER_12_197 VPWR VGND sg13g2_decap_8
XFILLER_5_820 VPWR VGND sg13g2_decap_8
XFILLER_5_897 VPWR VGND sg13g2_decap_8
XFILLER_4_374 VPWR VGND sg13g2_decap_8
XFILLER_48_562 VPWR VGND sg13g2_decap_8
XFILLER_24_908 VPWR VGND sg13g2_decap_8
XFILLER_35_256 VPWR VGND sg13g2_decap_8
XFILLER_36_757 VPWR VGND sg13g2_decap_8
XFILLER_17_971 VPWR VGND sg13g2_decap_8
XFILLER_16_492 VPWR VGND sg13g2_decap_8
XFILLER_31_440 VPWR VGND sg13g2_decap_4
XFILLER_32_974 VPWR VGND sg13g2_decap_8
XFILLER_8_691 VPWR VGND sg13g2_decap_8
Xhold113 DP_3.matrix\[32\] VPWR VGND net163 sg13g2_dlygate4sd3_1
Xhold124 _011_ VPWR VGND net174 sg13g2_dlygate4sd3_1
Xhold102 mac2.sum_lvl2_ff\[0\] VPWR VGND net152 sg13g2_dlygate4sd3_1
Xhold135 _020_ VPWR VGND net185 sg13g2_dlygate4sd3_1
Xhold157 mac2.sum_lvl3_ff\[0\] VPWR VGND net207 sg13g2_dlygate4sd3_1
Xhold146 mac2.sum_lvl2_ff\[4\] VPWR VGND net196 sg13g2_dlygate4sd3_1
XFILLER_2_1005 VPWR VGND sg13g2_decap_8
XFILLER_37_49 VPWR VGND sg13g2_decap_8
XFILLER_27_735 VPWR VGND sg13g2_decap_8
XFILLER_26_245 VPWR VGND sg13g2_decap_8
XFILLER_42_738 VPWR VGND sg13g2_decap_8
XFILLER_41_237 VPWR VGND sg13g2_decap_8
XFILLER_22_451 VPWR VGND sg13g2_decap_8
XFILLER_23_985 VPWR VGND sg13g2_decap_8
XFILLER_10_657 VPWR VGND sg13g2_decap_8
XFILLER_6_628 VPWR VGND sg13g2_decap_8
XFILLER_5_149 VPWR VGND sg13g2_decap_8
XFILLER_2_823 VPWR VGND sg13g2_decap_8
XFILLER_1_311 VPWR VGND sg13g2_decap_8
XFILLER_49_315 VPWR VGND sg13g2_decap_8
XFILLER_1_388 VPWR VGND sg13g2_decap_8
XFILLER_18_702 VPWR VGND sg13g2_decap_8
XFILLER_45_521 VPWR VGND sg13g2_decap_8
XFILLER_17_223 VPWR VGND sg13g2_decap_8
XFILLER_18_779 VPWR VGND sg13g2_decap_8
X_535_ net70 VGND VPWR net195 mac1.sum_lvl1_ff\[25\] clknet_5_25__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_716 VPWR VGND sg13g2_decap_8
XFILLER_45_598 VPWR VGND sg13g2_decap_8
X_466_ net72 VGND VPWR _088_ DP_2.matrix\[0\] clknet_5_21__leaf_clk sg13g2_dfrbpq_1
XFILLER_43_70 VPWR VGND sg13g2_decap_8
XFILLER_14_996 VPWR VGND sg13g2_decap_8
X_397_ net49 _091_ VPWR VGND sg13g2_buf_1
XFILLER_41_793 VPWR VGND sg13g2_decap_8
XFILLER_9_477 VPWR VGND sg13g2_fill_1
XFILLER_9_466 VPWR VGND sg13g2_decap_8
Xheichips25_template_5 VPWR VGND uio_out[0] sg13g2_tielo
XFILLER_5_694 VPWR VGND sg13g2_decap_8
XFILLER_4_64 VPWR VGND sg13g2_decap_8
XFILLER_49_860 VPWR VGND sg13g2_decap_8
XFILLER_36_554 VPWR VGND sg13g2_decap_8
XFILLER_23_204 VPWR VGND sg13g2_decap_8
XFILLER_24_705 VPWR VGND sg13g2_decap_8
XFILLER_17_1013 VPWR VGND sg13g2_decap_8
XFILLER_20_922 VPWR VGND sg13g2_decap_8
XFILLER_32_771 VPWR VGND sg13g2_decap_8
XFILLER_31_292 VPWR VGND sg13g2_decap_8
XFILLER_20_999 VPWR VGND sg13g2_decap_8
XFILLER_24_1006 VPWR VGND sg13g2_decap_8
XFILLER_46_307 VPWR VGND sg13g2_fill_1
XFILLER_27_532 VPWR VGND sg13g2_decap_8
XFILLER_15_727 VPWR VGND sg13g2_decap_8
XFILLER_42_535 VPWR VGND sg13g2_decap_8
X_320_ _187_ net125 net41 VPWR VGND sg13g2_nand2_1
XFILLER_11_900 VPWR VGND sg13g2_decap_8
X_251_ _150_ net178 net126 VPWR VGND sg13g2_nand2_1
Xfanout74 net75 net74 VPWR VGND sg13g2_buf_8
XFILLER_23_782 VPWR VGND sg13g2_decap_8
Xfanout63 net64 net63 VPWR VGND sg13g2_buf_8
XFILLER_7_926 VPWR VGND sg13g2_decap_8
XFILLER_11_977 VPWR VGND sg13g2_decap_8
XFILLER_6_414 VPWR VGND sg13g2_decap_8
XFILLER_2_620 VPWR VGND sg13g2_decap_8
XFILLER_1_130 VPWR VGND sg13g2_fill_2
XFILLER_49_112 VPWR VGND sg13g2_decap_8
XFILLER_1_185 VPWR VGND sg13g2_decap_8
XFILLER_2_697 VPWR VGND sg13g2_decap_8
XFILLER_49_189 VPWR VGND sg13g2_decap_8
XFILLER_46_841 VPWR VGND sg13g2_decap_8
XFILLER_18_554 VPWR VGND sg13g2_decap_8
XFILLER_33_513 VPWR VGND sg13g2_decap_8
XFILLER_45_395 VPWR VGND sg13g2_decap_8
XFILLER_18_598 VPWR VGND sg13g2_decap_8
X_518_ net57 VGND VPWR _140_ DP_4.matrix\[128\] clknet_5_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_21_708 VPWR VGND sg13g2_decap_8
X_449_ net72 VGND VPWR _071_ DP_1.matrix\[1\] clknet_5_21__leaf_clk sg13g2_dfrbpq_1
XFILLER_14_793 VPWR VGND sg13g2_decap_8
XFILLER_41_590 VPWR VGND sg13g2_decap_8
XFILLER_47_1028 VPWR VGND sg13g2_fill_1
XFILLER_47_1017 VPWR VGND sg13g2_decap_8
XFILLER_6_992 VPWR VGND sg13g2_decap_8
XFILLER_29_819 VPWR VGND sg13g2_decap_8
XFILLER_18_18 VPWR VGND sg13g2_decap_8
XFILLER_24_502 VPWR VGND sg13g2_decap_8
XFILLER_36_362 VPWR VGND sg13g2_decap_8
XFILLER_37_896 VPWR VGND sg13g2_decap_8
XFILLER_12_719 VPWR VGND sg13g2_decap_8
Xclkload5 clknet_5_19__leaf_clk clkload5/X VPWR VGND sg13g2_buf_1
XFILLER_30_1010 VPWR VGND sg13g2_decap_8
XFILLER_20_796 VPWR VGND sg13g2_decap_8
XFILLER_3_406 VPWR VGND sg13g2_decap_4
Xclkbuf_5_30__f_clk clknet_4_15_0_clk clknet_5_30__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_46_148 VPWR VGND sg13g2_decap_8
XFILLER_28_841 VPWR VGND sg13g2_decap_8
XFILLER_43_833 VPWR VGND sg13g2_decap_8
XFILLER_42_343 VPWR VGND sg13g2_decap_8
XFILLER_42_387 VPWR VGND sg13g2_decap_8
XFILLER_24_50 VPWR VGND sg13g2_decap_8
X_303_ _024_ _176_ _177_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_527 VPWR VGND sg13g2_decap_8
X_234_ net119 net150 _058_ VPWR VGND sg13g2_and2_1
XFILLER_7_723 VPWR VGND sg13g2_decap_8
XFILLER_11_774 VPWR VGND sg13g2_decap_8
XFILLER_6_211 VPWR VGND sg13g2_decap_8
XFILLER_40_60 VPWR VGND sg13g2_decap_8
XFILLER_6_288 VPWR VGND sg13g2_decap_8
XFILLER_34_7 VPWR VGND sg13g2_decap_8
XFILLER_49_91 VPWR VGND sg13g2_decap_8
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_37_126 VPWR VGND sg13g2_decap_8
XFILLER_38_649 VPWR VGND sg13g2_decap_8
XFILLER_1_98 VPWR VGND sg13g2_decap_8
XFILLER_18_340 VPWR VGND sg13g2_decap_4
XFILLER_19_896 VPWR VGND sg13g2_decap_8
XFILLER_34_855 VPWR VGND sg13g2_decap_8
XFILLER_33_398 VPWR VGND sg13g2_decap_8
Xhold28 DP_3.matrix\[81\] VPWR VGND net52 sg13g2_dlygate4sd3_1
Xhold17 DP_4.matrix\[113\] VPWR VGND net41 sg13g2_dlygate4sd3_1
XFILLER_29_28 VPWR VGND sg13g2_decap_8
XFILLER_21_1009 VPWR VGND sg13g2_decap_8
XFILLER_29_616 VPWR VGND sg13g2_decap_8
Xhold39 DP_1.matrix\[81\] VPWR VGND net89 sg13g2_dlygate4sd3_1
XFILLER_44_619 VPWR VGND sg13g2_decap_8
XFILLER_25_811 VPWR VGND sg13g2_decap_8
XFILLER_37_693 VPWR VGND sg13g2_decap_8
XFILLER_40_803 VPWR VGND sg13g2_decap_8
XFILLER_24_376 VPWR VGND sg13g2_decap_8
XFILLER_25_888 VPWR VGND sg13g2_decap_8
XFILLER_20_560 VPWR VGND sg13g2_decap_8
XFILLER_20_593 VPWR VGND sg13g2_decap_8
XFILLER_4_748 VPWR VGND sg13g2_decap_8
XFILLER_3_236 VPWR VGND sg13g2_decap_8
XFILLER_0_910 VPWR VGND sg13g2_decap_8
XFILLER_0_987 VPWR VGND sg13g2_decap_8
XFILLER_48_947 VPWR VGND sg13g2_decap_8
XFILLER_19_137 VPWR VGND sg13g2_decap_8
XFILLER_47_457 VPWR VGND sg13g2_decap_8
XFILLER_43_630 VPWR VGND sg13g2_decap_8
XFILLER_16_866 VPWR VGND sg13g2_decap_8
XFILLER_42_140 VPWR VGND sg13g2_decap_8
XFILLER_42_184 VPWR VGND sg13g2_decap_8
XFILLER_15_398 VPWR VGND sg13g2_decap_8
XFILLER_30_335 VPWR VGND sg13g2_decap_8
XFILLER_31_869 VPWR VGND sg13g2_decap_8
XFILLER_30_368 VPWR VGND sg13g2_decap_8
XFILLER_7_520 VPWR VGND sg13g2_decap_8
XFILLER_7_597 VPWR VGND sg13g2_decap_8
Xheichips25_template_19 VPWR VGND uio_oe[2] sg13g2_tiehi
XFILLER_39_914 VPWR VGND sg13g2_decap_8
XFILLER_20_1020 VPWR VGND sg13g2_decap_8
XFILLER_19_693 VPWR VGND sg13g2_decap_8
XFILLER_34_652 VPWR VGND sg13g2_decap_8
XFILLER_22_814 VPWR VGND sg13g2_decap_8
XFILLER_30_891 VPWR VGND sg13g2_decap_8
XFILLER_0_217 VPWR VGND sg13g2_decap_8
XFILLER_45_906 VPWR VGND sg13g2_decap_8
XFILLER_44_416 VPWR VGND sg13g2_decap_8
XFILLER_37_490 VPWR VGND sg13g2_decap_8
XFILLER_25_685 VPWR VGND sg13g2_decap_8
XFILLER_40_600 VPWR VGND sg13g2_decap_8
XFILLER_9_807 VPWR VGND sg13g2_decap_8
XFILLER_13_858 VPWR VGND sg13g2_decap_8
XFILLER_12_368 VPWR VGND sg13g2_decap_8
XFILLER_40_677 VPWR VGND sg13g2_decap_8
XFILLER_4_512 VPWR VGND sg13g2_decap_8
XFILLER_21_51 VPWR VGND sg13g2_decap_8
XFILLER_4_545 VPWR VGND sg13g2_decap_8
XFILLER_48_744 VPWR VGND sg13g2_decap_8
XFILLER_0_784 VPWR VGND sg13g2_decap_8
XFILLER_47_232 VPWR VGND sg13g2_decap_8
XFILLER_47_276 VPWR VGND sg13g2_decap_8
XFILLER_29_980 VPWR VGND sg13g2_decap_8
XFILLER_36_939 VPWR VGND sg13g2_decap_8
XFILLER_35_449 VPWR VGND sg13g2_decap_8
XFILLER_44_983 VPWR VGND sg13g2_decap_8
XFILLER_43_471 VPWR VGND sg13g2_decap_8
XFILLER_15_151 VPWR VGND sg13g2_decap_8
XFILLER_16_663 VPWR VGND sg13g2_decap_8
XFILLER_31_666 VPWR VGND sg13g2_decap_8
XFILLER_12_880 VPWR VGND sg13g2_decap_8
XFILLER_8_873 VPWR VGND sg13g2_decap_8
XFILLER_7_42 VPWR VGND sg13g2_decap_8
XFILLER_11_1019 VPWR VGND sg13g2_decap_8
XFILLER_39_711 VPWR VGND sg13g2_decap_8
XFILLER_27_917 VPWR VGND sg13g2_decap_8
XFILLER_39_788 VPWR VGND sg13g2_decap_8
XFILLER_26_18 VPWR VGND sg13g2_decap_8
XFILLER_19_490 VPWR VGND sg13g2_decap_8
XFILLER_22_611 VPWR VGND sg13g2_decap_8
XFILLER_42_28 VPWR VGND sg13g2_decap_8
XFILLER_10_839 VPWR VGND sg13g2_decap_8
XFILLER_22_688 VPWR VGND sg13g2_decap_8
XFILLER_5_309 VPWR VGND sg13g2_decap_8
XFILLER_27_1015 VPWR VGND sg13g2_decap_8
XFILLER_45_703 VPWR VGND sg13g2_decap_8
XFILLER_44_213 VPWR VGND sg13g2_decap_8
X_551_ net72 VGND VPWR _043_ mac1.products_ff\[1\] clknet_5_23__leaf_clk sg13g2_dfrbpq_1
XFILLER_29_265 VPWR VGND sg13g2_decap_8
XFILLER_17_438 VPWR VGND sg13g2_decap_8
XFILLER_26_950 VPWR VGND sg13g2_decap_8
X_482_ net59 VGND VPWR _104_ DP_2.matrix\[128\] clknet_5_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_13_600 VPWR VGND sg13g2_decap_4
XFILLER_16_62 VPWR VGND sg13g2_decap_8
XFILLER_25_471 VPWR VGND sg13g2_fill_2
XFILLER_25_482 VPWR VGND sg13g2_decap_8
XFILLER_9_604 VPWR VGND sg13g2_decap_8
XFILLER_13_655 VPWR VGND sg13g2_decap_8
XFILLER_40_430 VPWR VGND sg13g2_decap_8
XFILLER_41_975 VPWR VGND sg13g2_decap_8
XFILLER_12_176 VPWR VGND sg13g2_decap_8
XFILLER_40_474 VPWR VGND sg13g2_decap_8
XFILLER_5_876 VPWR VGND sg13g2_decap_8
XFILLER_4_353 VPWR VGND sg13g2_decap_8
XFILLER_0_581 VPWR VGND sg13g2_decap_8
XFILLER_48_541 VPWR VGND sg13g2_decap_8
XFILLER_36_736 VPWR VGND sg13g2_decap_8
XFILLER_17_950 VPWR VGND sg13g2_decap_8
XFILLER_35_235 VPWR VGND sg13g2_decap_8
XFILLER_44_780 VPWR VGND sg13g2_decap_8
XFILLER_16_471 VPWR VGND sg13g2_decap_8
XFILLER_32_953 VPWR VGND sg13g2_decap_8
XFILLER_8_670 VPWR VGND sg13g2_decap_8
Xhold114 DP_1.matrix\[48\] VPWR VGND net164 sg13g2_dlygate4sd3_1
Xhold103 _029_ VPWR VGND net153 sg13g2_dlygate4sd3_1
Xhold125 mac2.products_ff\[81\] VPWR VGND net175 sg13g2_dlygate4sd3_1
Xhold158 _033_ VPWR VGND net208 sg13g2_dlygate4sd3_1
Xhold147 _030_ VPWR VGND net197 sg13g2_dlygate4sd3_1
Xhold136 mac2.sum_lvl1_ff\[24\] VPWR VGND net186 sg13g2_dlygate4sd3_1
XFILLER_2_1028 VPWR VGND sg13g2_fill_1
XFILLER_27_714 VPWR VGND sg13g2_decap_8
XFILLER_39_585 VPWR VGND sg13g2_decap_8
XFILLER_15_909 VPWR VGND sg13g2_decap_8
XFILLER_26_224 VPWR VGND sg13g2_decap_8
XFILLER_42_717 VPWR VGND sg13g2_decap_8
XFILLER_26_268 VPWR VGND sg13g2_fill_1
XFILLER_41_216 VPWR VGND sg13g2_decap_8
XFILLER_23_964 VPWR VGND sg13g2_decap_8
XFILLER_10_636 VPWR VGND sg13g2_decap_8
XFILLER_6_607 VPWR VGND sg13g2_decap_8
XFILLER_5_128 VPWR VGND sg13g2_decap_8
XFILLER_2_802 VPWR VGND sg13g2_decap_8
XFILLER_2_879 VPWR VGND sg13g2_decap_8
XFILLER_1_367 VPWR VGND sg13g2_decap_8
XFILLER_45_500 VPWR VGND sg13g2_decap_8
XFILLER_17_202 VPWR VGND sg13g2_decap_8
XFILLER_18_758 VPWR VGND sg13g2_decap_8
XFILLER_27_72 VPWR VGND sg13g2_decap_4
XFILLER_45_577 VPWR VGND sg13g2_decap_8
X_534_ net70 VGND VPWR net38 mac1.sum_lvl1_ff\[24\] clknet_5_18__leaf_clk sg13g2_dfrbpq_1
X_465_ net56 VGND VPWR _087_ DP_1.matrix\[129\] clknet_5_4__leaf_clk sg13g2_dfrbpq_1
XFILLER_14_975 VPWR VGND sg13g2_decap_8
XFILLER_13_485 VPWR VGND sg13g2_decap_8
X_396_ net135 _090_ VPWR VGND sg13g2_buf_1
XFILLER_40_271 VPWR VGND sg13g2_fill_2
XFILLER_41_772 VPWR VGND sg13g2_decap_8
XFILLER_9_445 VPWR VGND sg13g2_decap_8
Xheichips25_template_6 VPWR VGND uio_out[1] sg13g2_tielo
XFILLER_5_673 VPWR VGND sg13g2_decap_8
XFILLER_4_172 VPWR VGND sg13g2_decap_4
XFILLER_4_43 VPWR VGND sg13g2_decap_8
XFILLER_4_32 VPWR VGND sg13g2_decap_8
XFILLER_36_533 VPWR VGND sg13g2_decap_8
XFILLER_20_901 VPWR VGND sg13g2_decap_8
XFILLER_32_750 VPWR VGND sg13g2_decap_8
XFILLER_20_978 VPWR VGND sg13g2_decap_8
XFILLER_2_109 VPWR VGND sg13g2_decap_8
XFILLER_48_49 VPWR VGND sg13g2_decap_8
XFILLER_27_511 VPWR VGND sg13g2_decap_8
XFILLER_15_706 VPWR VGND sg13g2_decap_8
XFILLER_42_514 VPWR VGND sg13g2_decap_8
XFILLER_14_216 VPWR VGND sg13g2_decap_8
XFILLER_27_588 VPWR VGND sg13g2_decap_8
XFILLER_30_709 VPWR VGND sg13g2_decap_8
XFILLER_10_411 VPWR VGND sg13g2_decap_8
X_250_ mac2.total_sum\[0\] mac1.total_sum\[0\] net1 VPWR VGND sg13g2_xor2_1
XFILLER_23_761 VPWR VGND sg13g2_decap_8
Xfanout64 net68 net64 VPWR VGND sg13g2_buf_8
XFILLER_7_905 VPWR VGND sg13g2_decap_8
XFILLER_11_956 VPWR VGND sg13g2_decap_8
Xfanout75 net81 net75 VPWR VGND sg13g2_buf_8
XFILLER_10_466 VPWR VGND sg13g2_fill_2
XFILLER_13_74 VPWR VGND sg13g2_decap_8
XFILLER_2_676 VPWR VGND sg13g2_decap_8
XFILLER_1_164 VPWR VGND sg13g2_decap_8
XFILLER_49_168 VPWR VGND sg13g2_decap_8
XFILLER_46_820 VPWR VGND sg13g2_decap_8
XFILLER_38_71 VPWR VGND sg13g2_decap_8
XFILLER_18_544 VPWR VGND sg13g2_fill_1
XFILLER_45_363 VPWR VGND sg13g2_fill_2
XFILLER_46_897 VPWR VGND sg13g2_decap_8
XFILLER_45_374 VPWR VGND sg13g2_decap_8
X_517_ net64 VGND VPWR _139_ DP_4.matrix\[113\] clknet_5_3__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_569 VPWR VGND sg13g2_decap_8
X_448_ net72 VGND VPWR _070_ DP_1.matrix\[0\] clknet_5_21__leaf_clk sg13g2_dfrbpq_1
XFILLER_14_772 VPWR VGND sg13g2_decap_8
XFILLER_13_282 VPWR VGND sg13g2_decap_8
X_379_ net40 _073_ VPWR VGND sg13g2_buf_1
XFILLER_9_264 VPWR VGND sg13g2_decap_8
XFILLER_6_971 VPWR VGND sg13g2_decap_8
XFILLER_5_492 VPWR VGND sg13g2_decap_8
XFILLER_37_875 VPWR VGND sg13g2_decap_8
Xclkload6 VPWR clkload6/Y clknet_5_23__leaf_clk VGND sg13g2_inv_1
XFILLER_20_775 VPWR VGND sg13g2_decap_8
XFILLER_47_639 VPWR VGND sg13g2_decap_8
XFILLER_19_319 VPWR VGND sg13g2_decap_8
XFILLER_46_127 VPWR VGND sg13g2_decap_8
XFILLER_28_820 VPWR VGND sg13g2_decap_8
XFILLER_43_812 VPWR VGND sg13g2_decap_8
XFILLER_28_897 VPWR VGND sg13g2_decap_8
XFILLER_42_322 VPWR VGND sg13g2_decap_8
XFILLER_43_889 VPWR VGND sg13g2_decap_8
X_302_ mac2.products_ff\[113\] mac2.products_ff\[97\] _177_ VPWR VGND sg13g2_xor2_1
XFILLER_30_506 VPWR VGND sg13g2_decap_8
X_233_ net128 net135 _056_ VPWR VGND sg13g2_and2_1
XFILLER_7_702 VPWR VGND sg13g2_decap_8
XFILLER_11_753 VPWR VGND sg13g2_decap_8
XFILLER_7_779 VPWR VGND sg13g2_decap_8
XFILLER_6_267 VPWR VGND sg13g2_decap_8
XFILLER_3_985 VPWR VGND sg13g2_decap_8
XFILLER_2_451 VPWR VGND sg13g2_decap_8
XFILLER_49_70 VPWR VGND sg13g2_decap_8
XFILLER_27_7 VPWR VGND sg13g2_decap_8
XFILLER_38_628 VPWR VGND sg13g2_decap_8
XFILLER_1_77 VPWR VGND sg13g2_decap_8
XFILLER_18_352 VPWR VGND sg13g2_fill_1
XFILLER_19_875 VPWR VGND sg13g2_decap_8
XFILLER_37_149 VPWR VGND sg13g2_fill_1
XFILLER_46_694 VPWR VGND sg13g2_decap_8
XFILLER_34_834 VPWR VGND sg13g2_decap_8
XFILLER_33_377 VPWR VGND sg13g2_decap_8
XFILLER_14_591 VPWR VGND sg13g2_decap_8
XFILLER_21_539 VPWR VGND sg13g2_decap_4
XFILLER_14_1017 VPWR VGND sg13g2_decap_8
XFILLER_14_1028 VPWR VGND sg13g2_fill_1
Xhold29 DP_2.matrix\[33\] VPWR VGND net53 sg13g2_dlygate4sd3_1
Xhold18 DP_3.matrix\[49\] VPWR VGND net42 sg13g2_dlygate4sd3_1
XFILLER_45_28 VPWR VGND sg13g2_decap_8
XFILLER_37_672 VPWR VGND sg13g2_decap_8
XFILLER_24_344 VPWR VGND sg13g2_decap_8
XFILLER_25_867 VPWR VGND sg13g2_decap_8
XFILLER_24_355 VPWR VGND sg13g2_fill_1
XFILLER_40_859 VPWR VGND sg13g2_decap_8
XFILLER_4_727 VPWR VGND sg13g2_decap_8
XFILLER_10_86 VPWR VGND sg13g2_decap_8
XFILLER_0_966 VPWR VGND sg13g2_decap_8
XFILLER_48_926 VPWR VGND sg13g2_decap_8
XFILLER_47_436 VPWR VGND sg13g2_decap_8
XFILLER_19_116 VPWR VGND sg13g2_decap_8
XFILLER_19_95 VPWR VGND sg13g2_decap_8
XFILLER_28_694 VPWR VGND sg13g2_decap_8
XFILLER_34_119 VPWR VGND sg13g2_decap_8
XFILLER_16_845 VPWR VGND sg13g2_decap_8
XFILLER_43_686 VPWR VGND sg13g2_decap_8
XFILLER_42_163 VPWR VGND sg13g2_decap_8
XFILLER_15_377 VPWR VGND sg13g2_decap_8
XFILLER_35_72 VPWR VGND sg13g2_decap_8
XFILLER_35_83 VPWR VGND sg13g2_fill_2
XFILLER_31_848 VPWR VGND sg13g2_decap_8
XFILLER_11_561 VPWR VGND sg13g2_fill_2
XFILLER_7_576 VPWR VGND sg13g2_decap_8
XFILLER_3_782 VPWR VGND sg13g2_decap_8
XFILLER_25_4 VPWR VGND sg13g2_decap_8
XFILLER_38_436 VPWR VGND sg13g2_decap_8
XFILLER_19_672 VPWR VGND sg13g2_decap_8
XFILLER_25_108 VPWR VGND sg13g2_decap_8
XFILLER_46_491 VPWR VGND sg13g2_decap_8
XFILLER_34_631 VPWR VGND sg13g2_decap_8
XFILLER_33_163 VPWR VGND sg13g2_decap_8
XFILLER_21_314 VPWR VGND sg13g2_decap_8
XFILLER_30_870 VPWR VGND sg13g2_decap_8
XFILLER_29_469 VPWR VGND sg13g2_decap_8
XFILLER_38_992 VPWR VGND sg13g2_decap_8
XFILLER_25_664 VPWR VGND sg13g2_decap_8
XFILLER_13_837 VPWR VGND sg13g2_decap_8
XFILLER_24_185 VPWR VGND sg13g2_decap_8
XFILLER_12_347 VPWR VGND sg13g2_decap_8
XFILLER_40_656 VPWR VGND sg13g2_decap_8
XFILLER_4_502 VPWR VGND sg13g2_fill_2
XFILLER_0_763 VPWR VGND sg13g2_decap_8
XFILLER_48_723 VPWR VGND sg13g2_decap_8
XFILLER_36_918 VPWR VGND sg13g2_decap_8
XFILLER_35_428 VPWR VGND sg13g2_decap_8
XFILLER_16_642 VPWR VGND sg13g2_decap_8
XFILLER_28_480 VPWR VGND sg13g2_decap_8
XFILLER_44_962 VPWR VGND sg13g2_decap_8
XFILLER_43_450 VPWR VGND sg13g2_decap_8
XFILLER_15_130 VPWR VGND sg13g2_decap_8
XFILLER_31_645 VPWR VGND sg13g2_decap_8
XFILLER_30_133 VPWR VGND sg13g2_decap_8
XFILLER_7_21 VPWR VGND sg13g2_decap_8
XFILLER_8_852 VPWR VGND sg13g2_decap_8
XFILLER_38_244 VPWR VGND sg13g2_decap_8
XFILLER_38_255 VPWR VGND sg13g2_fill_2
XFILLER_39_767 VPWR VGND sg13g2_decap_8
XFILLER_35_995 VPWR VGND sg13g2_decap_8
XFILLER_10_818 VPWR VGND sg13g2_decap_8
XFILLER_22_667 VPWR VGND sg13g2_decap_8
XFILLER_1_549 VPWR VGND sg13g2_decap_8
XFILLER_29_244 VPWR VGND sg13g2_decap_8
X_550_ net72 VGND VPWR _042_ mac1.products_ff\[0\] clknet_5_23__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_417 VPWR VGND sg13g2_decap_8
XFILLER_45_759 VPWR VGND sg13g2_decap_8
XFILLER_44_269 VPWR VGND sg13g2_decap_8
X_481_ net60 VGND VPWR _103_ DP_2.matrix\[113\] clknet_5_6__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_409 VPWR VGND sg13g2_decap_8
XFILLER_34_1009 VPWR VGND sg13g2_decap_8
XFILLER_41_954 VPWR VGND sg13g2_decap_8
XFILLER_12_155 VPWR VGND sg13g2_decap_8
XFILLER_32_95 VPWR VGND sg13g2_decap_8
XFILLER_5_855 VPWR VGND sg13g2_decap_8
XFILLER_4_332 VPWR VGND sg13g2_decap_8
XFILLER_4_310 VPWR VGND sg13g2_decap_4
XFILLER_48_520 VPWR VGND sg13g2_decap_8
XFILLER_0_560 VPWR VGND sg13g2_decap_8
XFILLER_48_597 VPWR VGND sg13g2_decap_8
XFILLER_36_715 VPWR VGND sg13g2_decap_8
XFILLER_35_214 VPWR VGND sg13g2_decap_8
XFILLER_16_450 VPWR VGND sg13g2_decap_8
XFILLER_32_932 VPWR VGND sg13g2_decap_8
Xhold115 mac1.sum_lvl3_ff\[0\] VPWR VGND net165 sg13g2_dlygate4sd3_1
Xhold104 DP_1.matrix\[0\] VPWR VGND net154 sg13g2_dlygate4sd3_1
Xhold126 _179_ VPWR VGND net176 sg13g2_dlygate4sd3_1
Xhold137 _028_ VPWR VGND net187 sg13g2_dlygate4sd3_1
Xhold148 mac2.sum_lvl1_ff\[1\] VPWR VGND net198 sg13g2_dlygate4sd3_1
XFILLER_39_564 VPWR VGND sg13g2_decap_8
XFILLER_23_943 VPWR VGND sg13g2_decap_8
XFILLER_35_792 VPWR VGND sg13g2_decap_8
XFILLER_34_280 VPWR VGND sg13g2_decap_8
XFILLER_34_291 VPWR VGND sg13g2_fill_1
XFILLER_10_615 VPWR VGND sg13g2_decap_8
XFILLER_22_486 VPWR VGND sg13g2_decap_8
XFILLER_5_107 VPWR VGND sg13g2_decap_8
XFILLER_2_858 VPWR VGND sg13g2_decap_8
Xclkbuf_5_13__f_clk clknet_4_6_0_clk clknet_5_13__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_1_346 VPWR VGND sg13g2_decap_8
XFILLER_40_1013 VPWR VGND sg13g2_decap_8
XFILLER_18_737 VPWR VGND sg13g2_decap_8
XFILLER_27_51 VPWR VGND sg13g2_decap_8
XFILLER_45_556 VPWR VGND sg13g2_decap_8
X_533_ net71 VGND VPWR _053_ mac1.products_ff\[49\] clknet_5_20__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_258 VPWR VGND sg13g2_decap_8
X_464_ net56 VGND VPWR _086_ DP_1.matrix\[128\] clknet_5_4__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_228 VPWR VGND sg13g2_decap_8
XFILLER_14_954 VPWR VGND sg13g2_decap_8
XFILLER_41_751 VPWR VGND sg13g2_decap_8
XFILLER_9_424 VPWR VGND sg13g2_decap_8
X_395_ net55 _089_ VPWR VGND sg13g2_buf_1
XFILLER_13_464 VPWR VGND sg13g2_decap_8
XFILLER_40_250 VPWR VGND sg13g2_decap_8
XFILLER_40_283 VPWR VGND sg13g2_decap_8
Xheichips25_template_7 VPWR VGND uio_out[2] sg13g2_tielo
XFILLER_5_652 VPWR VGND sg13g2_decap_8
XFILLER_4_151 VPWR VGND sg13g2_decap_8
XFILLER_4_162 VPWR VGND sg13g2_fill_1
XFILLER_4_11 VPWR VGND sg13g2_decap_8
XFILLER_4_99 VPWR VGND sg13g2_decap_8
XFILLER_49_895 VPWR VGND sg13g2_decap_8
XFILLER_36_512 VPWR VGND sg13g2_decap_8
XFILLER_48_394 VPWR VGND sg13g2_decap_8
XFILLER_36_589 VPWR VGND sg13g2_decap_8
XFILLER_23_239 VPWR VGND sg13g2_decap_8
XFILLER_31_250 VPWR VGND sg13g2_fill_1
XFILLER_20_957 VPWR VGND sg13g2_decap_8
XFILLER_48_28 VPWR VGND sg13g2_decap_8
XFILLER_27_567 VPWR VGND sg13g2_decap_8
XFILLER_23_740 VPWR VGND sg13g2_decap_8
Xfanout65 net68 net65 VPWR VGND sg13g2_buf_8
XFILLER_11_935 VPWR VGND sg13g2_decap_8
Xfanout76 net77 net76 VPWR VGND sg13g2_buf_8
XFILLER_13_53 VPWR VGND sg13g2_decap_8
XFILLER_1_143 VPWR VGND sg13g2_decap_8
XFILLER_2_655 VPWR VGND sg13g2_decap_8
XFILLER_49_147 VPWR VGND sg13g2_decap_8
XFILLER_38_50 VPWR VGND sg13g2_decap_8
XFILLER_18_512 VPWR VGND sg13g2_decap_8
XFILLER_46_876 VPWR VGND sg13g2_decap_8
XFILLER_45_342 VPWR VGND sg13g2_decap_8
X_516_ net64 VGND VPWR _138_ DP_4.matrix\[112\] clknet_5_2__leaf_clk sg13g2_dfrbpq_1
XFILLER_14_751 VPWR VGND sg13g2_decap_8
XFILLER_33_548 VPWR VGND sg13g2_decap_8
X_447_ net83 _141_ VPWR VGND sg13g2_buf_1
XFILLER_9_221 VPWR VGND sg13g2_fill_1
X_378_ net128 _072_ VPWR VGND sg13g2_buf_1
XFILLER_6_950 VPWR VGND sg13g2_decap_8
XFILLER_5_471 VPWR VGND sg13g2_decap_8
XFILLER_28_309 VPWR VGND sg13g2_decap_8
XFILLER_49_692 VPWR VGND sg13g2_decap_8
XFILLER_48_180 VPWR VGND sg13g2_decap_4
XFILLER_37_854 VPWR VGND sg13g2_decap_8
XFILLER_24_537 VPWR VGND sg13g2_decap_8
XFILLER_36_397 VPWR VGND sg13g2_decap_8
XFILLER_20_754 VPWR VGND sg13g2_decap_8
Xclkload7 VPWR clkload7/Y clknet_5_27__leaf_clk VGND sg13g2_inv_1
XFILLER_4_909 VPWR VGND sg13g2_decap_8
XFILLER_8_1013 VPWR VGND sg13g2_decap_8
XFILLER_47_618 VPWR VGND sg13g2_decap_8
XFILLER_28_876 VPWR VGND sg13g2_decap_8
XFILLER_42_301 VPWR VGND sg13g2_decap_8
XFILLER_15_504 VPWR VGND sg13g2_fill_2
XFILLER_15_526 VPWR VGND sg13g2_decap_8
XFILLER_43_868 VPWR VGND sg13g2_decap_8
XFILLER_15_559 VPWR VGND sg13g2_fill_1
X_301_ _176_ net180 net113 VPWR VGND sg13g2_nand2_1
X_232_ net160 net123 _054_ VPWR VGND sg13g2_and2_1
XFILLER_11_732 VPWR VGND sg13g2_decap_8
XFILLER_7_758 VPWR VGND sg13g2_decap_8
XFILLER_6_246 VPWR VGND sg13g2_decap_8
XFILLER_40_95 VPWR VGND sg13g2_decap_8
XFILLER_3_964 VPWR VGND sg13g2_decap_8
XFILLER_38_607 VPWR VGND sg13g2_decap_8
XFILLER_1_56 VPWR VGND sg13g2_decap_8
XFILLER_19_854 VPWR VGND sg13g2_decap_8
XFILLER_46_673 VPWR VGND sg13g2_decap_8
XFILLER_34_813 VPWR VGND sg13g2_decap_8
XFILLER_45_194 VPWR VGND sg13g2_decap_8
XFILLER_33_334 VPWR VGND sg13g2_decap_8
XFILLER_33_345 VPWR VGND sg13g2_fill_2
XFILLER_21_518 VPWR VGND sg13g2_decap_8
XFILLER_14_570 VPWR VGND sg13g2_decap_8
XFILLER_46_0 VPWR VGND sg13g2_decap_8
Xhold19 DP_3.matrix\[113\] VPWR VGND net43 sg13g2_dlygate4sd3_1
XFILLER_28_128 VPWR VGND sg13g2_decap_8
XFILLER_37_651 VPWR VGND sg13g2_decap_8
XFILLER_36_161 VPWR VGND sg13g2_fill_1
XFILLER_25_846 VPWR VGND sg13g2_decap_8
XFILLER_12_529 VPWR VGND sg13g2_decap_8
XFILLER_40_838 VPWR VGND sg13g2_decap_8
XFILLER_4_706 VPWR VGND sg13g2_decap_8
XFILLER_10_65 VPWR VGND sg13g2_decap_8
XFILLER_0_945 VPWR VGND sg13g2_decap_8
XFILLER_48_905 VPWR VGND sg13g2_decap_8
XFILLER_47_415 VPWR VGND sg13g2_decap_8
XFILLER_19_74 VPWR VGND sg13g2_decap_8
XFILLER_16_824 VPWR VGND sg13g2_decap_8
XFILLER_28_673 VPWR VGND sg13g2_decap_8
XFILLER_27_194 VPWR VGND sg13g2_decap_8
XFILLER_43_665 VPWR VGND sg13g2_decap_8
XFILLER_15_356 VPWR VGND sg13g2_fill_1
XFILLER_30_304 VPWR VGND sg13g2_decap_4
XFILLER_31_827 VPWR VGND sg13g2_decap_8
XFILLER_7_555 VPWR VGND sg13g2_decap_8
XFILLER_3_761 VPWR VGND sg13g2_decap_8
XFILLER_18_4 VPWR VGND sg13g2_decap_8
XFILLER_38_415 VPWR VGND sg13g2_decap_8
XFILLER_39_949 VPWR VGND sg13g2_decap_8
XFILLER_19_651 VPWR VGND sg13g2_decap_8
XFILLER_47_982 VPWR VGND sg13g2_decap_8
XFILLER_46_470 VPWR VGND sg13g2_decap_8
XFILLER_34_610 VPWR VGND sg13g2_decap_8
XFILLER_18_183 VPWR VGND sg13g2_decap_8
XFILLER_33_142 VPWR VGND sg13g2_decap_8
XFILLER_34_687 VPWR VGND sg13g2_decap_8
XFILLER_22_849 VPWR VGND sg13g2_decap_8
XFILLER_5_1027 VPWR VGND sg13g2_fill_2
XFILLER_5_1016 VPWR VGND sg13g2_decap_8
XFILLER_29_404 VPWR VGND sg13g2_decap_8
XFILLER_29_448 VPWR VGND sg13g2_decap_8
XFILLER_38_971 VPWR VGND sg13g2_decap_8
XFILLER_25_643 VPWR VGND sg13g2_decap_8
XFILLER_13_816 VPWR VGND sg13g2_decap_8
XFILLER_12_326 VPWR VGND sg13g2_decap_8
XFILLER_24_164 VPWR VGND sg13g2_decap_8
XFILLER_40_635 VPWR VGND sg13g2_decap_8
XFILLER_20_381 VPWR VGND sg13g2_decap_8
XFILLER_21_86 VPWR VGND sg13g2_decap_8
XFILLER_48_702 VPWR VGND sg13g2_decap_8
XFILLER_43_1022 VPWR VGND sg13g2_decap_8
XFILLER_0_742 VPWR VGND sg13g2_decap_8
XFILLER_48_779 VPWR VGND sg13g2_decap_8
XFILLER_46_83 VPWR VGND sg13g2_decap_4
XFILLER_44_941 VPWR VGND sg13g2_decap_8
XFILLER_16_621 VPWR VGND sg13g2_decap_8
XFILLER_16_698 VPWR VGND sg13g2_decap_8
XFILLER_30_112 VPWR VGND sg13g2_decap_8
XFILLER_31_624 VPWR VGND sg13g2_decap_8
XFILLER_8_831 VPWR VGND sg13g2_decap_8
XFILLER_7_77 VPWR VGND sg13g2_decap_8
XFILLER_7_385 VPWR VGND sg13g2_fill_2
XFILLER_39_746 VPWR VGND sg13g2_decap_8
XFILLER_35_974 VPWR VGND sg13g2_decap_8
XFILLER_34_484 VPWR VGND sg13g2_decap_8
XFILLER_21_134 VPWR VGND sg13g2_decap_8
XFILLER_22_646 VPWR VGND sg13g2_decap_8
XFILLER_21_189 VPWR VGND sg13g2_decap_8
XFILLER_1_528 VPWR VGND sg13g2_decap_8
XFILLER_29_223 VPWR VGND sg13g2_decap_8
XFILLER_18_919 VPWR VGND sg13g2_decap_8
XFILLER_45_738 VPWR VGND sg13g2_decap_8
XFILLER_29_289 VPWR VGND sg13g2_decap_8
XFILLER_44_248 VPWR VGND sg13g2_decap_8
X_480_ net60 VGND VPWR _102_ DP_2.matrix\[112\] clknet_5_7__leaf_clk sg13g2_dfrbpq_1
XFILLER_26_985 VPWR VGND sg13g2_decap_8
XFILLER_13_613 VPWR VGND sg13g2_fill_1
XFILLER_41_933 VPWR VGND sg13g2_decap_8
XFILLER_12_112 VPWR VGND sg13g2_decap_8
XFILLER_9_639 VPWR VGND sg13g2_decap_8
XFILLER_8_149 VPWR VGND sg13g2_decap_8
XFILLER_32_52 VPWR VGND sg13g2_fill_2
XFILLER_32_74 VPWR VGND sg13g2_decap_8
XFILLER_5_834 VPWR VGND sg13g2_decap_8
XFILLER_10_1021 VPWR VGND sg13g2_decap_8
XFILLER_4_388 VPWR VGND sg13g2_decap_8
XFILLER_48_576 VPWR VGND sg13g2_decap_8
XFILLER_17_985 VPWR VGND sg13g2_decap_8
XFILLER_32_911 VPWR VGND sg13g2_decap_8
XFILLER_32_988 VPWR VGND sg13g2_decap_8
Xhold116 _015_ VPWR VGND net166 sg13g2_dlygate4sd3_1
Xhold105 DP_4.matrix\[112\] VPWR VGND net155 sg13g2_dlygate4sd3_1
Xhold138 mac1.products_ff\[65\] VPWR VGND net188 sg13g2_dlygate4sd3_1
Xhold127 _022_ VPWR VGND net177 sg13g2_dlygate4sd3_1
Xhold149 _175_ VPWR VGND net199 sg13g2_dlygate4sd3_1
XFILLER_39_543 VPWR VGND sg13g2_decap_8
XFILLER_2_1019 VPWR VGND sg13g2_decap_8
XFILLER_27_749 VPWR VGND sg13g2_decap_8
XFILLER_26_259 VPWR VGND sg13g2_decap_8
XFILLER_23_922 VPWR VGND sg13g2_decap_8
XFILLER_35_771 VPWR VGND sg13g2_decap_8
XFILLER_22_432 VPWR VGND sg13g2_decap_4
XFILLER_22_465 VPWR VGND sg13g2_decap_8
XFILLER_23_999 VPWR VGND sg13g2_decap_8
XFILLER_33_1010 VPWR VGND sg13g2_decap_8
XFILLER_2_837 VPWR VGND sg13g2_decap_8
XFILLER_1_325 VPWR VGND sg13g2_decap_8
XFILLER_49_329 VPWR VGND sg13g2_decap_8
X_601_ net58 VGND VPWR net33 mac2.sum_lvl3_ff\[3\] clknet_5_6__leaf_clk sg13g2_dfrbpq_1
XFILLER_18_716 VPWR VGND sg13g2_decap_8
XFILLER_45_535 VPWR VGND sg13g2_decap_8
XFILLER_17_237 VPWR VGND sg13g2_decap_8
X_532_ net71 VGND VPWR _052_ mac1.products_ff\[48\] clknet_5_20__leaf_clk sg13g2_dfrbpq_1
XFILLER_14_933 VPWR VGND sg13g2_decap_8
X_463_ net60 VGND VPWR _085_ DP_1.matrix\[113\] clknet_5_6__leaf_clk sg13g2_dfrbpq_1
XFILLER_26_782 VPWR VGND sg13g2_decap_8
XFILLER_32_207 VPWR VGND sg13g2_decap_8
XFILLER_32_218 VPWR VGND sg13g2_fill_2
XFILLER_25_292 VPWR VGND sg13g2_decap_8
XFILLER_41_730 VPWR VGND sg13g2_decap_8
X_394_ net156 _088_ VPWR VGND sg13g2_buf_1
XFILLER_9_403 VPWR VGND sg13g2_decap_8
XFILLER_43_84 VPWR VGND sg13g2_decap_8
XFILLER_40_273 VPWR VGND sg13g2_fill_1
Xheichips25_template_8 VPWR VGND uio_out[3] sg13g2_tielo
XFILLER_5_631 VPWR VGND sg13g2_decap_8
XFILLER_4_130 VPWR VGND sg13g2_decap_8
XFILLER_4_78 VPWR VGND sg13g2_decap_8
XFILLER_1_892 VPWR VGND sg13g2_decap_8
XFILLER_49_874 VPWR VGND sg13g2_decap_8
XFILLER_48_351 VPWR VGND sg13g2_decap_8
XFILLER_24_719 VPWR VGND sg13g2_decap_8
XFILLER_36_568 VPWR VGND sg13g2_decap_8
XFILLER_17_782 VPWR VGND sg13g2_decap_8
XFILLER_23_218 VPWR VGND sg13g2_decap_8
XFILLER_16_281 VPWR VGND sg13g2_decap_8
XFILLER_17_1027 VPWR VGND sg13g2_fill_2
XFILLER_32_785 VPWR VGND sg13g2_decap_8
XFILLER_20_936 VPWR VGND sg13g2_decap_8
XFILLER_39_362 VPWR VGND sg13g2_fill_2
XFILLER_39_395 VPWR VGND sg13g2_decap_8
XFILLER_27_546 VPWR VGND sg13g2_decap_8
XFILLER_42_549 VPWR VGND sg13g2_decap_8
XFILLER_11_914 VPWR VGND sg13g2_decap_8
XFILLER_22_240 VPWR VGND sg13g2_decap_8
XFILLER_13_32 VPWR VGND sg13g2_decap_8
XFILLER_23_796 VPWR VGND sg13g2_decap_8
Xfanout77 net81 net77 VPWR VGND sg13g2_buf_8
Xfanout66 net68 net66 VPWR VGND sg13g2_buf_1
XFILLER_10_468 VPWR VGND sg13g2_fill_1
XFILLER_6_428 VPWR VGND sg13g2_decap_4
XFILLER_2_634 VPWR VGND sg13g2_decap_8
XFILLER_49_126 VPWR VGND sg13g2_decap_8
XFILLER_1_199 VPWR VGND sg13g2_decap_8
XFILLER_38_40 VPWR VGND sg13g2_fill_1
XFILLER_45_310 VPWR VGND sg13g2_decap_8
XFILLER_46_855 VPWR VGND sg13g2_decap_8
XFILLER_18_568 VPWR VGND sg13g2_fill_2
XFILLER_45_365 VPWR VGND sg13g2_fill_1
X_515_ net63 VGND VPWR _137_ DP_4.matrix\[97\] clknet_5_8__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_527 VPWR VGND sg13g2_decap_8
XFILLER_14_730 VPWR VGND sg13g2_decap_8
XFILLER_9_200 VPWR VGND sg13g2_decap_8
X_446_ net124 _140_ VPWR VGND sg13g2_buf_1
X_377_ net46 _071_ VPWR VGND sg13g2_buf_1
XFILLER_5_450 VPWR VGND sg13g2_decap_8
XFILLER_23_1020 VPWR VGND sg13g2_decap_8
XFILLER_49_671 VPWR VGND sg13g2_decap_8
XFILLER_37_833 VPWR VGND sg13g2_decap_8
XFILLER_24_516 VPWR VGND sg13g2_decap_8
XFILLER_36_376 VPWR VGND sg13g2_decap_8
XFILLER_20_733 VPWR VGND sg13g2_decap_8
XFILLER_32_582 VPWR VGND sg13g2_decap_8
Xclkload8 VPWR clkload8/Y clknet_5_31__leaf_clk VGND sg13g2_inv_1
XFILLER_30_1024 VPWR VGND sg13g2_decap_4
XFILLER_28_855 VPWR VGND sg13g2_decap_8
XFILLER_27_365 VPWR VGND sg13g2_decap_4
XFILLER_43_847 VPWR VGND sg13g2_decap_8
XFILLER_27_398 VPWR VGND sg13g2_fill_1
X_300_ mac2.sum_lvl1_ff\[0\] net121 _025_ VPWR VGND sg13g2_xor2_1
XFILLER_42_357 VPWR VGND sg13g2_decap_8
X_231_ net164 net132 _052_ VPWR VGND sg13g2_and2_1
XFILLER_11_711 VPWR VGND sg13g2_decap_8
XFILLER_23_593 VPWR VGND sg13g2_decap_8
XFILLER_24_64 VPWR VGND sg13g2_decap_4
XFILLER_24_97 VPWR VGND sg13g2_decap_8
XFILLER_7_737 VPWR VGND sg13g2_decap_8
XFILLER_6_225 VPWR VGND sg13g2_decap_8
XFILLER_11_788 VPWR VGND sg13g2_decap_8
XFILLER_40_74 VPWR VGND sg13g2_decap_8
XFILLER_3_943 VPWR VGND sg13g2_decap_8
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_19_833 VPWR VGND sg13g2_decap_8
XFILLER_46_652 VPWR VGND sg13g2_decap_8
XFILLER_45_173 VPWR VGND sg13g2_decap_8
XFILLER_33_313 VPWR VGND sg13g2_decap_8
XFILLER_34_869 VPWR VGND sg13g2_decap_8
X_429_ net87 _123_ VPWR VGND sg13g2_buf_1
XFILLER_39_0 VPWR VGND sg13g2_decap_8
XFILLER_28_107 VPWR VGND sg13g2_decap_8
XFILLER_37_630 VPWR VGND sg13g2_decap_8
XFILLER_24_302 VPWR VGND sg13g2_decap_8
XFILLER_25_825 VPWR VGND sg13g2_decap_8
XFILLER_36_140 VPWR VGND sg13g2_decap_8
XFILLER_36_173 VPWR VGND sg13g2_decap_8
XFILLER_12_508 VPWR VGND sg13g2_decap_8
XFILLER_40_817 VPWR VGND sg13g2_decap_8
XFILLER_33_891 VPWR VGND sg13g2_decap_8
XFILLER_10_11 VPWR VGND sg13g2_decap_8
XFILLER_10_22 VPWR VGND sg13g2_fill_2
XFILLER_0_924 VPWR VGND sg13g2_decap_8
XFILLER_19_53 VPWR VGND sg13g2_decap_8
XFILLER_28_652 VPWR VGND sg13g2_decap_8
XFILLER_16_803 VPWR VGND sg13g2_decap_8
XFILLER_43_644 VPWR VGND sg13g2_decap_8
XFILLER_15_335 VPWR VGND sg13g2_decap_8
XFILLER_27_173 VPWR VGND sg13g2_decap_8
XFILLER_31_806 VPWR VGND sg13g2_decap_8
XFILLER_37_1008 VPWR VGND sg13g2_decap_8
XFILLER_24_880 VPWR VGND sg13g2_decap_8
XFILLER_42_198 VPWR VGND sg13g2_decap_8
XFILLER_30_349 VPWR VGND sg13g2_decap_8
XFILLER_7_534 VPWR VGND sg13g2_decap_8
XFILLER_11_596 VPWR VGND sg13g2_decap_8
XFILLER_3_740 VPWR VGND sg13g2_decap_8
XFILLER_32_7 VPWR VGND sg13g2_decap_8
XFILLER_39_928 VPWR VGND sg13g2_decap_8
XFILLER_38_405 VPWR VGND sg13g2_fill_1
XFILLER_19_630 VPWR VGND sg13g2_decap_8
XFILLER_47_961 VPWR VGND sg13g2_decap_8
XFILLER_18_162 VPWR VGND sg13g2_decap_8
XFILLER_34_666 VPWR VGND sg13g2_decap_8
XFILLER_22_828 VPWR VGND sg13g2_decap_8
XFILLER_29_427 VPWR VGND sg13g2_decap_8
XFILLER_38_950 VPWR VGND sg13g2_decap_8
XFILLER_25_622 VPWR VGND sg13g2_decap_8
XFILLER_24_143 VPWR VGND sg13g2_decap_8
XFILLER_12_305 VPWR VGND sg13g2_decap_8
XFILLER_25_699 VPWR VGND sg13g2_decap_8
XFILLER_40_614 VPWR VGND sg13g2_decap_8
XFILLER_8_309 VPWR VGND sg13g2_decap_8
XFILLER_20_360 VPWR VGND sg13g2_decap_8
XFILLER_21_883 VPWR VGND sg13g2_decap_8
XFILLER_4_559 VPWR VGND sg13g2_decap_8
XFILLER_4_526 VPWR VGND sg13g2_decap_8
XFILLER_21_65 VPWR VGND sg13g2_decap_8
XFILLER_0_721 VPWR VGND sg13g2_decap_8
XFILLER_43_1001 VPWR VGND sg13g2_decap_8
XFILLER_0_798 VPWR VGND sg13g2_decap_8
XFILLER_48_758 VPWR VGND sg13g2_decap_8
XFILLER_47_246 VPWR VGND sg13g2_fill_2
XFILLER_16_600 VPWR VGND sg13g2_decap_8
XFILLER_28_460 VPWR VGND sg13g2_fill_1
XFILLER_44_920 VPWR VGND sg13g2_decap_8
XFILLER_29_994 VPWR VGND sg13g2_decap_8
XFILLER_16_677 VPWR VGND sg13g2_decap_8
XFILLER_44_997 VPWR VGND sg13g2_decap_8
Xclkbuf_5_0__f_clk clknet_4_0_0_clk clknet_5_0__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_15_165 VPWR VGND sg13g2_decap_8
XFILLER_31_603 VPWR VGND sg13g2_decap_8
XFILLER_8_810 VPWR VGND sg13g2_decap_8
XFILLER_12_894 VPWR VGND sg13g2_decap_8
XFILLER_8_887 VPWR VGND sg13g2_decap_8
XFILLER_7_364 VPWR VGND sg13g2_decap_8
XFILLER_7_56 VPWR VGND sg13g2_decap_8
XFILLER_39_725 VPWR VGND sg13g2_decap_8
XFILLER_26_419 VPWR VGND sg13g2_decap_8
XFILLER_35_953 VPWR VGND sg13g2_decap_8
XFILLER_22_625 VPWR VGND sg13g2_decap_8
XFILLER_34_463 VPWR VGND sg13g2_decap_8
XFILLER_1_507 VPWR VGND sg13g2_decap_8
XFILLER_45_717 VPWR VGND sg13g2_decap_8
XFILLER_29_279 VPWR VGND sg13g2_fill_1
XFILLER_44_227 VPWR VGND sg13g2_decap_8
XFILLER_16_32 VPWR VGND sg13g2_fill_2
XFILLER_25_441 VPWR VGND sg13g2_decap_8
XFILLER_26_964 VPWR VGND sg13g2_decap_8
XFILLER_16_76 VPWR VGND sg13g2_decap_8
XFILLER_16_87 VPWR VGND sg13g2_fill_1
XFILLER_41_912 VPWR VGND sg13g2_decap_8
XFILLER_25_496 VPWR VGND sg13g2_decap_8
XFILLER_40_444 VPWR VGND sg13g2_decap_8
XFILLER_9_618 VPWR VGND sg13g2_decap_8
XFILLER_13_669 VPWR VGND sg13g2_decap_8
XFILLER_41_989 VPWR VGND sg13g2_decap_8
XFILLER_21_680 VPWR VGND sg13g2_decap_8
XFILLER_40_488 VPWR VGND sg13g2_decap_8
XFILLER_5_813 VPWR VGND sg13g2_decap_8
XFILLER_10_1000 VPWR VGND sg13g2_decap_8
XFILLER_4_367 VPWR VGND sg13g2_decap_8
XFILLER_0_595 VPWR VGND sg13g2_decap_8
XFILLER_48_555 VPWR VGND sg13g2_decap_8
XFILLER_29_791 VPWR VGND sg13g2_decap_8
XFILLER_17_964 VPWR VGND sg13g2_decap_8
XFILLER_35_249 VPWR VGND sg13g2_decap_8
XFILLER_44_794 VPWR VGND sg13g2_decap_8
XFILLER_16_485 VPWR VGND sg13g2_decap_8
XFILLER_43_282 VPWR VGND sg13g2_decap_8
XFILLER_31_433 VPWR VGND sg13g2_decap_8
XFILLER_31_444 VPWR VGND sg13g2_fill_1
XFILLER_32_967 VPWR VGND sg13g2_decap_8
XFILLER_12_691 VPWR VGND sg13g2_decap_8
Xhold106 DP_2.matrix\[0\] VPWR VGND net156 sg13g2_dlygate4sd3_1
XFILLER_8_684 VPWR VGND sg13g2_decap_8
Xhold117 mac1.sum_lvl3_ff\[3\] VPWR VGND net167 sg13g2_dlygate4sd3_1
XFILLER_7_161 VPWR VGND sg13g2_decap_8
Xhold128 mac1.products_ff\[0\] VPWR VGND net178 sg13g2_dlygate4sd3_1
Xhold139 _161_ VPWR VGND net189 sg13g2_dlygate4sd3_1
XFILLER_39_522 VPWR VGND sg13g2_decap_8
XFILLER_27_728 VPWR VGND sg13g2_decap_8
XFILLER_39_599 VPWR VGND sg13g2_decap_8
XFILLER_26_238 VPWR VGND sg13g2_decap_8
XFILLER_35_750 VPWR VGND sg13g2_decap_8
XFILLER_23_901 VPWR VGND sg13g2_decap_8
XFILLER_22_411 VPWR VGND sg13g2_decap_8
XFILLER_23_978 VPWR VGND sg13g2_decap_8
XFILLER_2_816 VPWR VGND sg13g2_decap_8
XFILLER_1_304 VPWR VGND sg13g2_decap_8
XFILLER_49_308 VPWR VGND sg13g2_decap_8
X_600_ net58 VGND VPWR net36 mac2.sum_lvl3_ff\[2\] clknet_5_4__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_514 VPWR VGND sg13g2_decap_8
XFILLER_17_216 VPWR VGND sg13g2_decap_8
X_531_ net70 VGND VPWR net190 mac1.sum_lvl1_ff\[17\] clknet_5_28__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_709 VPWR VGND sg13g2_decap_8
XFILLER_14_912 VPWR VGND sg13g2_decap_8
X_462_ net62 VGND VPWR _084_ DP_1.matrix\[112\] clknet_5_7__leaf_clk sg13g2_dfrbpq_1
XFILLER_26_761 VPWR VGND sg13g2_decap_8
X_393_ net104 _087_ VPWR VGND sg13g2_buf_1
XFILLER_25_282 VPWR VGND sg13g2_fill_2
XFILLER_43_63 VPWR VGND sg13g2_decap_8
XFILLER_14_989 VPWR VGND sg13g2_decap_8
XFILLER_40_241 VPWR VGND sg13g2_fill_1
XFILLER_41_786 VPWR VGND sg13g2_decap_8
XFILLER_9_459 VPWR VGND sg13g2_decap_8
XFILLER_13_499 VPWR VGND sg13g2_decap_8
Xheichips25_template_9 VPWR VGND uio_out[4] sg13g2_tielo
XFILLER_5_610 VPWR VGND sg13g2_decap_8
XFILLER_4_120 VPWR VGND sg13g2_decap_4
XFILLER_5_687 VPWR VGND sg13g2_decap_8
XFILLER_4_197 VPWR VGND sg13g2_decap_8
XFILLER_4_57 VPWR VGND sg13g2_decap_8
XFILLER_1_871 VPWR VGND sg13g2_decap_8
XFILLER_49_853 VPWR VGND sg13g2_decap_8
XFILLER_48_330 VPWR VGND sg13g2_decap_8
XFILLER_0_392 VPWR VGND sg13g2_decap_8
XFILLER_36_547 VPWR VGND sg13g2_decap_8
XFILLER_17_761 VPWR VGND sg13g2_decap_8
XFILLER_44_591 VPWR VGND sg13g2_decap_8
XFILLER_17_1006 VPWR VGND sg13g2_decap_8
XFILLER_20_915 VPWR VGND sg13g2_decap_8
XFILLER_31_241 VPWR VGND sg13g2_decap_8
XFILLER_32_764 VPWR VGND sg13g2_decap_8
XFILLER_31_285 VPWR VGND sg13g2_decap_8
XFILLER_9_982 VPWR VGND sg13g2_decap_8
XFILLER_27_525 VPWR VGND sg13g2_decap_8
XFILLER_42_528 VPWR VGND sg13g2_decap_8
Xfanout56 net59 net56 VPWR VGND sg13g2_buf_8
XFILLER_23_775 VPWR VGND sg13g2_decap_8
XFILLER_10_425 VPWR VGND sg13g2_decap_8
XFILLER_13_11 VPWR VGND sg13g2_decap_8
Xfanout67 net68 net67 VPWR VGND sg13g2_buf_8
Xfanout78 net80 net78 VPWR VGND sg13g2_buf_8
XFILLER_7_919 VPWR VGND sg13g2_decap_8
XFILLER_6_407 VPWR VGND sg13g2_decap_8
XFILLER_13_88 VPWR VGND sg13g2_fill_2
XFILLER_2_613 VPWR VGND sg13g2_decap_8
XFILLER_8_4 VPWR VGND sg13g2_decap_8
XFILLER_1_112 VPWR VGND sg13g2_decap_8
XFILLER_49_105 VPWR VGND sg13g2_decap_8
XFILLER_1_178 VPWR VGND sg13g2_decap_8
XFILLER_46_834 VPWR VGND sg13g2_decap_8
XFILLER_38_85 VPWR VGND sg13g2_decap_4
XFILLER_45_388 VPWR VGND sg13g2_decap_8
X_514_ net63 VGND VPWR _136_ DP_4.matrix\[96\] clknet_5_2__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_506 VPWR VGND sg13g2_decap_8
X_445_ net41 _139_ VPWR VGND sg13g2_buf_1
X_376_ net154 _070_ VPWR VGND sg13g2_buf_1
XFILLER_14_786 VPWR VGND sg13g2_decap_8
XFILLER_41_583 VPWR VGND sg13g2_decap_8
XFILLER_13_296 VPWR VGND sg13g2_decap_8
XFILLER_9_278 VPWR VGND sg13g2_fill_2
XFILLER_6_985 VPWR VGND sg13g2_decap_8
XFILLER_49_650 VPWR VGND sg13g2_decap_8
XFILLER_37_812 VPWR VGND sg13g2_decap_8
XFILLER_36_322 VPWR VGND sg13g2_decap_8
XFILLER_36_333 VPWR VGND sg13g2_fill_2
XFILLER_36_355 VPWR VGND sg13g2_decap_8
XFILLER_37_889 VPWR VGND sg13g2_decap_8
XFILLER_20_712 VPWR VGND sg13g2_decap_8
XFILLER_32_561 VPWR VGND sg13g2_decap_8
XFILLER_20_789 VPWR VGND sg13g2_decap_8
XFILLER_30_1003 VPWR VGND sg13g2_decap_8
XFILLER_28_834 VPWR VGND sg13g2_decap_8
XFILLER_39_160 VPWR VGND sg13g2_fill_2
XFILLER_43_826 VPWR VGND sg13g2_decap_8
XFILLER_15_506 VPWR VGND sg13g2_fill_1
XFILLER_42_336 VPWR VGND sg13g2_decap_8
XFILLER_23_572 VPWR VGND sg13g2_decap_8
X_230_ net131 net157 _050_ VPWR VGND sg13g2_and2_1
XFILLER_10_222 VPWR VGND sg13g2_decap_8
XFILLER_7_716 VPWR VGND sg13g2_decap_8
XFILLER_11_767 VPWR VGND sg13g2_decap_8
XFILLER_10_299 VPWR VGND sg13g2_fill_2
XFILLER_40_53 VPWR VGND sg13g2_decap_8
XFILLER_3_922 VPWR VGND sg13g2_decap_8
XFILLER_3_999 VPWR VGND sg13g2_decap_8
XFILLER_49_84 VPWR VGND sg13g2_decap_8
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_19_812 VPWR VGND sg13g2_decap_8
XFILLER_37_119 VPWR VGND sg13g2_decap_8
XFILLER_46_631 VPWR VGND sg13g2_decap_8
XFILLER_18_333 VPWR VGND sg13g2_decap_8
XFILLER_45_152 VPWR VGND sg13g2_decap_8
XFILLER_19_889 VPWR VGND sg13g2_decap_8
XFILLER_34_848 VPWR VGND sg13g2_decap_8
XFILLER_33_347 VPWR VGND sg13g2_fill_1
XFILLER_42_892 VPWR VGND sg13g2_decap_8
X_428_ net142 _122_ VPWR VGND sg13g2_buf_1
XFILLER_41_380 VPWR VGND sg13g2_fill_1
X_359_ _211_ _210_ _059_ VPWR VGND sg13g2_xor2_1
XFILLER_6_782 VPWR VGND sg13g2_decap_8
XFILLER_29_609 VPWR VGND sg13g2_decap_8
XFILLER_25_804 VPWR VGND sg13g2_decap_8
XFILLER_37_686 VPWR VGND sg13g2_decap_8
XFILLER_24_369 VPWR VGND sg13g2_decap_8
XFILLER_33_870 VPWR VGND sg13g2_decap_8
XFILLER_20_553 VPWR VGND sg13g2_decap_8
XFILLER_20_586 VPWR VGND sg13g2_decap_8
XFILLER_3_229 VPWR VGND sg13g2_decap_8
XFILLER_0_903 VPWR VGND sg13g2_decap_8
XFILLER_19_32 VPWR VGND sg13g2_decap_8
XFILLER_28_631 VPWR VGND sg13g2_decap_8
XFILLER_43_623 VPWR VGND sg13g2_decap_8
XFILLER_16_859 VPWR VGND sg13g2_decap_8
XFILLER_42_133 VPWR VGND sg13g2_decap_8
XFILLER_42_177 VPWR VGND sg13g2_decap_8
Xclkbuf_5_19__f_clk clknet_4_9_0_clk clknet_5_19__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_7_513 VPWR VGND sg13g2_decap_8
XFILLER_2_240 VPWR VGND sg13g2_fill_1
XFILLER_3_796 VPWR VGND sg13g2_decap_8
XFILLER_39_907 VPWR VGND sg13g2_decap_8
XFILLER_47_940 VPWR VGND sg13g2_decap_8
XFILLER_20_1013 VPWR VGND sg13g2_decap_8
XFILLER_18_141 VPWR VGND sg13g2_decap_8
XFILLER_19_686 VPWR VGND sg13g2_decap_8
XFILLER_22_807 VPWR VGND sg13g2_decap_8
XFILLER_34_645 VPWR VGND sg13g2_decap_8
XFILLER_15_881 VPWR VGND sg13g2_decap_8
XFILLER_21_328 VPWR VGND sg13g2_decap_4
XFILLER_33_177 VPWR VGND sg13g2_fill_2
XFILLER_30_884 VPWR VGND sg13g2_decap_8
XFILLER_44_409 VPWR VGND sg13g2_decap_8
XFILLER_25_601 VPWR VGND sg13g2_decap_8
XFILLER_24_111 VPWR VGND sg13g2_decap_8
XFILLER_37_483 VPWR VGND sg13g2_decap_8
XFILLER_25_678 VPWR VGND sg13g2_decap_8
XFILLER_24_199 VPWR VGND sg13g2_fill_2
XFILLER_21_862 VPWR VGND sg13g2_decap_8
XFILLER_21_11 VPWR VGND sg13g2_decap_8
XFILLER_21_33 VPWR VGND sg13g2_fill_2
XFILLER_21_44 VPWR VGND sg13g2_decap_8
XFILLER_4_538 VPWR VGND sg13g2_decap_8
XFILLER_0_700 VPWR VGND sg13g2_decap_8
XFILLER_48_737 VPWR VGND sg13g2_decap_8
XFILLER_0_777 VPWR VGND sg13g2_decap_8
XFILLER_47_225 VPWR VGND sg13g2_decap_8
XFILLER_29_973 VPWR VGND sg13g2_decap_8
XFILLER_28_494 VPWR VGND sg13g2_decap_8
XFILLER_44_976 VPWR VGND sg13g2_decap_8
XFILLER_15_144 VPWR VGND sg13g2_decap_8
XFILLER_16_656 VPWR VGND sg13g2_decap_8
XFILLER_43_464 VPWR VGND sg13g2_decap_8
XFILLER_43_497 VPWR VGND sg13g2_decap_8
XFILLER_15_199 VPWR VGND sg13g2_decap_8
XFILLER_31_659 VPWR VGND sg13g2_decap_8
XFILLER_12_873 VPWR VGND sg13g2_decap_8
XFILLER_30_147 VPWR VGND sg13g2_decap_8
XFILLER_7_321 VPWR VGND sg13g2_decap_8
XFILLER_7_35 VPWR VGND sg13g2_decap_8
XFILLER_8_866 VPWR VGND sg13g2_decap_8
XFILLER_7_387 VPWR VGND sg13g2_fill_1
XFILLER_3_593 VPWR VGND sg13g2_decap_8
XFILLER_23_4 VPWR VGND sg13g2_decap_8
XFILLER_38_203 VPWR VGND sg13g2_decap_8
XFILLER_39_704 VPWR VGND sg13g2_decap_8
XFILLER_19_483 VPWR VGND sg13g2_decap_8
XFILLER_35_932 VPWR VGND sg13g2_decap_8
XFILLER_22_604 VPWR VGND sg13g2_decap_8
XFILLER_30_681 VPWR VGND sg13g2_decap_8
XFILLER_27_1008 VPWR VGND sg13g2_decap_8
XFILLER_29_258 VPWR VGND sg13g2_decap_8
XFILLER_16_11 VPWR VGND sg13g2_decap_8
XFILLER_26_943 VPWR VGND sg13g2_decap_8
XFILLER_13_604 VPWR VGND sg13g2_fill_1
XFILLER_25_464 VPWR VGND sg13g2_decap_8
XFILLER_13_648 VPWR VGND sg13g2_decap_8
XFILLER_40_423 VPWR VGND sg13g2_decap_8
XFILLER_41_968 VPWR VGND sg13g2_decap_8
XFILLER_12_169 VPWR VGND sg13g2_decap_8
XFILLER_40_467 VPWR VGND sg13g2_decap_8
XFILLER_5_869 VPWR VGND sg13g2_decap_8
XFILLER_4_346 VPWR VGND sg13g2_decap_8
XFILLER_0_574 VPWR VGND sg13g2_decap_8
XFILLER_48_534 VPWR VGND sg13g2_decap_8
XFILLER_29_770 VPWR VGND sg13g2_decap_8
XFILLER_35_228 VPWR VGND sg13g2_decap_8
XFILLER_36_729 VPWR VGND sg13g2_decap_8
XFILLER_17_943 VPWR VGND sg13g2_decap_8
XFILLER_44_773 VPWR VGND sg13g2_decap_8
XFILLER_43_261 VPWR VGND sg13g2_decap_8
XFILLER_16_464 VPWR VGND sg13g2_decap_8
XFILLER_31_412 VPWR VGND sg13g2_decap_8
XFILLER_32_946 VPWR VGND sg13g2_decap_8
XFILLER_31_456 VPWR VGND sg13g2_decap_4
XFILLER_12_670 VPWR VGND sg13g2_decap_8
XFILLER_8_663 VPWR VGND sg13g2_decap_8
XFILLER_7_140 VPWR VGND sg13g2_decap_8
XFILLER_11_191 VPWR VGND sg13g2_decap_8
Xhold107 DP_2.matrix\[64\] VPWR VGND net157 sg13g2_dlygate4sd3_1
XFILLER_7_195 VPWR VGND sg13g2_decap_8
Xhold118 _167_ VPWR VGND net168 sg13g2_dlygate4sd3_1
Xhold129 _001_ VPWR VGND net179 sg13g2_dlygate4sd3_1
XFILLER_27_707 VPWR VGND sg13g2_decap_8
XFILLER_39_578 VPWR VGND sg13g2_decap_8
XFILLER_19_291 VPWR VGND sg13g2_decap_8
XFILLER_41_209 VPWR VGND sg13g2_decap_8
XFILLER_23_957 VPWR VGND sg13g2_decap_8
XFILLER_10_629 VPWR VGND sg13g2_decap_8
XFILLER_40_1027 VPWR VGND sg13g2_fill_2
X_530_ net70 VGND VPWR net98 mac1.sum_lvl1_ff\[16\] clknet_5_25__leaf_clk sg13g2_dfrbpq_1
XFILLER_27_21 VPWR VGND sg13g2_decap_8
XFILLER_26_740 VPWR VGND sg13g2_decap_8
XFILLER_27_65 VPWR VGND sg13g2_decap_8
XFILLER_27_76 VPWR VGND sg13g2_fill_1
XFILLER_13_401 VPWR VGND sg13g2_decap_8
X_461_ net67 VGND VPWR _083_ DP_1.matrix\[97\] clknet_5_24__leaf_clk sg13g2_dfrbpq_1
X_392_ net119 _086_ VPWR VGND sg13g2_buf_1
XFILLER_25_261 VPWR VGND sg13g2_decap_8
XFILLER_43_42 VPWR VGND sg13g2_decap_8
XFILLER_14_968 VPWR VGND sg13g2_decap_8
XFILLER_41_765 VPWR VGND sg13g2_decap_8
XFILLER_9_438 VPWR VGND sg13g2_decap_8
XFILLER_13_478 VPWR VGND sg13g2_decap_8
XFILLER_40_264 VPWR VGND sg13g2_decap_8
XFILLER_40_297 VPWR VGND sg13g2_decap_8
XFILLER_5_666 VPWR VGND sg13g2_decap_8
XFILLER_4_25 VPWR VGND sg13g2_decap_8
XFILLER_1_850 VPWR VGND sg13g2_decap_8
XFILLER_49_832 VPWR VGND sg13g2_decap_8
XFILLER_0_371 VPWR VGND sg13g2_decap_8
XFILLER_36_526 VPWR VGND sg13g2_decap_8
XFILLER_17_740 VPWR VGND sg13g2_decap_8
XFILLER_44_570 VPWR VGND sg13g2_decap_8
XFILLER_16_261 VPWR VGND sg13g2_decap_4
XFILLER_32_743 VPWR VGND sg13g2_decap_8
XFILLER_31_231 VPWR VGND sg13g2_fill_1
XFILLER_9_961 VPWR VGND sg13g2_decap_8
XFILLER_8_493 VPWR VGND sg13g2_decap_8
XFILLER_27_504 VPWR VGND sg13g2_decap_8
XFILLER_39_364 VPWR VGND sg13g2_fill_1
XFILLER_42_507 VPWR VGND sg13g2_decap_8
XFILLER_14_209 VPWR VGND sg13g2_decap_8
XFILLER_23_754 VPWR VGND sg13g2_decap_8
XFILLER_10_404 VPWR VGND sg13g2_decap_8
Xfanout57 net59 net57 VPWR VGND sg13g2_buf_8
XFILLER_11_949 VPWR VGND sg13g2_decap_8
Xfanout68 rst_n net68 VPWR VGND sg13g2_buf_8
Xfanout79 net80 net79 VPWR VGND sg13g2_buf_8
XFILLER_10_459 VPWR VGND sg13g2_decap_8
XFILLER_13_67 VPWR VGND sg13g2_decap_8
XFILLER_1_157 VPWR VGND sg13g2_decap_8
XFILLER_2_669 VPWR VGND sg13g2_decap_8
XFILLER_46_813 VPWR VGND sg13g2_decap_8
XFILLER_18_526 VPWR VGND sg13g2_fill_1
XFILLER_38_64 VPWR VGND sg13g2_decap_8
XFILLER_45_323 VPWR VGND sg13g2_decap_4
X_513_ net65 VGND VPWR _135_ DP_4.matrix\[81\] clknet_5_11__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_356 VPWR VGND sg13g2_decap_8
X_444_ net155 _138_ VPWR VGND sg13g2_buf_1
XFILLER_14_765 VPWR VGND sg13g2_decap_8
XFILLER_13_275 VPWR VGND sg13g2_decap_8
X_375_ net171 VPWR _031_ VGND _182_ _184_ sg13g2_o21ai_1
XFILLER_41_562 VPWR VGND sg13g2_decap_8
XFILLER_6_964 VPWR VGND sg13g2_decap_8
XFILLER_10_993 VPWR VGND sg13g2_decap_8
XFILLER_5_485 VPWR VGND sg13g2_decap_8
XFILLER_36_301 VPWR VGND sg13g2_decap_8
XFILLER_37_868 VPWR VGND sg13g2_decap_8
XFILLER_32_540 VPWR VGND sg13g2_decap_8
XFILLER_20_768 VPWR VGND sg13g2_decap_8
XFILLER_8_1027 VPWR VGND sg13g2_fill_2
XFILLER_28_813 VPWR VGND sg13g2_decap_8
XFILLER_39_150 VPWR VGND sg13g2_fill_2
XFILLER_27_312 VPWR VGND sg13g2_decap_4
XFILLER_43_805 VPWR VGND sg13g2_decap_8
XFILLER_42_315 VPWR VGND sg13g2_decap_8
XFILLER_36_890 VPWR VGND sg13g2_decap_8
XFILLER_23_551 VPWR VGND sg13g2_decap_8
XFILLER_24_11 VPWR VGND sg13g2_decap_8
XFILLER_24_22 VPWR VGND sg13g2_fill_2
XFILLER_10_201 VPWR VGND sg13g2_decap_8
XFILLER_11_746 VPWR VGND sg13g2_decap_8
XFILLER_10_267 VPWR VGND sg13g2_decap_8
XFILLER_40_21 VPWR VGND sg13g2_decap_8
XFILLER_40_32 VPWR VGND sg13g2_fill_1
XFILLER_3_901 VPWR VGND sg13g2_decap_8
XFILLER_3_978 VPWR VGND sg13g2_decap_8
XFILLER_2_444 VPWR VGND sg13g2_decap_8
XFILLER_49_63 VPWR VGND sg13g2_decap_8
XFILLER_46_610 VPWR VGND sg13g2_decap_8
XFILLER_37_109 VPWR VGND sg13g2_fill_1
XFILLER_18_312 VPWR VGND sg13g2_decap_8
XFILLER_45_131 VPWR VGND sg13g2_decap_8
XFILLER_19_868 VPWR VGND sg13g2_decap_8
XFILLER_34_827 VPWR VGND sg13g2_decap_8
XFILLER_46_687 VPWR VGND sg13g2_decap_8
XFILLER_18_389 VPWR VGND sg13g2_fill_2
XFILLER_42_871 VPWR VGND sg13g2_decap_8
XFILLER_14_584 VPWR VGND sg13g2_decap_8
X_427_ net43 _121_ VPWR VGND sg13g2_buf_1
X_358_ _211_ net119 net96 VPWR VGND sg13g2_nand2_1
XFILLER_10_790 VPWR VGND sg13g2_decap_8
X_289_ _170_ net196 net152 VPWR VGND sg13g2_nand2_1
XFILLER_6_761 VPWR VGND sg13g2_decap_8
XFILLER_37_665 VPWR VGND sg13g2_decap_8
XFILLER_20_532 VPWR VGND sg13g2_decap_8
XFILLER_32_381 VPWR VGND sg13g2_decap_8
XFILLER_10_79 VPWR VGND sg13g2_decap_8
XFILLER_48_919 VPWR VGND sg13g2_decap_8
XFILLER_0_959 VPWR VGND sg13g2_decap_8
XFILLER_19_11 VPWR VGND sg13g2_decap_8
XFILLER_47_429 VPWR VGND sg13g2_decap_8
XFILLER_19_109 VPWR VGND sg13g2_decap_8
XFILLER_19_88 VPWR VGND sg13g2_decap_8
XFILLER_28_610 VPWR VGND sg13g2_decap_8
XFILLER_43_602 VPWR VGND sg13g2_decap_8
XFILLER_42_112 VPWR VGND sg13g2_decap_8
XFILLER_16_838 VPWR VGND sg13g2_decap_8
XFILLER_28_687 VPWR VGND sg13g2_decap_8
XFILLER_35_21 VPWR VGND sg13g2_decap_8
XFILLER_35_65 VPWR VGND sg13g2_decap_8
XFILLER_43_679 VPWR VGND sg13g2_decap_8
XFILLER_35_98 VPWR VGND sg13g2_decap_8
XFILLER_11_521 VPWR VGND sg13g2_decap_8
XFILLER_11_554 VPWR VGND sg13g2_decap_8
XFILLER_7_569 VPWR VGND sg13g2_decap_8
XFILLER_3_775 VPWR VGND sg13g2_decap_8
XFILLER_38_429 VPWR VGND sg13g2_decap_8
XFILLER_18_120 VPWR VGND sg13g2_decap_8
XFILLER_19_665 VPWR VGND sg13g2_decap_8
XFILLER_47_996 VPWR VGND sg13g2_decap_8
XFILLER_46_484 VPWR VGND sg13g2_decap_8
XFILLER_34_624 VPWR VGND sg13g2_decap_8
XFILLER_18_197 VPWR VGND sg13g2_decap_8
XFILLER_15_860 VPWR VGND sg13g2_decap_8
XFILLER_21_307 VPWR VGND sg13g2_decap_8
XFILLER_33_156 VPWR VGND sg13g2_decap_8
XFILLER_14_392 VPWR VGND sg13g2_decap_8
XFILLER_30_863 VPWR VGND sg13g2_decap_8
XFILLER_44_0 VPWR VGND sg13g2_decap_8
Xclkbuf_5_25__f_clk clknet_4_12_0_clk clknet_5_25__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_38_985 VPWR VGND sg13g2_decap_8
XFILLER_25_657 VPWR VGND sg13g2_decap_8
XFILLER_24_178 VPWR VGND sg13g2_decap_8
XFILLER_21_841 VPWR VGND sg13g2_decap_8
XFILLER_40_649 VPWR VGND sg13g2_decap_8
XFILLER_20_395 VPWR VGND sg13g2_decap_8
XFILLER_0_756 VPWR VGND sg13g2_decap_8
XFILLER_48_716 VPWR VGND sg13g2_decap_8
XFILLER_47_248 VPWR VGND sg13g2_fill_1
XFILLER_28_451 VPWR VGND sg13g2_decap_8
XFILLER_29_952 VPWR VGND sg13g2_decap_8
XFILLER_28_473 VPWR VGND sg13g2_decap_8
XFILLER_44_955 VPWR VGND sg13g2_decap_8
XFILLER_43_443 VPWR VGND sg13g2_decap_8
XFILLER_15_123 VPWR VGND sg13g2_decap_8
XFILLER_16_635 VPWR VGND sg13g2_decap_8
XFILLER_30_126 VPWR VGND sg13g2_decap_8
XFILLER_31_638 VPWR VGND sg13g2_decap_8
XFILLER_12_852 VPWR VGND sg13g2_decap_8
XFILLER_8_845 VPWR VGND sg13g2_decap_8
XFILLER_7_300 VPWR VGND sg13g2_decap_8
XFILLER_7_14 VPWR VGND sg13g2_decap_8
XFILLER_11_351 VPWR VGND sg13g2_decap_8
XFILLER_3_572 VPWR VGND sg13g2_decap_8
XFILLER_16_4 VPWR VGND sg13g2_decap_8
XFILLER_38_237 VPWR VGND sg13g2_decap_8
XFILLER_47_793 VPWR VGND sg13g2_decap_8
XFILLER_19_462 VPWR VGND sg13g2_decap_8
XFILLER_34_410 VPWR VGND sg13g2_fill_2
XFILLER_35_911 VPWR VGND sg13g2_decap_8
XFILLER_35_988 VPWR VGND sg13g2_decap_8
XFILLER_34_498 VPWR VGND sg13g2_decap_8
XFILLER_30_660 VPWR VGND sg13g2_decap_8
XFILLER_29_237 VPWR VGND sg13g2_decap_8
XFILLER_26_922 VPWR VGND sg13g2_decap_8
XFILLER_38_782 VPWR VGND sg13g2_decap_8
XFILLER_16_34 VPWR VGND sg13g2_fill_1
XFILLER_37_281 VPWR VGND sg13g2_decap_8
XFILLER_26_999 VPWR VGND sg13g2_decap_8
XFILLER_40_402 VPWR VGND sg13g2_decap_8
XFILLER_41_947 VPWR VGND sg13g2_decap_8
XFILLER_20_181 VPWR VGND sg13g2_decap_4
XFILLER_32_88 VPWR VGND sg13g2_decap_8
XFILLER_5_848 VPWR VGND sg13g2_decap_8
XFILLER_4_325 VPWR VGND sg13g2_decap_8
XFILLER_4_314 VPWR VGND sg13g2_fill_2
XFILLER_4_303 VPWR VGND sg13g2_decap_8
XFILLER_0_553 VPWR VGND sg13g2_decap_8
XFILLER_48_513 VPWR VGND sg13g2_decap_8
XFILLER_36_708 VPWR VGND sg13g2_decap_8
XFILLER_17_922 VPWR VGND sg13g2_decap_8
XFILLER_35_207 VPWR VGND sg13g2_decap_8
XFILLER_16_421 VPWR VGND sg13g2_decap_4
XFILLER_44_752 VPWR VGND sg13g2_decap_8
XFILLER_16_443 VPWR VGND sg13g2_decap_8
XFILLER_17_999 VPWR VGND sg13g2_decap_8
XFILLER_32_925 VPWR VGND sg13g2_decap_8
XFILLER_8_642 VPWR VGND sg13g2_decap_8
XFILLER_11_170 VPWR VGND sg13g2_decap_8
Xhold108 DP_2.matrix\[80\] VPWR VGND net158 sg13g2_dlygate4sd3_1
Xhold119 _014_ VPWR VGND net169 sg13g2_dlygate4sd3_1
XFILLER_4_881 VPWR VGND sg13g2_decap_8
XFILLER_3_380 VPWR VGND sg13g2_decap_8
XFILLER_26_1020 VPWR VGND sg13g2_decap_8
XFILLER_39_557 VPWR VGND sg13g2_decap_8
XFILLER_47_590 VPWR VGND sg13g2_decap_8
XFILLER_23_936 VPWR VGND sg13g2_decap_8
XFILLER_34_273 VPWR VGND sg13g2_decap_8
XFILLER_35_785 VPWR VGND sg13g2_decap_8
XFILLER_10_608 VPWR VGND sg13g2_decap_8
XFILLER_22_479 VPWR VGND sg13g2_decap_8
XFILLER_33_1024 VPWR VGND sg13g2_decap_4
XFILLER_1_339 VPWR VGND sg13g2_decap_8
XFILLER_40_1006 VPWR VGND sg13g2_decap_8
XFILLER_27_44 VPWR VGND sg13g2_decap_8
XFILLER_45_549 VPWR VGND sg13g2_decap_8
X_460_ net60 VGND VPWR _082_ DP_1.matrix\[96\] clknet_5_24__leaf_clk sg13g2_dfrbpq_1
XFILLER_25_240 VPWR VGND sg13g2_decap_8
XFILLER_43_21 VPWR VGND sg13g2_decap_8
XFILLER_13_424 VPWR VGND sg13g2_decap_4
XFILLER_14_947 VPWR VGND sg13g2_decap_8
X_391_ net47 _085_ VPWR VGND sg13g2_buf_1
XFILLER_26_796 VPWR VGND sg13g2_decap_8
XFILLER_9_417 VPWR VGND sg13g2_decap_8
XFILLER_13_457 VPWR VGND sg13g2_decap_8
XFILLER_40_232 VPWR VGND sg13g2_decap_8
XFILLER_41_744 VPWR VGND sg13g2_decap_8
XFILLER_43_98 VPWR VGND sg13g2_decap_8
XFILLER_5_645 VPWR VGND sg13g2_decap_8
XFILLER_4_144 VPWR VGND sg13g2_decap_8
XFILLER_49_811 VPWR VGND sg13g2_decap_8
XFILLER_0_350 VPWR VGND sg13g2_decap_8
XFILLER_49_888 VPWR VGND sg13g2_decap_8
XFILLER_48_387 VPWR VGND sg13g2_decap_8
XFILLER_36_505 VPWR VGND sg13g2_decap_8
XFILLER_1_1011 VPWR VGND sg13g2_decap_8
X_589_ net57 VGND VPWR net30 mac2.sum_lvl2_ff\[8\] clknet_5_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_796 VPWR VGND sg13g2_decap_8
XFILLER_31_210 VPWR VGND sg13g2_fill_1
XFILLER_32_722 VPWR VGND sg13g2_decap_8
XFILLER_16_295 VPWR VGND sg13g2_decap_8
XFILLER_32_799 VPWR VGND sg13g2_decap_8
XFILLER_9_940 VPWR VGND sg13g2_decap_8
XFILLER_13_991 VPWR VGND sg13g2_decap_8
XFILLER_8_472 VPWR VGND sg13g2_decap_8
XFILLER_23_733 VPWR VGND sg13g2_decap_8
XFILLER_35_582 VPWR VGND sg13g2_decap_8
XFILLER_11_928 VPWR VGND sg13g2_decap_8
Xfanout58 net59 net58 VPWR VGND sg13g2_buf_2
Xfanout69 net70 net69 VPWR VGND sg13g2_buf_8
XFILLER_22_254 VPWR VGND sg13g2_decap_8
XFILLER_13_46 VPWR VGND sg13g2_decap_8
XFILLER_2_648 VPWR VGND sg13g2_decap_8
XFILLER_1_136 VPWR VGND sg13g2_decap_8
XFILLER_38_21 VPWR VGND sg13g2_decap_8
XFILLER_18_505 VPWR VGND sg13g2_decap_8
XFILLER_46_869 VPWR VGND sg13g2_decap_8
X_512_ net65 VGND VPWR _134_ DP_4.matrix\[80\] clknet_5_10__leaf_clk sg13g2_dfrbpq_1
X_443_ net94 _137_ VPWR VGND sg13g2_buf_1
XFILLER_13_243 VPWR VGND sg13g2_decap_4
XFILLER_14_744 VPWR VGND sg13g2_decap_8
XFILLER_26_593 VPWR VGND sg13g2_decap_8
XFILLER_41_541 VPWR VGND sg13g2_decap_8
X_374_ _221_ _220_ _069_ VPWR VGND sg13g2_xor2_1
XFILLER_9_214 VPWR VGND sg13g2_decap_8
XFILLER_10_972 VPWR VGND sg13g2_decap_8
XFILLER_6_943 VPWR VGND sg13g2_decap_8
XFILLER_5_464 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
Xclkbuf_5_6__f_clk clknet_4_3_0_clk clknet_5_6__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_49_685 VPWR VGND sg13g2_decap_8
XFILLER_48_173 VPWR VGND sg13g2_decap_8
XFILLER_37_847 VPWR VGND sg13g2_decap_8
XFILLER_20_747 VPWR VGND sg13g2_decap_8
XFILLER_32_596 VPWR VGND sg13g2_decap_8
XFILLER_8_1006 VPWR VGND sg13g2_decap_8
XFILLER_39_195 VPWR VGND sg13g2_decap_8
XFILLER_28_869 VPWR VGND sg13g2_decap_8
XFILLER_11_725 VPWR VGND sg13g2_decap_8
XFILLER_10_257 VPWR VGND sg13g2_decap_4
XFILLER_6_239 VPWR VGND sg13g2_decap_8
XFILLER_40_88 VPWR VGND sg13g2_decap_8
XFILLER_46_1023 VPWR VGND sg13g2_decap_4
XFILLER_3_957 VPWR VGND sg13g2_decap_8
XFILLER_49_42 VPWR VGND sg13g2_decap_8
XFILLER_45_110 VPWR VGND sg13g2_decap_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_19_847 VPWR VGND sg13g2_decap_8
XFILLER_46_666 VPWR VGND sg13g2_decap_8
XFILLER_34_806 VPWR VGND sg13g2_decap_8
XFILLER_45_187 VPWR VGND sg13g2_decap_8
XFILLER_33_327 VPWR VGND sg13g2_decap_8
XFILLER_42_850 VPWR VGND sg13g2_decap_8
XFILLER_14_563 VPWR VGND sg13g2_decap_8
X_426_ net125 _120_ VPWR VGND sg13g2_buf_1
X_357_ _210_ net104 net150 VPWR VGND sg13g2_nand2_1
XFILLER_41_393 VPWR VGND sg13g2_decap_8
X_288_ net165 mac1.sum_lvl3_ff\[2\] _015_ VPWR VGND sg13g2_xor2_1
XFILLER_6_740 VPWR VGND sg13g2_decap_8
XFILLER_5_272 VPWR VGND sg13g2_fill_1
XFILLER_5_261 VPWR VGND sg13g2_decap_8
XFILLER_49_482 VPWR VGND sg13g2_decap_8
XFILLER_37_644 VPWR VGND sg13g2_decap_8
XFILLER_24_316 VPWR VGND sg13g2_fill_1
XFILLER_25_839 VPWR VGND sg13g2_decap_8
XFILLER_36_154 VPWR VGND sg13g2_decap_8
XFILLER_36_187 VPWR VGND sg13g2_decap_8
XFILLER_18_891 VPWR VGND sg13g2_decap_8
XFILLER_32_360 VPWR VGND sg13g2_decap_8
XFILLER_20_511 VPWR VGND sg13g2_decap_8
XFILLER_10_58 VPWR VGND sg13g2_decap_8
XFILLER_0_938 VPWR VGND sg13g2_decap_8
XFILLER_47_408 VPWR VGND sg13g2_decap_8
XFILLER_19_67 VPWR VGND sg13g2_decap_8
XFILLER_16_817 VPWR VGND sg13g2_decap_8
XFILLER_28_666 VPWR VGND sg13g2_decap_8
XFILLER_43_658 VPWR VGND sg13g2_decap_8
XFILLER_15_349 VPWR VGND sg13g2_decap_8
XFILLER_27_187 VPWR VGND sg13g2_decap_8
XFILLER_23_371 VPWR VGND sg13g2_decap_8
XFILLER_24_894 VPWR VGND sg13g2_decap_8
XFILLER_7_548 VPWR VGND sg13g2_decap_8
XFILLER_3_754 VPWR VGND sg13g2_decap_8
XFILLER_47_975 VPWR VGND sg13g2_decap_8
XFILLER_19_644 VPWR VGND sg13g2_decap_8
XFILLER_46_463 VPWR VGND sg13g2_decap_8
XFILLER_18_176 VPWR VGND sg13g2_decap_8
XFILLER_34_603 VPWR VGND sg13g2_decap_8
XFILLER_14_371 VPWR VGND sg13g2_decap_8
X_409_ net88 _103_ VPWR VGND sg13g2_buf_1
XFILLER_30_842 VPWR VGND sg13g2_decap_8
XFILLER_37_0 VPWR VGND sg13g2_decap_8
XFILLER_5_1009 VPWR VGND sg13g2_decap_8
XFILLER_2_81 VPWR VGND sg13g2_decap_8
XFILLER_38_964 VPWR VGND sg13g2_decap_8
XFILLER_25_636 VPWR VGND sg13g2_decap_8
XFILLER_13_809 VPWR VGND sg13g2_decap_8
XFILLER_24_157 VPWR VGND sg13g2_decap_8
XFILLER_12_319 VPWR VGND sg13g2_decap_8
XFILLER_21_820 VPWR VGND sg13g2_decap_8
XFILLER_40_628 VPWR VGND sg13g2_decap_8
XFILLER_20_374 VPWR VGND sg13g2_decap_8
XFILLER_21_897 VPWR VGND sg13g2_decap_8
XFILLER_21_79 VPWR VGND sg13g2_decap_8
XFILLER_43_1015 VPWR VGND sg13g2_decap_8
XFILLER_0_735 VPWR VGND sg13g2_decap_8
XFILLER_29_931 VPWR VGND sg13g2_decap_8
XFILLER_46_21 VPWR VGND sg13g2_decap_8
XFILLER_28_430 VPWR VGND sg13g2_decap_8
XFILLER_46_76 VPWR VGND sg13g2_decap_8
XFILLER_44_934 VPWR VGND sg13g2_decap_8
XFILLER_16_614 VPWR VGND sg13g2_decap_8
XFILLER_46_87 VPWR VGND sg13g2_fill_2
XFILLER_43_422 VPWR VGND sg13g2_decap_8
XFILLER_15_102 VPWR VGND sg13g2_decap_8
XFILLER_31_617 VPWR VGND sg13g2_decap_8
XFILLER_12_831 VPWR VGND sg13g2_decap_8
XFILLER_15_179 VPWR VGND sg13g2_decap_8
XFILLER_24_691 VPWR VGND sg13g2_decap_8
XFILLER_30_105 VPWR VGND sg13g2_decap_8
XFILLER_23_190 VPWR VGND sg13g2_decap_8
XFILLER_8_824 VPWR VGND sg13g2_decap_8
XFILLER_11_374 VPWR VGND sg13g2_decap_4
XFILLER_7_378 VPWR VGND sg13g2_decap_8
Xclkbuf_5_31__f_clk clknet_4_15_0_clk clknet_5_31__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_30_7 VPWR VGND sg13g2_decap_8
XFILLER_39_739 VPWR VGND sg13g2_decap_8
XFILLER_47_772 VPWR VGND sg13g2_decap_8
XFILLER_46_282 VPWR VGND sg13g2_decap_8
XFILLER_35_967 VPWR VGND sg13g2_decap_8
XFILLER_34_477 VPWR VGND sg13g2_decap_8
XFILLER_21_127 VPWR VGND sg13g2_decap_8
XFILLER_22_639 VPWR VGND sg13g2_decap_8
XFILLER_29_216 VPWR VGND sg13g2_decap_8
XFILLER_26_901 VPWR VGND sg13g2_decap_8
XFILLER_38_761 VPWR VGND sg13g2_decap_8
XFILLER_25_455 VPWR VGND sg13g2_decap_4
XFILLER_26_978 VPWR VGND sg13g2_decap_8
XFILLER_41_926 VPWR VGND sg13g2_decap_8
XFILLER_12_105 VPWR VGND sg13g2_decap_8
XFILLER_32_45 VPWR VGND sg13g2_decap_8
XFILLER_21_694 VPWR VGND sg13g2_decap_8
XFILLER_32_67 VPWR VGND sg13g2_decap_8
XFILLER_5_827 VPWR VGND sg13g2_decap_8
XFILLER_10_1014 VPWR VGND sg13g2_decap_8
XFILLER_0_532 VPWR VGND sg13g2_decap_8
XFILLER_48_569 VPWR VGND sg13g2_decap_8
XFILLER_17_901 VPWR VGND sg13g2_decap_8
XFILLER_44_731 VPWR VGND sg13g2_decap_8
XFILLER_43_241 VPWR VGND sg13g2_decap_4
XFILLER_17_978 VPWR VGND sg13g2_decap_8
XFILLER_32_904 VPWR VGND sg13g2_decap_8
XFILLER_16_499 VPWR VGND sg13g2_fill_1
XFILLER_43_296 VPWR VGND sg13g2_decap_8
XFILLER_8_621 VPWR VGND sg13g2_decap_8
XFILLER_40_992 VPWR VGND sg13g2_decap_8
XFILLER_8_698 VPWR VGND sg13g2_decap_8
Xhold109 DP_1.matrix\[112\] VPWR VGND net159 sg13g2_dlygate4sd3_1
XFILLER_4_860 VPWR VGND sg13g2_decap_8
XFILLER_39_536 VPWR VGND sg13g2_decap_8
XFILLER_23_915 VPWR VGND sg13g2_decap_8
XFILLER_34_252 VPWR VGND sg13g2_decap_8
XFILLER_35_764 VPWR VGND sg13g2_decap_8
XFILLER_22_425 VPWR VGND sg13g2_decap_8
XFILLER_22_436 VPWR VGND sg13g2_fill_2
XFILLER_22_458 VPWR VGND sg13g2_decap_8
XFILLER_34_296 VPWR VGND sg13g2_decap_8
XFILLER_31_981 VPWR VGND sg13g2_decap_8
XFILLER_33_1003 VPWR VGND sg13g2_decap_8
XFILLER_1_318 VPWR VGND sg13g2_decap_8
XFILLER_18_709 VPWR VGND sg13g2_decap_8
XFILLER_45_528 VPWR VGND sg13g2_decap_8
XFILLER_26_775 VPWR VGND sg13g2_decap_8
XFILLER_14_926 VPWR VGND sg13g2_decap_8
X_390_ net159 _084_ VPWR VGND sg13g2_buf_1
XFILLER_41_723 VPWR VGND sg13g2_decap_8
XFILLER_43_77 VPWR VGND sg13g2_decap_8
XFILLER_5_624 VPWR VGND sg13g2_decap_8
XFILLER_49_1021 VPWR VGND sg13g2_decap_8
XFILLER_1_885 VPWR VGND sg13g2_decap_8
XFILLER_49_867 VPWR VGND sg13g2_decap_8
XFILLER_48_344 VPWR VGND sg13g2_decap_8
XFILLER_16_274 VPWR VGND sg13g2_decap_8
XFILLER_17_775 VPWR VGND sg13g2_decap_8
XFILLER_32_701 VPWR VGND sg13g2_decap_8
X_588_ net67 VGND VPWR net187 mac2.sum_lvl2_ff\[5\] clknet_5_12__leaf_clk sg13g2_dfrbpq_1
XFILLER_31_222 VPWR VGND sg13g2_decap_8
XFILLER_13_970 VPWR VGND sg13g2_decap_8
XFILLER_20_929 VPWR VGND sg13g2_decap_8
XFILLER_32_778 VPWR VGND sg13g2_decap_8
XFILLER_31_299 VPWR VGND sg13g2_decap_8
XFILLER_8_451 VPWR VGND sg13g2_decap_8
XFILLER_9_996 VPWR VGND sg13g2_decap_8
XFILLER_39_344 VPWR VGND sg13g2_decap_4
XFILLER_27_539 VPWR VGND sg13g2_decap_8
XFILLER_23_712 VPWR VGND sg13g2_decap_8
XFILLER_35_561 VPWR VGND sg13g2_decap_8
XFILLER_11_907 VPWR VGND sg13g2_decap_8
XFILLER_22_233 VPWR VGND sg13g2_decap_8
Xfanout59 net62 net59 VPWR VGND sg13g2_buf_8
XFILLER_23_789 VPWR VGND sg13g2_decap_8
XFILLER_13_25 VPWR VGND sg13g2_decap_8
XFILLER_2_627 VPWR VGND sg13g2_decap_8
XFILLER_1_126 VPWR VGND sg13g2_decap_4
XFILLER_49_119 VPWR VGND sg13g2_decap_8
XFILLER_45_303 VPWR VGND sg13g2_decap_8
XFILLER_46_848 VPWR VGND sg13g2_decap_8
X_511_ net63 VGND VPWR _133_ DP_4.matrix\[65\] clknet_5_8__leaf_clk sg13g2_dfrbpq_1
XFILLER_14_723 VPWR VGND sg13g2_decap_8
X_442_ net136 _136_ VPWR VGND sg13g2_buf_1
XFILLER_26_572 VPWR VGND sg13g2_decap_8
XFILLER_13_222 VPWR VGND sg13g2_decap_8
XFILLER_41_520 VPWR VGND sg13g2_decap_8
X_373_ _221_ net161 net39 VPWR VGND sg13g2_nand2_1
XFILLER_16_1020 VPWR VGND sg13g2_decap_8
XFILLER_41_597 VPWR VGND sg13g2_decap_8
XFILLER_6_922 VPWR VGND sg13g2_decap_8
XFILLER_10_951 VPWR VGND sg13g2_decap_8
XFILLER_5_443 VPWR VGND sg13g2_decap_8
XFILLER_6_999 VPWR VGND sg13g2_decap_8
XFILLER_1_682 VPWR VGND sg13g2_decap_8
XFILLER_23_1013 VPWR VGND sg13g2_decap_8
XFILLER_49_664 VPWR VGND sg13g2_decap_8
XFILLER_48_152 VPWR VGND sg13g2_decap_8
XFILLER_37_826 VPWR VGND sg13g2_decap_8
XFILLER_24_509 VPWR VGND sg13g2_decap_8
XFILLER_36_369 VPWR VGND sg13g2_decap_8
XFILLER_45_892 VPWR VGND sg13g2_decap_8
XFILLER_17_550 VPWR VGND sg13g2_decap_8
XFILLER_32_575 VPWR VGND sg13g2_decap_8
XFILLER_20_726 VPWR VGND sg13g2_decap_8
XFILLER_30_1017 VPWR VGND sg13g2_decap_8
XFILLER_9_793 VPWR VGND sg13g2_decap_8
XFILLER_8_281 VPWR VGND sg13g2_decap_8
XFILLER_30_1028 VPWR VGND sg13g2_fill_1
XFILLER_28_848 VPWR VGND sg13g2_decap_8
XFILLER_27_358 VPWR VGND sg13g2_decap_8
XFILLER_27_369 VPWR VGND sg13g2_fill_2
XFILLER_35_380 VPWR VGND sg13g2_decap_8
XFILLER_35_391 VPWR VGND sg13g2_fill_2
XFILLER_11_704 VPWR VGND sg13g2_decap_8
XFILLER_24_57 VPWR VGND sg13g2_decap_8
XFILLER_23_586 VPWR VGND sg13g2_decap_8
XFILLER_24_68 VPWR VGND sg13g2_fill_2
XFILLER_10_236 VPWR VGND sg13g2_fill_1
XFILLER_6_218 VPWR VGND sg13g2_decap_8
XFILLER_40_67 VPWR VGND sg13g2_decap_8
XFILLER_3_936 VPWR VGND sg13g2_decap_8
XFILLER_49_21 VPWR VGND sg13g2_decap_8
XFILLER_46_1002 VPWR VGND sg13g2_decap_8
XFILLER_6_4 VPWR VGND sg13g2_decap_8
XFILLER_49_98 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_19_826 VPWR VGND sg13g2_decap_8
XFILLER_46_645 VPWR VGND sg13g2_decap_8
XFILLER_45_166 VPWR VGND sg13g2_decap_8
XFILLER_33_306 VPWR VGND sg13g2_decap_8
X_425_ net85 _119_ VPWR VGND sg13g2_buf_1
X_356_ net168 VPWR _014_ VGND _166_ _168_ sg13g2_o21ai_1
X_287_ _016_ _166_ _169_ VPWR VGND sg13g2_xnor2_1
XFILLER_5_240 VPWR VGND sg13g2_decap_8
XFILLER_6_796 VPWR VGND sg13g2_decap_8
XFILLER_2_991 VPWR VGND sg13g2_decap_8
XFILLER_49_461 VPWR VGND sg13g2_decap_8
XFILLER_37_623 VPWR VGND sg13g2_decap_8
XFILLER_36_133 VPWR VGND sg13g2_decap_8
XFILLER_18_870 VPWR VGND sg13g2_decap_8
XFILLER_25_818 VPWR VGND sg13g2_decap_8
XFILLER_36_166 VPWR VGND sg13g2_decap_8
XFILLER_17_391 VPWR VGND sg13g2_fill_2
XFILLER_33_884 VPWR VGND sg13g2_decap_8
XFILLER_20_567 VPWR VGND sg13g2_fill_2
XFILLER_9_590 VPWR VGND sg13g2_decap_8
XFILLER_0_917 VPWR VGND sg13g2_decap_8
XFILLER_19_46 VPWR VGND sg13g2_decap_8
XFILLER_28_645 VPWR VGND sg13g2_decap_8
XFILLER_27_166 VPWR VGND sg13g2_decap_8
XFILLER_43_637 VPWR VGND sg13g2_decap_8
XFILLER_15_328 VPWR VGND sg13g2_decap_8
XFILLER_42_158 VPWR VGND sg13g2_fill_1
XFILLER_42_147 VPWR VGND sg13g2_decap_8
XFILLER_23_350 VPWR VGND sg13g2_decap_8
XFILLER_24_873 VPWR VGND sg13g2_decap_8
XFILLER_11_567 VPWR VGND sg13g2_fill_2
XFILLER_7_527 VPWR VGND sg13g2_decap_8
XFILLER_13_1012 VPWR VGND sg13g2_decap_8
XFILLER_3_733 VPWR VGND sg13g2_decap_8
XFILLER_2_210 VPWR VGND sg13g2_fill_1
XFILLER_19_623 VPWR VGND sg13g2_decap_8
XFILLER_47_954 VPWR VGND sg13g2_decap_8
XFILLER_46_442 VPWR VGND sg13g2_decap_8
XFILLER_20_1027 VPWR VGND sg13g2_fill_2
XFILLER_18_155 VPWR VGND sg13g2_decap_8
XFILLER_34_659 VPWR VGND sg13g2_decap_8
XFILLER_14_350 VPWR VGND sg13g2_decap_8
XFILLER_15_895 VPWR VGND sg13g2_decap_8
X_408_ net120 _102_ VPWR VGND sg13g2_buf_1
XFILLER_30_821 VPWR VGND sg13g2_decap_8
X_339_ _199_ net151 net95 VPWR VGND sg13g2_nand2_1
XFILLER_30_898 VPWR VGND sg13g2_decap_8
XFILLER_6_593 VPWR VGND sg13g2_decap_8
XFILLER_2_60 VPWR VGND sg13g2_decap_8
XFILLER_49_280 VPWR VGND sg13g2_decap_8
XFILLER_37_442 VPWR VGND sg13g2_decap_8
XFILLER_38_943 VPWR VGND sg13g2_decap_8
XFILLER_25_615 VPWR VGND sg13g2_decap_8
XFILLER_37_497 VPWR VGND sg13g2_decap_8
XFILLER_24_136 VPWR VGND sg13g2_decap_8
XFILLER_40_607 VPWR VGND sg13g2_decap_8
XFILLER_33_681 VPWR VGND sg13g2_decap_8
XFILLER_36_1023 VPWR VGND sg13g2_decap_4
XFILLER_20_353 VPWR VGND sg13g2_decap_8
XFILLER_21_876 VPWR VGND sg13g2_decap_8
XFILLER_4_519 VPWR VGND sg13g2_decap_8
XFILLER_21_58 VPWR VGND sg13g2_decap_8
XFILLER_0_714 VPWR VGND sg13g2_decap_8
XFILLER_29_910 VPWR VGND sg13g2_decap_8
XFILLER_47_239 VPWR VGND sg13g2_decap_8
XFILLER_44_913 VPWR VGND sg13g2_decap_8
XFILLER_43_401 VPWR VGND sg13g2_decap_8
XFILLER_29_987 VPWR VGND sg13g2_decap_8
XFILLER_15_158 VPWR VGND sg13g2_decap_8
XFILLER_43_478 VPWR VGND sg13g2_fill_2
XFILLER_12_810 VPWR VGND sg13g2_decap_8
XFILLER_24_670 VPWR VGND sg13g2_decap_8
XFILLER_8_803 VPWR VGND sg13g2_decap_8
XFILLER_12_887 VPWR VGND sg13g2_decap_8
XFILLER_7_335 VPWR VGND sg13g2_decap_8
XFILLER_7_49 VPWR VGND sg13g2_decap_8
XFILLER_11_91 VPWR VGND sg13g2_decap_8
Xclkbuf_4_9_0_clk clknet_0_clk clknet_4_9_0_clk VPWR VGND sg13g2_buf_8
XFILLER_39_718 VPWR VGND sg13g2_decap_8
XFILLER_47_751 VPWR VGND sg13g2_decap_8
XFILLER_4_1021 VPWR VGND sg13g2_decap_8
XFILLER_19_497 VPWR VGND sg13g2_decap_8
XFILLER_34_412 VPWR VGND sg13g2_fill_1
XFILLER_35_946 VPWR VGND sg13g2_decap_8
XFILLER_34_456 VPWR VGND sg13g2_decap_8
XFILLER_22_618 VPWR VGND sg13g2_decap_8
XFILLER_15_692 VPWR VGND sg13g2_decap_8
XFILLER_30_695 VPWR VGND sg13g2_decap_8
XFILLER_7_891 VPWR VGND sg13g2_decap_8
XFILLER_29_206 VPWR VGND sg13g2_fill_2
XFILLER_38_740 VPWR VGND sg13g2_decap_8
XFILLER_16_25 VPWR VGND sg13g2_decap_8
XFILLER_25_434 VPWR VGND sg13g2_decap_8
XFILLER_26_957 VPWR VGND sg13g2_decap_8
XFILLER_16_69 VPWR VGND sg13g2_decap_8
XFILLER_41_905 VPWR VGND sg13g2_decap_8
XFILLER_25_489 VPWR VGND sg13g2_decap_8
XFILLER_40_437 VPWR VGND sg13g2_decap_8
XFILLER_21_673 VPWR VGND sg13g2_decap_8
XFILLER_5_806 VPWR VGND sg13g2_decap_8
XFILLER_0_511 VPWR VGND sg13g2_decap_8
XFILLER_0_588 VPWR VGND sg13g2_decap_8
XFILLER_48_548 VPWR VGND sg13g2_decap_8
XFILLER_44_710 VPWR VGND sg13g2_decap_8
XFILLER_17_957 VPWR VGND sg13g2_decap_8
XFILLER_29_784 VPWR VGND sg13g2_decap_8
XFILLER_43_220 VPWR VGND sg13g2_decap_8
XFILLER_44_787 VPWR VGND sg13g2_decap_8
XFILLER_43_275 VPWR VGND sg13g2_decap_8
XFILLER_16_478 VPWR VGND sg13g2_decap_8
XFILLER_31_426 VPWR VGND sg13g2_decap_8
XFILLER_8_600 VPWR VGND sg13g2_decap_8
XFILLER_40_971 VPWR VGND sg13g2_decap_8
XFILLER_7_110 VPWR VGND sg13g2_decap_8
XFILLER_12_684 VPWR VGND sg13g2_decap_8
XFILLER_8_677 VPWR VGND sg13g2_decap_8
XFILLER_7_154 VPWR VGND sg13g2_decap_8
XFILLER_21_4 VPWR VGND sg13g2_decap_8
XFILLER_39_515 VPWR VGND sg13g2_decap_8
XFILLER_34_231 VPWR VGND sg13g2_decap_8
XFILLER_35_743 VPWR VGND sg13g2_decap_8
XFILLER_22_404 VPWR VGND sg13g2_decap_8
XFILLER_31_960 VPWR VGND sg13g2_decap_8
XFILLER_8_81 VPWR VGND sg13g2_decap_8
XFILLER_2_809 VPWR VGND sg13g2_decap_8
XFILLER_45_507 VPWR VGND sg13g2_decap_8
XFILLER_17_209 VPWR VGND sg13g2_decap_8
XFILLER_27_35 VPWR VGND sg13g2_decap_4
XFILLER_14_905 VPWR VGND sg13g2_decap_8
XFILLER_26_754 VPWR VGND sg13g2_decap_8
XFILLER_25_275 VPWR VGND sg13g2_decap_8
XFILLER_41_702 VPWR VGND sg13g2_decap_8
XFILLER_43_56 VPWR VGND sg13g2_decap_8
XFILLER_41_779 VPWR VGND sg13g2_decap_8
XFILLER_22_982 VPWR VGND sg13g2_decap_8
XFILLER_5_603 VPWR VGND sg13g2_decap_8
XFILLER_49_1000 VPWR VGND sg13g2_decap_8
XFILLER_4_124 VPWR VGND sg13g2_fill_2
XFILLER_4_113 VPWR VGND sg13g2_decap_8
XFILLER_1_864 VPWR VGND sg13g2_decap_8
XFILLER_49_846 VPWR VGND sg13g2_decap_8
XFILLER_48_323 VPWR VGND sg13g2_decap_8
XFILLER_0_385 VPWR VGND sg13g2_decap_8
XFILLER_29_581 VPWR VGND sg13g2_decap_8
XFILLER_16_231 VPWR VGND sg13g2_fill_2
XFILLER_17_754 VPWR VGND sg13g2_decap_8
XFILLER_44_584 VPWR VGND sg13g2_decap_8
X_587_ net67 VGND VPWR net106 mac2.sum_lvl2_ff\[4\] clknet_5_12__leaf_clk sg13g2_dfrbpq_1
XFILLER_31_201 VPWR VGND sg13g2_decap_8
XFILLER_20_908 VPWR VGND sg13g2_decap_8
XFILLER_32_757 VPWR VGND sg13g2_decap_8
XFILLER_8_430 VPWR VGND sg13g2_decap_8
XFILLER_31_278 VPWR VGND sg13g2_decap_8
XFILLER_9_975 VPWR VGND sg13g2_decap_8
XFILLER_3_190 VPWR VGND sg13g2_decap_4
XFILLER_27_518 VPWR VGND sg13g2_decap_8
XFILLER_35_540 VPWR VGND sg13g2_decap_8
XFILLER_22_212 VPWR VGND sg13g2_decap_8
XFILLER_23_768 VPWR VGND sg13g2_decap_8
XFILLER_10_418 VPWR VGND sg13g2_decap_8
XFILLER_2_606 VPWR VGND sg13g2_decap_8
XFILLER_1_105 VPWR VGND sg13g2_decap_8
XFILLER_38_78 VPWR VGND sg13g2_decap_8
XFILLER_46_827 VPWR VGND sg13g2_decap_8
X_510_ net68 VGND VPWR _132_ DP_4.matrix\[64\] clknet_5_10__leaf_clk sg13g2_dfrbpq_1
X_441_ net50 _135_ VPWR VGND sg13g2_buf_1
XFILLER_14_702 VPWR VGND sg13g2_decap_8
XFILLER_26_551 VPWR VGND sg13g2_decap_8
X_372_ _220_ net133 net82 VPWR VGND sg13g2_nand2_1
XFILLER_14_779 VPWR VGND sg13g2_decap_8
XFILLER_41_576 VPWR VGND sg13g2_decap_8
XFILLER_9_249 VPWR VGND sg13g2_decap_8
XFILLER_10_930 VPWR VGND sg13g2_decap_8
XFILLER_13_289 VPWR VGND sg13g2_decap_8
XFILLER_6_901 VPWR VGND sg13g2_decap_8
XFILLER_6_978 VPWR VGND sg13g2_decap_8
XFILLER_5_499 VPWR VGND sg13g2_decap_8
XFILLER_1_661 VPWR VGND sg13g2_decap_8
XFILLER_49_643 VPWR VGND sg13g2_decap_8
XFILLER_48_131 VPWR VGND sg13g2_decap_8
XFILLER_0_182 VPWR VGND sg13g2_decap_8
XFILLER_37_805 VPWR VGND sg13g2_decap_8
XFILLER_36_315 VPWR VGND sg13g2_decap_8
XFILLER_36_348 VPWR VGND sg13g2_decap_8
XFILLER_45_871 VPWR VGND sg13g2_decap_8
XFILLER_20_705 VPWR VGND sg13g2_decap_8
XFILLER_32_554 VPWR VGND sg13g2_decap_8
XFILLER_9_772 VPWR VGND sg13g2_decap_8
XFILLER_8_260 VPWR VGND sg13g2_decap_8
XFILLER_5_93 VPWR VGND sg13g2_decap_8
XFILLER_28_827 VPWR VGND sg13g2_decap_8
XFILLER_43_819 VPWR VGND sg13g2_decap_8
XFILLER_42_329 VPWR VGND sg13g2_decap_8
XFILLER_23_565 VPWR VGND sg13g2_fill_2
XFILLER_10_215 VPWR VGND sg13g2_decap_8
XFILLER_7_709 VPWR VGND sg13g2_decap_8
XFILLER_40_46 VPWR VGND sg13g2_decap_8
XFILLER_3_915 VPWR VGND sg13g2_decap_8
XFILLER_2_458 VPWR VGND sg13g2_decap_4
XFILLER_49_77 VPWR VGND sg13g2_decap_8
XFILLER_19_805 VPWR VGND sg13g2_decap_8
XFILLER_46_624 VPWR VGND sg13g2_decap_8
XFILLER_18_326 VPWR VGND sg13g2_decap_8
XFILLER_45_145 VPWR VGND sg13g2_decap_8
XFILLER_27_882 VPWR VGND sg13g2_decap_8
XFILLER_14_532 VPWR VGND sg13g2_decap_8
X_424_ net137 _118_ VPWR VGND sg13g2_buf_1
XFILLER_42_885 VPWR VGND sg13g2_decap_8
XFILLER_14_598 VPWR VGND sg13g2_decap_8
X_355_ _209_ _208_ _057_ VPWR VGND sg13g2_xor2_1
XFILLER_41_373 VPWR VGND sg13g2_decap_8
X_286_ mac1.sum_lvl3_ff\[1\] net167 _169_ VPWR VGND sg13g2_xor2_1
XFILLER_6_775 VPWR VGND sg13g2_decap_8
Xclkbuf_5_14__f_clk clknet_4_7_0_clk clknet_5_14__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_2_970 VPWR VGND sg13g2_decap_8
XFILLER_49_440 VPWR VGND sg13g2_decap_8
XFILLER_37_602 VPWR VGND sg13g2_decap_8
XFILLER_36_112 VPWR VGND sg13g2_decap_8
XFILLER_37_679 VPWR VGND sg13g2_decap_8
XFILLER_17_370 VPWR VGND sg13g2_decap_8
XFILLER_33_863 VPWR VGND sg13g2_decap_8
XFILLER_20_546 VPWR VGND sg13g2_decap_8
XFILLER_32_395 VPWR VGND sg13g2_decap_8
XFILLER_20_579 VPWR VGND sg13g2_decap_8
XFILLER_19_25 VPWR VGND sg13g2_decap_8
XFILLER_28_624 VPWR VGND sg13g2_decap_8
XFILLER_43_616 VPWR VGND sg13g2_decap_8
XFILLER_27_145 VPWR VGND sg13g2_fill_1
XFILLER_42_126 VPWR VGND sg13g2_decap_8
XFILLER_35_35 VPWR VGND sg13g2_fill_2
XFILLER_24_852 VPWR VGND sg13g2_decap_8
XFILLER_35_79 VPWR VGND sg13g2_decap_4
XFILLER_7_506 VPWR VGND sg13g2_decap_8
XFILLER_11_535 VPWR VGND sg13g2_decap_4
XFILLER_3_712 VPWR VGND sg13g2_decap_8
XFILLER_3_789 VPWR VGND sg13g2_decap_8
XFILLER_2_277 VPWR VGND sg13g2_fill_1
XFILLER_47_933 VPWR VGND sg13g2_decap_8
XFILLER_19_602 VPWR VGND sg13g2_decap_8
XFILLER_46_421 VPWR VGND sg13g2_decap_8
XFILLER_18_134 VPWR VGND sg13g2_decap_8
XFILLER_20_1006 VPWR VGND sg13g2_decap_8
XFILLER_19_679 VPWR VGND sg13g2_decap_8
XFILLER_46_498 VPWR VGND sg13g2_decap_8
XFILLER_34_638 VPWR VGND sg13g2_decap_8
XFILLER_42_682 VPWR VGND sg13g2_decap_8
XFILLER_15_874 VPWR VGND sg13g2_decap_8
X_407_ net95 _101_ VPWR VGND sg13g2_buf_1
XFILLER_30_800 VPWR VGND sg13g2_decap_8
X_338_ _198_ net48 net140 VPWR VGND sg13g2_nand2_1
XFILLER_41_181 VPWR VGND sg13g2_decap_8
XFILLER_30_877 VPWR VGND sg13g2_decap_8
X_269_ _007_ _158_ net194 VPWR VGND sg13g2_xnor2_1
XFILLER_6_572 VPWR VGND sg13g2_decap_8
XFILLER_38_922 VPWR VGND sg13g2_decap_8
XFILLER_37_421 VPWR VGND sg13g2_decap_8
XFILLER_37_476 VPWR VGND sg13g2_decap_8
XFILLER_38_999 VPWR VGND sg13g2_decap_8
XFILLER_24_104 VPWR VGND sg13g2_decap_8
XFILLER_36_1002 VPWR VGND sg13g2_decap_8
XFILLER_33_660 VPWR VGND sg13g2_decap_8
XFILLER_21_855 VPWR VGND sg13g2_decap_8
XFILLER_29_966 VPWR VGND sg13g2_decap_8
XFILLER_16_649 VPWR VGND sg13g2_decap_8
XFILLER_28_487 VPWR VGND sg13g2_decap_8
XFILLER_44_969 VPWR VGND sg13g2_decap_8
XFILLER_43_457 VPWR VGND sg13g2_decap_8
XFILLER_15_137 VPWR VGND sg13g2_decap_8
XFILLER_11_321 VPWR VGND sg13g2_decap_8
XFILLER_7_314 VPWR VGND sg13g2_decap_8
XFILLER_7_28 VPWR VGND sg13g2_decap_8
XFILLER_12_866 VPWR VGND sg13g2_decap_8
XFILLER_8_859 VPWR VGND sg13g2_decap_8
XFILLER_3_586 VPWR VGND sg13g2_decap_8
XFILLER_4_1000 VPWR VGND sg13g2_decap_8
XFILLER_47_730 VPWR VGND sg13g2_decap_8
XFILLER_19_476 VPWR VGND sg13g2_decap_8
XFILLER_35_925 VPWR VGND sg13g2_decap_8
XFILLER_43_980 VPWR VGND sg13g2_decap_8
XFILLER_15_671 VPWR VGND sg13g2_decap_8
XFILLER_14_181 VPWR VGND sg13g2_fill_1
XFILLER_30_674 VPWR VGND sg13g2_decap_8
XFILLER_7_870 VPWR VGND sg13g2_decap_8
XFILLER_42_0 VPWR VGND sg13g2_decap_8
XFILLER_37_251 VPWR VGND sg13g2_decap_8
XFILLER_25_413 VPWR VGND sg13g2_decap_4
XFILLER_26_936 VPWR VGND sg13g2_decap_8
XFILLER_38_796 VPWR VGND sg13g2_decap_8
XFILLER_37_295 VPWR VGND sg13g2_decap_8
XFILLER_40_416 VPWR VGND sg13g2_decap_8
XFILLER_20_140 VPWR VGND sg13g2_decap_4
XFILLER_21_652 VPWR VGND sg13g2_decap_8
XFILLER_32_14 VPWR VGND sg13g2_decap_4
XFILLER_4_339 VPWR VGND sg13g2_decap_8
XFILLER_48_527 VPWR VGND sg13g2_decap_8
XFILLER_0_567 VPWR VGND sg13g2_decap_8
XFILLER_29_763 VPWR VGND sg13g2_decap_8
XFILLER_17_936 VPWR VGND sg13g2_decap_8
XFILLER_44_766 VPWR VGND sg13g2_decap_8
XFILLER_16_457 VPWR VGND sg13g2_decap_8
XFILLER_28_295 VPWR VGND sg13g2_decap_8
XFILLER_31_405 VPWR VGND sg13g2_decap_8
XFILLER_32_939 VPWR VGND sg13g2_decap_8
XFILLER_31_449 VPWR VGND sg13g2_decap_8
XFILLER_12_663 VPWR VGND sg13g2_decap_8
XFILLER_40_950 VPWR VGND sg13g2_decap_8
XFILLER_8_656 VPWR VGND sg13g2_decap_8
XFILLER_7_133 VPWR VGND sg13g2_decap_8
XFILLER_11_184 VPWR VGND sg13g2_decap_8
XFILLER_4_895 VPWR VGND sg13g2_decap_8
XFILLER_3_394 VPWR VGND sg13g2_decap_8
XFILLER_14_4 VPWR VGND sg13g2_decap_8
XFILLER_19_284 VPWR VGND sg13g2_decap_8
XFILLER_35_722 VPWR VGND sg13g2_decap_8
XFILLER_34_210 VPWR VGND sg13g2_decap_8
XFILLER_35_799 VPWR VGND sg13g2_decap_8
XFILLER_15_490 VPWR VGND sg13g2_decap_8
XFILLER_34_287 VPWR VGND sg13g2_decap_4
XFILLER_8_60 VPWR VGND sg13g2_decap_8
XFILLER_30_471 VPWR VGND sg13g2_fill_2
XFILLER_27_14 VPWR VGND sg13g2_decap_8
XFILLER_27_58 VPWR VGND sg13g2_decap_8
XFILLER_26_733 VPWR VGND sg13g2_decap_8
XFILLER_38_593 VPWR VGND sg13g2_decap_8
XFILLER_25_254 VPWR VGND sg13g2_decap_8
XFILLER_40_202 VPWR VGND sg13g2_decap_8
XFILLER_43_35 VPWR VGND sg13g2_decap_8
Xclkbuf_4_8_0_clk clknet_0_clk clknet_4_8_0_clk VPWR VGND sg13g2_buf_8
XFILLER_41_758 VPWR VGND sg13g2_decap_8
XFILLER_22_961 VPWR VGND sg13g2_decap_8
XFILLER_40_257 VPWR VGND sg13g2_decap_8
XFILLER_21_482 VPWR VGND sg13g2_decap_8
XFILLER_5_659 VPWR VGND sg13g2_decap_8
XFILLER_4_158 VPWR VGND sg13g2_decap_4
XFILLER_4_18 VPWR VGND sg13g2_decap_8
XFILLER_1_843 VPWR VGND sg13g2_decap_8
XFILLER_49_825 VPWR VGND sg13g2_decap_8
XFILLER_48_302 VPWR VGND sg13g2_decap_8
XFILLER_0_364 VPWR VGND sg13g2_decap_8
XFILLER_1_1025 VPWR VGND sg13g2_decap_4
XFILLER_29_560 VPWR VGND sg13g2_decap_8
XFILLER_36_519 VPWR VGND sg13g2_decap_8
XFILLER_16_210 VPWR VGND sg13g2_decap_8
XFILLER_17_733 VPWR VGND sg13g2_decap_8
XFILLER_44_563 VPWR VGND sg13g2_decap_8
X_586_ net79 VGND VPWR _069_ mac2.products_ff\[17\] clknet_5_27__leaf_clk sg13g2_dfrbpq_1
XFILLER_16_254 VPWR VGND sg13g2_decap_8
XFILLER_32_736 VPWR VGND sg13g2_decap_8
XFILLER_9_954 VPWR VGND sg13g2_decap_8
XFILLER_8_486 VPWR VGND sg13g2_decap_8
XFILLER_4_692 VPWR VGND sg13g2_decap_8
XFILLER_39_302 VPWR VGND sg13g2_decap_8
XFILLER_48_891 VPWR VGND sg13g2_decap_8
XFILLER_23_747 VPWR VGND sg13g2_decap_8
XFILLER_35_596 VPWR VGND sg13g2_decap_8
XFILLER_30_290 VPWR VGND sg13g2_decap_8
XFILLER_46_806 VPWR VGND sg13g2_decap_8
XFILLER_38_57 VPWR VGND sg13g2_decap_8
XFILLER_45_327 VPWR VGND sg13g2_fill_2
XFILLER_18_519 VPWR VGND sg13g2_decap_8
XFILLER_45_349 VPWR VGND sg13g2_decap_8
X_440_ net144 _134_ VPWR VGND sg13g2_buf_1
X_371_ _219_ _218_ _067_ VPWR VGND sg13g2_xor2_1
XFILLER_14_758 VPWR VGND sg13g2_decap_8
XFILLER_41_555 VPWR VGND sg13g2_decap_8
XFILLER_10_986 VPWR VGND sg13g2_decap_8
XFILLER_6_957 VPWR VGND sg13g2_decap_8
XFILLER_5_478 VPWR VGND sg13g2_decap_8
XFILLER_1_640 VPWR VGND sg13g2_decap_8
XFILLER_49_622 VPWR VGND sg13g2_decap_8
XFILLER_48_110 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_49_699 VPWR VGND sg13g2_decap_8
XFILLER_45_850 VPWR VGND sg13g2_decap_8
XFILLER_44_371 VPWR VGND sg13g2_decap_8
XFILLER_32_533 VPWR VGND sg13g2_decap_8
X_569_ net57 VGND VPWR _036_ mac2.products_ff\[128\] clknet_5_0__leaf_clk sg13g2_dfrbpq_1
XFILLER_9_751 VPWR VGND sg13g2_decap_8
XFILLER_5_61 VPWR VGND sg13g2_decap_4
XFILLER_28_806 VPWR VGND sg13g2_decap_8
XFILLER_39_143 VPWR VGND sg13g2_decap_8
XFILLER_27_305 VPWR VGND sg13g2_decap_8
XFILLER_27_316 VPWR VGND sg13g2_fill_2
XFILLER_42_308 VPWR VGND sg13g2_decap_8
XFILLER_23_500 VPWR VGND sg13g2_fill_1
XFILLER_36_883 VPWR VGND sg13g2_decap_8
XFILLER_23_544 VPWR VGND sg13g2_decap_8
XFILLER_11_739 VPWR VGND sg13g2_decap_8
XFILLER_40_14 VPWR VGND sg13g2_decap_8
XFILLER_49_56 VPWR VGND sg13g2_decap_8
XFILLER_46_603 VPWR VGND sg13g2_decap_8
XFILLER_18_305 VPWR VGND sg13g2_decap_8
XFILLER_45_124 VPWR VGND sg13g2_decap_8
XFILLER_27_861 VPWR VGND sg13g2_decap_8
X_423_ net52 _117_ VPWR VGND sg13g2_buf_1
XFILLER_26_382 VPWR VGND sg13g2_decap_8
XFILLER_42_864 VPWR VGND sg13g2_decap_8
XFILLER_14_577 VPWR VGND sg13g2_decap_8
X_354_ _209_ net128 net49 VPWR VGND sg13g2_nand2_1
X_285_ net167 mac1.sum_lvl3_ff\[1\] _168_ VPWR VGND sg13g2_nor2_1
XFILLER_14_81 VPWR VGND sg13g2_decap_8
XFILLER_10_783 VPWR VGND sg13g2_decap_8
XFILLER_6_754 VPWR VGND sg13g2_decap_8
XFILLER_46_7 VPWR VGND sg13g2_decap_8
XFILLER_30_91 VPWR VGND sg13g2_decap_8
XFILLER_49_496 VPWR VGND sg13g2_decap_8
XFILLER_37_658 VPWR VGND sg13g2_decap_8
XFILLER_17_393 VPWR VGND sg13g2_fill_1
XFILLER_33_842 VPWR VGND sg13g2_decap_8
XFILLER_32_374 VPWR VGND sg13g2_decap_8
XFILLER_20_525 VPWR VGND sg13g2_decap_8
XFILLER_20_569 VPWR VGND sg13g2_fill_1
XFILLER_28_603 VPWR VGND sg13g2_decap_8
XFILLER_27_124 VPWR VGND sg13g2_decap_4
XFILLER_35_14 VPWR VGND sg13g2_decap_8
XFILLER_24_831 VPWR VGND sg13g2_decap_8
XFILLER_35_58 VPWR VGND sg13g2_decap_8
XFILLER_36_680 VPWR VGND sg13g2_decap_8
Xclkbuf_5_20__f_clk clknet_4_10_0_clk clknet_5_20__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_3_768 VPWR VGND sg13g2_decap_8
XFILLER_47_912 VPWR VGND sg13g2_decap_8
XFILLER_46_400 VPWR VGND sg13g2_decap_8
XFILLER_18_113 VPWR VGND sg13g2_decap_8
XFILLER_19_658 VPWR VGND sg13g2_decap_8
XFILLER_47_989 VPWR VGND sg13g2_decap_8
XFILLER_46_477 VPWR VGND sg13g2_decap_8
XFILLER_34_617 VPWR VGND sg13g2_decap_8
XFILLER_15_853 VPWR VGND sg13g2_decap_8
XFILLER_26_190 VPWR VGND sg13g2_decap_8
XFILLER_33_149 VPWR VGND sg13g2_decap_8
XFILLER_42_661 VPWR VGND sg13g2_decap_8
X_406_ net140 _100_ VPWR VGND sg13g2_buf_1
XFILLER_25_80 VPWR VGND sg13g2_decap_8
XFILLER_14_385 VPWR VGND sg13g2_decap_8
XFILLER_30_856 VPWR VGND sg13g2_decap_8
X_337_ _197_ _196_ _045_ VPWR VGND sg13g2_xor2_1
X_268_ net193 mac1.products_ff\[113\] _159_ VPWR VGND sg13g2_xor2_1
XFILLER_38_901 VPWR VGND sg13g2_decap_8
XFILLER_2_95 VPWR VGND sg13g2_decap_8
XFILLER_38_978 VPWR VGND sg13g2_decap_8
XFILLER_21_834 VPWR VGND sg13g2_decap_8
XFILLER_32_160 VPWR VGND sg13g2_decap_4
XFILLER_32_193 VPWR VGND sg13g2_decap_8
XFILLER_20_344 VPWR VGND sg13g2_fill_1
XFILLER_20_388 VPWR VGND sg13g2_decap_8
XFILLER_48_709 VPWR VGND sg13g2_decap_8
XFILLER_0_749 VPWR VGND sg13g2_decap_8
XFILLER_29_945 VPWR VGND sg13g2_decap_8
XFILLER_46_35 VPWR VGND sg13g2_decap_8
XFILLER_28_444 VPWR VGND sg13g2_decap_8
XFILLER_28_466 VPWR VGND sg13g2_decap_8
XFILLER_44_948 VPWR VGND sg13g2_decap_8
XFILLER_15_116 VPWR VGND sg13g2_decap_8
XFILLER_16_628 VPWR VGND sg13g2_decap_8
XFILLER_43_436 VPWR VGND sg13g2_decap_8
XFILLER_30_119 VPWR VGND sg13g2_decap_8
XFILLER_11_300 VPWR VGND sg13g2_decap_8
XFILLER_12_845 VPWR VGND sg13g2_decap_8
XFILLER_8_838 VPWR VGND sg13g2_decap_8
XFILLER_3_543 VPWR VGND sg13g2_decap_4
XFILLER_3_565 VPWR VGND sg13g2_decap_8
XFILLER_19_422 VPWR VGND sg13g2_decap_4
XFILLER_19_455 VPWR VGND sg13g2_decap_8
XFILLER_35_904 VPWR VGND sg13g2_decap_8
XFILLER_47_786 VPWR VGND sg13g2_decap_8
XFILLER_34_403 VPWR VGND sg13g2_decap_8
XFILLER_46_296 VPWR VGND sg13g2_decap_8
XFILLER_15_650 VPWR VGND sg13g2_decap_8
XFILLER_30_653 VPWR VGND sg13g2_decap_8
XFILLER_35_0 VPWR VGND sg13g2_decap_8
XFILLER_26_915 VPWR VGND sg13g2_decap_8
XFILLER_38_775 VPWR VGND sg13g2_decap_8
XFILLER_37_274 VPWR VGND sg13g2_decap_8
XFILLER_34_981 VPWR VGND sg13g2_decap_8
XFILLER_12_119 VPWR VGND sg13g2_decap_4
XFILLER_21_631 VPWR VGND sg13g2_decap_8
XFILLER_20_185 VPWR VGND sg13g2_fill_1
XFILLER_10_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_546 VPWR VGND sg13g2_decap_8
XFILLER_48_506 VPWR VGND sg13g2_decap_8
XFILLER_29_742 VPWR VGND sg13g2_decap_8
XFILLER_17_915 VPWR VGND sg13g2_decap_8
XFILLER_28_252 VPWR VGND sg13g2_decap_8
XFILLER_44_745 VPWR VGND sg13g2_decap_8
XFILLER_16_425 VPWR VGND sg13g2_fill_2
XFILLER_16_436 VPWR VGND sg13g2_decap_8
XFILLER_32_918 VPWR VGND sg13g2_decap_8
XFILLER_12_620 VPWR VGND sg13g2_decap_4
XFILLER_12_642 VPWR VGND sg13g2_decap_8
XFILLER_8_635 VPWR VGND sg13g2_decap_8
XFILLER_11_163 VPWR VGND sg13g2_decap_8
XFILLER_4_874 VPWR VGND sg13g2_decap_8
XFILLER_3_373 VPWR VGND sg13g2_decap_8
XFILLER_26_1013 VPWR VGND sg13g2_decap_8
XFILLER_19_241 VPWR VGND sg13g2_decap_8
XFILLER_47_583 VPWR VGND sg13g2_decap_8
XFILLER_35_701 VPWR VGND sg13g2_decap_8
XFILLER_23_929 VPWR VGND sg13g2_decap_8
XFILLER_34_266 VPWR VGND sg13g2_decap_8
XFILLER_35_778 VPWR VGND sg13g2_decap_8
XFILLER_16_992 VPWR VGND sg13g2_decap_8
XFILLER_33_1017 VPWR VGND sg13g2_decap_8
XFILLER_30_461 VPWR VGND sg13g2_decap_4
XFILLER_31_995 VPWR VGND sg13g2_decap_8
XFILLER_33_1028 VPWR VGND sg13g2_fill_1
XFILLER_26_712 VPWR VGND sg13g2_decap_8
XFILLER_38_572 VPWR VGND sg13g2_decap_8
XFILLER_43_14 VPWR VGND sg13g2_decap_8
XFILLER_26_789 VPWR VGND sg13g2_decap_8
XFILLER_13_428 VPWR VGND sg13g2_fill_2
XFILLER_25_299 VPWR VGND sg13g2_decap_8
XFILLER_41_737 VPWR VGND sg13g2_decap_8
XFILLER_22_940 VPWR VGND sg13g2_decap_8
XFILLER_21_450 VPWR VGND sg13g2_decap_8
XFILLER_21_461 VPWR VGND sg13g2_fill_1
XFILLER_5_638 VPWR VGND sg13g2_decap_8
XFILLER_4_137 VPWR VGND sg13g2_decap_8
XFILLER_1_822 VPWR VGND sg13g2_decap_8
XFILLER_49_804 VPWR VGND sg13g2_decap_8
XFILLER_0_343 VPWR VGND sg13g2_decap_8
XFILLER_1_899 VPWR VGND sg13g2_decap_8
XFILLER_48_358 VPWR VGND sg13g2_fill_2
XFILLER_1_1004 VPWR VGND sg13g2_decap_8
XFILLER_17_712 VPWR VGND sg13g2_decap_8
XFILLER_44_542 VPWR VGND sg13g2_decap_8
XFILLER_17_789 VPWR VGND sg13g2_decap_8
XFILLER_32_715 VPWR VGND sg13g2_decap_8
X_585_ net79 VGND VPWR _068_ mac2.products_ff\[16\] clknet_5_26__leaf_clk sg13g2_dfrbpq_1
XFILLER_16_288 VPWR VGND sg13g2_decap_8
XFILLER_9_933 VPWR VGND sg13g2_decap_8
XFILLER_12_472 VPWR VGND sg13g2_decap_8
XFILLER_13_984 VPWR VGND sg13g2_decap_8
XFILLER_8_465 VPWR VGND sg13g2_decap_8
XFILLER_4_671 VPWR VGND sg13g2_decap_8
XFILLER_48_870 VPWR VGND sg13g2_decap_8
XFILLER_35_575 VPWR VGND sg13g2_decap_8
Xclkbuf_5_1__f_clk clknet_4_0_0_clk clknet_5_1__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_23_726 VPWR VGND sg13g2_decap_8
XFILLER_22_247 VPWR VGND sg13g2_decap_8
XFILLER_13_39 VPWR VGND sg13g2_decap_8
XFILLER_31_792 VPWR VGND sg13g2_decap_8
XFILLER_38_14 VPWR VGND sg13g2_decap_8
XFILLER_45_317 VPWR VGND sg13g2_fill_2
XFILLER_38_391 VPWR VGND sg13g2_decap_8
X_370_ _219_ net163 net54 VPWR VGND sg13g2_nand2_1
XFILLER_14_737 VPWR VGND sg13g2_decap_8
XFILLER_26_586 VPWR VGND sg13g2_decap_8
XFILLER_41_534 VPWR VGND sg13g2_decap_8
XFILLER_9_207 VPWR VGND sg13g2_decap_8
XFILLER_13_236 VPWR VGND sg13g2_decap_8
XFILLER_13_247 VPWR VGND sg13g2_fill_1
XFILLER_6_936 VPWR VGND sg13g2_decap_8
XFILLER_5_402 VPWR VGND sg13g2_fill_2
XFILLER_10_965 VPWR VGND sg13g2_decap_8
XFILLER_5_457 VPWR VGND sg13g2_decap_8
XFILLER_49_601 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_1_696 VPWR VGND sg13g2_decap_8
XFILLER_23_1027 VPWR VGND sg13g2_fill_2
XFILLER_49_678 VPWR VGND sg13g2_decap_8
XFILLER_48_166 VPWR VGND sg13g2_decap_8
XFILLER_44_350 VPWR VGND sg13g2_decap_8
XFILLER_17_564 VPWR VGND sg13g2_fill_2
XFILLER_17_575 VPWR VGND sg13g2_fill_2
XFILLER_32_512 VPWR VGND sg13g2_decap_8
X_568_ net77 VGND VPWR net185 mac2.sum_lvl1_ff\[9\] clknet_5_15__leaf_clk sg13g2_dfrbpq_1
X_499_ net64 VGND VPWR _121_ DP_3.matrix\[113\] clknet_5_2__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_589 VPWR VGND sg13g2_decap_8
XFILLER_9_730 VPWR VGND sg13g2_decap_8
XFILLER_13_781 VPWR VGND sg13g2_decap_8
XFILLER_12_291 VPWR VGND sg13g2_decap_8
XFILLER_8_295 VPWR VGND sg13g2_decap_8
Xclkbuf_4_7_0_clk clknet_0_clk clknet_4_7_0_clk VPWR VGND sg13g2_buf_8
XFILLER_39_122 VPWR VGND sg13g2_decap_8
XFILLER_39_188 VPWR VGND sg13g2_decap_8
XFILLER_36_862 VPWR VGND sg13g2_decap_8
XFILLER_39_1012 VPWR VGND sg13g2_decap_8
XFILLER_11_718 VPWR VGND sg13g2_decap_8
XFILLER_23_567 VPWR VGND sg13g2_fill_1
XFILLER_49_35 VPWR VGND sg13g2_decap_8
XFILLER_46_1027 VPWR VGND sg13g2_fill_2
XFILLER_46_1016 VPWR VGND sg13g2_decap_8
XFILLER_46_659 VPWR VGND sg13g2_decap_8
XFILLER_45_103 VPWR VGND sg13g2_decap_8
XFILLER_27_840 VPWR VGND sg13g2_decap_8
X_422_ net138 _116_ VPWR VGND sg13g2_buf_1
XFILLER_26_361 VPWR VGND sg13g2_decap_8
XFILLER_42_843 VPWR VGND sg13g2_decap_8
XFILLER_41_342 VPWR VGND sg13g2_decap_4
X_353_ _208_ net40 net135 VPWR VGND sg13g2_nand2_1
X_284_ _167_ net167 mac1.sum_lvl3_ff\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_14_60 VPWR VGND sg13g2_decap_8
XFILLER_10_762 VPWR VGND sg13g2_decap_8
XFILLER_6_733 VPWR VGND sg13g2_decap_8
XFILLER_5_254 VPWR VGND sg13g2_decap_8
XFILLER_30_70 VPWR VGND sg13g2_decap_8
XFILLER_7_1010 VPWR VGND sg13g2_decap_8
XFILLER_39_7 VPWR VGND sg13g2_decap_8
XFILLER_1_493 VPWR VGND sg13g2_decap_8
XFILLER_49_475 VPWR VGND sg13g2_decap_8
XFILLER_37_637 VPWR VGND sg13g2_decap_8
XFILLER_24_309 VPWR VGND sg13g2_decap_8
XFILLER_36_147 VPWR VGND sg13g2_decap_8
XFILLER_18_884 VPWR VGND sg13g2_decap_8
XFILLER_33_821 VPWR VGND sg13g2_decap_8
XFILLER_44_180 VPWR VGND sg13g2_decap_8
XFILLER_20_504 VPWR VGND sg13g2_decap_8
XFILLER_32_353 VPWR VGND sg13g2_decap_8
XFILLER_33_898 VPWR VGND sg13g2_decap_8
XFILLER_9_571 VPWR VGND sg13g2_fill_1
XFILLER_10_18 VPWR VGND sg13g2_decap_4
XFILLER_28_659 VPWR VGND sg13g2_decap_8
XFILLER_24_810 VPWR VGND sg13g2_decap_8
XFILLER_23_364 VPWR VGND sg13g2_decap_8
XFILLER_24_887 VPWR VGND sg13g2_decap_8
XFILLER_13_1026 VPWR VGND sg13g2_fill_2
XFILLER_4_4 VPWR VGND sg13g2_decap_8
XFILLER_3_747 VPWR VGND sg13g2_decap_8
XFILLER_19_637 VPWR VGND sg13g2_decap_8
XFILLER_47_968 VPWR VGND sg13g2_decap_8
XFILLER_46_456 VPWR VGND sg13g2_decap_8
XFILLER_18_169 VPWR VGND sg13g2_decap_8
XFILLER_42_640 VPWR VGND sg13g2_decap_8
XFILLER_15_832 VPWR VGND sg13g2_decap_8
XFILLER_14_364 VPWR VGND sg13g2_decap_8
X_405_ net84 _099_ VPWR VGND sg13g2_buf_1
XFILLER_30_835 VPWR VGND sg13g2_decap_8
X_336_ _197_ net146 net51 VPWR VGND sg13g2_nand2_1
XFILLER_41_161 VPWR VGND sg13g2_decap_8
X_267_ _158_ mac1.products_ff\[112\] net37 VPWR VGND sg13g2_nand2_1
XFILLER_29_1022 VPWR VGND sg13g2_decap_8
XFILLER_1_290 VPWR VGND sg13g2_decap_8
XFILLER_2_74 VPWR VGND sg13g2_decap_8
XFILLER_38_957 VPWR VGND sg13g2_decap_8
XFILLER_49_294 VPWR VGND sg13g2_decap_8
XFILLER_18_681 VPWR VGND sg13g2_decap_8
XFILLER_25_629 VPWR VGND sg13g2_decap_8
XFILLER_21_813 VPWR VGND sg13g2_decap_8
XFILLER_20_301 VPWR VGND sg13g2_decap_8
XFILLER_32_172 VPWR VGND sg13g2_decap_8
XFILLER_33_695 VPWR VGND sg13g2_decap_8
XFILLER_20_367 VPWR VGND sg13g2_decap_8
XFILLER_0_728 VPWR VGND sg13g2_decap_8
XFILLER_43_1008 VPWR VGND sg13g2_decap_8
XFILLER_46_14 VPWR VGND sg13g2_decap_8
XFILLER_28_423 VPWR VGND sg13g2_decap_8
XFILLER_29_924 VPWR VGND sg13g2_decap_8
XFILLER_16_607 VPWR VGND sg13g2_decap_8
XFILLER_46_69 VPWR VGND sg13g2_decap_8
XFILLER_44_927 VPWR VGND sg13g2_decap_8
XFILLER_43_415 VPWR VGND sg13g2_decap_8
XFILLER_12_824 VPWR VGND sg13g2_decap_8
XFILLER_23_183 VPWR VGND sg13g2_decap_8
XFILLER_24_684 VPWR VGND sg13g2_decap_8
XFILLER_8_817 VPWR VGND sg13g2_decap_8
XFILLER_11_378 VPWR VGND sg13g2_fill_2
XFILLER_3_522 VPWR VGND sg13g2_decap_8
XFILLER_47_765 VPWR VGND sg13g2_decap_8
XFILLER_46_275 VPWR VGND sg13g2_decap_8
XFILLER_36_91 VPWR VGND sg13g2_decap_8
XFILLER_14_172 VPWR VGND sg13g2_decap_8
XFILLER_30_632 VPWR VGND sg13g2_decap_8
X_319_ _186_ net155 net43 VPWR VGND sg13g2_nand2_1
XFILLER_38_754 VPWR VGND sg13g2_decap_8
XFILLER_25_448 VPWR VGND sg13g2_decap_8
XFILLER_25_459 VPWR VGND sg13g2_fill_1
XFILLER_34_960 VPWR VGND sg13g2_decap_8
XFILLER_41_919 VPWR VGND sg13g2_decap_8
XFILLER_21_610 VPWR VGND sg13g2_decap_8
XFILLER_33_492 VPWR VGND sg13g2_decap_8
XFILLER_21_687 VPWR VGND sg13g2_decap_8
XFILLER_10_1007 VPWR VGND sg13g2_decap_8
XFILLER_0_525 VPWR VGND sg13g2_decap_8
XFILLER_29_721 VPWR VGND sg13g2_decap_8
XFILLER_28_231 VPWR VGND sg13g2_decap_8
XFILLER_44_724 VPWR VGND sg13g2_decap_8
XFILLER_29_798 VPWR VGND sg13g2_decap_8
XFILLER_43_234 VPWR VGND sg13g2_decap_8
XFILLER_43_289 VPWR VGND sg13g2_decap_8
XFILLER_12_610 VPWR VGND sg13g2_decap_4
XFILLER_24_481 VPWR VGND sg13g2_decap_8
XFILLER_25_993 VPWR VGND sg13g2_decap_8
XFILLER_8_614 VPWR VGND sg13g2_decap_8
XFILLER_11_142 VPWR VGND sg13g2_decap_8
XFILLER_12_698 VPWR VGND sg13g2_decap_8
XFILLER_40_985 VPWR VGND sg13g2_decap_8
XFILLER_7_179 VPWR VGND sg13g2_decap_8
XFILLER_7_168 VPWR VGND sg13g2_decap_8
XFILLER_22_71 VPWR VGND sg13g2_decap_8
XFILLER_22_82 VPWR VGND sg13g2_fill_1
XFILLER_4_853 VPWR VGND sg13g2_decap_8
XFILLER_3_352 VPWR VGND sg13g2_decap_8
XFILLER_39_529 VPWR VGND sg13g2_decap_8
XFILLER_47_562 VPWR VGND sg13g2_decap_8
XFILLER_35_757 VPWR VGND sg13g2_decap_8
XFILLER_16_971 VPWR VGND sg13g2_decap_8
XFILLER_23_908 VPWR VGND sg13g2_decap_8
XFILLER_34_245 VPWR VGND sg13g2_decap_8
XFILLER_22_418 VPWR VGND sg13g2_decap_8
XFILLER_30_473 VPWR VGND sg13g2_fill_1
XFILLER_31_974 VPWR VGND sg13g2_decap_8
XFILLER_8_95 VPWR VGND sg13g2_decap_8
XFILLER_38_551 VPWR VGND sg13g2_decap_8
XFILLER_14_919 VPWR VGND sg13g2_decap_8
XFILLER_26_768 VPWR VGND sg13g2_decap_8
XFILLER_41_716 VPWR VGND sg13g2_decap_8
XFILLER_22_996 VPWR VGND sg13g2_decap_8
XFILLER_5_617 VPWR VGND sg13g2_decap_8
XFILLER_49_1014 VPWR VGND sg13g2_decap_8
XFILLER_1_801 VPWR VGND sg13g2_decap_8
XFILLER_0_322 VPWR VGND sg13g2_decap_8
XFILLER_1_878 VPWR VGND sg13g2_decap_8
XFILLER_48_337 VPWR VGND sg13g2_decap_8
XFILLER_0_399 VPWR VGND sg13g2_decap_8
XFILLER_44_521 VPWR VGND sg13g2_decap_8
XFILLER_29_595 VPWR VGND sg13g2_decap_8
XFILLER_17_71 VPWR VGND sg13g2_decap_8
XFILLER_17_768 VPWR VGND sg13g2_decap_8
X_584_ net67 VGND VPWR net200 mac2.sum_lvl2_ff\[1\] clknet_5_13__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_598 VPWR VGND sg13g2_decap_8
XFILLER_31_215 VPWR VGND sg13g2_decap_8
XFILLER_9_912 VPWR VGND sg13g2_decap_8
XFILLER_13_963 VPWR VGND sg13g2_decap_8
XFILLER_25_790 VPWR VGND sg13g2_decap_8
XFILLER_31_248 VPWR VGND sg13g2_fill_2
XFILLER_8_400 VPWR VGND sg13g2_decap_8
XFILLER_12_451 VPWR VGND sg13g2_decap_8
XFILLER_40_782 VPWR VGND sg13g2_decap_8
XFILLER_8_444 VPWR VGND sg13g2_decap_8
XFILLER_9_989 VPWR VGND sg13g2_decap_8
XFILLER_4_650 VPWR VGND sg13g2_decap_8
XFILLER_39_337 VPWR VGND sg13g2_decap_8
XFILLER_39_348 VPWR VGND sg13g2_fill_1
XFILLER_23_705 VPWR VGND sg13g2_decap_8
XFILLER_35_554 VPWR VGND sg13g2_decap_8
XFILLER_22_226 VPWR VGND sg13g2_decap_8
XFILLER_13_18 VPWR VGND sg13g2_decap_8
XFILLER_31_771 VPWR VGND sg13g2_decap_8
XFILLER_1_119 VPWR VGND sg13g2_decap_8
XFILLER_26_532 VPWR VGND sg13g2_decap_8
XFILLER_38_370 VPWR VGND sg13g2_decap_8
XFILLER_39_893 VPWR VGND sg13g2_decap_8
XFILLER_26_565 VPWR VGND sg13g2_decap_8
XFILLER_13_204 VPWR VGND sg13g2_decap_4
XFILLER_14_716 VPWR VGND sg13g2_decap_8
XFILLER_41_513 VPWR VGND sg13g2_decap_8
XFILLER_16_1013 VPWR VGND sg13g2_decap_8
XFILLER_10_944 VPWR VGND sg13g2_decap_8
XFILLER_22_793 VPWR VGND sg13g2_decap_8
XFILLER_6_915 VPWR VGND sg13g2_decap_8
XFILLER_5_436 VPWR VGND sg13g2_decap_8
XFILLER_1_675 VPWR VGND sg13g2_decap_8
XFILLER_49_657 VPWR VGND sg13g2_decap_8
XFILLER_0_196 VPWR VGND sg13g2_decap_8
XFILLER_23_1006 VPWR VGND sg13g2_decap_8
XFILLER_48_145 VPWR VGND sg13g2_decap_8
XFILLER_37_819 VPWR VGND sg13g2_decap_8
XFILLER_28_81 VPWR VGND sg13g2_decap_4
XFILLER_36_329 VPWR VGND sg13g2_decap_4
XFILLER_17_543 VPWR VGND sg13g2_decap_8
XFILLER_45_885 VPWR VGND sg13g2_decap_8
X_567_ net81 VGND VPWR net118 mac2.sum_lvl1_ff\[8\] clknet_5_13__leaf_clk sg13g2_dfrbpq_1
XFILLER_13_760 VPWR VGND sg13g2_decap_8
X_498_ net64 VGND VPWR _120_ DP_3.matrix\[112\] clknet_5_3__leaf_clk sg13g2_dfrbpq_1
XFILLER_20_719 VPWR VGND sg13g2_decap_8
XFILLER_32_568 VPWR VGND sg13g2_decap_8
XFILLER_12_281 VPWR VGND sg13g2_fill_2
XFILLER_9_786 VPWR VGND sg13g2_decap_8
XFILLER_8_274 VPWR VGND sg13g2_decap_8
XFILLER_5_981 VPWR VGND sg13g2_decap_8
XFILLER_39_101 VPWR VGND sg13g2_decap_8
XFILLER_39_156 VPWR VGND sg13g2_decap_4
XFILLER_36_841 VPWR VGND sg13g2_decap_8
XFILLER_35_373 VPWR VGND sg13g2_decap_8
XFILLER_23_579 VPWR VGND sg13g2_decap_8
XFILLER_10_229 VPWR VGND sg13g2_decap_8
XFILLER_3_929 VPWR VGND sg13g2_decap_8
XFILLER_49_14 VPWR VGND sg13g2_decap_8
XFILLER_19_819 VPWR VGND sg13g2_decap_8
XFILLER_46_638 VPWR VGND sg13g2_decap_8
XFILLER_39_690 VPWR VGND sg13g2_decap_8
XFILLER_45_159 VPWR VGND sg13g2_decap_8
XFILLER_26_340 VPWR VGND sg13g2_decap_8
XFILLER_42_822 VPWR VGND sg13g2_decap_8
XFILLER_27_896 VPWR VGND sg13g2_decap_8
X_421_ net93 _115_ VPWR VGND sg13g2_buf_1
X_352_ _207_ _206_ _055_ VPWR VGND sg13g2_xor2_1
XFILLER_14_546 VPWR VGND sg13g2_decap_4
XFILLER_41_321 VPWR VGND sg13g2_decap_8
XFILLER_42_899 VPWR VGND sg13g2_decap_8
X_283_ _166_ net205 net165 VPWR VGND sg13g2_nand2_1
XFILLER_10_741 VPWR VGND sg13g2_decap_8
XFILLER_6_712 VPWR VGND sg13g2_decap_8
XFILLER_22_590 VPWR VGND sg13g2_decap_8
XFILLER_5_233 VPWR VGND sg13g2_decap_8
XFILLER_6_789 VPWR VGND sg13g2_decap_8
XFILLER_2_984 VPWR VGND sg13g2_decap_8
XFILLER_1_472 VPWR VGND sg13g2_decap_8
XFILLER_49_454 VPWR VGND sg13g2_decap_8
XFILLER_37_616 VPWR VGND sg13g2_decap_8
XFILLER_39_80 VPWR VGND sg13g2_decap_8
XFILLER_36_126 VPWR VGND sg13g2_decap_8
XFILLER_18_863 VPWR VGND sg13g2_decap_8
XFILLER_45_682 VPWR VGND sg13g2_decap_8
XFILLER_33_800 VPWR VGND sg13g2_decap_8
XFILLER_17_384 VPWR VGND sg13g2_decap_8
XFILLER_32_332 VPWR VGND sg13g2_decap_8
XFILLER_33_877 VPWR VGND sg13g2_decap_8
XFILLER_9_550 VPWR VGND sg13g2_decap_8
XFILLER_9_583 VPWR VGND sg13g2_decap_8
XFILLER_19_39 VPWR VGND sg13g2_decap_8
XFILLER_27_104 VPWR VGND sg13g2_decap_4
XFILLER_28_638 VPWR VGND sg13g2_decap_8
XFILLER_27_159 VPWR VGND sg13g2_decap_8
XFILLER_23_332 VPWR VGND sg13g2_decap_8
XFILLER_24_866 VPWR VGND sg13g2_decap_8
XFILLER_13_1005 VPWR VGND sg13g2_decap_8
XFILLER_3_726 VPWR VGND sg13g2_decap_8
XFILLER_2_203 VPWR VGND sg13g2_decap_8
XFILLER_47_947 VPWR VGND sg13g2_decap_8
XFILLER_19_616 VPWR VGND sg13g2_decap_8
XFILLER_46_435 VPWR VGND sg13g2_decap_8
XFILLER_18_148 VPWR VGND sg13g2_decap_8
XFILLER_15_811 VPWR VGND sg13g2_decap_8
XFILLER_27_693 VPWR VGND sg13g2_decap_8
XFILLER_14_343 VPWR VGND sg13g2_decap_8
XFILLER_15_888 VPWR VGND sg13g2_decap_8
XFILLER_30_814 VPWR VGND sg13g2_decap_8
X_404_ net158 _098_ VPWR VGND sg13g2_buf_1
XFILLER_41_140 VPWR VGND sg13g2_decap_8
XFILLER_42_696 VPWR VGND sg13g2_decap_8
X_335_ _196_ net143 net45 VPWR VGND sg13g2_nand2_1
X_266_ net129 mac1.sum_lvl1_ff\[8\] _008_ VPWR VGND sg13g2_xor2_1
Xclkbuf_4_6_0_clk clknet_0_clk clknet_4_6_0_clk VPWR VGND sg13g2_buf_8
XFILLER_41_195 VPWR VGND sg13g2_decap_8
XFILLER_6_531 VPWR VGND sg13g2_decap_8
XFILLER_41_70 VPWR VGND sg13g2_decap_8
XFILLER_6_586 VPWR VGND sg13g2_decap_8
XFILLER_29_1001 VPWR VGND sg13g2_decap_8
XFILLER_2_781 VPWR VGND sg13g2_decap_8
XFILLER_2_53 VPWR VGND sg13g2_decap_8
XFILLER_49_273 VPWR VGND sg13g2_decap_8
XFILLER_38_936 VPWR VGND sg13g2_decap_8
XFILLER_37_435 VPWR VGND sg13g2_decap_8
XFILLER_18_660 VPWR VGND sg13g2_decap_8
XFILLER_25_608 VPWR VGND sg13g2_decap_8
XFILLER_17_170 VPWR VGND sg13g2_decap_4
XFILLER_24_118 VPWR VGND sg13g2_fill_2
XFILLER_24_129 VPWR VGND sg13g2_decap_8
XFILLER_33_674 VPWR VGND sg13g2_decap_8
XFILLER_36_1016 VPWR VGND sg13g2_decap_8
XFILLER_36_1027 VPWR VGND sg13g2_fill_2
XFILLER_21_869 VPWR VGND sg13g2_decap_8
XFILLER_21_18 VPWR VGND sg13g2_decap_8
XFILLER_21_29 VPWR VGND sg13g2_decap_4
XFILLER_0_707 VPWR VGND sg13g2_decap_8
XFILLER_29_903 VPWR VGND sg13g2_decap_8
XFILLER_28_413 VPWR VGND sg13g2_fill_1
XFILLER_44_906 VPWR VGND sg13g2_decap_8
XFILLER_37_980 VPWR VGND sg13g2_decap_8
XFILLER_12_803 VPWR VGND sg13g2_decap_8
XFILLER_24_663 VPWR VGND sg13g2_decap_8
XFILLER_23_162 VPWR VGND sg13g2_decap_8
XFILLER_11_335 VPWR VGND sg13g2_fill_2
XFILLER_7_328 VPWR VGND sg13g2_decap_8
XFILLER_20_880 VPWR VGND sg13g2_decap_8
XFILLER_11_51 VPWR VGND sg13g2_decap_8
XFILLER_11_62 VPWR VGND sg13g2_fill_2
XFILLER_4_1014 VPWR VGND sg13g2_decap_8
XFILLER_19_413 VPWR VGND sg13g2_fill_1
XFILLER_47_744 VPWR VGND sg13g2_decap_8
XFILLER_35_939 VPWR VGND sg13g2_decap_8
XFILLER_27_490 VPWR VGND sg13g2_decap_8
XFILLER_34_449 VPWR VGND sg13g2_decap_8
XFILLER_36_70 VPWR VGND sg13g2_decap_8
XFILLER_43_994 VPWR VGND sg13g2_decap_8
XFILLER_14_151 VPWR VGND sg13g2_decap_8
XFILLER_15_685 VPWR VGND sg13g2_decap_8
XFILLER_30_611 VPWR VGND sg13g2_decap_8
XFILLER_42_493 VPWR VGND sg13g2_decap_8
XFILLER_14_195 VPWR VGND sg13g2_decap_8
X_318_ net107 mac2.sum_lvl3_ff\[0\] _032_ VPWR VGND sg13g2_xor2_1
XFILLER_30_688 VPWR VGND sg13g2_decap_8
X_249_ net3 _146_ _149_ VPWR VGND sg13g2_xnor2_1
XFILLER_7_884 VPWR VGND sg13g2_decap_8
XFILLER_6_394 VPWR VGND sg13g2_decap_8
XFILLER_6_372 VPWR VGND sg13g2_fill_2
XFILLER_38_733 VPWR VGND sg13g2_decap_8
XFILLER_16_18 VPWR VGND sg13g2_decap_8
XFILLER_19_980 VPWR VGND sg13g2_decap_8
XFILLER_25_427 VPWR VGND sg13g2_decap_8
XFILLER_21_666 VPWR VGND sg13g2_decap_8
XFILLER_0_504 VPWR VGND sg13g2_decap_8
XFILLER_29_700 VPWR VGND sg13g2_decap_8
XFILLER_44_703 VPWR VGND sg13g2_decap_8
XFILLER_29_777 VPWR VGND sg13g2_decap_8
XFILLER_43_213 VPWR VGND sg13g2_decap_8
XFILLER_43_268 VPWR VGND sg13g2_decap_8
XFILLER_19_1022 VPWR VGND sg13g2_decap_8
XFILLER_24_460 VPWR VGND sg13g2_decap_8
XFILLER_25_972 VPWR VGND sg13g2_decap_8
XFILLER_31_419 VPWR VGND sg13g2_decap_8
XFILLER_40_964 VPWR VGND sg13g2_decap_8
XFILLER_7_103 VPWR VGND sg13g2_decap_8
XFILLER_12_677 VPWR VGND sg13g2_decap_8
XFILLER_7_147 VPWR VGND sg13g2_decap_8
XFILLER_11_198 VPWR VGND sg13g2_decap_8
XFILLER_22_50 VPWR VGND sg13g2_decap_8
XFILLER_4_832 VPWR VGND sg13g2_decap_8
XFILLER_39_508 VPWR VGND sg13g2_decap_8
XFILLER_47_541 VPWR VGND sg13g2_decap_8
XFILLER_19_298 VPWR VGND sg13g2_decap_8
XFILLER_34_224 VPWR VGND sg13g2_decap_8
XFILLER_35_736 VPWR VGND sg13g2_decap_8
XFILLER_16_950 VPWR VGND sg13g2_decap_8
XFILLER_43_791 VPWR VGND sg13g2_decap_8
XFILLER_31_953 VPWR VGND sg13g2_decap_8
XFILLER_8_74 VPWR VGND sg13g2_decap_8
XFILLER_30_485 VPWR VGND sg13g2_decap_4
XFILLER_7_681 VPWR VGND sg13g2_decap_8
XFILLER_40_0 VPWR VGND sg13g2_decap_8
XFILLER_38_530 VPWR VGND sg13g2_decap_8
XFILLER_27_28 VPWR VGND sg13g2_decap_8
XFILLER_27_39 VPWR VGND sg13g2_fill_1
XFILLER_26_747 VPWR VGND sg13g2_decap_8
XFILLER_13_408 VPWR VGND sg13g2_decap_8
XFILLER_25_268 VPWR VGND sg13g2_decap_8
XFILLER_40_216 VPWR VGND sg13g2_fill_2
XFILLER_43_49 VPWR VGND sg13g2_decap_8
XFILLER_22_975 VPWR VGND sg13g2_decap_8
XFILLER_4_106 VPWR VGND sg13g2_decap_8
XFILLER_0_301 VPWR VGND sg13g2_decap_8
XFILLER_1_857 VPWR VGND sg13g2_decap_8
XFILLER_49_839 VPWR VGND sg13g2_decap_8
XFILLER_48_316 VPWR VGND sg13g2_decap_8
XFILLER_0_378 VPWR VGND sg13g2_decap_8
Xclkbuf_5_26__f_clk clknet_4_13_0_clk clknet_5_26__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_44_500 VPWR VGND sg13g2_decap_8
XFILLER_16_224 VPWR VGND sg13g2_decap_8
XFILLER_17_747 VPWR VGND sg13g2_decap_8
XFILLER_29_574 VPWR VGND sg13g2_decap_8
X_583_ net67 VGND VPWR net122 mac2.sum_lvl2_ff\[0\] clknet_5_13__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_577 VPWR VGND sg13g2_decap_8
XFILLER_12_430 VPWR VGND sg13g2_decap_8
XFILLER_13_942 VPWR VGND sg13g2_decap_8
XFILLER_33_60 VPWR VGND sg13g2_decap_8
XFILLER_40_761 VPWR VGND sg13g2_decap_8
XFILLER_8_423 VPWR VGND sg13g2_decap_8
XFILLER_9_968 VPWR VGND sg13g2_decap_8
XFILLER_3_161 VPWR VGND sg13g2_fill_2
XFILLER_3_150 VPWR VGND sg13g2_decap_8
XFILLER_3_194 VPWR VGND sg13g2_fill_1
XFILLER_12_4 VPWR VGND sg13g2_decap_8
Xhold1 mac2.sum_lvl1_ff\[33\] VPWR VGND net25 sg13g2_dlygate4sd3_1
XFILLER_35_533 VPWR VGND sg13g2_decap_8
XFILLER_22_205 VPWR VGND sg13g2_decap_8
XFILLER_31_750 VPWR VGND sg13g2_decap_8
XFILLER_38_38 VPWR VGND sg13g2_fill_2
XFILLER_39_872 VPWR VGND sg13g2_decap_8
XFILLER_26_511 VPWR VGND sg13g2_decap_8
XFILLER_26_544 VPWR VGND sg13g2_decap_8
XFILLER_22_772 VPWR VGND sg13g2_decap_8
XFILLER_41_569 VPWR VGND sg13g2_decap_8
XFILLER_10_923 VPWR VGND sg13g2_decap_8
XFILLER_21_260 VPWR VGND sg13g2_decap_4
XFILLER_21_293 VPWR VGND sg13g2_decap_8
XFILLER_1_654 VPWR VGND sg13g2_decap_8
XFILLER_49_636 VPWR VGND sg13g2_decap_8
XFILLER_48_124 VPWR VGND sg13g2_decap_8
XFILLER_0_175 VPWR VGND sg13g2_decap_8
XFILLER_36_308 VPWR VGND sg13g2_decap_8
XFILLER_17_522 VPWR VGND sg13g2_decap_8
XFILLER_28_60 VPWR VGND sg13g2_decap_8
XFILLER_45_864 VPWR VGND sg13g2_decap_8
XFILLER_17_566 VPWR VGND sg13g2_fill_1
X_566_ net79 VGND VPWR net202 mac2.sum_lvl1_ff\[1\] clknet_5_26__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_599 VPWR VGND sg13g2_decap_8
XFILLER_32_547 VPWR VGND sg13g2_decap_8
X_497_ net63 VGND VPWR _119_ DP_3.matrix\[97\] clknet_5_2__leaf_clk sg13g2_dfrbpq_1
XFILLER_12_260 VPWR VGND sg13g2_decap_8
XFILLER_9_765 VPWR VGND sg13g2_decap_8
XFILLER_5_960 VPWR VGND sg13g2_decap_8
XFILLER_4_481 VPWR VGND sg13g2_decap_8
XFILLER_36_820 VPWR VGND sg13g2_decap_8
XFILLER_35_330 VPWR VGND sg13g2_fill_2
XFILLER_36_897 VPWR VGND sg13g2_decap_8
XFILLER_24_18 VPWR VGND sg13g2_decap_4
XFILLER_23_558 VPWR VGND sg13g2_decap_8
XFILLER_10_208 VPWR VGND sg13g2_decap_8
XFILLER_40_28 VPWR VGND sg13g2_decap_4
XFILLER_3_908 VPWR VGND sg13g2_decap_8
XFILLER_46_617 VPWR VGND sg13g2_decap_8
XFILLER_18_319 VPWR VGND sg13g2_decap_8
XFILLER_45_138 VPWR VGND sg13g2_decap_8
XFILLER_42_801 VPWR VGND sg13g2_decap_8
XFILLER_27_875 VPWR VGND sg13g2_decap_8
X_420_ net141 _114_ VPWR VGND sg13g2_buf_1
X_351_ _207_ net160 net53 VPWR VGND sg13g2_nand2_1
XFILLER_14_525 VPWR VGND sg13g2_decap_8
XFILLER_26_396 VPWR VGND sg13g2_decap_8
XFILLER_41_300 VPWR VGND sg13g2_decap_8
XFILLER_42_878 VPWR VGND sg13g2_decap_8
XFILLER_10_720 VPWR VGND sg13g2_decap_8
X_282_ net147 mac2.products_ff\[16\] _017_ VPWR VGND sg13g2_xor2_1
XFILLER_14_95 VPWR VGND sg13g2_decap_8
XFILLER_10_797 VPWR VGND sg13g2_decap_8
XFILLER_5_212 VPWR VGND sg13g2_decap_8
XFILLER_6_768 VPWR VGND sg13g2_decap_8
XFILLER_2_963 VPWR VGND sg13g2_decap_8
XFILLER_1_451 VPWR VGND sg13g2_decap_8
XFILLER_49_433 VPWR VGND sg13g2_decap_8
XFILLER_36_105 VPWR VGND sg13g2_decap_8
XFILLER_18_842 VPWR VGND sg13g2_decap_8
XFILLER_45_661 VPWR VGND sg13g2_decap_8
XFILLER_17_363 VPWR VGND sg13g2_decap_8
XFILLER_32_311 VPWR VGND sg13g2_decap_8
XFILLER_33_856 VPWR VGND sg13g2_decap_8
X_549_ net61 VGND VPWR net26 mac1.sum_lvl2_ff\[9\] clknet_5_16__leaf_clk sg13g2_dfrbpq_1
XFILLER_20_539 VPWR VGND sg13g2_decap_8
XFILLER_32_388 VPWR VGND sg13g2_decap_8
XFILLER_19_18 VPWR VGND sg13g2_decap_8
XFILLER_28_617 VPWR VGND sg13g2_decap_8
XFILLER_27_138 VPWR VGND sg13g2_decap_8
XFILLER_43_609 VPWR VGND sg13g2_decap_8
XFILLER_35_28 VPWR VGND sg13g2_decap_8
XFILLER_42_119 VPWR VGND sg13g2_decap_8
XFILLER_23_311 VPWR VGND sg13g2_decap_8
XFILLER_24_845 VPWR VGND sg13g2_decap_8
XFILLER_36_694 VPWR VGND sg13g2_decap_8
XFILLER_35_193 VPWR VGND sg13g2_decap_8
XFILLER_11_528 VPWR VGND sg13g2_decap_8
XFILLER_11_539 VPWR VGND sg13g2_fill_2
XFILLER_13_1028 VPWR VGND sg13g2_fill_1
XFILLER_3_705 VPWR VGND sg13g2_decap_8
XFILLER_47_926 VPWR VGND sg13g2_decap_8
XFILLER_46_414 VPWR VGND sg13g2_decap_8
XFILLER_18_127 VPWR VGND sg13g2_decap_8
XFILLER_27_672 VPWR VGND sg13g2_decap_8
X_403_ net91 _097_ VPWR VGND sg13g2_buf_1
XFILLER_15_867 VPWR VGND sg13g2_decap_8
XFILLER_42_675 VPWR VGND sg13g2_decap_8
X_334_ _195_ _194_ _043_ VPWR VGND sg13g2_xor2_1
XFILLER_14_399 VPWR VGND sg13g2_decap_8
XFILLER_25_94 VPWR VGND sg13g2_decap_8
XFILLER_41_174 VPWR VGND sg13g2_decap_8
X_265_ _009_ _156_ _157_ VPWR VGND sg13g2_xnor2_1
XFILLER_6_510 VPWR VGND sg13g2_decap_8
XFILLER_10_594 VPWR VGND sg13g2_decap_8
XFILLER_6_565 VPWR VGND sg13g2_decap_8
XFILLER_44_7 VPWR VGND sg13g2_decap_8
XFILLER_2_760 VPWR VGND sg13g2_decap_8
XFILLER_2_32 VPWR VGND sg13g2_decap_8
XFILLER_38_915 VPWR VGND sg13g2_decap_8
XFILLER_49_252 VPWR VGND sg13g2_decap_8
XFILLER_46_981 VPWR VGND sg13g2_decap_8
XFILLER_37_469 VPWR VGND sg13g2_decap_8
XFILLER_33_653 VPWR VGND sg13g2_decap_8
XFILLER_21_848 VPWR VGND sg13g2_decap_8
Xclkbuf_5_7__f_clk clknet_4_3_0_clk clknet_5_7__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_28_458 VPWR VGND sg13g2_fill_2
XFILLER_29_959 VPWR VGND sg13g2_decap_8
XFILLER_24_642 VPWR VGND sg13g2_decap_8
XFILLER_36_491 VPWR VGND sg13g2_decap_8
XFILLER_11_314 VPWR VGND sg13g2_decap_8
XFILLER_23_141 VPWR VGND sg13g2_decap_8
XFILLER_12_859 VPWR VGND sg13g2_decap_8
XFILLER_7_307 VPWR VGND sg13g2_decap_8
XFILLER_11_358 VPWR VGND sg13g2_decap_8
XFILLER_3_579 VPWR VGND sg13g2_decap_8
XFILLER_47_723 VPWR VGND sg13g2_decap_8
XFILLER_46_222 VPWR VGND sg13g2_fill_2
XFILLER_46_211 VPWR VGND sg13g2_decap_8
XFILLER_19_469 VPWR VGND sg13g2_decap_8
XFILLER_35_918 VPWR VGND sg13g2_decap_8
XFILLER_28_981 VPWR VGND sg13g2_decap_8
XFILLER_43_973 VPWR VGND sg13g2_decap_8
XFILLER_14_130 VPWR VGND sg13g2_decap_8
XFILLER_15_664 VPWR VGND sg13g2_decap_8
X_317_ _033_ _182_ _185_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_667 VPWR VGND sg13g2_decap_8
X_248_ _149_ _148_ _147_ VPWR VGND sg13g2_nand2b_1
XFILLER_7_863 VPWR VGND sg13g2_decap_8
XFILLER_6_351 VPWR VGND sg13g2_decap_8
XFILLER_38_712 VPWR VGND sg13g2_decap_8
XFILLER_26_929 VPWR VGND sg13g2_decap_8
XFILLER_37_244 VPWR VGND sg13g2_decap_8
XFILLER_38_789 VPWR VGND sg13g2_decap_8
XFILLER_25_417 VPWR VGND sg13g2_fill_1
XFILLER_37_288 VPWR VGND sg13g2_decap_8
XFILLER_18_491 VPWR VGND sg13g2_decap_8
XFILLER_40_409 VPWR VGND sg13g2_decap_8
XFILLER_34_995 VPWR VGND sg13g2_decap_8
XFILLER_21_645 VPWR VGND sg13g2_decap_8
XFILLER_20_133 VPWR VGND sg13g2_decap_8
XFILLER_20_144 VPWR VGND sg13g2_fill_1
Xclkbuf_4_5_0_clk clknet_0_clk clknet_4_5_0_clk VPWR VGND sg13g2_buf_8
XFILLER_28_211 VPWR VGND sg13g2_decap_4
XFILLER_29_756 VPWR VGND sg13g2_decap_8
XFILLER_17_929 VPWR VGND sg13g2_decap_8
XFILLER_28_288 VPWR VGND sg13g2_decap_8
XFILLER_44_759 VPWR VGND sg13g2_decap_8
XFILLER_19_1001 VPWR VGND sg13g2_decap_8
XFILLER_25_951 VPWR VGND sg13g2_decap_8
XFILLER_11_100 VPWR VGND sg13g2_fill_1
XFILLER_40_943 VPWR VGND sg13g2_decap_8
XFILLER_12_656 VPWR VGND sg13g2_decap_8
XFILLER_8_649 VPWR VGND sg13g2_decap_8
XFILLER_11_177 VPWR VGND sg13g2_decap_8
XFILLER_4_811 VPWR VGND sg13g2_decap_8
XFILLER_4_888 VPWR VGND sg13g2_decap_8
XFILLER_3_387 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_26_1027 VPWR VGND sg13g2_fill_2
XFILLER_47_520 VPWR VGND sg13g2_decap_8
XFILLER_19_200 VPWR VGND sg13g2_fill_1
XFILLER_19_255 VPWR VGND sg13g2_fill_2
XFILLER_35_715 VPWR VGND sg13g2_decap_8
XFILLER_47_597 VPWR VGND sg13g2_decap_8
XFILLER_34_203 VPWR VGND sg13g2_decap_8
XFILLER_43_770 VPWR VGND sg13g2_decap_8
XFILLER_15_483 VPWR VGND sg13g2_decap_8
XFILLER_31_932 VPWR VGND sg13g2_decap_8
XFILLER_8_53 VPWR VGND sg13g2_decap_8
XFILLER_7_660 VPWR VGND sg13g2_decap_8
XFILLER_33_0 VPWR VGND sg13g2_decap_8
XFILLER_26_726 VPWR VGND sg13g2_decap_8
XFILLER_38_586 VPWR VGND sg13g2_decap_8
XFILLER_25_247 VPWR VGND sg13g2_decap_8
XFILLER_43_28 VPWR VGND sg13g2_decap_8
XFILLER_22_954 VPWR VGND sg13g2_decap_8
XFILLER_33_280 VPWR VGND sg13g2_fill_2
XFILLER_34_792 VPWR VGND sg13g2_decap_8
XFILLER_40_239 VPWR VGND sg13g2_fill_2
XFILLER_21_475 VPWR VGND sg13g2_decap_8
XFILLER_1_836 VPWR VGND sg13g2_decap_8
XFILLER_49_818 VPWR VGND sg13g2_decap_8
XFILLER_0_357 VPWR VGND sg13g2_decap_8
XFILLER_29_553 VPWR VGND sg13g2_decap_8
X_582_ net76 VGND VPWR _067_ mac2.products_ff\[33\] clknet_5_14__leaf_clk sg13g2_dfrbpq_1
XFILLER_1_1018 VPWR VGND sg13g2_decap_8
XFILLER_16_203 VPWR VGND sg13g2_decap_8
XFILLER_17_726 VPWR VGND sg13g2_decap_8
XFILLER_44_556 VPWR VGND sg13g2_decap_8
XFILLER_16_247 VPWR VGND sg13g2_decap_8
XFILLER_32_729 VPWR VGND sg13g2_decap_8
XFILLER_13_921 VPWR VGND sg13g2_decap_8
XFILLER_40_740 VPWR VGND sg13g2_decap_8
XFILLER_9_947 VPWR VGND sg13g2_decap_8
XFILLER_13_998 VPWR VGND sg13g2_decap_8
XFILLER_33_94 VPWR VGND sg13g2_decap_4
XFILLER_8_479 VPWR VGND sg13g2_decap_8
XFILLER_4_685 VPWR VGND sg13g2_decap_8
Xhold2 mac1.sum_lvl1_ff\[33\] VPWR VGND net26 sg13g2_dlygate4sd3_1
XFILLER_48_884 VPWR VGND sg13g2_decap_8
XFILLER_47_372 VPWR VGND sg13g2_fill_2
XFILLER_35_512 VPWR VGND sg13g2_decap_8
XFILLER_35_589 VPWR VGND sg13g2_decap_8
XFILLER_30_283 VPWR VGND sg13g2_decap_8
XFILLER_38_28 VPWR VGND sg13g2_fill_2
XFILLER_39_851 VPWR VGND sg13g2_decap_8
XFILLER_41_548 VPWR VGND sg13g2_decap_8
XFILLER_10_902 VPWR VGND sg13g2_decap_8
XFILLER_22_751 VPWR VGND sg13g2_decap_8
XFILLER_10_979 VPWR VGND sg13g2_decap_8
XFILLER_1_633 VPWR VGND sg13g2_decap_8
XFILLER_49_615 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_48_103 VPWR VGND sg13g2_decap_8
XFILLER_29_361 VPWR VGND sg13g2_decap_8
XFILLER_45_843 VPWR VGND sg13g2_decap_8
XFILLER_44_364 VPWR VGND sg13g2_decap_8
X_565_ net78 VGND VPWR net148 mac2.sum_lvl1_ff\[0\] clknet_5_30__leaf_clk sg13g2_dfrbpq_2
X_496_ net63 VGND VPWR _118_ DP_3.matrix\[96\] clknet_5_8__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_526 VPWR VGND sg13g2_decap_8
XFILLER_9_744 VPWR VGND sg13g2_decap_8
XFILLER_13_795 VPWR VGND sg13g2_decap_8
XFILLER_4_460 VPWR VGND sg13g2_decap_8
XFILLER_5_65 VPWR VGND sg13g2_fill_1
XFILLER_39_136 VPWR VGND sg13g2_decap_8
XFILLER_48_681 VPWR VGND sg13g2_decap_8
XFILLER_36_876 VPWR VGND sg13g2_decap_8
XFILLER_39_1026 VPWR VGND sg13g2_fill_2
XFILLER_23_537 VPWR VGND sg13g2_decap_8
XFILLER_49_49 VPWR VGND sg13g2_decap_8
XFILLER_45_117 VPWR VGND sg13g2_decap_8
XFILLER_27_854 VPWR VGND sg13g2_decap_8
XFILLER_42_857 VPWR VGND sg13g2_decap_8
X_350_ _206_ net92 net123 VPWR VGND sg13g2_nand2_1
XFILLER_26_375 VPWR VGND sg13g2_decap_8
X_281_ _018_ _164_ _165_ VPWR VGND sg13g2_xnor2_1
XFILLER_14_74 VPWR VGND sg13g2_decap_8
XFILLER_10_776 VPWR VGND sg13g2_decap_8
XFILLER_6_747 VPWR VGND sg13g2_decap_8
XFILLER_5_268 VPWR VGND sg13g2_decap_4
XFILLER_2_942 VPWR VGND sg13g2_decap_8
XFILLER_30_84 VPWR VGND sg13g2_decap_8
XFILLER_1_430 VPWR VGND sg13g2_decap_8
XFILLER_49_412 VPWR VGND sg13g2_decap_8
XFILLER_7_1024 VPWR VGND sg13g2_decap_4
XFILLER_49_489 VPWR VGND sg13g2_decap_8
XFILLER_18_821 VPWR VGND sg13g2_decap_8
XFILLER_45_640 VPWR VGND sg13g2_decap_8
XFILLER_17_342 VPWR VGND sg13g2_decap_8
X_548_ net61 VGND VPWR net34 mac1.sum_lvl2_ff\[8\] clknet_5_16__leaf_clk sg13g2_dfrbpq_1
XFILLER_18_898 VPWR VGND sg13g2_decap_8
XFILLER_33_835 VPWR VGND sg13g2_decap_8
XFILLER_44_194 VPWR VGND sg13g2_decap_4
XFILLER_20_518 VPWR VGND sg13g2_decap_8
X_479_ net67 VGND VPWR _101_ DP_2.matrix\[97\] clknet_5_13__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_367 VPWR VGND sg13g2_decap_8
XFILLER_27_117 VPWR VGND sg13g2_decap_8
XFILLER_27_128 VPWR VGND sg13g2_fill_1
XFILLER_36_673 VPWR VGND sg13g2_decap_8
XFILLER_24_824 VPWR VGND sg13g2_decap_8
XFILLER_35_172 VPWR VGND sg13g2_decap_8
XFILLER_23_378 VPWR VGND sg13g2_fill_1
XFILLER_32_890 VPWR VGND sg13g2_decap_8
XFILLER_2_238 VPWR VGND sg13g2_fill_2
XFILLER_47_905 VPWR VGND sg13g2_decap_8
XFILLER_27_651 VPWR VGND sg13g2_decap_8
XFILLER_15_846 VPWR VGND sg13g2_decap_8
X_402_ net157 _096_ VPWR VGND sg13g2_buf_1
XFILLER_42_654 VPWR VGND sg13g2_decap_8
XFILLER_26_183 VPWR VGND sg13g2_decap_8
X_333_ _195_ net154 net55 VPWR VGND sg13g2_nand2_1
XFILLER_14_378 VPWR VGND sg13g2_decap_8
XFILLER_25_73 VPWR VGND sg13g2_decap_8
X_264_ mac1.sum_lvl1_ff\[1\] mac1.sum_lvl1_ff\[9\] _157_ VPWR VGND sg13g2_xor2_1
XFILLER_30_849 VPWR VGND sg13g2_decap_8
XFILLER_10_584 VPWR VGND sg13g2_fill_1
XFILLER_37_7 VPWR VGND sg13g2_decap_8
XFILLER_49_231 VPWR VGND sg13g2_decap_8
XFILLER_2_11 VPWR VGND sg13g2_decap_8
XFILLER_2_88 VPWR VGND sg13g2_decap_8
XFILLER_46_960 VPWR VGND sg13g2_decap_8
XFILLER_18_695 VPWR VGND sg13g2_decap_8
XFILLER_33_632 VPWR VGND sg13g2_decap_8
XFILLER_20_315 VPWR VGND sg13g2_fill_2
XFILLER_21_827 VPWR VGND sg13g2_decap_8
XFILLER_32_153 VPWR VGND sg13g2_decap_8
XFILLER_32_186 VPWR VGND sg13g2_decap_8
XFILLER_9_382 VPWR VGND sg13g2_decap_8
XFILLER_29_938 VPWR VGND sg13g2_decap_8
XFILLER_46_28 VPWR VGND sg13g2_decap_8
XFILLER_28_437 VPWR VGND sg13g2_decap_8
XFILLER_43_429 VPWR VGND sg13g2_decap_8
XFILLER_15_109 VPWR VGND sg13g2_decap_8
XFILLER_24_621 VPWR VGND sg13g2_decap_8
XFILLER_23_120 VPWR VGND sg13g2_decap_8
XFILLER_12_838 VPWR VGND sg13g2_decap_8
XFILLER_24_698 VPWR VGND sg13g2_decap_8
XFILLER_23_197 VPWR VGND sg13g2_decap_8
XFILLER_3_503 VPWR VGND sg13g2_fill_2
XFILLER_3_536 VPWR VGND sg13g2_decap_8
XFILLER_3_558 VPWR VGND sg13g2_decap_8
XFILLER_3_547 VPWR VGND sg13g2_fill_2
XFILLER_2_4 VPWR VGND sg13g2_decap_8
XFILLER_47_702 VPWR VGND sg13g2_decap_8
XFILLER_19_426 VPWR VGND sg13g2_fill_2
XFILLER_47_779 VPWR VGND sg13g2_decap_8
XFILLER_28_960 VPWR VGND sg13g2_decap_8
XFILLER_46_289 VPWR VGND sg13g2_decap_8
XFILLER_43_952 VPWR VGND sg13g2_decap_8
XFILLER_15_643 VPWR VGND sg13g2_decap_8
X_316_ mac2.sum_lvl3_ff\[3\] net170 _185_ VPWR VGND sg13g2_xor2_1
XFILLER_30_646 VPWR VGND sg13g2_decap_8
XFILLER_7_842 VPWR VGND sg13g2_decap_8
XFILLER_11_893 VPWR VGND sg13g2_decap_8
X_247_ VGND VPWR _148_ mac2.total_sum\[2\] mac1.total_sum\[2\] sg13g2_or2_1
XFILLER_42_1011 VPWR VGND sg13g2_decap_8
XFILLER_37_223 VPWR VGND sg13g2_fill_1
XFILLER_26_908 VPWR VGND sg13g2_decap_8
XFILLER_38_768 VPWR VGND sg13g2_decap_8
XFILLER_18_470 VPWR VGND sg13g2_decap_8
XFILLER_33_473 VPWR VGND sg13g2_fill_2
XFILLER_34_974 VPWR VGND sg13g2_decap_8
XFILLER_20_112 VPWR VGND sg13g2_decap_8
XFILLER_21_624 VPWR VGND sg13g2_decap_8
XFILLER_0_539 VPWR VGND sg13g2_decap_8
XFILLER_29_735 VPWR VGND sg13g2_decap_8
XFILLER_17_908 VPWR VGND sg13g2_decap_8
XFILLER_28_245 VPWR VGND sg13g2_decap_8
XFILLER_44_738 VPWR VGND sg13g2_decap_8
XFILLER_25_930 VPWR VGND sg13g2_decap_8
XFILLER_40_922 VPWR VGND sg13g2_decap_8
XFILLER_12_624 VPWR VGND sg13g2_fill_2
XFILLER_12_635 VPWR VGND sg13g2_decap_8
XFILLER_24_495 VPWR VGND sg13g2_decap_8
XFILLER_8_628 VPWR VGND sg13g2_decap_8
XFILLER_11_156 VPWR VGND sg13g2_decap_8
XFILLER_40_999 VPWR VGND sg13g2_decap_8
XFILLER_4_867 VPWR VGND sg13g2_decap_8
XFILLER_3_366 VPWR VGND sg13g2_decap_8
XFILLER_26_1006 VPWR VGND sg13g2_decap_8
XFILLER_19_223 VPWR VGND sg13g2_fill_2
XFILLER_47_71 VPWR VGND sg13g2_decap_8
XFILLER_47_60 VPWR VGND sg13g2_fill_2
XFILLER_19_234 VPWR VGND sg13g2_decap_8
XFILLER_47_576 VPWR VGND sg13g2_decap_8
XFILLER_15_462 VPWR VGND sg13g2_decap_8
XFILLER_16_985 VPWR VGND sg13g2_decap_8
XFILLER_31_911 VPWR VGND sg13g2_decap_8
XFILLER_34_259 VPWR VGND sg13g2_decap_8
XFILLER_8_32 VPWR VGND sg13g2_decap_8
XFILLER_30_454 VPWR VGND sg13g2_decap_8
XFILLER_30_465 VPWR VGND sg13g2_fill_2
XFILLER_31_988 VPWR VGND sg13g2_decap_8
XFILLER_11_690 VPWR VGND sg13g2_decap_8
XFILLER_26_705 VPWR VGND sg13g2_decap_8
XFILLER_38_565 VPWR VGND sg13g2_decap_8
XFILLER_34_771 VPWR VGND sg13g2_decap_8
XFILLER_22_933 VPWR VGND sg13g2_decap_8
XFILLER_40_218 VPWR VGND sg13g2_fill_1
XFILLER_21_443 VPWR VGND sg13g2_decap_8
XFILLER_49_1028 VPWR VGND sg13g2_fill_1
XFILLER_1_815 VPWR VGND sg13g2_decap_8
XFILLER_0_336 VPWR VGND sg13g2_decap_8
XFILLER_17_705 VPWR VGND sg13g2_decap_8
XFILLER_29_532 VPWR VGND sg13g2_decap_8
X_581_ net76 VGND VPWR _066_ mac2.products_ff\[32\] clknet_5_15__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_535 VPWR VGND sg13g2_decap_8
XFILLER_16_237 VPWR VGND sg13g2_fill_1
XFILLER_13_900 VPWR VGND sg13g2_decap_8
XFILLER_17_85 VPWR VGND sg13g2_fill_2
XFILLER_32_708 VPWR VGND sg13g2_decap_8
XFILLER_31_229 VPWR VGND sg13g2_fill_2
XFILLER_9_926 VPWR VGND sg13g2_decap_8
XFILLER_13_977 VPWR VGND sg13g2_decap_8
XFILLER_24_292 VPWR VGND sg13g2_fill_2
XFILLER_12_465 VPWR VGND sg13g2_decap_8
XFILLER_40_796 VPWR VGND sg13g2_decap_8
XFILLER_8_458 VPWR VGND sg13g2_decap_8
XFILLER_4_664 VPWR VGND sg13g2_decap_8
Xhold3 mac1.products_ff\[129\] VPWR VGND net27 sg13g2_dlygate4sd3_1
XFILLER_48_863 VPWR VGND sg13g2_decap_8
XFILLER_47_351 VPWR VGND sg13g2_decap_8
XFILLER_23_719 VPWR VGND sg13g2_decap_8
XFILLER_35_568 VPWR VGND sg13g2_decap_8
XFILLER_16_782 VPWR VGND sg13g2_decap_8
XFILLER_30_262 VPWR VGND sg13g2_decap_8
XFILLER_31_785 VPWR VGND sg13g2_decap_8
Xclkbuf_4_4_0_clk clknet_0_clk clknet_4_4_0_clk VPWR VGND sg13g2_buf_8
XFILLER_8_992 VPWR VGND sg13g2_decap_8
XFILLER_39_830 VPWR VGND sg13g2_decap_8
XFILLER_38_384 VPWR VGND sg13g2_decap_8
XFILLER_26_579 VPWR VGND sg13g2_decap_8
XFILLER_13_229 VPWR VGND sg13g2_decap_8
XFILLER_41_527 VPWR VGND sg13g2_decap_8
XFILLER_22_730 VPWR VGND sg13g2_decap_8
XFILLER_16_1027 VPWR VGND sg13g2_fill_2
XFILLER_10_958 VPWR VGND sg13g2_decap_8
XFILLER_6_929 VPWR VGND sg13g2_decap_8
XFILLER_1_612 VPWR VGND sg13g2_decap_8
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_1_689 VPWR VGND sg13g2_decap_8
XFILLER_48_159 VPWR VGND sg13g2_decap_8
XFILLER_45_822 VPWR VGND sg13g2_decap_8
XFILLER_44_343 VPWR VGND sg13g2_fill_2
XFILLER_17_557 VPWR VGND sg13g2_decap_8
XFILLER_32_505 VPWR VGND sg13g2_decap_8
X_564_ net68 VGND VPWR _061_ mac2.products_ff\[65\] clknet_5_9__leaf_clk sg13g2_dfrbpq_1
X_495_ net65 VGND VPWR _117_ DP_3.matrix\[81\] clknet_5_10__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_899 VPWR VGND sg13g2_decap_8
XFILLER_44_61 VPWR VGND sg13g2_decap_8
XFILLER_9_723 VPWR VGND sg13g2_decap_8
XFILLER_13_774 VPWR VGND sg13g2_decap_8
XFILLER_40_593 VPWR VGND sg13g2_decap_8
XFILLER_8_288 VPWR VGND sg13g2_decap_8
XFILLER_5_995 VPWR VGND sg13g2_decap_8
XFILLER_39_115 VPWR VGND sg13g2_decap_8
XFILLER_48_660 VPWR VGND sg13g2_decap_8
XFILLER_47_181 VPWR VGND sg13g2_decap_8
XFILLER_36_855 VPWR VGND sg13g2_decap_8
XFILLER_39_1005 VPWR VGND sg13g2_decap_8
XFILLER_35_387 VPWR VGND sg13g2_decap_4
XFILLER_31_582 VPWR VGND sg13g2_decap_8
XFILLER_49_28 VPWR VGND sg13g2_decap_8
XFILLER_46_1009 VPWR VGND sg13g2_decap_8
XFILLER_27_833 VPWR VGND sg13g2_decap_8
XFILLER_38_170 VPWR VGND sg13g2_fill_2
XFILLER_26_354 VPWR VGND sg13g2_decap_8
XFILLER_42_836 VPWR VGND sg13g2_decap_8
XFILLER_41_335 VPWR VGND sg13g2_decap_8
X_280_ mac2.products_ff\[1\] mac2.products_ff\[17\] _165_ VPWR VGND sg13g2_xor2_1
XFILLER_14_53 VPWR VGND sg13g2_decap_8
XFILLER_10_755 VPWR VGND sg13g2_decap_8
XFILLER_6_726 VPWR VGND sg13g2_decap_8
XFILLER_5_247 VPWR VGND sg13g2_decap_8
XFILLER_30_63 VPWR VGND sg13g2_decap_8
XFILLER_2_921 VPWR VGND sg13g2_decap_8
XFILLER_7_1003 VPWR VGND sg13g2_decap_8
XFILLER_2_998 VPWR VGND sg13g2_decap_8
XFILLER_1_486 VPWR VGND sg13g2_decap_8
XFILLER_49_468 VPWR VGND sg13g2_decap_8
XFILLER_18_800 VPWR VGND sg13g2_decap_8
XFILLER_39_94 VPWR VGND sg13g2_decap_8
XFILLER_17_321 VPWR VGND sg13g2_decap_8
XFILLER_18_877 VPWR VGND sg13g2_decap_8
XFILLER_29_192 VPWR VGND sg13g2_decap_8
XFILLER_33_814 VPWR VGND sg13g2_decap_8
XFILLER_45_696 VPWR VGND sg13g2_decap_8
X_547_ net70 VGND VPWR net174 mac1.sum_lvl2_ff\[5\] clknet_5_19__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_346 VPWR VGND sg13g2_decap_8
X_478_ net60 VGND VPWR _100_ DP_2.matrix\[96\] clknet_5_24__leaf_clk sg13g2_dfrbpq_1
XFILLER_13_593 VPWR VGND sg13g2_decap_8
XFILLER_41_891 VPWR VGND sg13g2_decap_8
XFILLER_9_564 VPWR VGND sg13g2_decap_8
XFILLER_9_597 VPWR VGND sg13g2_decap_8
XFILLER_5_792 VPWR VGND sg13g2_decap_8
XFILLER_24_803 VPWR VGND sg13g2_decap_8
XFILLER_36_652 VPWR VGND sg13g2_decap_8
XFILLER_35_151 VPWR VGND sg13g2_decap_8
XFILLER_23_357 VPWR VGND sg13g2_decap_8
XFILLER_13_1019 VPWR VGND sg13g2_decap_8
XFILLER_46_449 VPWR VGND sg13g2_decap_8
XFILLER_27_630 VPWR VGND sg13g2_decap_8
XFILLER_39_490 VPWR VGND sg13g2_decap_8
X_401_ net100 _095_ VPWR VGND sg13g2_buf_1
XFILLER_15_825 VPWR VGND sg13g2_decap_8
XFILLER_26_162 VPWR VGND sg13g2_decap_8
XFILLER_42_633 VPWR VGND sg13g2_decap_8
XFILLER_25_52 VPWR VGND sg13g2_decap_8
X_332_ _194_ net46 net156 VPWR VGND sg13g2_nand2_1
XFILLER_14_357 VPWR VGND sg13g2_decap_8
XFILLER_30_828 VPWR VGND sg13g2_decap_8
XFILLER_41_154 VPWR VGND sg13g2_decap_8
X_263_ _156_ net191 net129 VPWR VGND sg13g2_nand2_1
XFILLER_23_880 VPWR VGND sg13g2_decap_8
XFILLER_6_545 VPWR VGND sg13g2_decap_4
XFILLER_41_84 VPWR VGND sg13g2_fill_1
XFILLER_29_1015 VPWR VGND sg13g2_decap_8
XFILLER_49_210 VPWR VGND sg13g2_decap_8
XFILLER_2_795 VPWR VGND sg13g2_decap_8
XFILLER_1_283 VPWR VGND sg13g2_decap_8
XFILLER_2_67 VPWR VGND sg13g2_decap_8
XFILLER_37_405 VPWR VGND sg13g2_fill_2
XFILLER_49_287 VPWR VGND sg13g2_decap_8
XFILLER_37_449 VPWR VGND sg13g2_decap_8
XFILLER_18_674 VPWR VGND sg13g2_decap_8
XFILLER_33_611 VPWR VGND sg13g2_decap_8
XFILLER_45_493 VPWR VGND sg13g2_decap_8
XFILLER_17_195 VPWR VGND sg13g2_decap_8
XFILLER_21_806 VPWR VGND sg13g2_decap_8
XFILLER_33_688 VPWR VGND sg13g2_decap_8
XFILLER_14_891 VPWR VGND sg13g2_decap_8
XFILLER_9_361 VPWR VGND sg13g2_decap_8
XFILLER_29_917 VPWR VGND sg13g2_decap_8
XFILLER_43_408 VPWR VGND sg13g2_decap_8
XFILLER_24_600 VPWR VGND sg13g2_decap_8
XFILLER_37_994 VPWR VGND sg13g2_decap_8
XFILLER_12_817 VPWR VGND sg13g2_decap_8
XFILLER_24_677 VPWR VGND sg13g2_decap_8
XFILLER_23_176 VPWR VGND sg13g2_decap_8
XFILLER_20_894 VPWR VGND sg13g2_decap_8
XFILLER_11_98 VPWR VGND sg13g2_fill_2
XFILLER_4_1028 VPWR VGND sg13g2_fill_1
XFILLER_47_758 VPWR VGND sg13g2_decap_8
XFILLER_43_931 VPWR VGND sg13g2_decap_8
XFILLER_15_622 VPWR VGND sg13g2_decap_8
XFILLER_36_84 VPWR VGND sg13g2_decap_8
XFILLER_14_165 VPWR VGND sg13g2_decap_8
X_315_ net170 mac2.sum_lvl3_ff\[3\] _184_ VPWR VGND sg13g2_nor2_1
XFILLER_15_699 VPWR VGND sg13g2_decap_8
XFILLER_30_625 VPWR VGND sg13g2_decap_8
XFILLER_7_821 VPWR VGND sg13g2_decap_8
XFILLER_11_872 VPWR VGND sg13g2_decap_8
X_246_ mac1.total_sum\[2\] mac2.total_sum\[2\] _147_ VPWR VGND sg13g2_and2_1
XFILLER_7_898 VPWR VGND sg13g2_decap_8
XFILLER_2_592 VPWR VGND sg13g2_decap_8
XFILLER_28_4 VPWR VGND sg13g2_fill_2
XFILLER_37_202 VPWR VGND sg13g2_decap_8
XFILLER_38_747 VPWR VGND sg13g2_decap_8
XFILLER_19_994 VPWR VGND sg13g2_decap_8
XFILLER_34_953 VPWR VGND sg13g2_decap_8
XFILLER_33_485 VPWR VGND sg13g2_decap_8
Xclkbuf_5_15__f_clk clknet_4_7_0_clk clknet_5_15__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_0_518 VPWR VGND sg13g2_decap_8
XFILLER_29_714 VPWR VGND sg13g2_decap_8
XFILLER_28_224 VPWR VGND sg13g2_decap_8
XFILLER_44_717 VPWR VGND sg13g2_decap_8
XFILLER_43_227 VPWR VGND sg13g2_decap_8
XFILLER_37_791 VPWR VGND sg13g2_decap_8
XFILLER_25_986 VPWR VGND sg13g2_decap_8
XFILLER_40_901 VPWR VGND sg13g2_decap_8
XFILLER_12_614 VPWR VGND sg13g2_fill_2
XFILLER_24_474 VPWR VGND sg13g2_decap_8
XFILLER_8_607 VPWR VGND sg13g2_decap_8
XFILLER_11_135 VPWR VGND sg13g2_decap_8
XFILLER_40_978 VPWR VGND sg13g2_decap_8
XFILLER_7_117 VPWR VGND sg13g2_fill_2
XFILLER_20_691 VPWR VGND sg13g2_decap_8
XFILLER_22_64 VPWR VGND sg13g2_decap_8
XFILLER_4_846 VPWR VGND sg13g2_decap_8
XFILLER_3_345 VPWR VGND sg13g2_decap_8
XFILLER_47_555 VPWR VGND sg13g2_decap_8
XFILLER_34_238 VPWR VGND sg13g2_decap_8
XFILLER_15_441 VPWR VGND sg13g2_decap_8
XFILLER_16_964 VPWR VGND sg13g2_decap_8
XFILLER_8_11 VPWR VGND sg13g2_decap_8
XFILLER_31_967 VPWR VGND sg13g2_decap_8
XFILLER_8_88 VPWR VGND sg13g2_decap_8
X_229_ net162 net158 _048_ VPWR VGND sg13g2_and2_1
XFILLER_30_499 VPWR VGND sg13g2_decap_8
XFILLER_7_695 VPWR VGND sg13g2_decap_8
XFILLER_6_194 VPWR VGND sg13g2_decap_4
XFILLER_38_544 VPWR VGND sg13g2_decap_8
XFILLER_19_791 VPWR VGND sg13g2_decap_8
XFILLER_22_912 VPWR VGND sg13g2_decap_8
XFILLER_34_750 VPWR VGND sg13g2_decap_8
XFILLER_41_709 VPWR VGND sg13g2_decap_8
XFILLER_21_422 VPWR VGND sg13g2_decap_8
XFILLER_22_989 VPWR VGND sg13g2_decap_8
XFILLER_49_1007 VPWR VGND sg13g2_decap_8
XFILLER_0_315 VPWR VGND sg13g2_decap_8
XFILLER_29_511 VPWR VGND sg13g2_decap_8
XFILLER_44_514 VPWR VGND sg13g2_decap_8
X_580_ net64 VGND VPWR _035_ mac2.products_ff\[113\] clknet_5_3__leaf_clk sg13g2_dfrbpq_1
XFILLER_29_588 VPWR VGND sg13g2_decap_8
XFILLER_31_208 VPWR VGND sg13g2_fill_2
XFILLER_12_411 VPWR VGND sg13g2_decap_8
XFILLER_24_271 VPWR VGND sg13g2_decap_8
XFILLER_25_783 VPWR VGND sg13g2_decap_8
XFILLER_9_905 VPWR VGND sg13g2_decap_8
XFILLER_12_444 VPWR VGND sg13g2_decap_8
XFILLER_13_956 VPWR VGND sg13g2_decap_8
XFILLER_8_437 VPWR VGND sg13g2_decap_8
XFILLER_40_775 VPWR VGND sg13g2_decap_8
XFILLER_4_643 VPWR VGND sg13g2_decap_8
Xhold4 mac2.products_ff\[128\] VPWR VGND net28 sg13g2_dlygate4sd3_1
XFILLER_0_882 VPWR VGND sg13g2_decap_8
XFILLER_48_842 VPWR VGND sg13g2_decap_8
XFILLER_35_547 VPWR VGND sg13g2_decap_8
XFILLER_16_761 VPWR VGND sg13g2_decap_8
XFILLER_22_219 VPWR VGND sg13g2_decap_8
XFILLER_15_282 VPWR VGND sg13g2_decap_4
XFILLER_30_241 VPWR VGND sg13g2_decap_8
XFILLER_31_764 VPWR VGND sg13g2_decap_8
XFILLER_8_971 VPWR VGND sg13g2_decap_8
XFILLER_7_492 VPWR VGND sg13g2_decap_8
XFILLER_38_363 VPWR VGND sg13g2_decap_8
XFILLER_39_886 VPWR VGND sg13g2_decap_8
XFILLER_26_525 VPWR VGND sg13g2_decap_8
XFILLER_14_709 VPWR VGND sg13g2_decap_8
XFILLER_26_558 VPWR VGND sg13g2_decap_8
XFILLER_41_506 VPWR VGND sg13g2_decap_8
XFILLER_13_208 VPWR VGND sg13g2_fill_1
XFILLER_16_1006 VPWR VGND sg13g2_decap_8
XFILLER_10_937 VPWR VGND sg13g2_decap_8
XFILLER_22_786 VPWR VGND sg13g2_decap_8
XFILLER_6_908 VPWR VGND sg13g2_decap_8
XFILLER_5_429 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_1_668 VPWR VGND sg13g2_decap_8
XFILLER_48_138 VPWR VGND sg13g2_decap_8
XFILLER_0_189 VPWR VGND sg13g2_decap_8
XFILLER_45_801 VPWR VGND sg13g2_decap_8
XFILLER_28_74 VPWR VGND sg13g2_decap_8
XFILLER_17_536 VPWR VGND sg13g2_decap_8
XFILLER_28_85 VPWR VGND sg13g2_fill_2
XFILLER_45_878 VPWR VGND sg13g2_decap_8
X_563_ net63 VGND VPWR _060_ mac2.products_ff\[64\] clknet_5_8__leaf_clk sg13g2_dfrbpq_1
X_494_ net65 VGND VPWR _116_ DP_3.matrix\[80\] clknet_5_11__leaf_clk sg13g2_dfrbpq_1
XFILLER_9_702 VPWR VGND sg13g2_decap_8
XFILLER_13_753 VPWR VGND sg13g2_decap_8
XFILLER_8_212 VPWR VGND sg13g2_decap_8
XFILLER_40_572 VPWR VGND sg13g2_decap_8
XFILLER_12_274 VPWR VGND sg13g2_decap_8
XFILLER_9_779 VPWR VGND sg13g2_decap_8
XFILLER_8_267 VPWR VGND sg13g2_decap_8
XFILLER_5_974 VPWR VGND sg13g2_decap_8
XFILLER_4_495 VPWR VGND sg13g2_decap_8
XFILLER_10_4 VPWR VGND sg13g2_decap_8
XFILLER_47_160 VPWR VGND sg13g2_decap_8
XFILLER_36_834 VPWR VGND sg13g2_decap_8
XFILLER_39_1028 VPWR VGND sg13g2_fill_1
XFILLER_35_366 VPWR VGND sg13g2_decap_8
XFILLER_31_561 VPWR VGND sg13g2_decap_8
XFILLER_22_1010 VPWR VGND sg13g2_decap_8
XFILLER_27_812 VPWR VGND sg13g2_decap_8
XFILLER_38_182 VPWR VGND sg13g2_decap_8
XFILLER_39_683 VPWR VGND sg13g2_decap_8
XFILLER_26_333 VPWR VGND sg13g2_decap_8
XFILLER_42_815 VPWR VGND sg13g2_decap_8
XFILLER_14_539 VPWR VGND sg13g2_decap_8
XFILLER_27_889 VPWR VGND sg13g2_decap_8
XFILLER_41_314 VPWR VGND sg13g2_decap_8
XFILLER_14_32 VPWR VGND sg13g2_decap_8
XFILLER_22_550 VPWR VGND sg13g2_decap_8
XFILLER_10_734 VPWR VGND sg13g2_decap_8
XFILLER_22_583 VPWR VGND sg13g2_decap_8
XFILLER_6_705 VPWR VGND sg13g2_decap_8
XFILLER_5_226 VPWR VGND sg13g2_decap_8
XFILLER_2_900 VPWR VGND sg13g2_decap_8
XFILLER_30_42 VPWR VGND sg13g2_decap_8
XFILLER_2_977 VPWR VGND sg13g2_decap_8
XFILLER_1_465 VPWR VGND sg13g2_decap_8
XFILLER_49_447 VPWR VGND sg13g2_decap_8
XFILLER_39_73 VPWR VGND sg13g2_decap_8
Xclkbuf_4_3_0_clk clknet_0_clk clknet_4_3_0_clk VPWR VGND sg13g2_buf_8
XFILLER_37_609 VPWR VGND sg13g2_decap_8
XFILLER_17_300 VPWR VGND sg13g2_decap_8
XFILLER_29_171 VPWR VGND sg13g2_decap_8
XFILLER_36_119 VPWR VGND sg13g2_decap_8
XFILLER_18_856 VPWR VGND sg13g2_decap_8
XFILLER_45_675 VPWR VGND sg13g2_decap_8
X_546_ net70 VGND VPWR net103 mac1.sum_lvl2_ff\[4\] clknet_5_19__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_377 VPWR VGND sg13g2_decap_8
XFILLER_32_325 VPWR VGND sg13g2_decap_8
X_477_ net78 VGND VPWR _099_ DP_2.matrix\[81\] clknet_5_29__leaf_clk sg13g2_dfrbpq_1
XFILLER_41_870 VPWR VGND sg13g2_decap_8
XFILLER_9_543 VPWR VGND sg13g2_decap_8
XFILLER_13_572 VPWR VGND sg13g2_decap_8
XFILLER_9_576 VPWR VGND sg13g2_decap_8
XFILLER_5_771 VPWR VGND sg13g2_decap_8
XFILLER_35_130 VPWR VGND sg13g2_decap_8
XFILLER_36_631 VPWR VGND sg13g2_decap_8
XFILLER_23_325 VPWR VGND sg13g2_decap_8
XFILLER_24_859 VPWR VGND sg13g2_decap_8
XFILLER_31_391 VPWR VGND sg13g2_decap_8
XFILLER_3_719 VPWR VGND sg13g2_decap_8
XFILLER_19_609 VPWR VGND sg13g2_decap_8
XFILLER_46_428 VPWR VGND sg13g2_decap_8
XFILLER_42_612 VPWR VGND sg13g2_decap_8
X_400_ net132 _094_ VPWR VGND sg13g2_buf_1
XFILLER_14_303 VPWR VGND sg13g2_fill_1
XFILLER_15_804 VPWR VGND sg13g2_decap_8
XFILLER_27_686 VPWR VGND sg13g2_decap_8
XFILLER_14_336 VPWR VGND sg13g2_decap_8
X_331_ _193_ _192_ _041_ VPWR VGND sg13g2_xor2_1
XFILLER_42_689 VPWR VGND sg13g2_decap_8
XFILLER_30_807 VPWR VGND sg13g2_decap_8
XFILLER_41_133 VPWR VGND sg13g2_decap_8
X_262_ net102 mac1.sum_lvl1_ff\[24\] _010_ VPWR VGND sg13g2_xor2_1
XFILLER_41_188 VPWR VGND sg13g2_decap_8
XFILLER_10_542 VPWR VGND sg13g2_decap_8
XFILLER_6_524 VPWR VGND sg13g2_decap_8
XFILLER_41_63 VPWR VGND sg13g2_decap_8
XFILLER_6_579 VPWR VGND sg13g2_decap_8
XFILLER_2_774 VPWR VGND sg13g2_decap_8
XFILLER_1_262 VPWR VGND sg13g2_decap_8
XFILLER_49_266 VPWR VGND sg13g2_decap_8
XFILLER_2_46 VPWR VGND sg13g2_decap_8
XFILLER_38_929 VPWR VGND sg13g2_decap_8
XFILLER_37_428 VPWR VGND sg13g2_decap_8
XFILLER_18_653 VPWR VGND sg13g2_decap_8
XFILLER_46_995 VPWR VGND sg13g2_decap_8
XFILLER_45_472 VPWR VGND sg13g2_decap_8
XFILLER_17_163 VPWR VGND sg13g2_decap_8
XFILLER_17_185 VPWR VGND sg13g2_fill_1
XFILLER_32_111 VPWR VGND sg13g2_fill_1
XFILLER_36_1009 VPWR VGND sg13g2_decap_8
X_529_ net61 VGND VPWR _059_ mac1.products_ff\[129\] clknet_5_4__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_667 VPWR VGND sg13g2_decap_8
XFILLER_14_870 VPWR VGND sg13g2_decap_8
XFILLER_12_1020 VPWR VGND sg13g2_decap_8
XFILLER_49_0 VPWR VGND sg13g2_decap_8
XFILLER_28_406 VPWR VGND sg13g2_decap_8
XFILLER_37_973 VPWR VGND sg13g2_decap_8
XFILLER_23_100 VPWR VGND sg13g2_decap_4
XFILLER_23_155 VPWR VGND sg13g2_decap_8
XFILLER_24_656 VPWR VGND sg13g2_decap_8
XFILLER_11_328 VPWR VGND sg13g2_decap_8
XFILLER_20_873 VPWR VGND sg13g2_decap_8
XFILLER_11_11 VPWR VGND sg13g2_decap_4
XFILLER_11_44 VPWR VGND sg13g2_decap_8
XFILLER_4_1007 VPWR VGND sg13g2_decap_8
XFILLER_47_737 VPWR VGND sg13g2_decap_8
XFILLER_43_910 VPWR VGND sg13g2_decap_8
XFILLER_15_601 VPWR VGND sg13g2_decap_8
XFILLER_28_995 VPWR VGND sg13g2_decap_8
XFILLER_36_63 VPWR VGND sg13g2_decap_8
XFILLER_27_483 VPWR VGND sg13g2_decap_8
XFILLER_43_987 VPWR VGND sg13g2_decap_8
XFILLER_42_464 VPWR VGND sg13g2_fill_2
XFILLER_42_453 VPWR VGND sg13g2_fill_2
XFILLER_14_144 VPWR VGND sg13g2_decap_8
XFILLER_15_678 VPWR VGND sg13g2_decap_8
XFILLER_30_604 VPWR VGND sg13g2_decap_8
X_314_ _183_ net170 mac2.sum_lvl3_ff\[3\] VPWR VGND sg13g2_nand2_1
X_245_ _143_ VPWR _146_ VGND _142_ _144_ sg13g2_o21ai_1
XFILLER_7_800 VPWR VGND sg13g2_decap_8
XFILLER_11_851 VPWR VGND sg13g2_decap_8
XFILLER_10_383 VPWR VGND sg13g2_fill_1
XFILLER_7_877 VPWR VGND sg13g2_decap_8
XFILLER_6_387 VPWR VGND sg13g2_decap_8
XFILLER_6_365 VPWR VGND sg13g2_decap_8
XFILLER_42_7 VPWR VGND sg13g2_decap_8
XFILLER_2_571 VPWR VGND sg13g2_decap_8
XFILLER_38_726 VPWR VGND sg13g2_decap_8
XFILLER_19_973 VPWR VGND sg13g2_decap_8
XFILLER_37_258 VPWR VGND sg13g2_decap_8
XFILLER_46_792 VPWR VGND sg13g2_decap_8
XFILLER_34_932 VPWR VGND sg13g2_decap_8
XFILLER_33_475 VPWR VGND sg13g2_fill_1
XFILLER_21_659 VPWR VGND sg13g2_decap_8
XFILLER_43_206 VPWR VGND sg13g2_decap_8
XFILLER_37_770 VPWR VGND sg13g2_decap_8
XFILLER_19_1015 VPWR VGND sg13g2_decap_8
XFILLER_24_453 VPWR VGND sg13g2_decap_8
XFILLER_25_965 VPWR VGND sg13g2_decap_8
XFILLER_40_957 VPWR VGND sg13g2_decap_8
XFILLER_20_670 VPWR VGND sg13g2_decap_8
XFILLER_22_43 VPWR VGND sg13g2_decap_8
XFILLER_4_825 VPWR VGND sg13g2_decap_8
XFILLER_3_313 VPWR VGND sg13g2_decap_4
XFILLER_47_534 VPWR VGND sg13g2_decap_8
XFILLER_47_51 VPWR VGND sg13g2_fill_1
XFILLER_35_729 VPWR VGND sg13g2_decap_8
XFILLER_16_943 VPWR VGND sg13g2_decap_8
XFILLER_28_792 VPWR VGND sg13g2_decap_8
XFILLER_34_217 VPWR VGND sg13g2_decap_8
Xclkbuf_5_21__f_clk clknet_4_10_0_clk clknet_5_21__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_43_784 VPWR VGND sg13g2_decap_8
XFILLER_31_946 VPWR VGND sg13g2_decap_8
XFILLER_42_294 VPWR VGND sg13g2_decap_8
XFILLER_15_497 VPWR VGND sg13g2_decap_8
XFILLER_8_67 VPWR VGND sg13g2_decap_8
XFILLER_30_478 VPWR VGND sg13g2_decap_8
XFILLER_30_489 VPWR VGND sg13g2_fill_1
X_228_ net151 net140 _046_ VPWR VGND sg13g2_and2_1
XFILLER_7_674 VPWR VGND sg13g2_decap_8
XFILLER_3_880 VPWR VGND sg13g2_decap_8
XFILLER_38_523 VPWR VGND sg13g2_decap_8
XFILLER_19_770 VPWR VGND sg13g2_decap_8
XFILLER_18_291 VPWR VGND sg13g2_decap_8
XFILLER_21_412 VPWR VGND sg13g2_fill_2
XFILLER_40_209 VPWR VGND sg13g2_decap_8
XFILLER_22_968 VPWR VGND sg13g2_decap_8
XFILLER_21_489 VPWR VGND sg13g2_fill_2
XFILLER_48_309 VPWR VGND sg13g2_decap_8
XFILLER_17_21 VPWR VGND sg13g2_fill_2
XFILLER_29_567 VPWR VGND sg13g2_decap_8
XFILLER_16_217 VPWR VGND sg13g2_decap_8
XFILLER_17_87 VPWR VGND sg13g2_fill_1
XFILLER_25_762 VPWR VGND sg13g2_decap_8
XFILLER_13_935 VPWR VGND sg13g2_decap_8
XFILLER_24_250 VPWR VGND sg13g2_decap_8
XFILLER_40_754 VPWR VGND sg13g2_decap_8
XFILLER_8_416 VPWR VGND sg13g2_decap_8
XFILLER_33_53 VPWR VGND sg13g2_decap_8
XFILLER_32_1023 VPWR VGND sg13g2_decap_4
XFILLER_4_622 VPWR VGND sg13g2_decap_8
XFILLER_3_143 VPWR VGND sg13g2_decap_8
XFILLER_4_699 VPWR VGND sg13g2_decap_8
XFILLER_48_821 VPWR VGND sg13g2_decap_8
XFILLER_0_861 VPWR VGND sg13g2_decap_8
XFILLER_39_309 VPWR VGND sg13g2_fill_1
Xhold5 mac1.sum_lvl2_ff\[9\] VPWR VGND net29 sg13g2_dlygate4sd3_1
XFILLER_48_898 VPWR VGND sg13g2_decap_8
XFILLER_35_526 VPWR VGND sg13g2_decap_8
XFILLER_16_740 VPWR VGND sg13g2_decap_8
XFILLER_15_261 VPWR VGND sg13g2_decap_8
XFILLER_43_581 VPWR VGND sg13g2_decap_8
XFILLER_31_743 VPWR VGND sg13g2_decap_8
XFILLER_8_950 VPWR VGND sg13g2_decap_8
XFILLER_30_297 VPWR VGND sg13g2_decap_8
XFILLER_7_471 VPWR VGND sg13g2_decap_4
XFILLER_31_0 VPWR VGND sg13g2_decap_8
XFILLER_26_504 VPWR VGND sg13g2_decap_8
XFILLER_38_342 VPWR VGND sg13g2_decap_8
XFILLER_39_865 VPWR VGND sg13g2_decap_8
XFILLER_10_916 VPWR VGND sg13g2_decap_8
XFILLER_21_253 VPWR VGND sg13g2_decap_8
XFILLER_21_264 VPWR VGND sg13g2_fill_2
XFILLER_22_765 VPWR VGND sg13g2_decap_8
XFILLER_1_647 VPWR VGND sg13g2_decap_8
XFILLER_49_629 VPWR VGND sg13g2_decap_8
XFILLER_48_117 VPWR VGND sg13g2_decap_8
XFILLER_0_168 VPWR VGND sg13g2_decap_8
XFILLER_29_331 VPWR VGND sg13g2_decap_8
XFILLER_29_375 VPWR VGND sg13g2_fill_2
X_562_ net65 VGND VPWR _039_ mac2.products_ff\[81\] clknet_5_10__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_857 VPWR VGND sg13g2_decap_8
XFILLER_44_378 VPWR VGND sg13g2_decap_4
XFILLER_25_570 VPWR VGND sg13g2_decap_8
X_493_ net63 VGND VPWR _115_ DP_3.matrix\[65\] clknet_5_8__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_96 VPWR VGND sg13g2_decap_8
XFILLER_13_732 VPWR VGND sg13g2_decap_8
XFILLER_12_253 VPWR VGND sg13g2_decap_8
XFILLER_40_551 VPWR VGND sg13g2_decap_8
XFILLER_9_758 VPWR VGND sg13g2_decap_8
XFILLER_5_953 VPWR VGND sg13g2_decap_8
XFILLER_4_474 VPWR VGND sg13g2_decap_8
XFILLER_36_813 VPWR VGND sg13g2_decap_8
XFILLER_48_695 VPWR VGND sg13g2_decap_8
XFILLER_35_323 VPWR VGND sg13g2_decap_8
XFILLER_31_540 VPWR VGND sg13g2_decap_8
XFILLER_39_662 VPWR VGND sg13g2_decap_8
XFILLER_26_312 VPWR VGND sg13g2_decap_8
XFILLER_38_172 VPWR VGND sg13g2_fill_1
XFILLER_27_868 VPWR VGND sg13g2_decap_8
XFILLER_14_518 VPWR VGND sg13g2_decap_8
XFILLER_26_389 VPWR VGND sg13g2_decap_8
XFILLER_14_11 VPWR VGND sg13g2_decap_8
XFILLER_35_890 VPWR VGND sg13g2_decap_8
XFILLER_10_713 VPWR VGND sg13g2_decap_8
XFILLER_14_88 VPWR VGND sg13g2_decap_8
XFILLER_5_205 VPWR VGND sg13g2_decap_8
XFILLER_30_21 VPWR VGND sg13g2_decap_8
XFILLER_30_98 VPWR VGND sg13g2_decap_8
XFILLER_2_956 VPWR VGND sg13g2_decap_8
XFILLER_1_444 VPWR VGND sg13g2_decap_8
XFILLER_49_426 VPWR VGND sg13g2_decap_8
XFILLER_18_835 VPWR VGND sg13g2_decap_8
XFILLER_29_150 VPWR VGND sg13g2_decap_8
XFILLER_45_654 VPWR VGND sg13g2_decap_8
XFILLER_44_131 VPWR VGND sg13g2_decap_8
XFILLER_44_142 VPWR VGND sg13g2_fill_2
XFILLER_17_356 VPWR VGND sg13g2_decap_8
X_545_ net73 VGND VPWR _057_ mac1.products_ff\[17\] clknet_5_23__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_304 VPWR VGND sg13g2_decap_8
XFILLER_33_849 VPWR VGND sg13g2_decap_8
XFILLER_13_551 VPWR VGND sg13g2_decap_8
X_476_ net78 VGND VPWR _098_ DP_2.matrix\[80\] clknet_5_29__leaf_clk sg13g2_dfrbpq_1
XFILLER_9_522 VPWR VGND sg13g2_decap_8
XFILLER_5_750 VPWR VGND sg13g2_decap_8
XFILLER_45_1011 VPWR VGND sg13g2_decap_8
XFILLER_4_282 VPWR VGND sg13g2_decap_8
XFILLER_49_993 VPWR VGND sg13g2_decap_8
XFILLER_36_610 VPWR VGND sg13g2_decap_8
XFILLER_48_492 VPWR VGND sg13g2_decap_8
XFILLER_23_304 VPWR VGND sg13g2_decap_8
XFILLER_24_838 VPWR VGND sg13g2_decap_8
XFILLER_36_687 VPWR VGND sg13g2_decap_8
XFILLER_35_186 VPWR VGND sg13g2_decap_8
XFILLER_31_370 VPWR VGND sg13g2_decap_8
XFILLER_47_919 VPWR VGND sg13g2_decap_8
XFILLER_46_407 VPWR VGND sg13g2_decap_8
XFILLER_39_470 VPWR VGND sg13g2_decap_8
XFILLER_39_481 VPWR VGND sg13g2_decap_4
Xclkbuf_5_2__f_clk clknet_4_1_0_clk clknet_5_2__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_27_665 VPWR VGND sg13g2_decap_8
XFILLER_25_32 VPWR VGND sg13g2_decap_8
X_330_ _193_ net137 net94 VPWR VGND sg13g2_nand2_1
XFILLER_41_112 VPWR VGND sg13g2_decap_8
XFILLER_42_668 VPWR VGND sg13g2_decap_8
XFILLER_25_87 VPWR VGND sg13g2_decap_8
X_261_ _011_ _154_ _155_ VPWR VGND sg13g2_xnor2_1
XFILLER_10_521 VPWR VGND sg13g2_decap_8
XFILLER_6_503 VPWR VGND sg13g2_decap_8
XFILLER_41_42 VPWR VGND sg13g2_decap_8
XFILLER_6_558 VPWR VGND sg13g2_decap_8
XFILLER_2_753 VPWR VGND sg13g2_decap_8
XFILLER_1_241 VPWR VGND sg13g2_decap_8
XFILLER_2_25 VPWR VGND sg13g2_decap_8
XFILLER_49_245 VPWR VGND sg13g2_decap_8
XFILLER_38_908 VPWR VGND sg13g2_decap_8
XFILLER_37_407 VPWR VGND sg13g2_fill_1
XFILLER_18_632 VPWR VGND sg13g2_decap_8
XFILLER_46_974 VPWR VGND sg13g2_decap_8
XFILLER_45_451 VPWR VGND sg13g2_decap_8
XFILLER_17_142 VPWR VGND sg13g2_decap_8
XFILLER_33_646 VPWR VGND sg13g2_decap_8
X_528_ net59 VGND VPWR _058_ mac1.products_ff\[128\] clknet_5_4__leaf_clk sg13g2_dfrbpq_1
X_459_ net80 VGND VPWR _081_ DP_1.matrix\[81\] clknet_5_30__leaf_clk sg13g2_dfrbpq_1
XFILLER_9_396 VPWR VGND sg13g2_decap_8
XFILLER_49_790 VPWR VGND sg13g2_decap_8
XFILLER_37_952 VPWR VGND sg13g2_decap_8
XFILLER_36_451 VPWR VGND sg13g2_decap_4
XFILLER_24_635 VPWR VGND sg13g2_decap_8
XFILLER_36_484 VPWR VGND sg13g2_decap_8
XFILLER_23_134 VPWR VGND sg13g2_decap_8
XFILLER_11_307 VPWR VGND sg13g2_decap_8
XFILLER_20_852 VPWR VGND sg13g2_decap_8
Xclkbuf_4_2_0_clk clknet_0_clk clknet_4_2_0_clk VPWR VGND sg13g2_buf_8
XFILLER_47_716 VPWR VGND sg13g2_decap_8
XFILLER_46_204 VPWR VGND sg13g2_decap_8
XFILLER_27_440 VPWR VGND sg13g2_fill_2
XFILLER_28_974 VPWR VGND sg13g2_decap_8
XFILLER_36_42 VPWR VGND sg13g2_decap_8
XFILLER_43_966 VPWR VGND sg13g2_decap_8
XFILLER_42_443 VPWR VGND sg13g2_fill_2
XFILLER_14_123 VPWR VGND sg13g2_decap_8
XFILLER_15_657 VPWR VGND sg13g2_decap_8
X_313_ _182_ net207 net107 VPWR VGND sg13g2_nand2_1
X_244_ net2 _142_ _145_ VPWR VGND sg13g2_xnor2_1
XFILLER_11_830 VPWR VGND sg13g2_decap_8
XFILLER_10_362 VPWR VGND sg13g2_decap_8
XFILLER_7_856 VPWR VGND sg13g2_decap_8
XFILLER_6_344 VPWR VGND sg13g2_decap_8
XFILLER_35_7 VPWR VGND sg13g2_decap_8
XFILLER_42_1025 VPWR VGND sg13g2_decap_4
XFILLER_38_705 VPWR VGND sg13g2_decap_8
XFILLER_19_952 VPWR VGND sg13g2_decap_8
XFILLER_37_237 VPWR VGND sg13g2_decap_8
XFILLER_46_771 VPWR VGND sg13g2_decap_8
XFILLER_34_911 VPWR VGND sg13g2_decap_8
XFILLER_18_484 VPWR VGND sg13g2_decap_8
XFILLER_33_443 VPWR VGND sg13g2_fill_2
XFILLER_34_988 VPWR VGND sg13g2_decap_8
XFILLER_21_638 VPWR VGND sg13g2_decap_8
XFILLER_20_126 VPWR VGND sg13g2_decap_8
XFILLER_9_193 VPWR VGND sg13g2_decap_8
XFILLER_28_204 VPWR VGND sg13g2_decap_8
XFILLER_29_749 VPWR VGND sg13g2_decap_8
XFILLER_28_259 VPWR VGND sg13g2_fill_2
XFILLER_25_944 VPWR VGND sg13g2_decap_8
XFILLER_24_432 VPWR VGND sg13g2_decap_8
XFILLER_36_292 VPWR VGND sg13g2_fill_1
XFILLER_40_936 VPWR VGND sg13g2_decap_8
XFILLER_12_649 VPWR VGND sg13g2_decap_8
XFILLER_7_119 VPWR VGND sg13g2_fill_1
XFILLER_22_11 VPWR VGND sg13g2_decap_4
XFILLER_4_804 VPWR VGND sg13g2_decap_8
XFILLER_47_513 VPWR VGND sg13g2_decap_8
XFILLER_47_85 VPWR VGND sg13g2_decap_4
XFILLER_19_248 VPWR VGND sg13g2_decap_8
XFILLER_35_708 VPWR VGND sg13g2_decap_8
XFILLER_16_922 VPWR VGND sg13g2_decap_8
XFILLER_28_771 VPWR VGND sg13g2_decap_8
XFILLER_43_763 VPWR VGND sg13g2_decap_8
XFILLER_15_421 VPWR VGND sg13g2_fill_1
XFILLER_15_476 VPWR VGND sg13g2_decap_8
XFILLER_16_999 VPWR VGND sg13g2_decap_8
XFILLER_31_925 VPWR VGND sg13g2_decap_8
XFILLER_8_46 VPWR VGND sg13g2_decap_8
X_227_ net143 net146 _044_ VPWR VGND sg13g2_and2_1
XFILLER_7_653 VPWR VGND sg13g2_decap_8
XFILLER_6_152 VPWR VGND sg13g2_decap_8
XFILLER_26_719 VPWR VGND sg13g2_decap_8
XFILLER_38_579 VPWR VGND sg13g2_decap_8
XFILLER_18_270 VPWR VGND sg13g2_decap_8
XFILLER_34_785 VPWR VGND sg13g2_decap_8
XFILLER_22_947 VPWR VGND sg13g2_decap_8
XFILLER_33_273 VPWR VGND sg13g2_decap_8
XFILLER_21_457 VPWR VGND sg13g2_decap_4
XFILLER_1_829 VPWR VGND sg13g2_decap_8
XFILLER_29_546 VPWR VGND sg13g2_decap_8
XFILLER_17_719 VPWR VGND sg13g2_decap_8
XFILLER_17_55 VPWR VGND sg13g2_fill_2
XFILLER_44_549 VPWR VGND sg13g2_decap_8
XFILLER_25_741 VPWR VGND sg13g2_decap_8
XFILLER_13_914 VPWR VGND sg13g2_decap_8
XFILLER_40_733 VPWR VGND sg13g2_decap_8
XFILLER_12_479 VPWR VGND sg13g2_fill_2
XFILLER_32_1002 VPWR VGND sg13g2_decap_8
XFILLER_4_601 VPWR VGND sg13g2_decap_8
XFILLER_20_490 VPWR VGND sg13g2_decap_8
XFILLER_4_678 VPWR VGND sg13g2_decap_8
XFILLER_0_840 VPWR VGND sg13g2_decap_8
XFILLER_48_800 VPWR VGND sg13g2_decap_8
Xhold6 mac2.sum_lvl1_ff\[32\] VPWR VGND net30 sg13g2_dlygate4sd3_1
XFILLER_48_877 VPWR VGND sg13g2_decap_8
XFILLER_47_365 VPWR VGND sg13g2_decap_8
XFILLER_35_505 VPWR VGND sg13g2_decap_8
XFILLER_43_560 VPWR VGND sg13g2_decap_8
XFILLER_16_796 VPWR VGND sg13g2_decap_8
XFILLER_31_722 VPWR VGND sg13g2_decap_8
XFILLER_30_276 VPWR VGND sg13g2_decap_8
XFILLER_31_799 VPWR VGND sg13g2_decap_8
XFILLER_7_450 VPWR VGND sg13g2_decap_8
XFILLER_38_321 VPWR VGND sg13g2_decap_8
XFILLER_39_844 VPWR VGND sg13g2_decap_8
XFILLER_38_398 VPWR VGND sg13g2_decap_8
XFILLER_0_1022 VPWR VGND sg13g2_decap_8
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_22_744 VPWR VGND sg13g2_decap_8
XFILLER_34_582 VPWR VGND sg13g2_decap_8
XFILLER_21_232 VPWR VGND sg13g2_decap_4
XFILLER_1_626 VPWR VGND sg13g2_decap_8
XFILLER_49_608 VPWR VGND sg13g2_decap_8
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_29_310 VPWR VGND sg13g2_decap_8
XFILLER_29_354 VPWR VGND sg13g2_decap_8
XFILLER_45_836 VPWR VGND sg13g2_decap_8
X_561_ net65 VGND VPWR _038_ mac2.products_ff\[80\] clknet_5_11__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_357 VPWR VGND sg13g2_decap_8
XFILLER_13_711 VPWR VGND sg13g2_decap_8
XFILLER_32_519 VPWR VGND sg13g2_decap_8
X_492_ net68 VGND VPWR _114_ DP_3.matrix\[64\] clknet_5_10__leaf_clk sg13g2_dfrbpq_1
XFILLER_44_75 VPWR VGND sg13g2_fill_1
XFILLER_40_530 VPWR VGND sg13g2_decap_8
XFILLER_12_232 VPWR VGND sg13g2_decap_8
XFILLER_9_737 VPWR VGND sg13g2_decap_8
XFILLER_13_788 VPWR VGND sg13g2_decap_8
XFILLER_12_298 VPWR VGND sg13g2_decap_8
XFILLER_5_932 VPWR VGND sg13g2_decap_8
XFILLER_4_420 VPWR VGND sg13g2_fill_1
XFILLER_4_453 VPWR VGND sg13g2_decap_8
XFILLER_39_129 VPWR VGND sg13g2_decap_8
XFILLER_48_674 VPWR VGND sg13g2_decap_8
XFILLER_35_302 VPWR VGND sg13g2_decap_8
XFILLER_36_869 VPWR VGND sg13g2_decap_8
XFILLER_39_1019 VPWR VGND sg13g2_decap_8
XFILLER_16_593 VPWR VGND sg13g2_decap_8
XFILLER_31_596 VPWR VGND sg13g2_decap_8
XFILLER_39_641 VPWR VGND sg13g2_decap_8
XFILLER_27_847 VPWR VGND sg13g2_decap_8
XFILLER_26_368 VPWR VGND sg13g2_decap_8
XFILLER_22_530 VPWR VGND sg13g2_decap_8
XFILLER_14_67 VPWR VGND sg13g2_decap_8
XFILLER_10_769 VPWR VGND sg13g2_decap_8
XFILLER_30_77 VPWR VGND sg13g2_decap_8
XFILLER_2_935 VPWR VGND sg13g2_decap_8
XFILLER_1_423 VPWR VGND sg13g2_decap_8
XFILLER_49_405 VPWR VGND sg13g2_decap_8
XFILLER_7_1017 VPWR VGND sg13g2_decap_8
XFILLER_7_1028 VPWR VGND sg13g2_fill_1
XFILLER_18_814 VPWR VGND sg13g2_decap_8
XFILLER_45_633 VPWR VGND sg13g2_decap_8
XFILLER_44_110 VPWR VGND sg13g2_decap_8
XFILLER_17_335 VPWR VGND sg13g2_decap_8
X_544_ net74 VGND VPWR _056_ mac1.products_ff\[16\] clknet_5_22__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_828 VPWR VGND sg13g2_decap_8
XFILLER_44_198 VPWR VGND sg13g2_fill_2
XFILLER_44_187 VPWR VGND sg13g2_decap_8
XFILLER_26_880 VPWR VGND sg13g2_decap_8
X_475_ net77 VGND VPWR _097_ DP_2.matrix\[65\] clknet_5_30__leaf_clk sg13g2_dfrbpq_1
XFILLER_1_990 VPWR VGND sg13g2_decap_8
XFILLER_49_972 VPWR VGND sg13g2_decap_8
XFILLER_48_471 VPWR VGND sg13g2_decap_8
XFILLER_24_817 VPWR VGND sg13g2_decap_8
XFILLER_35_165 VPWR VGND sg13g2_decap_8
XFILLER_36_666 VPWR VGND sg13g2_decap_8
XFILLER_17_880 VPWR VGND sg13g2_decap_8
XFILLER_32_883 VPWR VGND sg13g2_decap_8
XFILLER_27_644 VPWR VGND sg13g2_decap_8
XFILLER_25_11 VPWR VGND sg13g2_decap_8
XFILLER_42_647 VPWR VGND sg13g2_decap_8
XFILLER_15_839 VPWR VGND sg13g2_decap_8
XFILLER_26_176 VPWR VGND sg13g2_decap_8
XFILLER_25_66 VPWR VGND sg13g2_decap_8
XFILLER_10_500 VPWR VGND sg13g2_decap_8
X_260_ mac1.sum_lvl1_ff\[17\] mac1.sum_lvl1_ff\[25\] _155_ VPWR VGND sg13g2_xor2_1
XFILLER_23_894 VPWR VGND sg13g2_decap_8
XFILLER_41_168 VPWR VGND sg13g2_fill_2
XFILLER_41_21 VPWR VGND sg13g2_decap_8
XFILLER_2_732 VPWR VGND sg13g2_decap_8
XFILLER_1_220 VPWR VGND sg13g2_decap_8
XFILLER_49_224 VPWR VGND sg13g2_decap_8
XFILLER_1_297 VPWR VGND sg13g2_decap_8
XFILLER_46_953 VPWR VGND sg13g2_decap_8
XFILLER_45_430 VPWR VGND sg13g2_decap_8
X_527_ net71 VGND VPWR net183 mac1.sum_lvl1_ff\[9\] clknet_5_20__leaf_clk sg13g2_dfrbpq_1
XFILLER_18_688 VPWR VGND sg13g2_decap_8
XFILLER_32_102 VPWR VGND sg13g2_decap_8
XFILLER_33_625 VPWR VGND sg13g2_decap_8
XFILLER_32_146 VPWR VGND sg13g2_decap_8
XFILLER_20_308 VPWR VGND sg13g2_decap_8
X_458_ net73 VGND VPWR _080_ DP_1.matrix\[80\] clknet_5_28__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_179 VPWR VGND sg13g2_decap_8
X_389_ net48 _083_ VPWR VGND sg13g2_buf_1
XFILLER_9_375 VPWR VGND sg13g2_decap_8
XFILLER_37_931 VPWR VGND sg13g2_decap_8
XFILLER_36_430 VPWR VGND sg13g2_decap_8
XFILLER_23_113 VPWR VGND sg13g2_decap_8
XFILLER_24_614 VPWR VGND sg13g2_decap_8
XFILLER_20_831 VPWR VGND sg13g2_decap_8
XFILLER_32_680 VPWR VGND sg13g2_decap_8
XFILLER_3_529 VPWR VGND sg13g2_decap_8
XFILLER_28_953 VPWR VGND sg13g2_decap_8
XFILLER_36_21 VPWR VGND sg13g2_decap_8
XFILLER_43_945 VPWR VGND sg13g2_decap_8
XFILLER_42_422 VPWR VGND sg13g2_decap_8
XFILLER_14_102 VPWR VGND sg13g2_decap_8
XFILLER_15_636 VPWR VGND sg13g2_decap_8
XFILLER_36_98 VPWR VGND sg13g2_decap_8
XFILLER_14_179 VPWR VGND sg13g2_fill_2
X_312_ net117 mac2.products_ff\[48\] _019_ VPWR VGND sg13g2_xor2_1
X_243_ mac2.total_sum\[1\] mac1.total_sum\[1\] _145_ VPWR VGND sg13g2_xor2_1
XFILLER_23_691 VPWR VGND sg13g2_decap_8
XFILLER_30_639 VPWR VGND sg13g2_decap_8
XFILLER_11_886 VPWR VGND sg13g2_decap_8
XFILLER_7_835 VPWR VGND sg13g2_decap_8
XFILLER_42_1004 VPWR VGND sg13g2_decap_8
XFILLER_19_931 VPWR VGND sg13g2_decap_8
XFILLER_37_216 VPWR VGND sg13g2_decap_8
XFILLER_46_750 VPWR VGND sg13g2_decap_8
XFILLER_18_463 VPWR VGND sg13g2_decap_8
XFILLER_45_282 VPWR VGND sg13g2_decap_8
XFILLER_34_967 VPWR VGND sg13g2_decap_8
XFILLER_21_617 VPWR VGND sg13g2_decap_8
XFILLER_33_466 VPWR VGND sg13g2_decap_8
XFILLER_33_499 VPWR VGND sg13g2_decap_8
XFILLER_13_190 VPWR VGND sg13g2_decap_8
XFILLER_29_728 VPWR VGND sg13g2_decap_8
XFILLER_3_1020 VPWR VGND sg13g2_decap_8
XFILLER_28_238 VPWR VGND sg13g2_decap_8
XFILLER_24_411 VPWR VGND sg13g2_decap_8
XFILLER_25_923 VPWR VGND sg13g2_decap_8
XFILLER_36_260 VPWR VGND sg13g2_decap_8
XFILLER_24_488 VPWR VGND sg13g2_decap_8
XFILLER_40_915 VPWR VGND sg13g2_decap_8
XFILLER_11_149 VPWR VGND sg13g2_decap_8
XFILLER_22_78 VPWR VGND sg13g2_decap_4
XFILLER_3_359 VPWR VGND sg13g2_decap_8
XFILLER_47_42 VPWR VGND sg13g2_decap_8
XFILLER_19_216 VPWR VGND sg13g2_decap_8
XFILLER_47_569 VPWR VGND sg13g2_decap_8
XFILLER_16_901 VPWR VGND sg13g2_decap_8
XFILLER_28_750 VPWR VGND sg13g2_decap_8
XFILLER_27_260 VPWR VGND sg13g2_fill_2
XFILLER_43_742 VPWR VGND sg13g2_decap_8
XFILLER_16_978 VPWR VGND sg13g2_decap_8
XFILLER_15_455 VPWR VGND sg13g2_decap_8
XFILLER_30_403 VPWR VGND sg13g2_decap_4
XFILLER_31_904 VPWR VGND sg13g2_decap_8
XFILLER_8_25 VPWR VGND sg13g2_decap_8
XFILLER_7_632 VPWR VGND sg13g2_decap_8
XFILLER_11_683 VPWR VGND sg13g2_decap_8
X_226_ net154 net156 _042_ VPWR VGND sg13g2_and2_1
XFILLER_6_131 VPWR VGND sg13g2_decap_8
XFILLER_2_370 VPWR VGND sg13g2_decap_8
XFILLER_26_4 VPWR VGND sg13g2_decap_8
Xclkbuf_4_1_0_clk clknet_0_clk clknet_4_1_0_clk VPWR VGND sg13g2_buf_8
XFILLER_38_558 VPWR VGND sg13g2_decap_8
XFILLER_22_926 VPWR VGND sg13g2_decap_8
XFILLER_33_252 VPWR VGND sg13g2_decap_8
XFILLER_34_764 VPWR VGND sg13g2_decap_8
XFILLER_21_436 VPWR VGND sg13g2_decap_8
XFILLER_1_808 VPWR VGND sg13g2_decap_8
XFILLER_0_329 VPWR VGND sg13g2_decap_8
XFILLER_25_1021 VPWR VGND sg13g2_decap_8
XFILLER_29_525 VPWR VGND sg13g2_decap_8
XFILLER_17_23 VPWR VGND sg13g2_fill_1
XFILLER_44_528 VPWR VGND sg13g2_decap_8
XFILLER_17_78 VPWR VGND sg13g2_decap_8
XFILLER_25_720 VPWR VGND sg13g2_decap_8
XFILLER_40_712 VPWR VGND sg13g2_decap_8
XFILLER_24_285 VPWR VGND sg13g2_decap_8
XFILLER_25_797 VPWR VGND sg13g2_decap_8
XFILLER_9_919 VPWR VGND sg13g2_decap_8
XFILLER_12_458 VPWR VGND sg13g2_decap_8
XFILLER_21_981 VPWR VGND sg13g2_decap_8
XFILLER_40_789 VPWR VGND sg13g2_decap_8
XFILLER_4_657 VPWR VGND sg13g2_decap_8
XFILLER_47_322 VPWR VGND sg13g2_decap_4
XFILLER_47_311 VPWR VGND sg13g2_decap_8
Xhold7 mac1.sum_lvl2_ff\[8\] VPWR VGND net31 sg13g2_dlygate4sd3_1
XFILLER_0_896 VPWR VGND sg13g2_decap_8
XFILLER_48_856 VPWR VGND sg13g2_decap_8
XFILLER_47_344 VPWR VGND sg13g2_decap_8
XFILLER_16_775 VPWR VGND sg13g2_decap_8
XFILLER_31_701 VPWR VGND sg13g2_decap_8
XFILLER_30_255 VPWR VGND sg13g2_decap_8
XFILLER_31_778 VPWR VGND sg13g2_decap_8
XFILLER_12_992 VPWR VGND sg13g2_decap_8
XFILLER_8_985 VPWR VGND sg13g2_decap_8
XFILLER_48_1010 VPWR VGND sg13g2_decap_8
XFILLER_39_823 VPWR VGND sg13g2_decap_8
XFILLER_17_0 VPWR VGND sg13g2_decap_8
XFILLER_0_1001 VPWR VGND sg13g2_decap_8
XFILLER_38_377 VPWR VGND sg13g2_decap_8
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_26_539 VPWR VGND sg13g2_fill_1
XFILLER_34_561 VPWR VGND sg13g2_decap_8
XFILLER_22_723 VPWR VGND sg13g2_decap_8
XFILLER_1_605 VPWR VGND sg13g2_decap_8
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_45_815 VPWR VGND sg13g2_decap_8
X_560_ net61 VGND VPWR net29 mac1.sum_lvl3_ff\[3\] clknet_5_16__leaf_clk sg13g2_dfrbpq_2
XFILLER_44_336 VPWR VGND sg13g2_decap_8
XFILLER_44_32 VPWR VGND sg13g2_fill_2
XFILLER_44_21 VPWR VGND sg13g2_decap_8
X_491_ net66 VGND VPWR _113_ DP_3.matrix\[49\] clknet_5_11__leaf_clk sg13g2_dfrbpq_1
XFILLER_12_211 VPWR VGND sg13g2_fill_2
XFILLER_25_594 VPWR VGND sg13g2_decap_8
XFILLER_9_716 VPWR VGND sg13g2_decap_8
XFILLER_13_767 VPWR VGND sg13g2_decap_8
XFILLER_8_226 VPWR VGND sg13g2_decap_8
XFILLER_40_586 VPWR VGND sg13g2_decap_8
XFILLER_5_911 VPWR VGND sg13g2_decap_8
XFILLER_4_432 VPWR VGND sg13g2_decap_8
XFILLER_5_988 VPWR VGND sg13g2_decap_8
XFILLER_39_108 VPWR VGND sg13g2_decap_8
XFILLER_48_653 VPWR VGND sg13g2_decap_8
XFILLER_0_693 VPWR VGND sg13g2_decap_8
XFILLER_47_174 VPWR VGND sg13g2_decap_8
XFILLER_36_848 VPWR VGND sg13g2_decap_8
XFILLER_44_892 VPWR VGND sg13g2_decap_8
XFILLER_43_380 VPWR VGND sg13g2_decap_8
XFILLER_31_575 VPWR VGND sg13g2_decap_8
XFILLER_8_782 VPWR VGND sg13g2_decap_8
XFILLER_39_620 VPWR VGND sg13g2_decap_8
XFILLER_22_1024 VPWR VGND sg13g2_decap_4
XFILLER_27_826 VPWR VGND sg13g2_decap_8
XFILLER_26_347 VPWR VGND sg13g2_decap_8
XFILLER_38_196 VPWR VGND sg13g2_decap_8
XFILLER_39_697 VPWR VGND sg13g2_decap_8
XFILLER_42_829 VPWR VGND sg13g2_decap_8
XFILLER_22_520 VPWR VGND sg13g2_decap_4
XFILLER_41_328 VPWR VGND sg13g2_decap_8
XFILLER_14_46 VPWR VGND sg13g2_decap_8
XFILLER_22_564 VPWR VGND sg13g2_decap_4
XFILLER_10_748 VPWR VGND sg13g2_decap_8
XFILLER_22_597 VPWR VGND sg13g2_decap_8
XFILLER_6_719 VPWR VGND sg13g2_decap_8
XFILLER_30_56 VPWR VGND sg13g2_decap_8
XFILLER_2_914 VPWR VGND sg13g2_decap_8
XFILLER_1_402 VPWR VGND sg13g2_decap_8
XFILLER_39_21 VPWR VGND sg13g2_fill_2
XFILLER_1_479 VPWR VGND sg13g2_decap_8
XFILLER_39_87 VPWR VGND sg13g2_decap_8
XFILLER_45_612 VPWR VGND sg13g2_decap_8
XFILLER_17_314 VPWR VGND sg13g2_decap_8
XFILLER_29_185 VPWR VGND sg13g2_decap_8
XFILLER_45_689 VPWR VGND sg13g2_decap_8
X_543_ net73 VGND VPWR net192 mac1.sum_lvl2_ff\[1\] clknet_5_22__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_807 VPWR VGND sg13g2_decap_8
X_474_ net77 VGND VPWR _096_ DP_2.matrix\[64\] clknet_5_24__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_339 VPWR VGND sg13g2_decap_8
XFILLER_38_1020 VPWR VGND sg13g2_decap_8
XFILLER_13_520 VPWR VGND sg13g2_decap_8
XFILLER_13_586 VPWR VGND sg13g2_decap_8
XFILLER_41_884 VPWR VGND sg13g2_decap_8
XFILLER_9_557 VPWR VGND sg13g2_decap_8
XFILLER_5_785 VPWR VGND sg13g2_decap_8
Xclkbuf_5_27__f_clk clknet_4_13_0_clk clknet_5_27__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_49_951 VPWR VGND sg13g2_decap_8
XFILLER_0_490 VPWR VGND sg13g2_decap_8
XFILLER_48_450 VPWR VGND sg13g2_decap_8
XFILLER_36_645 VPWR VGND sg13g2_decap_8
XFILLER_35_144 VPWR VGND sg13g2_decap_8
XFILLER_23_339 VPWR VGND sg13g2_fill_2
XFILLER_32_862 VPWR VGND sg13g2_decap_8
XFILLER_39_461 VPWR VGND sg13g2_fill_1
XFILLER_27_623 VPWR VGND sg13g2_decap_8
XFILLER_15_818 VPWR VGND sg13g2_decap_8
XFILLER_42_626 VPWR VGND sg13g2_decap_8
XFILLER_41_147 VPWR VGND sg13g2_decap_8
XFILLER_23_873 VPWR VGND sg13g2_decap_8
XFILLER_22_372 VPWR VGND sg13g2_decap_8
XFILLER_10_556 VPWR VGND sg13g2_fill_1
XFILLER_6_538 VPWR VGND sg13g2_decap_8
XFILLER_41_77 VPWR VGND sg13g2_decap_8
XFILLER_2_711 VPWR VGND sg13g2_decap_8
XFILLER_29_1008 VPWR VGND sg13g2_decap_8
XFILLER_49_203 VPWR VGND sg13g2_decap_8
XFILLER_2_788 VPWR VGND sg13g2_decap_8
XFILLER_1_276 VPWR VGND sg13g2_decap_8
XFILLER_46_932 VPWR VGND sg13g2_decap_8
XFILLER_18_667 VPWR VGND sg13g2_decap_8
XFILLER_33_604 VPWR VGND sg13g2_decap_8
XFILLER_45_486 VPWR VGND sg13g2_decap_8
X_526_ net71 VGND VPWR net110 mac1.sum_lvl1_ff\[8\] clknet_5_20__leaf_clk sg13g2_dfrbpq_1
XFILLER_13_361 VPWR VGND sg13g2_decap_4
XFILLER_14_884 VPWR VGND sg13g2_decap_8
X_457_ net77 VGND VPWR _079_ DP_1.matrix\[65\] clknet_5_26__leaf_clk sg13g2_dfrbpq_1
XFILLER_13_394 VPWR VGND sg13g2_decap_8
X_388_ net151 _082_ VPWR VGND sg13g2_buf_1
XFILLER_41_681 VPWR VGND sg13g2_decap_8
XFILLER_9_354 VPWR VGND sg13g2_decap_8
XFILLER_5_582 VPWR VGND sg13g2_decap_8
XFILLER_37_910 VPWR VGND sg13g2_decap_8
XFILLER_37_987 VPWR VGND sg13g2_decap_8
XFILLER_20_810 VPWR VGND sg13g2_decap_8
XFILLER_23_169 VPWR VGND sg13g2_decap_8
XFILLER_31_180 VPWR VGND sg13g2_decap_8
XFILLER_20_887 VPWR VGND sg13g2_decap_8
XFILLER_11_58 VPWR VGND sg13g2_decap_4
Xclkbuf_5_10__f_clk clknet_4_5_0_clk clknet_5_10__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_19_409 VPWR VGND sg13g2_decap_4
XFILLER_46_228 VPWR VGND sg13g2_decap_8
XFILLER_28_932 VPWR VGND sg13g2_decap_8
XFILLER_43_924 VPWR VGND sg13g2_decap_8
XFILLER_42_401 VPWR VGND sg13g2_decap_8
XFILLER_15_615 VPWR VGND sg13g2_decap_8
XFILLER_36_77 VPWR VGND sg13g2_decap_8
XFILLER_27_497 VPWR VGND sg13g2_decap_8
XFILLER_14_158 VPWR VGND sg13g2_decap_8
XFILLER_30_618 VPWR VGND sg13g2_decap_8
XFILLER_35_1023 VPWR VGND sg13g2_decap_4
X_311_ _020_ _180_ _181_ VPWR VGND sg13g2_xnor2_1
X_242_ mac1.total_sum\[1\] mac2.total_sum\[1\] _144_ VPWR VGND sg13g2_nor2_1
XFILLER_23_670 VPWR VGND sg13g2_decap_8
XFILLER_10_320 VPWR VGND sg13g2_fill_2
XFILLER_7_814 VPWR VGND sg13g2_decap_8
XFILLER_6_302 VPWR VGND sg13g2_decap_4
XFILLER_11_865 VPWR VGND sg13g2_decap_8
XFILLER_22_191 VPWR VGND sg13g2_decap_8
XFILLER_10_397 VPWR VGND sg13g2_decap_8
XFILLER_2_530 VPWR VGND sg13g2_fill_2
XFILLER_2_585 VPWR VGND sg13g2_decap_8
XFILLER_19_910 VPWR VGND sg13g2_decap_8
XFILLER_18_442 VPWR VGND sg13g2_decap_8
XFILLER_45_261 VPWR VGND sg13g2_decap_8
XFILLER_19_987 VPWR VGND sg13g2_decap_8
XFILLER_33_412 VPWR VGND sg13g2_decap_8
XFILLER_33_423 VPWR VGND sg13g2_fill_2
XFILLER_33_445 VPWR VGND sg13g2_fill_1
XFILLER_34_946 VPWR VGND sg13g2_decap_8
X_509_ net66 VGND VPWR _131_ DP_4.matrix\[49\] clknet_5_14__leaf_clk sg13g2_dfrbpq_1
XFILLER_42_990 VPWR VGND sg13g2_decap_8
XFILLER_14_681 VPWR VGND sg13g2_decap_8
XFILLER_6_880 VPWR VGND sg13g2_decap_8
XFILLER_47_0 VPWR VGND sg13g2_decap_8
XFILLER_3_81 VPWR VGND sg13g2_decap_8
XFILLER_29_707 VPWR VGND sg13g2_decap_8
XFILLER_25_902 VPWR VGND sg13g2_decap_8
XFILLER_37_784 VPWR VGND sg13g2_decap_8
XFILLER_24_467 VPWR VGND sg13g2_decap_8
XFILLER_25_979 VPWR VGND sg13g2_decap_8
XFILLER_11_128 VPWR VGND sg13g2_decap_8
XFILLER_20_684 VPWR VGND sg13g2_decap_8
XFILLER_22_57 VPWR VGND sg13g2_decap_8
XFILLER_4_839 VPWR VGND sg13g2_decap_8
XFILLER_47_21 VPWR VGND sg13g2_decap_8
XFILLER_47_548 VPWR VGND sg13g2_decap_8
XFILLER_43_721 VPWR VGND sg13g2_decap_8
XFILLER_15_412 VPWR VGND sg13g2_decap_8
XFILLER_16_957 VPWR VGND sg13g2_decap_8
XFILLER_43_798 VPWR VGND sg13g2_decap_8
XFILLER_7_611 VPWR VGND sg13g2_decap_8
XFILLER_11_662 VPWR VGND sg13g2_decap_8
X_225_ net136 net137 _040_ VPWR VGND sg13g2_and2_1
XFILLER_10_194 VPWR VGND sg13g2_decap_8
XFILLER_7_688 VPWR VGND sg13g2_decap_8
XFILLER_40_7 VPWR VGND sg13g2_decap_8
XFILLER_3_894 VPWR VGND sg13g2_decap_8
XFILLER_19_4 VPWR VGND sg13g2_decap_8
XFILLER_38_537 VPWR VGND sg13g2_decap_8
XFILLER_19_784 VPWR VGND sg13g2_decap_8
XFILLER_34_743 VPWR VGND sg13g2_decap_8
XFILLER_22_905 VPWR VGND sg13g2_decap_8
XFILLER_30_982 VPWR VGND sg13g2_decap_8
XFILLER_0_308 VPWR VGND sg13g2_decap_8
XFILLER_25_1000 VPWR VGND sg13g2_decap_8
XFILLER_29_504 VPWR VGND sg13g2_decap_8
XFILLER_44_507 VPWR VGND sg13g2_decap_8
XFILLER_17_57 VPWR VGND sg13g2_fill_1
XFILLER_37_581 VPWR VGND sg13g2_decap_8
XFILLER_25_776 VPWR VGND sg13g2_decap_8
XFILLER_12_404 VPWR VGND sg13g2_decap_8
XFILLER_12_437 VPWR VGND sg13g2_decap_8
XFILLER_13_949 VPWR VGND sg13g2_decap_8
XFILLER_24_264 VPWR VGND sg13g2_decap_8
XFILLER_40_768 VPWR VGND sg13g2_decap_8
XFILLER_21_960 VPWR VGND sg13g2_decap_8
XFILLER_3_102 VPWR VGND sg13g2_decap_8
XFILLER_4_636 VPWR VGND sg13g2_decap_8
XFILLER_3_157 VPWR VGND sg13g2_decap_4
Xclkbuf_5_8__f_clk clknet_4_4_0_clk clknet_5_8__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_0_875 VPWR VGND sg13g2_decap_8
XFILLER_48_835 VPWR VGND sg13g2_decap_8
Xhold8 mac2.products_ff\[129\] VPWR VGND net32 sg13g2_dlygate4sd3_1
XFILLER_16_754 VPWR VGND sg13g2_decap_8
XFILLER_43_595 VPWR VGND sg13g2_decap_8
XFILLER_15_275 VPWR VGND sg13g2_decap_8
XFILLER_15_286 VPWR VGND sg13g2_fill_2
XFILLER_30_234 VPWR VGND sg13g2_decap_8
XFILLER_31_757 VPWR VGND sg13g2_decap_8
XFILLER_12_971 VPWR VGND sg13g2_decap_8
XFILLER_8_964 VPWR VGND sg13g2_decap_8
XFILLER_11_470 VPWR VGND sg13g2_decap_4
XFILLER_7_485 VPWR VGND sg13g2_decap_8
XFILLER_3_691 VPWR VGND sg13g2_decap_8
XFILLER_39_802 VPWR VGND sg13g2_decap_8
XFILLER_39_879 VPWR VGND sg13g2_decap_8
XFILLER_26_518 VPWR VGND sg13g2_decap_8
XFILLER_38_356 VPWR VGND sg13g2_decap_8
XFILLER_19_581 VPWR VGND sg13g2_decap_8
XFILLER_22_702 VPWR VGND sg13g2_decap_8
XFILLER_34_540 VPWR VGND sg13g2_decap_8
XFILLER_22_779 VPWR VGND sg13g2_decap_8
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_44_304 VPWR VGND sg13g2_decap_4
XFILLER_17_529 VPWR VGND sg13g2_decap_8
XFILLER_28_67 VPWR VGND sg13g2_decap_8
X_490_ net66 VGND VPWR _112_ DP_3.matrix\[48\] clknet_5_14__leaf_clk sg13g2_dfrbpq_1
XFILLER_25_584 VPWR VGND sg13g2_fill_1
XFILLER_13_746 VPWR VGND sg13g2_decap_8
XFILLER_8_205 VPWR VGND sg13g2_decap_8
XFILLER_12_267 VPWR VGND sg13g2_decap_8
XFILLER_40_565 VPWR VGND sg13g2_decap_8
XFILLER_5_967 VPWR VGND sg13g2_decap_8
Xclkbuf_4_0_0_clk clknet_0_clk clknet_4_0_0_clk VPWR VGND sg13g2_buf_8
XFILLER_4_488 VPWR VGND sg13g2_decap_8
XFILLER_0_672 VPWR VGND sg13g2_decap_8
XFILLER_48_632 VPWR VGND sg13g2_decap_8
XFILLER_47_153 VPWR VGND sg13g2_decap_8
XFILLER_36_827 VPWR VGND sg13g2_decap_8
XFILLER_35_359 VPWR VGND sg13g2_decap_8
XFILLER_44_871 VPWR VGND sg13g2_decap_8
XFILLER_31_554 VPWR VGND sg13g2_decap_8
XFILLER_15_1021 VPWR VGND sg13g2_decap_8
XFILLER_8_761 VPWR VGND sg13g2_decap_8
XFILLER_7_293 VPWR VGND sg13g2_decap_8
XFILLER_22_1003 VPWR VGND sg13g2_decap_8
XFILLER_27_805 VPWR VGND sg13g2_decap_8
XFILLER_39_676 VPWR VGND sg13g2_decap_8
XFILLER_26_326 VPWR VGND sg13g2_decap_8
XFILLER_42_808 VPWR VGND sg13g2_decap_8
XFILLER_41_307 VPWR VGND sg13g2_decap_8
XFILLER_14_25 VPWR VGND sg13g2_decap_8
XFILLER_22_543 VPWR VGND sg13g2_decap_8
XFILLER_10_727 VPWR VGND sg13g2_decap_8
XFILLER_22_576 VPWR VGND sg13g2_decap_8
XFILLER_5_219 VPWR VGND sg13g2_decap_8
XFILLER_30_35 VPWR VGND sg13g2_decap_8
XFILLER_1_458 VPWR VGND sg13g2_decap_8
XFILLER_39_66 VPWR VGND sg13g2_decap_8
XFILLER_18_849 VPWR VGND sg13g2_decap_8
XFILLER_29_164 VPWR VGND sg13g2_decap_8
XFILLER_45_668 VPWR VGND sg13g2_decap_8
X_542_ net69 VGND VPWR net130 mac1.sum_lvl2_ff\[0\] clknet_5_19__leaf_clk sg13g2_dfrbpq_1
X_473_ net71 VGND VPWR _095_ DP_2.matrix\[49\] clknet_5_17__leaf_clk sg13g2_dfrbpq_1
XFILLER_32_318 VPWR VGND sg13g2_decap_8
XFILLER_25_392 VPWR VGND sg13g2_decap_4
XFILLER_13_565 VPWR VGND sg13g2_decap_8
XFILLER_40_351 VPWR VGND sg13g2_decap_8
XFILLER_40_362 VPWR VGND sg13g2_fill_1
XFILLER_41_863 VPWR VGND sg13g2_decap_8
XFILLER_9_536 VPWR VGND sg13g2_decap_8
XFILLER_5_764 VPWR VGND sg13g2_decap_8
XFILLER_45_1025 VPWR VGND sg13g2_decap_4
XFILLER_4_296 VPWR VGND sg13g2_decap_8
XFILLER_49_930 VPWR VGND sg13g2_decap_8
XFILLER_36_624 VPWR VGND sg13g2_decap_8
XFILLER_35_123 VPWR VGND sg13g2_decap_8
XFILLER_23_318 VPWR VGND sg13g2_decap_8
XFILLER_32_841 VPWR VGND sg13g2_decap_8
XFILLER_31_384 VPWR VGND sg13g2_decap_8
XFILLER_6_81 VPWR VGND sg13g2_decap_8
XFILLER_27_602 VPWR VGND sg13g2_decap_8
XFILLER_27_679 VPWR VGND sg13g2_decap_8
XFILLER_42_605 VPWR VGND sg13g2_decap_8
XFILLER_23_852 VPWR VGND sg13g2_decap_8
XFILLER_41_126 VPWR VGND sg13g2_decap_8
XFILLER_22_351 VPWR VGND sg13g2_decap_8
XFILLER_10_535 VPWR VGND sg13g2_decap_8
XFILLER_6_517 VPWR VGND sg13g2_decap_8
XFILLER_41_56 VPWR VGND sg13g2_decap_8
XFILLER_2_767 VPWR VGND sg13g2_decap_8
XFILLER_1_255 VPWR VGND sg13g2_decap_8
XFILLER_2_39 VPWR VGND sg13g2_decap_8
XFILLER_49_259 VPWR VGND sg13g2_decap_8
XFILLER_46_911 VPWR VGND sg13g2_decap_8
XFILLER_18_646 VPWR VGND sg13g2_decap_8
XFILLER_46_988 VPWR VGND sg13g2_decap_8
XFILLER_45_465 VPWR VGND sg13g2_decap_8
X_525_ net72 VGND VPWR net179 mac1.sum_lvl1_ff\[1\] clknet_5_22__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_156 VPWR VGND sg13g2_decap_8
XFILLER_17_178 VPWR VGND sg13g2_decap_8
XFILLER_14_863 VPWR VGND sg13g2_decap_8
X_456_ net77 VGND VPWR _078_ DP_1.matrix\[64\] clknet_5_25__leaf_clk sg13g2_dfrbpq_1
XFILLER_41_660 VPWR VGND sg13g2_decap_8
XFILLER_9_322 VPWR VGND sg13g2_decap_8
X_387_ net89 _081_ VPWR VGND sg13g2_buf_1
XFILLER_40_181 VPWR VGND sg13g2_decap_8
XFILLER_12_1013 VPWR VGND sg13g2_decap_8
XFILLER_5_561 VPWR VGND sg13g2_decap_8
XFILLER_48_281 VPWR VGND sg13g2_decap_8
XFILLER_37_966 VPWR VGND sg13g2_decap_8
XFILLER_23_104 VPWR VGND sg13g2_fill_1
XFILLER_24_649 VPWR VGND sg13g2_decap_8
XFILLER_36_498 VPWR VGND sg13g2_decap_8
XFILLER_23_148 VPWR VGND sg13g2_decap_8
XFILLER_20_866 VPWR VGND sg13g2_decap_8
XFILLER_11_15 VPWR VGND sg13g2_fill_2
XFILLER_46_218 VPWR VGND sg13g2_decap_4
XFILLER_28_911 VPWR VGND sg13g2_decap_8
XFILLER_43_903 VPWR VGND sg13g2_decap_8
XFILLER_39_281 VPWR VGND sg13g2_decap_8
XFILLER_28_988 VPWR VGND sg13g2_decap_8
XFILLER_36_56 VPWR VGND sg13g2_decap_8
XFILLER_14_137 VPWR VGND sg13g2_decap_8
X_310_ mac2.products_ff\[33\] mac2.products_ff\[49\] _181_ VPWR VGND sg13g2_xor2_1
XFILLER_35_1002 VPWR VGND sg13g2_decap_8
X_241_ _143_ mac1.total_sum\[1\] mac2.total_sum\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_10_332 VPWR VGND sg13g2_decap_8
XFILLER_11_844 VPWR VGND sg13g2_decap_8
XFILLER_10_376 VPWR VGND sg13g2_decap_8
XFILLER_6_358 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_2_564 VPWR VGND sg13g2_decap_8
XFILLER_38_719 VPWR VGND sg13g2_decap_8
XFILLER_18_421 VPWR VGND sg13g2_decap_8
XFILLER_19_966 VPWR VGND sg13g2_decap_8
XFILLER_46_785 VPWR VGND sg13g2_decap_8
XFILLER_34_925 VPWR VGND sg13g2_decap_8
XFILLER_18_498 VPWR VGND sg13g2_decap_8
X_508_ net66 VGND VPWR _130_ DP_4.matrix\[48\] clknet_5_12__leaf_clk sg13g2_dfrbpq_1
XFILLER_14_660 VPWR VGND sg13g2_decap_8
X_439_ net44 _133_ VPWR VGND sg13g2_buf_1
XFILLER_9_152 VPWR VGND sg13g2_decap_4
XFILLER_9_174 VPWR VGND sg13g2_decap_4
XFILLER_3_60 VPWR VGND sg13g2_decap_8
XFILLER_37_763 VPWR VGND sg13g2_decap_8
XFILLER_19_1008 VPWR VGND sg13g2_decap_8
XFILLER_25_958 VPWR VGND sg13g2_decap_8
XFILLER_24_446 VPWR VGND sg13g2_decap_8
XFILLER_20_663 VPWR VGND sg13g2_decap_8
XFILLER_4_818 VPWR VGND sg13g2_decap_8
XFILLER_3_306 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_47_527 VPWR VGND sg13g2_decap_8
XFILLER_43_700 VPWR VGND sg13g2_decap_8
XFILLER_28_785 VPWR VGND sg13g2_decap_8
XFILLER_16_936 VPWR VGND sg13g2_decap_8
XFILLER_43_777 VPWR VGND sg13g2_decap_8
XFILLER_42_254 VPWR VGND sg13g2_decap_4
XFILLER_42_287 VPWR VGND sg13g2_decap_8
XFILLER_31_939 VPWR VGND sg13g2_decap_8
X_224_ net144 net138 _038_ VPWR VGND sg13g2_and2_1
XFILLER_11_641 VPWR VGND sg13g2_decap_8
XFILLER_7_667 VPWR VGND sg13g2_decap_8
XFILLER_6_166 VPWR VGND sg13g2_fill_1
XFILLER_12_80 VPWR VGND sg13g2_decap_8
XFILLER_3_873 VPWR VGND sg13g2_decap_8
XFILLER_33_7 VPWR VGND sg13g2_decap_8
XFILLER_38_516 VPWR VGND sg13g2_decap_8
XFILLER_19_763 VPWR VGND sg13g2_decap_8
XFILLER_46_582 VPWR VGND sg13g2_decap_8
XFILLER_18_284 VPWR VGND sg13g2_decap_8
XFILLER_34_722 VPWR VGND sg13g2_decap_8
XFILLER_21_405 VPWR VGND sg13g2_decap_8
XFILLER_34_799 VPWR VGND sg13g2_decap_8
XFILLER_30_961 VPWR VGND sg13g2_decap_8
XFILLER_17_14 VPWR VGND sg13g2_decap_8
XFILLER_37_560 VPWR VGND sg13g2_decap_8
XFILLER_24_243 VPWR VGND sg13g2_decap_8
XFILLER_25_755 VPWR VGND sg13g2_decap_8
XFILLER_13_928 VPWR VGND sg13g2_decap_8
XFILLER_33_46 VPWR VGND sg13g2_decap_8
XFILLER_40_747 VPWR VGND sg13g2_decap_8
XFILLER_32_1016 VPWR VGND sg13g2_decap_8
XFILLER_32_1027 VPWR VGND sg13g2_fill_2
XFILLER_4_615 VPWR VGND sg13g2_decap_8
XFILLER_0_854 VPWR VGND sg13g2_decap_8
XFILLER_48_814 VPWR VGND sg13g2_decap_8
Xhold9 mac2.sum_lvl2_ff\[9\] VPWR VGND net33 sg13g2_dlygate4sd3_1
XFILLER_35_519 VPWR VGND sg13g2_decap_8
XFILLER_16_733 VPWR VGND sg13g2_decap_8
XFILLER_28_582 VPWR VGND sg13g2_decap_8
XFILLER_43_574 VPWR VGND sg13g2_decap_8
XFILLER_15_254 VPWR VGND sg13g2_decap_8
XFILLER_31_736 VPWR VGND sg13g2_decap_8
XFILLER_12_950 VPWR VGND sg13g2_decap_8
XFILLER_8_943 VPWR VGND sg13g2_decap_8
XFILLER_7_475 VPWR VGND sg13g2_fill_2
XFILLER_7_464 VPWR VGND sg13g2_decap_8
XFILLER_3_670 VPWR VGND sg13g2_decap_8
XFILLER_38_335 VPWR VGND sg13g2_decap_8
XFILLER_39_858 VPWR VGND sg13g2_decap_8
XFILLER_19_560 VPWR VGND sg13g2_decap_8
XFILLER_47_891 VPWR VGND sg13g2_decap_8
XFILLER_10_909 VPWR VGND sg13g2_decap_8
XFILLER_21_246 VPWR VGND sg13g2_decap_8
XFILLER_22_758 VPWR VGND sg13g2_decap_8
XFILLER_34_596 VPWR VGND sg13g2_decap_8
XFILLER_29_324 VPWR VGND sg13g2_decap_8
XFILLER_29_368 VPWR VGND sg13g2_decap_8
XFILLER_38_880 VPWR VGND sg13g2_decap_8
XFILLER_13_725 VPWR VGND sg13g2_decap_8
XFILLER_25_563 VPWR VGND sg13g2_decap_8
XFILLER_44_89 VPWR VGND sg13g2_decap_8
XFILLER_40_544 VPWR VGND sg13g2_decap_8
XFILLER_12_246 VPWR VGND sg13g2_decap_8
XFILLER_5_946 VPWR VGND sg13g2_decap_8
XFILLER_4_467 VPWR VGND sg13g2_decap_8
XFILLER_48_611 VPWR VGND sg13g2_decap_8
XFILLER_0_651 VPWR VGND sg13g2_decap_8
XFILLER_48_688 VPWR VGND sg13g2_decap_8
XFILLER_47_132 VPWR VGND sg13g2_decap_8
XFILLER_36_806 VPWR VGND sg13g2_decap_8
XFILLER_35_316 VPWR VGND sg13g2_decap_8
XFILLER_44_850 VPWR VGND sg13g2_decap_8
XFILLER_18_90 VPWR VGND sg13g2_decap_8
XFILLER_31_533 VPWR VGND sg13g2_decap_8
XFILLER_15_1000 VPWR VGND sg13g2_decap_8
XFILLER_8_740 VPWR VGND sg13g2_decap_8
XFILLER_7_272 VPWR VGND sg13g2_decap_8
XFILLER_38_132 VPWR VGND sg13g2_decap_8
XFILLER_39_655 VPWR VGND sg13g2_decap_8
XFILLER_26_305 VPWR VGND sg13g2_decap_8
XFILLER_19_390 VPWR VGND sg13g2_decap_4
XFILLER_22_500 VPWR VGND sg13g2_fill_2
XFILLER_35_883 VPWR VGND sg13g2_decap_8
XFILLER_34_382 VPWR VGND sg13g2_decap_8
XFILLER_10_706 VPWR VGND sg13g2_decap_8
XFILLER_30_14 VPWR VGND sg13g2_decap_8
XFILLER_2_949 VPWR VGND sg13g2_decap_8
XFILLER_1_437 VPWR VGND sg13g2_decap_8
XFILLER_49_419 VPWR VGND sg13g2_decap_8
XFILLER_29_143 VPWR VGND sg13g2_decap_8
X_541_ net69 VGND VPWR _055_ mac1.products_ff\[33\] clknet_5_17__leaf_clk sg13g2_dfrbpq_1
XFILLER_18_828 VPWR VGND sg13g2_decap_8
XFILLER_45_647 VPWR VGND sg13g2_decap_8
XFILLER_44_124 VPWR VGND sg13g2_decap_8
XFILLER_17_349 VPWR VGND sg13g2_decap_8
X_472_ net71 VGND VPWR _094_ DP_2.matrix\[48\] clknet_5_20__leaf_clk sg13g2_dfrbpq_1
XFILLER_13_544 VPWR VGND sg13g2_decap_8
XFILLER_25_371 VPWR VGND sg13g2_decap_8
XFILLER_26_894 VPWR VGND sg13g2_decap_8
XFILLER_41_842 VPWR VGND sg13g2_decap_8
XFILLER_9_515 VPWR VGND sg13g2_decap_8
XFILLER_5_743 VPWR VGND sg13g2_decap_8
XFILLER_4_275 VPWR VGND sg13g2_decap_8
XFILLER_45_1004 VPWR VGND sg13g2_decap_8
XFILLER_49_986 VPWR VGND sg13g2_decap_8
XFILLER_36_603 VPWR VGND sg13g2_decap_8
XFILLER_48_485 VPWR VGND sg13g2_decap_8
XFILLER_35_179 VPWR VGND sg13g2_decap_8
XFILLER_16_393 VPWR VGND sg13g2_fill_1
XFILLER_17_894 VPWR VGND sg13g2_decap_8
XFILLER_32_820 VPWR VGND sg13g2_decap_8
XFILLER_31_330 VPWR VGND sg13g2_decap_8
XFILLER_31_363 VPWR VGND sg13g2_decap_8
XFILLER_32_897 VPWR VGND sg13g2_decap_8
XFILLER_6_60 VPWR VGND sg13g2_decap_8
XFILLER_6_1020 VPWR VGND sg13g2_decap_8
XFILLER_39_452 VPWR VGND sg13g2_decap_8
XFILLER_39_485 VPWR VGND sg13g2_fill_1
XFILLER_26_124 VPWR VGND sg13g2_fill_2
XFILLER_27_658 VPWR VGND sg13g2_decap_8
XFILLER_25_25 VPWR VGND sg13g2_decap_8
XFILLER_23_831 VPWR VGND sg13g2_decap_8
XFILLER_35_680 VPWR VGND sg13g2_decap_8
XFILLER_22_330 VPWR VGND sg13g2_decap_8
XFILLER_10_514 VPWR VGND sg13g2_decap_8
XFILLER_41_35 VPWR VGND sg13g2_decap_8
XFILLER_9_4 VPWR VGND sg13g2_decap_8
XFILLER_2_746 VPWR VGND sg13g2_decap_8
XFILLER_1_234 VPWR VGND sg13g2_decap_8
XFILLER_49_238 VPWR VGND sg13g2_decap_8
XFILLER_2_18 VPWR VGND sg13g2_decap_8
XFILLER_18_625 VPWR VGND sg13g2_decap_8
XFILLER_46_967 VPWR VGND sg13g2_decap_8
XFILLER_45_444 VPWR VGND sg13g2_decap_8
XFILLER_17_135 VPWR VGND sg13g2_decap_8
X_524_ net73 VGND VPWR net127 mac1.sum_lvl1_ff\[0\] clknet_5_22__leaf_clk sg13g2_dfrbpq_1
X_455_ net71 VGND VPWR _077_ DP_1.matrix\[49\] clknet_5_21__leaf_clk sg13g2_dfrbpq_1
XFILLER_14_842 VPWR VGND sg13g2_decap_8
XFILLER_26_691 VPWR VGND sg13g2_decap_8
XFILLER_33_639 VPWR VGND sg13g2_decap_8
X_386_ net162 _080_ VPWR VGND sg13g2_buf_1
XFILLER_40_160 VPWR VGND sg13g2_decap_8
XFILLER_9_389 VPWR VGND sg13g2_decap_8
XFILLER_49_783 VPWR VGND sg13g2_decap_8
XFILLER_48_260 VPWR VGND sg13g2_decap_8
XFILLER_36_444 VPWR VGND sg13g2_decap_8
XFILLER_37_945 VPWR VGND sg13g2_decap_8
XFILLER_24_628 VPWR VGND sg13g2_decap_8
XFILLER_36_455 VPWR VGND sg13g2_fill_2
XFILLER_17_691 VPWR VGND sg13g2_decap_8
XFILLER_23_127 VPWR VGND sg13g2_decap_8
XFILLER_32_694 VPWR VGND sg13g2_decap_8
XFILLER_20_845 VPWR VGND sg13g2_decap_8
XFILLER_47_709 VPWR VGND sg13g2_decap_8
XFILLER_39_271 VPWR VGND sg13g2_fill_1
XFILLER_27_422 VPWR VGND sg13g2_decap_8
XFILLER_28_967 VPWR VGND sg13g2_decap_8
XFILLER_36_35 VPWR VGND sg13g2_decap_8
XFILLER_27_455 VPWR VGND sg13g2_fill_1
XFILLER_43_959 VPWR VGND sg13g2_decap_8
XFILLER_42_436 VPWR VGND sg13g2_decap_8
XFILLER_14_116 VPWR VGND sg13g2_decap_8
X_240_ _142_ mac1.total_sum\[0\] mac2.total_sum\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_11_823 VPWR VGND sg13g2_decap_8
XFILLER_10_322 VPWR VGND sg13g2_fill_1
XFILLER_10_355 VPWR VGND sg13g2_decap_8
XFILLER_7_849 VPWR VGND sg13g2_decap_8
XFILLER_2_532 VPWR VGND sg13g2_fill_1
XFILLER_42_1018 VPWR VGND sg13g2_decap_8
XFILLER_18_400 VPWR VGND sg13g2_decap_8
XFILLER_19_945 VPWR VGND sg13g2_decap_8
XFILLER_46_764 VPWR VGND sg13g2_decap_8
XFILLER_45_241 VPWR VGND sg13g2_decap_8
XFILLER_18_477 VPWR VGND sg13g2_decap_8
XFILLER_34_904 VPWR VGND sg13g2_decap_8
XFILLER_45_296 VPWR VGND sg13g2_decap_8
XFILLER_33_436 VPWR VGND sg13g2_decap_8
X_507_ net76 VGND VPWR _129_ DP_4.matrix\[33\] clknet_5_14__leaf_clk sg13g2_dfrbpq_1
XFILLER_20_119 VPWR VGND sg13g2_decap_8
X_438_ net134 _132_ VPWR VGND sg13g2_buf_1
X_369_ _218_ net139 net99 VPWR VGND sg13g2_nand2_1
XFILLER_9_131 VPWR VGND sg13g2_decap_8
XFILLER_49_580 VPWR VGND sg13g2_decap_8
XFILLER_37_742 VPWR VGND sg13g2_decap_8
XFILLER_24_425 VPWR VGND sg13g2_decap_8
XFILLER_25_937 VPWR VGND sg13g2_decap_8
XFILLER_36_285 VPWR VGND sg13g2_decap_8
XFILLER_40_929 VPWR VGND sg13g2_decap_8
XFILLER_20_642 VPWR VGND sg13g2_decap_8
XFILLER_22_15 VPWR VGND sg13g2_fill_1
XFILLER_32_491 VPWR VGND sg13g2_decap_8
XFILLER_47_506 VPWR VGND sg13g2_decap_8
XFILLER_47_89 VPWR VGND sg13g2_fill_2
XFILLER_47_78 VPWR VGND sg13g2_decap_8
XFILLER_47_56 VPWR VGND sg13g2_decap_4
XFILLER_16_915 VPWR VGND sg13g2_decap_8
XFILLER_28_764 VPWR VGND sg13g2_decap_8
XFILLER_43_756 VPWR VGND sg13g2_decap_8
XFILLER_15_469 VPWR VGND sg13g2_decap_8
XFILLER_31_918 VPWR VGND sg13g2_decap_8
XFILLER_24_992 VPWR VGND sg13g2_decap_8
XFILLER_8_39 VPWR VGND sg13g2_decap_8
X_223_ net124 net142 _036_ VPWR VGND sg13g2_and2_1
XFILLER_10_163 VPWR VGND sg13g2_decap_4
XFILLER_7_646 VPWR VGND sg13g2_decap_8
XFILLER_11_697 VPWR VGND sg13g2_decap_8
XFILLER_6_145 VPWR VGND sg13g2_decap_8
XFILLER_3_852 VPWR VGND sg13g2_decap_8
XFILLER_2_384 VPWR VGND sg13g2_decap_4
XFILLER_19_742 VPWR VGND sg13g2_decap_8
XFILLER_46_561 VPWR VGND sg13g2_decap_8
XFILLER_34_701 VPWR VGND sg13g2_decap_8
XFILLER_18_263 VPWR VGND sg13g2_decap_8
XFILLER_34_778 VPWR VGND sg13g2_decap_8
XFILLER_33_266 VPWR VGND sg13g2_decap_8
XFILLER_30_940 VPWR VGND sg13g2_decap_8
XFILLER_33_299 VPWR VGND sg13g2_decap_8
XFILLER_29_539 VPWR VGND sg13g2_decap_8
XFILLER_25_734 VPWR VGND sg13g2_decap_8
XFILLER_13_907 VPWR VGND sg13g2_decap_8
XFILLER_33_14 VPWR VGND sg13g2_decap_4
XFILLER_40_726 VPWR VGND sg13g2_decap_8
XFILLER_20_483 VPWR VGND sg13g2_decap_8
XFILLER_21_995 VPWR VGND sg13g2_decap_8
XFILLER_0_833 VPWR VGND sg13g2_decap_8
XFILLER_47_358 VPWR VGND sg13g2_decap_8
XFILLER_16_712 VPWR VGND sg13g2_decap_8
XFILLER_28_561 VPWR VGND sg13g2_decap_8
XFILLER_43_553 VPWR VGND sg13g2_decap_8
XFILLER_16_789 VPWR VGND sg13g2_decap_8
XFILLER_31_715 VPWR VGND sg13g2_decap_8
XFILLER_8_922 VPWR VGND sg13g2_decap_8
XFILLER_30_269 VPWR VGND sg13g2_decap_8
XFILLER_8_999 VPWR VGND sg13g2_decap_8
XFILLER_7_443 VPWR VGND sg13g2_decap_8
XFILLER_48_1024 VPWR VGND sg13g2_decap_4
XFILLER_24_4 VPWR VGND sg13g2_decap_8
XFILLER_38_314 VPWR VGND sg13g2_decap_8
XFILLER_39_837 VPWR VGND sg13g2_decap_8
XFILLER_47_870 VPWR VGND sg13g2_decap_8
XFILLER_0_1015 VPWR VGND sg13g2_decap_8
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_34_575 VPWR VGND sg13g2_decap_8
XFILLER_21_225 VPWR VGND sg13g2_decap_8
XFILLER_21_236 VPWR VGND sg13g2_fill_1
XFILLER_22_737 VPWR VGND sg13g2_decap_8
XFILLER_9_60 VPWR VGND sg13g2_fill_2
XFILLER_9_82 VPWR VGND sg13g2_decap_8
XFILLER_1_619 VPWR VGND sg13g2_decap_8
XFILLER_29_303 VPWR VGND sg13g2_decap_8
XFILLER_45_829 VPWR VGND sg13g2_decap_8
XFILLER_25_531 VPWR VGND sg13g2_decap_4
XFILLER_37_391 VPWR VGND sg13g2_decap_8
XFILLER_44_68 VPWR VGND sg13g2_decap_8
XFILLER_13_704 VPWR VGND sg13g2_decap_8
XFILLER_12_225 VPWR VGND sg13g2_decap_8
XFILLER_40_523 VPWR VGND sg13g2_decap_8
XFILLER_21_792 VPWR VGND sg13g2_decap_8
Xclkbuf_5_16__f_clk clknet_4_8_0_clk clknet_5_16__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_20_280 VPWR VGND sg13g2_decap_8
XFILLER_5_925 VPWR VGND sg13g2_decap_8
XFILLER_4_402 VPWR VGND sg13g2_decap_8
XFILLER_4_446 VPWR VGND sg13g2_decap_8
XFILLER_0_630 VPWR VGND sg13g2_decap_8
XFILLER_48_667 VPWR VGND sg13g2_decap_8
XFILLER_47_188 VPWR VGND sg13g2_fill_1
XFILLER_16_531 VPWR VGND sg13g2_decap_8
XFILLER_43_394 VPWR VGND sg13g2_decap_8
XFILLER_16_586 VPWR VGND sg13g2_decap_8
XFILLER_31_512 VPWR VGND sg13g2_decap_8
XFILLER_34_90 VPWR VGND sg13g2_decap_8
XFILLER_31_589 VPWR VGND sg13g2_decap_8
XFILLER_8_796 VPWR VGND sg13g2_decap_8
XFILLER_7_251 VPWR VGND sg13g2_decap_8
XFILLER_3_490 VPWR VGND sg13g2_decap_8
XFILLER_38_111 VPWR VGND sg13g2_decap_8
XFILLER_39_634 VPWR VGND sg13g2_decap_8
XFILLER_35_862 VPWR VGND sg13g2_decap_8
XFILLER_2_928 VPWR VGND sg13g2_decap_8
XFILLER_1_416 VPWR VGND sg13g2_decap_8
XFILLER_18_807 VPWR VGND sg13g2_decap_8
XFILLER_29_122 VPWR VGND sg13g2_decap_8
XFILLER_45_626 VPWR VGND sg13g2_decap_8
XFILLER_44_103 VPWR VGND sg13g2_decap_8
X_540_ net70 VGND VPWR _054_ mac1.products_ff\[32\] clknet_5_19__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_328 VPWR VGND sg13g2_decap_8
XFILLER_29_199 VPWR VGND sg13g2_decap_8
X_471_ net69 VGND VPWR _093_ DP_2.matrix\[33\] clknet_5_17__leaf_clk sg13g2_dfrbpq_1
XFILLER_25_350 VPWR VGND sg13g2_decap_8
XFILLER_26_873 VPWR VGND sg13g2_decap_8
XFILLER_40_320 VPWR VGND sg13g2_decap_8
XFILLER_41_821 VPWR VGND sg13g2_decap_8
XFILLER_41_898 VPWR VGND sg13g2_decap_8
XFILLER_5_722 VPWR VGND sg13g2_decap_8
XFILLER_5_799 VPWR VGND sg13g2_decap_8
XFILLER_20_81 VPWR VGND sg13g2_decap_8
XFILLER_1_983 VPWR VGND sg13g2_decap_8
XFILLER_49_965 VPWR VGND sg13g2_decap_8
XFILLER_48_464 VPWR VGND sg13g2_decap_8
Xhold90 DP_2.matrix\[96\] VPWR VGND net140 sg13g2_dlygate4sd3_1
XFILLER_36_659 VPWR VGND sg13g2_decap_8
XFILLER_17_873 VPWR VGND sg13g2_decap_8
XFILLER_35_158 VPWR VGND sg13g2_decap_8
XFILLER_16_372 VPWR VGND sg13g2_decap_8
XFILLER_32_876 VPWR VGND sg13g2_decap_8
XFILLER_8_593 VPWR VGND sg13g2_decap_8
XFILLER_39_431 VPWR VGND sg13g2_decap_8
XFILLER_27_637 VPWR VGND sg13g2_decap_8
XFILLER_39_497 VPWR VGND sg13g2_fill_2
XFILLER_26_169 VPWR VGND sg13g2_decap_8
XFILLER_23_810 VPWR VGND sg13g2_decap_8
XFILLER_25_59 VPWR VGND sg13g2_decap_8
XFILLER_22_386 VPWR VGND sg13g2_fill_2
XFILLER_23_887 VPWR VGND sg13g2_decap_8
XFILLER_41_14 VPWR VGND sg13g2_decap_8
XFILLER_22_397 VPWR VGND sg13g2_decap_8
XFILLER_2_725 VPWR VGND sg13g2_decap_8
XFILLER_1_213 VPWR VGND sg13g2_decap_8
XFILLER_49_217 VPWR VGND sg13g2_decap_8
XFILLER_46_946 VPWR VGND sg13g2_decap_8
XFILLER_45_423 VPWR VGND sg13g2_decap_8
X_523_ net77 VGND VPWR _051_ mac1.products_ff\[65\] clknet_5_28__leaf_clk sg13g2_dfrbpq_1
XFILLER_33_618 VPWR VGND sg13g2_decap_8
X_454_ net71 VGND VPWR _076_ DP_1.matrix\[48\] clknet_5_21__leaf_clk sg13g2_dfrbpq_1
XFILLER_14_821 VPWR VGND sg13g2_decap_8
XFILLER_26_670 VPWR VGND sg13g2_decap_8
XFILLER_13_331 VPWR VGND sg13g2_decap_8
XFILLER_32_139 VPWR VGND sg13g2_decap_8
XFILLER_14_898 VPWR VGND sg13g2_decap_8
XFILLER_15_81 VPWR VGND sg13g2_fill_1
X_385_ net101 _079_ VPWR VGND sg13g2_buf_1
XFILLER_41_695 VPWR VGND sg13g2_decap_8
XFILLER_9_368 VPWR VGND sg13g2_decap_8
XFILLER_31_91 VPWR VGND sg13g2_decap_8
XFILLER_5_596 VPWR VGND sg13g2_decap_8
Xoutput1 net1 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_1_780 VPWR VGND sg13g2_decap_8
XFILLER_49_762 VPWR VGND sg13g2_decap_8
XFILLER_48_250 VPWR VGND sg13g2_fill_1
XFILLER_37_924 VPWR VGND sg13g2_decap_8
XFILLER_36_423 VPWR VGND sg13g2_decap_8
XFILLER_24_607 VPWR VGND sg13g2_decap_8
XFILLER_45_990 VPWR VGND sg13g2_decap_8
XFILLER_17_670 VPWR VGND sg13g2_decap_8
XFILLER_20_824 VPWR VGND sg13g2_decap_8
XFILLER_31_150 VPWR VGND sg13g2_fill_2
XFILLER_32_673 VPWR VGND sg13g2_decap_8
XFILLER_31_194 VPWR VGND sg13g2_decap_8
XFILLER_9_891 VPWR VGND sg13g2_decap_8
XFILLER_28_946 VPWR VGND sg13g2_decap_8
XFILLER_36_14 VPWR VGND sg13g2_decap_8
XFILLER_43_938 VPWR VGND sg13g2_decap_8
XFILLER_42_415 VPWR VGND sg13g2_decap_8
XFILLER_15_629 VPWR VGND sg13g2_decap_8
XFILLER_11_802 VPWR VGND sg13g2_decap_8
XFILLER_23_684 VPWR VGND sg13g2_decap_8
XFILLER_7_828 VPWR VGND sg13g2_decap_8
XFILLER_11_879 VPWR VGND sg13g2_decap_8
XFILLER_2_599 VPWR VGND sg13g2_decap_8
XFILLER_19_924 VPWR VGND sg13g2_decap_8
XFILLER_37_209 VPWR VGND sg13g2_decap_8
XFILLER_46_743 VPWR VGND sg13g2_decap_8
XFILLER_18_456 VPWR VGND sg13g2_decap_8
X_506_ net76 VGND VPWR _128_ DP_4.matrix\[32\] clknet_5_15__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_275 VPWR VGND sg13g2_decap_8
XFILLER_26_91 VPWR VGND sg13g2_decap_8
XFILLER_33_459 VPWR VGND sg13g2_decap_8
X_437_ net90 _131_ VPWR VGND sg13g2_buf_1
XFILLER_9_110 VPWR VGND sg13g2_decap_8
XFILLER_14_695 VPWR VGND sg13g2_decap_8
X_368_ _217_ _216_ _065_ VPWR VGND sg13g2_xor2_1
XFILLER_41_492 VPWR VGND sg13g2_decap_8
X_299_ _026_ _174_ net199 VPWR VGND sg13g2_xnor2_1
XFILLER_6_894 VPWR VGND sg13g2_decap_8
XFILLER_3_95 VPWR VGND sg13g2_decap_8
XFILLER_3_1013 VPWR VGND sg13g2_decap_8
XFILLER_37_721 VPWR VGND sg13g2_decap_8
XFILLER_25_916 VPWR VGND sg13g2_decap_8
XFILLER_36_253 VPWR VGND sg13g2_decap_8
XFILLER_24_404 VPWR VGND sg13g2_decap_8
XFILLER_37_798 VPWR VGND sg13g2_decap_8
XFILLER_40_908 VPWR VGND sg13g2_decap_8
XFILLER_33_982 VPWR VGND sg13g2_decap_8
XFILLER_20_621 VPWR VGND sg13g2_decap_8
XFILLER_20_698 VPWR VGND sg13g2_decap_8
XFILLER_47_35 VPWR VGND sg13g2_decap_8
XFILLER_19_209 VPWR VGND sg13g2_decap_8
XFILLER_28_743 VPWR VGND sg13g2_decap_8
XFILLER_27_242 VPWR VGND sg13g2_decap_8
XFILLER_43_735 VPWR VGND sg13g2_decap_8
XFILLER_42_212 VPWR VGND sg13g2_decap_8
XFILLER_15_426 VPWR VGND sg13g2_fill_2
XFILLER_15_448 VPWR VGND sg13g2_decap_8
XFILLER_24_971 VPWR VGND sg13g2_decap_8
XFILLER_30_407 VPWR VGND sg13g2_fill_2
XFILLER_30_418 VPWR VGND sg13g2_fill_1
XFILLER_8_18 VPWR VGND sg13g2_decap_8
X_222_ net155 net125 _034_ VPWR VGND sg13g2_and2_1
XFILLER_10_142 VPWR VGND sg13g2_decap_8
XFILLER_7_625 VPWR VGND sg13g2_decap_8
XFILLER_11_676 VPWR VGND sg13g2_decap_8
XFILLER_3_831 VPWR VGND sg13g2_decap_8
XFILLER_2_363 VPWR VGND sg13g2_decap_8
XFILLER_19_721 VPWR VGND sg13g2_decap_8
XFILLER_46_540 VPWR VGND sg13g2_decap_8
XFILLER_18_242 VPWR VGND sg13g2_decap_8
XFILLER_19_798 VPWR VGND sg13g2_decap_8
XFILLER_33_245 VPWR VGND sg13g2_decap_8
XFILLER_34_757 VPWR VGND sg13g2_decap_8
XFILLER_18_1010 VPWR VGND sg13g2_decap_8
XFILLER_22_919 VPWR VGND sg13g2_decap_8
XFILLER_15_993 VPWR VGND sg13g2_decap_8
XFILLER_21_429 VPWR VGND sg13g2_decap_8
XFILLER_30_996 VPWR VGND sg13g2_decap_8
XFILLER_45_0 VPWR VGND sg13g2_decap_8
XFILLER_6_691 VPWR VGND sg13g2_decap_8
XFILLER_25_1014 VPWR VGND sg13g2_decap_8
XFILLER_29_518 VPWR VGND sg13g2_decap_8
XFILLER_25_713 VPWR VGND sg13g2_decap_8
XFILLER_37_595 VPWR VGND sg13g2_decap_8
XFILLER_12_418 VPWR VGND sg13g2_decap_4
XFILLER_24_278 VPWR VGND sg13g2_decap_8
XFILLER_40_705 VPWR VGND sg13g2_decap_8
XFILLER_21_974 VPWR VGND sg13g2_decap_8
XFILLER_20_462 VPWR VGND sg13g2_decap_8
XFILLER_0_812 VPWR VGND sg13g2_decap_8
XFILLER_47_304 VPWR VGND sg13g2_decap_8
XFILLER_0_889 VPWR VGND sg13g2_decap_8
XFILLER_48_849 VPWR VGND sg13g2_decap_8
XFILLER_47_337 VPWR VGND sg13g2_decap_8
XFILLER_47_326 VPWR VGND sg13g2_fill_2
XFILLER_28_540 VPWR VGND sg13g2_decap_8
XFILLER_43_532 VPWR VGND sg13g2_decap_8
XFILLER_16_768 VPWR VGND sg13g2_decap_8
XFILLER_8_901 VPWR VGND sg13g2_decap_8
XFILLER_30_248 VPWR VGND sg13g2_decap_8
XFILLER_7_422 VPWR VGND sg13g2_decap_8
XFILLER_12_985 VPWR VGND sg13g2_decap_8
XFILLER_8_978 VPWR VGND sg13g2_decap_8
XFILLER_7_499 VPWR VGND sg13g2_decap_8
XFILLER_48_1003 VPWR VGND sg13g2_decap_8
XFILLER_39_816 VPWR VGND sg13g2_decap_8
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_19_595 VPWR VGND sg13g2_decap_8
XFILLER_22_716 VPWR VGND sg13g2_decap_8
XFILLER_34_554 VPWR VGND sg13g2_decap_8
XFILLER_15_790 VPWR VGND sg13g2_decap_8
XFILLER_30_793 VPWR VGND sg13g2_decap_8
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_45_808 VPWR VGND sg13g2_decap_8
XFILLER_25_510 VPWR VGND sg13g2_decap_8
XFILLER_44_14 VPWR VGND sg13g2_decap_8
XFILLER_37_370 VPWR VGND sg13g2_decap_8
XFILLER_40_502 VPWR VGND sg13g2_decap_8
XFILLER_9_709 VPWR VGND sg13g2_decap_8
XFILLER_12_204 VPWR VGND sg13g2_decap_8
XFILLER_40_579 VPWR VGND sg13g2_decap_8
XFILLER_8_219 VPWR VGND sg13g2_decap_8
XFILLER_21_771 VPWR VGND sg13g2_decap_8
XFILLER_5_904 VPWR VGND sg13g2_decap_8
XFILLER_4_425 VPWR VGND sg13g2_decap_8
XFILLER_0_686 VPWR VGND sg13g2_decap_8
XFILLER_48_646 VPWR VGND sg13g2_decap_8
XFILLER_47_167 VPWR VGND sg13g2_decap_8
XFILLER_29_882 VPWR VGND sg13g2_decap_8
XFILLER_28_392 VPWR VGND sg13g2_decap_8
XFILLER_44_885 VPWR VGND sg13g2_decap_8
XFILLER_43_373 VPWR VGND sg13g2_decap_8
XFILLER_31_568 VPWR VGND sg13g2_decap_8
XFILLER_12_782 VPWR VGND sg13g2_decap_8
XFILLER_7_230 VPWR VGND sg13g2_decap_8
XFILLER_8_775 VPWR VGND sg13g2_decap_8
XFILLER_39_613 VPWR VGND sg13g2_decap_8
XFILLER_22_1017 VPWR VGND sg13g2_decap_8
XFILLER_22_1028 VPWR VGND sg13g2_fill_1
XFILLER_27_819 VPWR VGND sg13g2_decap_8
XFILLER_35_841 VPWR VGND sg13g2_decap_8
XFILLER_38_189 VPWR VGND sg13g2_decap_8
Xclkbuf_5_22__f_clk clknet_4_11_0_clk clknet_5_22__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_22_524 VPWR VGND sg13g2_fill_2
XFILLER_14_39 VPWR VGND sg13g2_decap_8
XFILLER_22_557 VPWR VGND sg13g2_decap_8
XFILLER_30_590 VPWR VGND sg13g2_decap_8
XFILLER_2_907 VPWR VGND sg13g2_decap_8
XFILLER_30_49 VPWR VGND sg13g2_decap_8
XFILLER_39_14 VPWR VGND sg13g2_decap_8
XFILLER_29_101 VPWR VGND sg13g2_decap_8
XFILLER_45_605 VPWR VGND sg13g2_decap_8
XFILLER_17_307 VPWR VGND sg13g2_decap_8
XFILLER_29_178 VPWR VGND sg13g2_decap_8
X_470_ net69 VGND VPWR _092_ DP_2.matrix\[32\] clknet_5_19__leaf_clk sg13g2_dfrbpq_1
XFILLER_26_852 VPWR VGND sg13g2_decap_8
XFILLER_38_1013 VPWR VGND sg13g2_decap_8
XFILLER_41_800 VPWR VGND sg13g2_decap_8
XFILLER_13_513 VPWR VGND sg13g2_decap_8
XFILLER_41_877 VPWR VGND sg13g2_decap_8
XFILLER_13_579 VPWR VGND sg13g2_decap_8
XFILLER_5_701 VPWR VGND sg13g2_decap_8
XFILLER_4_211 VPWR VGND sg13g2_decap_8
XFILLER_5_778 VPWR VGND sg13g2_decap_8
XFILLER_20_60 VPWR VGND sg13g2_decap_8
XFILLER_1_962 VPWR VGND sg13g2_decap_8
XFILLER_49_944 VPWR VGND sg13g2_decap_8
XFILLER_48_443 VPWR VGND sg13g2_decap_8
XFILLER_0_483 VPWR VGND sg13g2_decap_8
XFILLER_29_80 VPWR VGND sg13g2_decap_8
Xhold80 _008_ VPWR VGND net130 sg13g2_dlygate4sd3_1
Xhold91 DP_3.matrix\[64\] VPWR VGND net141 sg13g2_dlygate4sd3_1
XFILLER_35_137 VPWR VGND sg13g2_decap_8
XFILLER_36_638 VPWR VGND sg13g2_decap_8
XFILLER_16_351 VPWR VGND sg13g2_decap_8
XFILLER_17_852 VPWR VGND sg13g2_decap_8
XFILLER_44_682 VPWR VGND sg13g2_decap_8
X_599_ net60 VGND VPWR net197 mac2.sum_lvl3_ff\[1\] clknet_5_13__leaf_clk sg13g2_dfrbpq_2
XFILLER_43_192 VPWR VGND sg13g2_decap_8
XFILLER_32_855 VPWR VGND sg13g2_decap_8
XFILLER_31_398 VPWR VGND sg13g2_decap_8
XFILLER_27_616 VPWR VGND sg13g2_decap_8
XFILLER_42_619 VPWR VGND sg13g2_decap_8
XFILLER_23_866 VPWR VGND sg13g2_decap_8
XFILLER_22_365 VPWR VGND sg13g2_decap_8
XFILLER_10_549 VPWR VGND sg13g2_decap_8
XFILLER_2_704 VPWR VGND sg13g2_decap_8
XFILLER_1_269 VPWR VGND sg13g2_decap_8
XFILLER_46_925 VPWR VGND sg13g2_decap_8
XFILLER_45_402 VPWR VGND sg13g2_decap_8
XFILLER_18_605 VPWR VGND sg13g2_decap_4
XFILLER_45_479 VPWR VGND sg13g2_decap_8
X_522_ net77 VGND VPWR _050_ mac1.products_ff\[64\] clknet_5_28__leaf_clk sg13g2_dfrbpq_1
X_453_ net69 VGND VPWR _075_ DP_1.matrix\[33\] clknet_5_17__leaf_clk sg13g2_dfrbpq_1
XFILLER_14_800 VPWR VGND sg13g2_decap_8
XFILLER_13_310 VPWR VGND sg13g2_decap_4
XFILLER_25_181 VPWR VGND sg13g2_decap_8
XFILLER_13_354 VPWR VGND sg13g2_decap_8
XFILLER_13_365 VPWR VGND sg13g2_fill_1
XFILLER_14_877 VPWR VGND sg13g2_decap_8
XFILLER_15_60 VPWR VGND sg13g2_decap_8
X_384_ net131 _078_ VPWR VGND sg13g2_buf_1
XFILLER_41_674 VPWR VGND sg13g2_decap_8
XFILLER_9_336 VPWR VGND sg13g2_fill_2
XFILLER_40_195 VPWR VGND sg13g2_decap_8
XFILLER_12_1027 VPWR VGND sg13g2_fill_2
XFILLER_5_520 VPWR VGND sg13g2_decap_8
XFILLER_31_70 VPWR VGND sg13g2_decap_8
XFILLER_49_7 VPWR VGND sg13g2_decap_8
XFILLER_5_575 VPWR VGND sg13g2_decap_8
Xoutput2 net2 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_49_741 VPWR VGND sg13g2_decap_8
XFILLER_0_280 VPWR VGND sg13g2_decap_8
XFILLER_37_903 VPWR VGND sg13g2_decap_8
XFILLER_48_295 VPWR VGND sg13g2_decap_8
XFILLER_20_803 VPWR VGND sg13g2_decap_8
XFILLER_32_652 VPWR VGND sg13g2_decap_8
XFILLER_31_173 VPWR VGND sg13g2_decap_8
XFILLER_9_870 VPWR VGND sg13g2_decap_8
XFILLER_8_380 VPWR VGND sg13g2_decap_8
XFILLER_28_1023 VPWR VGND sg13g2_decap_4
XFILLER_28_925 VPWR VGND sg13g2_decap_8
XFILLER_39_295 VPWR VGND sg13g2_decap_8
XFILLER_43_917 VPWR VGND sg13g2_decap_8
XFILLER_15_608 VPWR VGND sg13g2_decap_8
XFILLER_42_449 VPWR VGND sg13g2_decap_4
XFILLER_23_663 VPWR VGND sg13g2_decap_8
XFILLER_35_1016 VPWR VGND sg13g2_decap_8
XFILLER_35_1027 VPWR VGND sg13g2_fill_2
XFILLER_10_313 VPWR VGND sg13g2_decap_8
XFILLER_7_807 VPWR VGND sg13g2_decap_8
XFILLER_11_858 VPWR VGND sg13g2_decap_8
XFILLER_22_162 VPWR VGND sg13g2_decap_4
XFILLER_22_184 VPWR VGND sg13g2_decap_8
XFILLER_6_306 VPWR VGND sg13g2_fill_2
XFILLER_2_523 VPWR VGND sg13g2_decap_8
XFILLER_2_578 VPWR VGND sg13g2_decap_8
XFILLER_19_903 VPWR VGND sg13g2_decap_8
XFILLER_46_722 VPWR VGND sg13g2_decap_8
XFILLER_18_435 VPWR VGND sg13g2_decap_8
XFILLER_45_254 VPWR VGND sg13g2_fill_2
X_505_ net79 VGND VPWR _127_ DP_4.matrix\[17\] clknet_5_27__leaf_clk sg13g2_dfrbpq_1
XFILLER_46_799 VPWR VGND sg13g2_decap_8
XFILLER_27_980 VPWR VGND sg13g2_decap_8
XFILLER_33_405 VPWR VGND sg13g2_decap_8
XFILLER_34_939 VPWR VGND sg13g2_decap_8
XFILLER_26_70 VPWR VGND sg13g2_decap_8
XFILLER_26_490 VPWR VGND sg13g2_decap_8
XFILLER_42_983 VPWR VGND sg13g2_decap_8
XFILLER_13_151 VPWR VGND sg13g2_fill_2
XFILLER_14_674 VPWR VGND sg13g2_decap_8
X_436_ net145 _130_ VPWR VGND sg13g2_buf_1
X_367_ _217_ net149 net90 VPWR VGND sg13g2_nand2_1
XFILLER_41_471 VPWR VGND sg13g2_decap_8
X_298_ net198 mac2.sum_lvl1_ff\[9\] _175_ VPWR VGND sg13g2_xor2_1
XFILLER_6_873 VPWR VGND sg13g2_decap_8
XFILLER_3_74 VPWR VGND sg13g2_decap_8
XFILLER_37_700 VPWR VGND sg13g2_decap_8
XFILLER_36_232 VPWR VGND sg13g2_decap_8
XFILLER_37_777 VPWR VGND sg13g2_decap_8
XFILLER_20_600 VPWR VGND sg13g2_decap_8
XFILLER_33_961 VPWR VGND sg13g2_decap_8
XFILLER_20_677 VPWR VGND sg13g2_decap_8
XFILLER_47_14 VPWR VGND sg13g2_decap_8
XFILLER_28_722 VPWR VGND sg13g2_decap_8
XFILLER_27_221 VPWR VGND sg13g2_decap_8
XFILLER_43_714 VPWR VGND sg13g2_decap_8
XFILLER_15_405 VPWR VGND sg13g2_decap_8
XFILLER_28_799 VPWR VGND sg13g2_decap_8
XFILLER_27_298 VPWR VGND sg13g2_decap_8
XFILLER_24_950 VPWR VGND sg13g2_decap_8
XFILLER_23_493 VPWR VGND sg13g2_decap_8
XFILLER_10_121 VPWR VGND sg13g2_decap_8
XFILLER_7_604 VPWR VGND sg13g2_decap_8
XFILLER_11_655 VPWR VGND sg13g2_decap_8
XFILLER_3_810 VPWR VGND sg13g2_decap_8
XFILLER_12_94 VPWR VGND sg13g2_fill_2
XFILLER_3_887 VPWR VGND sg13g2_decap_8
XFILLER_2_342 VPWR VGND sg13g2_decap_8
XFILLER_19_700 VPWR VGND sg13g2_decap_8
Xclkbuf_5_3__f_clk clknet_4_1_0_clk clknet_5_3__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_19_777 VPWR VGND sg13g2_decap_8
XFILLER_46_596 VPWR VGND sg13g2_decap_8
XFILLER_18_298 VPWR VGND sg13g2_decap_8
XFILLER_34_736 VPWR VGND sg13g2_decap_8
XFILLER_15_972 VPWR VGND sg13g2_decap_8
XFILLER_42_780 VPWR VGND sg13g2_decap_8
X_419_ net42 _113_ VPWR VGND sg13g2_buf_1
XFILLER_30_975 VPWR VGND sg13g2_decap_8
XFILLER_6_670 VPWR VGND sg13g2_decap_8
XFILLER_5_191 VPWR VGND sg13g2_decap_8
XFILLER_38_0 VPWR VGND sg13g2_decap_8
XFILLER_37_574 VPWR VGND sg13g2_decap_8
XFILLER_24_257 VPWR VGND sg13g2_decap_8
XFILLER_25_769 VPWR VGND sg13g2_decap_8
XFILLER_20_441 VPWR VGND sg13g2_decap_8
XFILLER_21_953 VPWR VGND sg13g2_decap_8
XFILLER_32_290 VPWR VGND sg13g2_fill_1
XFILLER_4_629 VPWR VGND sg13g2_decap_8
XFILLER_48_828 VPWR VGND sg13g2_decap_8
XFILLER_0_868 VPWR VGND sg13g2_decap_8
XFILLER_43_511 VPWR VGND sg13g2_decap_8
XFILLER_15_213 VPWR VGND sg13g2_fill_1
XFILLER_16_747 VPWR VGND sg13g2_decap_8
XFILLER_28_596 VPWR VGND sg13g2_decap_8
XFILLER_15_268 VPWR VGND sg13g2_decap_8
XFILLER_43_588 VPWR VGND sg13g2_decap_8
XFILLER_30_227 VPWR VGND sg13g2_decap_8
XFILLER_12_964 VPWR VGND sg13g2_decap_8
XFILLER_23_290 VPWR VGND sg13g2_decap_8
XFILLER_8_957 VPWR VGND sg13g2_decap_8
XFILLER_11_463 VPWR VGND sg13g2_decap_8
XFILLER_11_474 VPWR VGND sg13g2_fill_2
XFILLER_23_93 VPWR VGND sg13g2_decap_8
XFILLER_3_684 VPWR VGND sg13g2_decap_8
XFILLER_31_7 VPWR VGND sg13g2_decap_8
XFILLER_38_305 VPWR VGND sg13g2_fill_1
XFILLER_38_349 VPWR VGND sg13g2_decap_8
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_19_574 VPWR VGND sg13g2_decap_8
XFILLER_46_393 VPWR VGND sg13g2_decap_8
XFILLER_34_533 VPWR VGND sg13g2_decap_8
XFILLER_30_772 VPWR VGND sg13g2_decap_8
Xclkbuf_4_15_0_clk clknet_0_clk clknet_4_15_0_clk VPWR VGND sg13g2_buf_8
XFILLER_29_338 VPWR VGND sg13g2_decap_8
XFILLER_44_308 VPWR VGND sg13g2_fill_1
XFILLER_38_894 VPWR VGND sg13g2_decap_8
XFILLER_25_577 VPWR VGND sg13g2_decap_8
XFILLER_13_739 VPWR VGND sg13g2_decap_8
XFILLER_21_750 VPWR VGND sg13g2_decap_8
XFILLER_40_558 VPWR VGND sg13g2_decap_8
XFILLER_0_665 VPWR VGND sg13g2_decap_8
XFILLER_48_625 VPWR VGND sg13g2_decap_8
XFILLER_47_146 VPWR VGND sg13g2_decap_8
XFILLER_29_861 VPWR VGND sg13g2_decap_8
XFILLER_28_371 VPWR VGND sg13g2_decap_8
XFILLER_44_864 VPWR VGND sg13g2_decap_8
XFILLER_43_352 VPWR VGND sg13g2_decap_8
XFILLER_31_547 VPWR VGND sg13g2_decap_8
XFILLER_12_761 VPWR VGND sg13g2_decap_8
XFILLER_15_1014 VPWR VGND sg13g2_decap_8
XFILLER_8_754 VPWR VGND sg13g2_decap_8
XFILLER_11_293 VPWR VGND sg13g2_decap_8
XFILLER_7_286 VPWR VGND sg13g2_decap_8
XFILLER_4_993 VPWR VGND sg13g2_decap_8
XFILLER_38_102 VPWR VGND sg13g2_fill_1
XFILLER_39_669 VPWR VGND sg13g2_decap_8
XFILLER_26_319 VPWR VGND sg13g2_decap_8
XFILLER_35_820 VPWR VGND sg13g2_decap_8
XFILLER_46_190 VPWR VGND sg13g2_decap_4
XFILLER_14_18 VPWR VGND sg13g2_decap_8
XFILLER_35_897 VPWR VGND sg13g2_decap_8
XFILLER_34_396 VPWR VGND sg13g2_decap_8
XFILLER_30_28 VPWR VGND sg13g2_decap_8
XFILLER_39_59 VPWR VGND sg13g2_decap_8
XFILLER_29_157 VPWR VGND sg13g2_decap_8
XFILLER_44_138 VPWR VGND sg13g2_decap_4
XFILLER_26_831 VPWR VGND sg13g2_decap_8
XFILLER_38_691 VPWR VGND sg13g2_decap_8
XFILLER_25_385 VPWR VGND sg13g2_decap_8
XFILLER_13_558 VPWR VGND sg13g2_decap_8
XFILLER_41_856 VPWR VGND sg13g2_decap_8
XFILLER_9_529 VPWR VGND sg13g2_decap_8
XFILLER_5_757 VPWR VGND sg13g2_decap_8
XFILLER_4_289 VPWR VGND sg13g2_decap_8
XFILLER_45_1018 VPWR VGND sg13g2_decap_8
XFILLER_1_941 VPWR VGND sg13g2_decap_8
XFILLER_49_923 VPWR VGND sg13g2_decap_8
XFILLER_0_462 VPWR VGND sg13g2_decap_8
XFILLER_48_422 VPWR VGND sg13g2_decap_8
Xhold92 DP_3.matrix\[128\] VPWR VGND net142 sg13g2_dlygate4sd3_1
Xhold70 DP_2.matrix\[112\] VPWR VGND net120 sg13g2_dlygate4sd3_1
Xhold81 DP_1.matrix\[64\] VPWR VGND net131 sg13g2_dlygate4sd3_1
XFILLER_36_617 VPWR VGND sg13g2_decap_8
XFILLER_48_499 VPWR VGND sg13g2_decap_8
XFILLER_17_831 VPWR VGND sg13g2_decap_8
XFILLER_35_105 VPWR VGND sg13g2_fill_1
XFILLER_16_330 VPWR VGND sg13g2_decap_8
XFILLER_28_190 VPWR VGND sg13g2_decap_8
XFILLER_45_80 VPWR VGND sg13g2_decap_8
XFILLER_44_661 VPWR VGND sg13g2_decap_8
X_598_ net60 VGND VPWR net153 mac2.sum_lvl3_ff\[0\] clknet_5_7__leaf_clk sg13g2_dfrbpq_2
XFILLER_32_834 VPWR VGND sg13g2_decap_8
XFILLER_31_344 VPWR VGND sg13g2_fill_2
XFILLER_31_377 VPWR VGND sg13g2_decap_8
XFILLER_12_591 VPWR VGND sg13g2_decap_8
XFILLER_8_573 VPWR VGND sg13g2_decap_8
XFILLER_6_74 VPWR VGND sg13g2_decap_8
XFILLER_4_790 VPWR VGND sg13g2_decap_8
XFILLER_26_105 VPWR VGND sg13g2_decap_8
XFILLER_25_39 VPWR VGND sg13g2_fill_1
XFILLER_41_119 VPWR VGND sg13g2_decap_8
XFILLER_23_845 VPWR VGND sg13g2_decap_8
XFILLER_34_182 VPWR VGND sg13g2_decap_8
XFILLER_35_694 VPWR VGND sg13g2_decap_8
XFILLER_22_344 VPWR VGND sg13g2_decap_8
XFILLER_10_528 VPWR VGND sg13g2_decap_8
XFILLER_41_49 VPWR VGND sg13g2_decap_8
XFILLER_1_248 VPWR VGND sg13g2_decap_8
XFILLER_46_904 VPWR VGND sg13g2_decap_8
XFILLER_18_639 VPWR VGND sg13g2_decap_8
XFILLER_45_458 VPWR VGND sg13g2_decap_8
XFILLER_17_149 VPWR VGND sg13g2_decap_8
X_521_ net78 VGND VPWR _049_ mac1.products_ff\[81\] clknet_5_30__leaf_clk sg13g2_dfrbpq_1
X_452_ net69 VGND VPWR _074_ DP_1.matrix\[32\] clknet_5_17__leaf_clk sg13g2_dfrbpq_1
XFILLER_25_160 VPWR VGND sg13g2_decap_8
X_383_ net86 _077_ VPWR VGND sg13g2_buf_1
XFILLER_13_322 VPWR VGND sg13g2_decap_4
XFILLER_14_856 VPWR VGND sg13g2_decap_8
XFILLER_9_315 VPWR VGND sg13g2_decap_8
XFILLER_41_653 VPWR VGND sg13g2_decap_8
XFILLER_40_174 VPWR VGND sg13g2_decap_8
XFILLER_12_1006 VPWR VGND sg13g2_decap_8
Xoutput3 net3 uo_out[2] VPWR VGND sg13g2_buf_1
XFILLER_49_720 VPWR VGND sg13g2_decap_8
XFILLER_48_241 VPWR VGND sg13g2_decap_8
XFILLER_49_797 VPWR VGND sg13g2_decap_8
XFILLER_48_274 VPWR VGND sg13g2_decap_8
XFILLER_37_959 VPWR VGND sg13g2_decap_8
XFILLER_32_631 VPWR VGND sg13g2_decap_8
XFILLER_20_859 VPWR VGND sg13g2_decap_8
XFILLER_28_1002 VPWR VGND sg13g2_decap_8
XFILLER_28_904 VPWR VGND sg13g2_decap_8
XFILLER_39_230 VPWR VGND sg13g2_decap_8
XFILLER_27_436 VPWR VGND sg13g2_decap_4
XFILLER_36_49 VPWR VGND sg13g2_decap_8
XFILLER_36_981 VPWR VGND sg13g2_decap_8
XFILLER_23_642 VPWR VGND sg13g2_decap_8
XFILLER_35_491 VPWR VGND sg13g2_decap_8
XFILLER_22_152 VPWR VGND sg13g2_decap_4
XFILLER_11_837 VPWR VGND sg13g2_decap_8
XFILLER_10_369 VPWR VGND sg13g2_decap_8
XFILLER_46_701 VPWR VGND sg13g2_decap_8
XFILLER_18_414 VPWR VGND sg13g2_decap_8
XFILLER_19_959 VPWR VGND sg13g2_decap_8
XFILLER_46_778 VPWR VGND sg13g2_decap_8
XFILLER_34_918 VPWR VGND sg13g2_decap_8
X_504_ net79 VGND VPWR _126_ DP_4.matrix\[16\] clknet_5_26__leaf_clk sg13g2_dfrbpq_1
X_435_ net54 _129_ VPWR VGND sg13g2_buf_1
XFILLER_42_962 VPWR VGND sg13g2_decap_8
XFILLER_14_653 VPWR VGND sg13g2_decap_8
X_366_ _216_ net145 net42 VPWR VGND sg13g2_nand2_1
XFILLER_9_156 VPWR VGND sg13g2_fill_2
XFILLER_9_167 VPWR VGND sg13g2_decap_8
XFILLER_9_145 VPWR VGND sg13g2_decap_8
X_297_ _174_ net121 mac2.sum_lvl1_ff\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_42_81 VPWR VGND sg13g2_decap_4
XFILLER_9_178 VPWR VGND sg13g2_fill_2
XFILLER_10_881 VPWR VGND sg13g2_decap_8
XFILLER_6_852 VPWR VGND sg13g2_decap_8
XFILLER_5_351 VPWR VGND sg13g2_decap_8
XFILLER_5_395 VPWR VGND sg13g2_decap_8
XFILLER_3_53 VPWR VGND sg13g2_decap_8
XFILLER_49_594 VPWR VGND sg13g2_decap_8
XFILLER_36_211 VPWR VGND sg13g2_decap_8
XFILLER_37_756 VPWR VGND sg13g2_decap_8
XFILLER_24_439 VPWR VGND sg13g2_decap_8
XFILLER_33_940 VPWR VGND sg13g2_decap_8
XFILLER_20_656 VPWR VGND sg13g2_decap_8
XFILLER_41_1010 VPWR VGND sg13g2_decap_8
XFILLER_28_701 VPWR VGND sg13g2_decap_8
XFILLER_16_929 VPWR VGND sg13g2_decap_8
XFILLER_28_778 VPWR VGND sg13g2_decap_8
XFILLER_42_258 VPWR VGND sg13g2_fill_2
XFILLER_42_247 VPWR VGND sg13g2_decap_8
XFILLER_10_100 VPWR VGND sg13g2_decap_8
XFILLER_23_472 VPWR VGND sg13g2_decap_8
XFILLER_6_159 VPWR VGND sg13g2_decap_8
XFILLER_12_73 VPWR VGND sg13g2_decap_8
XFILLER_2_321 VPWR VGND sg13g2_decap_8
XFILLER_3_866 VPWR VGND sg13g2_decap_8
XFILLER_38_509 VPWR VGND sg13g2_decap_8
XFILLER_18_211 VPWR VGND sg13g2_decap_4
XFILLER_19_756 VPWR VGND sg13g2_decap_8
XFILLER_46_575 VPWR VGND sg13g2_decap_8
XFILLER_18_277 VPWR VGND sg13g2_decap_8
XFILLER_34_715 VPWR VGND sg13g2_decap_8
XFILLER_37_70 VPWR VGND sg13g2_decap_4
XFILLER_15_951 VPWR VGND sg13g2_decap_8
X_418_ net149 _112_ VPWR VGND sg13g2_buf_1
XFILLER_14_461 VPWR VGND sg13g2_decap_8
XFILLER_30_954 VPWR VGND sg13g2_decap_8
X_349_ _205_ _204_ _053_ VPWR VGND sg13g2_xor2_1
XFILLER_5_170 VPWR VGND sg13g2_decap_8
XFILLER_49_391 VPWR VGND sg13g2_decap_8
XFILLER_37_553 VPWR VGND sg13g2_decap_8
XFILLER_24_236 VPWR VGND sg13g2_decap_8
XFILLER_25_748 VPWR VGND sg13g2_decap_8
XFILLER_21_932 VPWR VGND sg13g2_decap_8
XFILLER_32_1009 VPWR VGND sg13g2_decap_8
XFILLER_20_497 VPWR VGND sg13g2_decap_8
XFILLER_4_608 VPWR VGND sg13g2_decap_8
XFILLER_0_847 VPWR VGND sg13g2_decap_8
XFILLER_48_807 VPWR VGND sg13g2_decap_8
XFILLER_28_575 VPWR VGND sg13g2_decap_8
XFILLER_16_726 VPWR VGND sg13g2_decap_8
XFILLER_43_567 VPWR VGND sg13g2_decap_8
XFILLER_15_247 VPWR VGND sg13g2_decap_8
XFILLER_31_729 VPWR VGND sg13g2_decap_8
XFILLER_11_442 VPWR VGND sg13g2_decap_8
XFILLER_12_943 VPWR VGND sg13g2_decap_8
XFILLER_8_936 VPWR VGND sg13g2_decap_8
XFILLER_23_72 VPWR VGND sg13g2_decap_8
XFILLER_7_457 VPWR VGND sg13g2_decap_8
XFILLER_3_663 VPWR VGND sg13g2_decap_8
XFILLER_2_173 VPWR VGND sg13g2_fill_2
XFILLER_38_328 VPWR VGND sg13g2_decap_8
XFILLER_47_884 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_19_553 VPWR VGND sg13g2_decap_8
XFILLER_34_512 VPWR VGND sg13g2_decap_8
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_34_589 VPWR VGND sg13g2_decap_8
XFILLER_9_96 VPWR VGND sg13g2_decap_8
XFILLER_30_751 VPWR VGND sg13g2_decap_8
XFILLER_9_1010 VPWR VGND sg13g2_decap_8
XFILLER_29_317 VPWR VGND sg13g2_decap_8
XFILLER_38_873 VPWR VGND sg13g2_decap_8
XFILLER_13_718 VPWR VGND sg13g2_decap_8
XFILLER_12_239 VPWR VGND sg13g2_decap_8
XFILLER_40_537 VPWR VGND sg13g2_decap_8
XFILLER_5_939 VPWR VGND sg13g2_decap_8
XFILLER_4_416 VPWR VGND sg13g2_decap_4
XFILLER_20_294 VPWR VGND sg13g2_decap_8
XFILLER_0_644 VPWR VGND sg13g2_decap_8
XFILLER_48_604 VPWR VGND sg13g2_decap_8
XFILLER_47_125 VPWR VGND sg13g2_decap_8
XFILLER_29_840 VPWR VGND sg13g2_decap_8
XFILLER_35_309 VPWR VGND sg13g2_decap_8
XFILLER_44_843 VPWR VGND sg13g2_decap_8
XFILLER_43_331 VPWR VGND sg13g2_decap_8
XFILLER_16_545 VPWR VGND sg13g2_decap_8
XFILLER_31_526 VPWR VGND sg13g2_decap_8
XFILLER_12_740 VPWR VGND sg13g2_decap_8
XFILLER_8_733 VPWR VGND sg13g2_decap_8
XFILLER_11_272 VPWR VGND sg13g2_decap_8
XFILLER_7_265 VPWR VGND sg13g2_decap_8
XFILLER_4_972 VPWR VGND sg13g2_decap_8
XFILLER_22_4 VPWR VGND sg13g2_decap_8
XFILLER_38_125 VPWR VGND sg13g2_decap_8
XFILLER_39_648 VPWR VGND sg13g2_decap_8
XFILLER_47_681 VPWR VGND sg13g2_decap_8
XFILLER_19_383 VPWR VGND sg13g2_decap_8
XFILLER_19_394 VPWR VGND sg13g2_fill_2
XFILLER_34_331 VPWR VGND sg13g2_decap_8
XFILLER_35_876 VPWR VGND sg13g2_decap_8
XFILLER_34_375 VPWR VGND sg13g2_decap_8
XFILLER_22_537 VPWR VGND sg13g2_fill_1
XFILLER_29_136 VPWR VGND sg13g2_decap_8
XFILLER_44_117 VPWR VGND sg13g2_decap_8
XFILLER_26_810 VPWR VGND sg13g2_decap_8
XFILLER_38_670 VPWR VGND sg13g2_decap_8
XFILLER_25_364 VPWR VGND sg13g2_decap_8
XFILLER_26_887 VPWR VGND sg13g2_decap_8
XFILLER_41_835 VPWR VGND sg13g2_decap_8
XFILLER_9_508 VPWR VGND sg13g2_decap_8
XFILLER_40_334 VPWR VGND sg13g2_decap_4
XFILLER_21_570 VPWR VGND sg13g2_decap_8
XFILLER_21_581 VPWR VGND sg13g2_fill_2
XFILLER_5_736 VPWR VGND sg13g2_decap_8
XFILLER_4_268 VPWR VGND sg13g2_decap_8
XFILLER_1_920 VPWR VGND sg13g2_decap_8
XFILLER_20_95 VPWR VGND sg13g2_decap_4
XFILLER_49_902 VPWR VGND sg13g2_decap_8
XFILLER_48_401 VPWR VGND sg13g2_decap_8
XFILLER_0_441 VPWR VGND sg13g2_decap_8
XFILLER_1_997 VPWR VGND sg13g2_decap_8
XFILLER_49_979 VPWR VGND sg13g2_decap_8
XFILLER_48_478 VPWR VGND sg13g2_decap_8
Xhold82 DP_2.matrix\[48\] VPWR VGND net132 sg13g2_dlygate4sd3_1
Xhold60 _002_ VPWR VGND net110 sg13g2_dlygate4sd3_1
Xhold71 mac2.sum_lvl1_ff\[8\] VPWR VGND net121 sg13g2_dlygate4sd3_1
Xhold93 DP_4.matrix\[0\] VPWR VGND net143 sg13g2_dlygate4sd3_1
XFILLER_17_810 VPWR VGND sg13g2_decap_8
XFILLER_44_640 VPWR VGND sg13g2_decap_8
X_597_ net56 VGND VPWR net172 mac2.total_sum\[2\] clknet_5_18__leaf_clk sg13g2_dfrbpq_1
XFILLER_17_887 VPWR VGND sg13g2_decap_8
XFILLER_32_813 VPWR VGND sg13g2_decap_8
XFILLER_16_386 VPWR VGND sg13g2_decap_8
XFILLER_31_323 VPWR VGND sg13g2_decap_8
Xclkbuf_4_14_0_clk clknet_0_clk clknet_4_14_0_clk VPWR VGND sg13g2_buf_8
XFILLER_8_552 VPWR VGND sg13g2_decap_8
XFILLER_6_1013 VPWR VGND sg13g2_decap_8
XFILLER_39_445 VPWR VGND sg13g2_decap_8
XFILLER_19_191 VPWR VGND sg13g2_decap_8
XFILLER_25_18 VPWR VGND sg13g2_decap_8
XFILLER_23_824 VPWR VGND sg13g2_decap_8
XFILLER_34_161 VPWR VGND sg13g2_decap_8
XFILLER_35_673 VPWR VGND sg13g2_decap_8
XFILLER_22_323 VPWR VGND sg13g2_decap_8
XFILLER_10_507 VPWR VGND sg13g2_decap_8
XFILLER_31_890 VPWR VGND sg13g2_decap_8
XFILLER_41_28 VPWR VGND sg13g2_decap_8
XFILLER_2_739 VPWR VGND sg13g2_decap_8
XFILLER_1_227 VPWR VGND sg13g2_decap_8
XFILLER_18_618 VPWR VGND sg13g2_decap_8
X_520_ net73 VGND VPWR _048_ mac1.products_ff\[80\] clknet_5_28__leaf_clk sg13g2_dfrbpq_1
XFILLER_45_437 VPWR VGND sg13g2_decap_8
XFILLER_17_128 VPWR VGND sg13g2_decap_8
X_451_ net73 VGND VPWR _073_ DP_1.matrix\[17\] clknet_5_29__leaf_clk sg13g2_dfrbpq_1
XFILLER_26_684 VPWR VGND sg13g2_decap_8
XFILLER_32_109 VPWR VGND sg13g2_fill_2
X_382_ net164 _076_ VPWR VGND sg13g2_buf_1
XFILLER_14_835 VPWR VGND sg13g2_decap_8
XFILLER_41_632 VPWR VGND sg13g2_decap_8
XFILLER_40_153 VPWR VGND sg13g2_decap_8
XFILLER_15_95 VPWR VGND sg13g2_decap_8
Xoutput4 net4 uo_out[3] VPWR VGND sg13g2_buf_1
XFILLER_1_794 VPWR VGND sg13g2_decap_8
XFILLER_49_776 VPWR VGND sg13g2_decap_8
XFILLER_48_220 VPWR VGND sg13g2_decap_8
XFILLER_36_404 VPWR VGND sg13g2_decap_4
XFILLER_37_938 VPWR VGND sg13g2_decap_8
XFILLER_36_437 VPWR VGND sg13g2_decap_8
XFILLER_17_684 VPWR VGND sg13g2_decap_8
XFILLER_32_610 VPWR VGND sg13g2_decap_8
XFILLER_20_838 VPWR VGND sg13g2_decap_8
XFILLER_32_687 VPWR VGND sg13g2_decap_8
XFILLER_27_415 VPWR VGND sg13g2_decap_8
XFILLER_36_28 VPWR VGND sg13g2_decap_8
XFILLER_14_109 VPWR VGND sg13g2_decap_8
XFILLER_36_960 VPWR VGND sg13g2_decap_8
XFILLER_42_429 VPWR VGND sg13g2_decap_8
XFILLER_23_621 VPWR VGND sg13g2_decap_8
XFILLER_35_470 VPWR VGND sg13g2_decap_8
XFILLER_11_816 VPWR VGND sg13g2_decap_8
XFILLER_22_131 VPWR VGND sg13g2_decap_8
XFILLER_23_698 VPWR VGND sg13g2_decap_8
XFILLER_45_201 VPWR VGND sg13g2_decap_8
XFILLER_19_938 VPWR VGND sg13g2_decap_8
XFILLER_46_757 VPWR VGND sg13g2_decap_8
XFILLER_45_234 VPWR VGND sg13g2_decap_8
XFILLER_26_50 VPWR VGND sg13g2_fill_1
X_503_ net78 VGND VPWR _125_ DP_4.matrix\[1\] clknet_5_31__leaf_clk sg13g2_dfrbpq_1
X_434_ net139 _128_ VPWR VGND sg13g2_buf_1
XFILLER_45_289 VPWR VGND sg13g2_decap_8
XFILLER_42_941 VPWR VGND sg13g2_decap_8
XFILLER_33_429 VPWR VGND sg13g2_decap_8
XFILLER_9_124 VPWR VGND sg13g2_decap_8
XFILLER_13_153 VPWR VGND sg13g2_fill_1
X_365_ _215_ _214_ _063_ VPWR VGND sg13g2_xor2_1
XFILLER_42_60 VPWR VGND sg13g2_fill_1
XFILLER_13_197 VPWR VGND sg13g2_decap_8
X_296_ net105 mac2.sum_lvl1_ff\[24\] _027_ VPWR VGND sg13g2_xor2_1
XFILLER_10_860 VPWR VGND sg13g2_decap_8
XFILLER_6_831 VPWR VGND sg13g2_decap_8
XFILLER_5_330 VPWR VGND sg13g2_decap_8
XFILLER_3_32 VPWR VGND sg13g2_decap_8
XFILLER_1_591 VPWR VGND sg13g2_decap_8
XFILLER_49_573 VPWR VGND sg13g2_decap_8
XFILLER_3_1027 VPWR VGND sg13g2_fill_2
XFILLER_37_735 VPWR VGND sg13g2_decap_8
XFILLER_18_982 VPWR VGND sg13g2_decap_8
XFILLER_24_418 VPWR VGND sg13g2_decap_8
XFILLER_36_267 VPWR VGND sg13g2_fill_2
XFILLER_36_278 VPWR VGND sg13g2_decap_8
XFILLER_17_481 VPWR VGND sg13g2_decap_4
XFILLER_32_451 VPWR VGND sg13g2_decap_8
XFILLER_32_462 VPWR VGND sg13g2_fill_2
XFILLER_33_996 VPWR VGND sg13g2_decap_8
XFILLER_20_635 VPWR VGND sg13g2_decap_8
Xclkbuf_5_28__f_clk clknet_4_14_0_clk clknet_5_28__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_47_49 VPWR VGND sg13g2_fill_2
XFILLER_27_201 VPWR VGND sg13g2_decap_4
XFILLER_16_908 VPWR VGND sg13g2_decap_8
XFILLER_28_757 VPWR VGND sg13g2_decap_8
XFILLER_27_256 VPWR VGND sg13g2_decap_4
XFILLER_43_749 VPWR VGND sg13g2_decap_8
XFILLER_23_451 VPWR VGND sg13g2_decap_8
XFILLER_24_985 VPWR VGND sg13g2_decap_8
XFILLER_10_156 VPWR VGND sg13g2_decap_8
XFILLER_7_639 VPWR VGND sg13g2_decap_8
XFILLER_12_30 VPWR VGND sg13g2_decap_4
XFILLER_6_138 VPWR VGND sg13g2_decap_8
XFILLER_12_52 VPWR VGND sg13g2_decap_8
XFILLER_3_845 VPWR VGND sg13g2_decap_8
XFILLER_2_377 VPWR VGND sg13g2_decap_8
XFILLER_2_388 VPWR VGND sg13g2_fill_2
XFILLER_19_735 VPWR VGND sg13g2_decap_8
XFILLER_46_554 VPWR VGND sg13g2_decap_8
XFILLER_18_256 VPWR VGND sg13g2_decap_8
XFILLER_15_930 VPWR VGND sg13g2_decap_8
XFILLER_33_215 VPWR VGND sg13g2_fill_2
XFILLER_33_259 VPWR VGND sg13g2_decap_8
X_417_ net99 _111_ VPWR VGND sg13g2_buf_1
XFILLER_18_1024 VPWR VGND sg13g2_decap_4
XFILLER_30_933 VPWR VGND sg13g2_decap_8
X_348_ _205_ net164 net100 VPWR VGND sg13g2_nand2_1
XFILLER_14_495 VPWR VGND sg13g2_decap_4
X_279_ _164_ net201 net147 VPWR VGND sg13g2_nand2_1
XFILLER_25_1028 VPWR VGND sg13g2_fill_1
XFILLER_37_532 VPWR VGND sg13g2_decap_8
XFILLER_25_727 VPWR VGND sg13g2_decap_8
XFILLER_40_719 VPWR VGND sg13g2_decap_8
XFILLER_21_911 VPWR VGND sg13g2_decap_8
XFILLER_33_18 VPWR VGND sg13g2_fill_1
XFILLER_33_793 VPWR VGND sg13g2_decap_8
XFILLER_21_988 VPWR VGND sg13g2_decap_8
XFILLER_0_826 VPWR VGND sg13g2_decap_8
XFILLER_16_705 VPWR VGND sg13g2_decap_8
XFILLER_28_554 VPWR VGND sg13g2_decap_8
XFILLER_43_546 VPWR VGND sg13g2_decap_8
XFILLER_31_708 VPWR VGND sg13g2_decap_8
XFILLER_12_922 VPWR VGND sg13g2_decap_8
XFILLER_24_782 VPWR VGND sg13g2_decap_8
XFILLER_30_207 VPWR VGND sg13g2_fill_2
XFILLER_11_421 VPWR VGND sg13g2_decap_8
XFILLER_8_915 VPWR VGND sg13g2_decap_8
XFILLER_12_999 VPWR VGND sg13g2_decap_8
XFILLER_23_51 VPWR VGND sg13g2_decap_8
XFILLER_7_436 VPWR VGND sg13g2_decap_8
XFILLER_48_1017 VPWR VGND sg13g2_decap_8
XFILLER_48_1028 VPWR VGND sg13g2_fill_1
XFILLER_3_642 VPWR VGND sg13g2_decap_8
Xclkbuf_5_11__f_clk clknet_4_5_0_clk clknet_5_11__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_2_185 VPWR VGND sg13g2_fill_2
XFILLER_2_196 VPWR VGND sg13g2_decap_8
XFILLER_48_70 VPWR VGND sg13g2_decap_8
XFILLER_17_7 VPWR VGND sg13g2_decap_8
XFILLER_19_532 VPWR VGND sg13g2_decap_8
XFILLER_47_863 VPWR VGND sg13g2_decap_8
XFILLER_0_1008 VPWR VGND sg13g2_decap_8
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_34_568 VPWR VGND sg13g2_decap_8
XFILLER_21_218 VPWR VGND sg13g2_decap_8
XFILLER_30_730 VPWR VGND sg13g2_decap_8
XFILLER_9_75 VPWR VGND sg13g2_decap_8
XFILLER_43_0 VPWR VGND sg13g2_decap_8
XFILLER_38_852 VPWR VGND sg13g2_decap_8
XFILLER_25_524 VPWR VGND sg13g2_decap_8
XFILLER_37_384 VPWR VGND sg13g2_decap_8
XFILLER_44_28 VPWR VGND sg13g2_decap_4
XFILLER_25_535 VPWR VGND sg13g2_fill_1
XFILLER_40_516 VPWR VGND sg13g2_decap_8
XFILLER_33_590 VPWR VGND sg13g2_decap_8
XFILLER_20_273 VPWR VGND sg13g2_decap_8
XFILLER_21_785 VPWR VGND sg13g2_decap_8
XFILLER_5_918 VPWR VGND sg13g2_decap_8
XFILLER_4_439 VPWR VGND sg13g2_decap_8
XFILLER_0_623 VPWR VGND sg13g2_decap_8
XFILLER_18_62 VPWR VGND sg13g2_decap_8
XFILLER_44_822 VPWR VGND sg13g2_decap_8
XFILLER_43_310 VPWR VGND sg13g2_decap_8
XFILLER_16_524 VPWR VGND sg13g2_decap_8
XFILLER_29_896 VPWR VGND sg13g2_decap_8
XFILLER_44_899 VPWR VGND sg13g2_decap_8
XFILLER_16_579 VPWR VGND sg13g2_decap_4
XFILLER_31_505 VPWR VGND sg13g2_decap_8
XFILLER_43_387 VPWR VGND sg13g2_decap_8
XFILLER_8_712 VPWR VGND sg13g2_decap_8
XFILLER_34_83 VPWR VGND sg13g2_decap_8
XFILLER_11_251 VPWR VGND sg13g2_decap_8
XFILLER_12_796 VPWR VGND sg13g2_decap_8
XFILLER_8_789 VPWR VGND sg13g2_decap_8
XFILLER_7_244 VPWR VGND sg13g2_decap_8
XFILLER_4_951 VPWR VGND sg13g2_decap_8
XFILLER_3_461 VPWR VGND sg13g2_decap_8
XFILLER_3_483 VPWR VGND sg13g2_decap_8
XFILLER_39_627 VPWR VGND sg13g2_decap_8
XFILLER_15_4 VPWR VGND sg13g2_decap_8
XFILLER_19_340 VPWR VGND sg13g2_fill_2
XFILLER_47_660 VPWR VGND sg13g2_decap_8
XFILLER_19_362 VPWR VGND sg13g2_decap_8
XFILLER_34_310 VPWR VGND sg13g2_decap_8
XFILLER_35_855 VPWR VGND sg13g2_decap_8
XFILLER_1_409 VPWR VGND sg13g2_decap_8
XFILLER_29_115 VPWR VGND sg13g2_decap_8
XFILLER_45_619 VPWR VGND sg13g2_decap_8
XFILLER_25_343 VPWR VGND sg13g2_decap_8
XFILLER_26_866 VPWR VGND sg13g2_decap_8
XFILLER_37_181 VPWR VGND sg13g2_decap_8
XFILLER_38_1027 VPWR VGND sg13g2_fill_2
XFILLER_41_814 VPWR VGND sg13g2_decap_8
XFILLER_13_527 VPWR VGND sg13g2_decap_4
XFILLER_5_715 VPWR VGND sg13g2_decap_8
XFILLER_4_225 VPWR VGND sg13g2_decap_8
XFILLER_20_74 VPWR VGND sg13g2_decap_8
XFILLER_0_420 VPWR VGND sg13g2_decap_8
XFILLER_1_976 VPWR VGND sg13g2_decap_8
XFILLER_49_958 VPWR VGND sg13g2_decap_8
Xhold50 DP_2.matrix\[49\] VPWR VGND net100 sg13g2_dlygate4sd3_1
XFILLER_0_497 VPWR VGND sg13g2_decap_8
XFILLER_48_457 VPWR VGND sg13g2_decap_8
Xhold83 DP_4.matrix\[16\] VPWR VGND net133 sg13g2_dlygate4sd3_1
XFILLER_29_94 VPWR VGND sg13g2_decap_8
Xhold72 _025_ VPWR VGND net122 sg13g2_dlygate4sd3_1
Xhold61 mac2.products_ff\[64\] VPWR VGND net111 sg13g2_dlygate4sd3_1
Xhold94 DP_4.matrix\[80\] VPWR VGND net144 sg13g2_dlygate4sd3_1
XFILLER_17_866 VPWR VGND sg13g2_decap_8
XFILLER_29_693 VPWR VGND sg13g2_decap_8
X_596_ net56 VGND VPWR net208 mac2.total_sum\[1\] clknet_5_5__leaf_clk sg13g2_dfrbpq_1
XFILLER_16_365 VPWR VGND sg13g2_decap_8
XFILLER_44_696 VPWR VGND sg13g2_decap_8
XFILLER_31_313 VPWR VGND sg13g2_decap_4
XFILLER_32_869 VPWR VGND sg13g2_decap_8
XFILLER_40_880 VPWR VGND sg13g2_decap_8
Xclkbuf_5_9__f_clk clknet_4_4_0_clk clknet_5_9__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_39_402 VPWR VGND sg13g2_fill_2
XFILLER_23_803 VPWR VGND sg13g2_decap_8
XFILLER_34_140 VPWR VGND sg13g2_decap_8
XFILLER_35_652 VPWR VGND sg13g2_decap_8
XFILLER_22_302 VPWR VGND sg13g2_decap_8
XFILLER_22_379 VPWR VGND sg13g2_decap_8
XFILLER_2_718 VPWR VGND sg13g2_decap_8
XFILLER_1_206 VPWR VGND sg13g2_decap_8
XFILLER_46_939 VPWR VGND sg13g2_decap_8
XFILLER_45_416 VPWR VGND sg13g2_decap_8
XFILLER_39_991 VPWR VGND sg13g2_decap_8
XFILLER_14_814 VPWR VGND sg13g2_decap_8
X_450_ net73 VGND VPWR _072_ DP_1.matrix\[16\] clknet_5_29__leaf_clk sg13g2_dfrbpq_1
XFILLER_26_663 VPWR VGND sg13g2_decap_8
X_381_ net92 _075_ VPWR VGND sg13g2_buf_1
XFILLER_41_611 VPWR VGND sg13g2_decap_8
XFILLER_15_74 VPWR VGND sg13g2_decap_8
XFILLER_25_195 VPWR VGND sg13g2_decap_4
XFILLER_40_132 VPWR VGND sg13g2_decap_8
XFILLER_41_688 VPWR VGND sg13g2_decap_8
XFILLER_22_891 VPWR VGND sg13g2_decap_8
XFILLER_31_84 VPWR VGND sg13g2_decap_8
XFILLER_5_589 VPWR VGND sg13g2_decap_8
XFILLER_1_773 VPWR VGND sg13g2_decap_8
XFILLER_49_755 VPWR VGND sg13g2_decap_8
XFILLER_0_294 VPWR VGND sg13g2_decap_8
XFILLER_37_917 VPWR VGND sg13g2_decap_8
XFILLER_29_490 VPWR VGND sg13g2_decap_8
XFILLER_45_983 VPWR VGND sg13g2_decap_8
XFILLER_17_663 VPWR VGND sg13g2_decap_8
XFILLER_44_493 VPWR VGND sg13g2_decap_8
XFILLER_16_151 VPWR VGND sg13g2_decap_8
X_579_ net64 VGND VPWR _034_ mac2.products_ff\[112\] clknet_5_3__leaf_clk sg13g2_dfrbpq_1
XFILLER_31_143 VPWR VGND sg13g2_decap_8
XFILLER_32_666 VPWR VGND sg13g2_decap_8
XFILLER_20_817 VPWR VGND sg13g2_decap_8
XFILLER_31_187 VPWR VGND sg13g2_decap_8
XFILLER_9_884 VPWR VGND sg13g2_decap_8
XFILLER_8_394 VPWR VGND sg13g2_fill_2
XFILLER_28_939 VPWR VGND sg13g2_decap_8
XFILLER_42_408 VPWR VGND sg13g2_decap_8
XFILLER_23_600 VPWR VGND sg13g2_decap_8
XFILLER_22_110 VPWR VGND sg13g2_decap_8
XFILLER_23_677 VPWR VGND sg13g2_decap_8
XFILLER_22_198 VPWR VGND sg13g2_decap_8
Xclkbuf_4_13_0_clk clknet_0_clk clknet_4_13_0_clk VPWR VGND sg13g2_buf_8
XFILLER_19_917 VPWR VGND sg13g2_decap_8
XFILLER_46_736 VPWR VGND sg13g2_decap_8
XFILLER_18_449 VPWR VGND sg13g2_decap_8
XFILLER_45_268 VPWR VGND sg13g2_decap_8
XFILLER_33_419 VPWR VGND sg13g2_decap_4
X_502_ net78 VGND VPWR _124_ DP_4.matrix\[0\] clknet_5_31__leaf_clk sg13g2_dfrbpq_1
X_433_ net39 _127_ VPWR VGND sg13g2_buf_1
XFILLER_42_920 VPWR VGND sg13g2_decap_8
XFILLER_26_84 VPWR VGND sg13g2_decap_8
XFILLER_27_994 VPWR VGND sg13g2_decap_8
XFILLER_13_110 VPWR VGND sg13g2_decap_8
XFILLER_41_430 VPWR VGND sg13g2_decap_4
XFILLER_42_997 VPWR VGND sg13g2_decap_8
XFILLER_9_103 VPWR VGND sg13g2_decap_8
XFILLER_14_688 VPWR VGND sg13g2_decap_8
X_364_ _215_ net159 net88 VPWR VGND sg13g2_nand2_1
XFILLER_41_463 VPWR VGND sg13g2_decap_4
XFILLER_41_485 VPWR VGND sg13g2_decap_8
X_295_ _028_ _172_ _173_ VPWR VGND sg13g2_xnor2_1
XFILLER_6_810 VPWR VGND sg13g2_decap_8
XFILLER_6_887 VPWR VGND sg13g2_decap_8
XFILLER_47_7 VPWR VGND sg13g2_decap_8
XFILLER_3_11 VPWR VGND sg13g2_decap_8
XFILLER_1_570 VPWR VGND sg13g2_decap_8
XFILLER_3_88 VPWR VGND sg13g2_decap_8
XFILLER_49_552 VPWR VGND sg13g2_decap_8
XFILLER_3_1006 VPWR VGND sg13g2_decap_8
XFILLER_37_714 VPWR VGND sg13g2_decap_8
XFILLER_18_961 VPWR VGND sg13g2_decap_8
XFILLER_25_909 VPWR VGND sg13g2_decap_8
XFILLER_36_246 VPWR VGND sg13g2_decap_8
XFILLER_45_780 VPWR VGND sg13g2_decap_8
XFILLER_44_290 VPWR VGND sg13g2_decap_8
XFILLER_32_430 VPWR VGND sg13g2_decap_8
XFILLER_20_614 VPWR VGND sg13g2_decap_8
XFILLER_33_975 VPWR VGND sg13g2_decap_8
XFILLER_9_681 VPWR VGND sg13g2_decap_8
XFILLER_8_191 VPWR VGND sg13g2_decap_8
XFILLER_47_28 VPWR VGND sg13g2_decap_8
XFILLER_27_235 VPWR VGND sg13g2_decap_8
XFILLER_28_736 VPWR VGND sg13g2_decap_8
XFILLER_43_728 VPWR VGND sg13g2_decap_8
XFILLER_42_205 VPWR VGND sg13g2_decap_8
XFILLER_15_419 VPWR VGND sg13g2_fill_2
XFILLER_24_964 VPWR VGND sg13g2_decap_8
XFILLER_11_603 VPWR VGND sg13g2_decap_8
XFILLER_10_135 VPWR VGND sg13g2_decap_8
XFILLER_7_618 VPWR VGND sg13g2_decap_8
XFILLER_11_669 VPWR VGND sg13g2_decap_8
XFILLER_3_824 VPWR VGND sg13g2_decap_8
XFILLER_2_356 VPWR VGND sg13g2_decap_8
XFILLER_19_714 VPWR VGND sg13g2_decap_8
XFILLER_46_533 VPWR VGND sg13g2_decap_8
XFILLER_27_791 VPWR VGND sg13g2_decap_8
XFILLER_18_1003 VPWR VGND sg13g2_decap_8
X_416_ net163 _110_ VPWR VGND sg13g2_buf_1
XFILLER_15_986 VPWR VGND sg13g2_decap_8
XFILLER_30_912 VPWR VGND sg13g2_decap_8
XFILLER_42_794 VPWR VGND sg13g2_decap_8
X_347_ _204_ net86 net132 VPWR VGND sg13g2_nand2_1
XFILLER_41_293 VPWR VGND sg13g2_decap_8
XFILLER_30_989 VPWR VGND sg13g2_decap_8
X_278_ net109 mac1.products_ff\[32\] _002_ VPWR VGND sg13g2_xor2_1
XFILLER_6_684 VPWR VGND sg13g2_decap_8
XFILLER_25_1007 VPWR VGND sg13g2_decap_8
XFILLER_49_371 VPWR VGND sg13g2_decap_4
XFILLER_37_511 VPWR VGND sg13g2_decap_8
XFILLER_25_706 VPWR VGND sg13g2_decap_8
XFILLER_37_588 VPWR VGND sg13g2_decap_8
XFILLER_33_772 VPWR VGND sg13g2_decap_8
XFILLER_20_455 VPWR VGND sg13g2_decap_8
XFILLER_21_967 VPWR VGND sg13g2_decap_8
XFILLER_3_109 VPWR VGND sg13g2_decap_8
XFILLER_0_805 VPWR VGND sg13g2_decap_8
XFILLER_28_533 VPWR VGND sg13g2_decap_8
XFILLER_43_525 VPWR VGND sg13g2_decap_8
XFILLER_15_227 VPWR VGND sg13g2_fill_2
XFILLER_12_901 VPWR VGND sg13g2_decap_8
XFILLER_24_761 VPWR VGND sg13g2_decap_8
XFILLER_23_260 VPWR VGND sg13g2_decap_8
XFILLER_7_415 VPWR VGND sg13g2_fill_2
XFILLER_12_978 VPWR VGND sg13g2_decap_8
XFILLER_3_621 VPWR VGND sg13g2_decap_8
XFILLER_2_120 VPWR VGND sg13g2_fill_1
XFILLER_3_698 VPWR VGND sg13g2_decap_8
XFILLER_2_164 VPWR VGND sg13g2_decap_4
XFILLER_39_809 VPWR VGND sg13g2_decap_8
XFILLER_47_842 VPWR VGND sg13g2_decap_8
XFILLER_19_511 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_19_588 VPWR VGND sg13g2_decap_8
XFILLER_22_709 VPWR VGND sg13g2_decap_8
XFILLER_34_547 VPWR VGND sg13g2_decap_8
XFILLER_42_591 VPWR VGND sg13g2_decap_8
XFILLER_14_282 VPWR VGND sg13g2_decap_8
XFILLER_15_783 VPWR VGND sg13g2_decap_8
XFILLER_30_786 VPWR VGND sg13g2_decap_8
XFILLER_7_982 VPWR VGND sg13g2_decap_8
XFILLER_36_0 VPWR VGND sg13g2_decap_8
XFILLER_38_831 VPWR VGND sg13g2_decap_8
XFILLER_25_503 VPWR VGND sg13g2_decap_8
XFILLER_37_363 VPWR VGND sg13g2_decap_8
XFILLER_21_764 VPWR VGND sg13g2_decap_8
XFILLER_20_252 VPWR VGND sg13g2_decap_8
XFILLER_0_602 VPWR VGND sg13g2_decap_8
XFILLER_0_679 VPWR VGND sg13g2_decap_8
XFILLER_48_639 VPWR VGND sg13g2_decap_8
XFILLER_28_330 VPWR VGND sg13g2_decap_8
XFILLER_44_801 VPWR VGND sg13g2_decap_8
XFILLER_29_875 VPWR VGND sg13g2_decap_8
XFILLER_28_385 VPWR VGND sg13g2_decap_8
XFILLER_44_878 VPWR VGND sg13g2_decap_8
XFILLER_43_366 VPWR VGND sg13g2_decap_8
XFILLER_34_62 VPWR VGND sg13g2_decap_8
XFILLER_11_230 VPWR VGND sg13g2_decap_8
XFILLER_15_1028 VPWR VGND sg13g2_fill_1
XFILLER_7_223 VPWR VGND sg13g2_decap_8
XFILLER_12_775 VPWR VGND sg13g2_decap_8
XFILLER_8_768 VPWR VGND sg13g2_decap_8
XFILLER_4_930 VPWR VGND sg13g2_decap_8
XFILLER_3_440 VPWR VGND sg13g2_decap_8
XFILLER_39_606 VPWR VGND sg13g2_decap_8
XFILLER_35_834 VPWR VGND sg13g2_decap_8
XFILLER_22_506 VPWR VGND sg13g2_fill_1
XFILLER_30_583 VPWR VGND sg13g2_decap_8
XFILLER_26_845 VPWR VGND sg13g2_decap_8
XFILLER_13_506 VPWR VGND sg13g2_decap_8
XFILLER_38_1006 VPWR VGND sg13g2_decap_8
XFILLER_40_358 VPWR VGND sg13g2_decap_4
XFILLER_4_204 VPWR VGND sg13g2_decap_8
XFILLER_20_53 VPWR VGND sg13g2_decap_8
XFILLER_1_955 VPWR VGND sg13g2_decap_8
XFILLER_49_937 VPWR VGND sg13g2_decap_8
XFILLER_48_436 VPWR VGND sg13g2_decap_8
Xhold40 DP_4.matrix\[49\] VPWR VGND net90 sg13g2_dlygate4sd3_1
XFILLER_0_476 VPWR VGND sg13g2_decap_8
Xhold73 DP_2.matrix\[32\] VPWR VGND net123 sg13g2_dlygate4sd3_1
XFILLER_29_73 VPWR VGND sg13g2_decap_8
Xhold62 _021_ VPWR VGND net112 sg13g2_dlygate4sd3_1
Xhold51 DP_1.matrix\[65\] VPWR VGND net101 sg13g2_dlygate4sd3_1
XFILLER_29_672 VPWR VGND sg13g2_decap_8
Xhold84 DP_4.matrix\[64\] VPWR VGND net134 sg13g2_dlygate4sd3_1
Xhold95 DP_4.matrix\[48\] VPWR VGND net145 sg13g2_dlygate4sd3_1
XFILLER_17_845 VPWR VGND sg13g2_decap_8
XFILLER_44_675 VPWR VGND sg13g2_decap_8
X_595_ net56 VGND VPWR net108 mac2.total_sum\[0\] clknet_5_5__leaf_clk sg13g2_dfrbpq_1
XFILLER_16_344 VPWR VGND sg13g2_decap_8
XFILLER_43_185 VPWR VGND sg13g2_decap_8
XFILLER_32_848 VPWR VGND sg13g2_decap_8
XFILLER_12_550 VPWR VGND sg13g2_decap_8
XFILLER_6_11 VPWR VGND sg13g2_decap_4
XFILLER_6_44 VPWR VGND sg13g2_fill_2
XFILLER_6_88 VPWR VGND sg13g2_decap_8
XFILLER_3_292 VPWR VGND sg13g2_decap_8
XFILLER_27_609 VPWR VGND sg13g2_decap_8
XFILLER_35_631 VPWR VGND sg13g2_decap_8
XFILLER_22_358 VPWR VGND sg13g2_decap_8
XFILLER_23_859 VPWR VGND sg13g2_decap_8
XFILLER_34_196 VPWR VGND sg13g2_decap_8
XFILLER_46_918 VPWR VGND sg13g2_decap_8
XFILLER_18_609 VPWR VGND sg13g2_fill_1
Xheichips25_template_20 VPWR VGND uio_oe[3] sg13g2_tiehi
XFILLER_39_970 VPWR VGND sg13g2_decap_8
XFILLER_26_642 VPWR VGND sg13g2_decap_8
X_380_ net160 _074_ VPWR VGND sg13g2_buf_1
XFILLER_13_303 VPWR VGND sg13g2_decap_8
XFILLER_25_174 VPWR VGND sg13g2_decap_8
XFILLER_13_347 VPWR VGND sg13g2_decap_8
XFILLER_15_53 VPWR VGND sg13g2_decap_8
XFILLER_41_667 VPWR VGND sg13g2_decap_8
XFILLER_9_329 VPWR VGND sg13g2_decap_8
XFILLER_22_870 VPWR VGND sg13g2_decap_8
XFILLER_40_188 VPWR VGND sg13g2_decap_8
XFILLER_5_513 VPWR VGND sg13g2_fill_2
XFILLER_31_63 VPWR VGND sg13g2_decap_8
XFILLER_5_568 VPWR VGND sg13g2_decap_8
XFILLER_1_752 VPWR VGND sg13g2_decap_8
XFILLER_49_734 VPWR VGND sg13g2_decap_8
XFILLER_0_273 VPWR VGND sg13g2_decap_8
XFILLER_48_288 VPWR VGND sg13g2_decap_8
XFILLER_45_962 VPWR VGND sg13g2_decap_8
XFILLER_16_130 VPWR VGND sg13g2_decap_8
XFILLER_17_642 VPWR VGND sg13g2_decap_8
XFILLER_44_472 VPWR VGND sg13g2_decap_8
X_578_ net58 VGND VPWR net32 mac2.sum_lvl1_ff\[33\] clknet_5_1__leaf_clk sg13g2_dfrbpq_1
XFILLER_16_196 VPWR VGND sg13g2_decap_8
XFILLER_32_645 VPWR VGND sg13g2_decap_8
XFILLER_9_863 VPWR VGND sg13g2_decap_8
XFILLER_8_373 VPWR VGND sg13g2_decap_8
XFILLER_28_1016 VPWR VGND sg13g2_decap_8
XFILLER_28_1027 VPWR VGND sg13g2_fill_2
.ends

